magic
tech sky130A
magscale 1 2
timestamp 1668718364
<< nmos >>
rect -505 -6917 -385 6917
rect -327 -6917 -207 6917
rect -149 -6917 -29 6917
rect 29 -6917 149 6917
rect 207 -6917 327 6917
rect 385 -6917 505 6917
<< ndiff >>
rect -563 6905 -505 6917
rect -563 -6905 -551 6905
rect -517 -6905 -505 6905
rect -563 -6917 -505 -6905
rect -385 6905 -327 6917
rect -385 -6905 -373 6905
rect -339 -6905 -327 6905
rect -385 -6917 -327 -6905
rect -207 6905 -149 6917
rect -207 -6905 -195 6905
rect -161 -6905 -149 6905
rect -207 -6917 -149 -6905
rect -29 6905 29 6917
rect -29 -6905 -17 6905
rect 17 -6905 29 6905
rect -29 -6917 29 -6905
rect 149 6905 207 6917
rect 149 -6905 161 6905
rect 195 -6905 207 6905
rect 149 -6917 207 -6905
rect 327 6905 385 6917
rect 327 -6905 339 6905
rect 373 -6905 385 6905
rect 327 -6917 385 -6905
rect 505 6905 563 6917
rect 505 -6905 517 6905
rect 551 -6905 563 6905
rect 505 -6917 563 -6905
<< ndiffc >>
rect -551 -6905 -517 6905
rect -373 -6905 -339 6905
rect -195 -6905 -161 6905
rect -17 -6905 17 6905
rect 161 -6905 195 6905
rect 339 -6905 373 6905
rect 517 -6905 551 6905
<< poly >>
rect -505 6917 -385 7005
rect -327 6995 -207 7005
rect -149 6995 -29 7005
rect -327 6949 -29 6995
rect -327 6917 -207 6949
rect -149 6917 -29 6949
rect 29 6995 149 7005
rect 207 6995 327 7005
rect 29 6949 327 6995
rect 29 6917 149 6949
rect 207 6917 327 6949
rect 385 6917 505 7005
rect -505 -6949 -385 -6917
rect -327 -6949 -207 -6917
rect -505 -6995 -207 -6949
rect -505 -7005 -385 -6995
rect -327 -7005 -207 -6995
rect -149 -6949 -29 -6917
rect 29 -6949 149 -6917
rect -149 -6995 149 -6949
rect -149 -7005 -29 -6995
rect 29 -7005 149 -6995
rect 207 -6949 327 -6917
rect 385 -6949 505 -6917
rect 207 -6995 505 -6949
rect 207 -7005 327 -6995
rect 385 -7005 505 -6995
<< locali >>
rect -551 6905 -517 6921
rect -551 -6921 -517 -6905
rect -373 6905 -339 6921
rect -373 -6921 -339 -6905
rect -195 6905 -161 6921
rect -195 -6921 -161 -6905
rect -17 6905 17 6921
rect -17 -6921 17 -6905
rect 161 6905 195 6921
rect 161 -6921 195 -6905
rect 339 6905 373 6921
rect 339 -6921 373 -6905
rect 517 6905 551 6921
rect 517 -6921 551 -6905
<< viali >>
rect -551 -6905 -517 6905
rect -373 -6905 -339 6905
rect -195 -6905 -161 6905
rect -17 -6905 17 6905
rect 161 -6905 195 6905
rect 339 -6905 373 6905
rect 517 -6905 551 6905
<< metal1 >>
rect -557 6905 -511 6917
rect -557 -6905 -551 6905
rect -517 -6905 -511 6905
rect -557 -6917 -511 -6905
rect -379 6905 -333 6917
rect -379 -6905 -373 6905
rect -339 -6905 -333 6905
rect -379 -6917 -333 -6905
rect -201 6905 -155 6917
rect -201 -6905 -195 6905
rect -161 -6905 -155 6905
rect -201 -6917 -155 -6905
rect -23 6905 23 6917
rect -23 -6905 -17 6905
rect 17 -6905 23 6905
rect -23 -6917 23 -6905
rect 155 6905 201 6917
rect 155 -6905 161 6905
rect 195 -6905 201 6905
rect 155 -6917 201 -6905
rect 333 6905 379 6917
rect 333 -6905 339 6905
rect 373 -6905 379 6905
rect 333 -6917 379 -6905
rect 511 6905 557 6917
rect 511 -6905 517 6905
rect 551 -6905 557 6905
rect 511 -6917 557 -6905
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 69.17 l 0.6 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
