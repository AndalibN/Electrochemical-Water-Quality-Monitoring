magic
tech sky130A
magscale 1 2
timestamp 1662641497
<< error_p >>
rect -31 -186 31 -180
rect -31 -220 -19 -186
rect -31 -226 31 -220
<< nwell >>
rect -129 -239 129 273
<< pmos >>
rect -35 -139 35 211
<< pdiff >>
rect -93 199 -35 211
rect -93 -127 -81 199
rect -47 -127 -35 199
rect -93 -139 -35 -127
rect 35 199 93 211
rect 35 -127 47 199
rect 81 -127 93 199
rect 35 -139 93 -127
<< pdiffc >>
rect -81 -127 -47 199
rect 47 -127 81 199
<< poly >>
rect -35 211 35 237
rect -35 -186 35 -139
rect -35 -220 -19 -186
rect 19 -220 35 -186
rect -35 -236 35 -220
<< polycont >>
rect -19 -220 19 -186
<< locali >>
rect -81 199 -47 215
rect -81 -143 -47 -127
rect 47 199 81 215
rect 47 -143 81 -127
rect -35 -220 -19 -186
rect 19 -220 35 -186
<< viali >>
rect -81 -127 -47 199
rect 47 -127 81 199
rect -19 -220 19 -186
<< metal1 >>
rect -87 199 -41 211
rect -87 -127 -81 199
rect -47 -127 -41 199
rect -87 -139 -41 -127
rect 41 199 87 211
rect 41 -127 47 199
rect 81 -127 87 199
rect 41 -139 87 -127
rect -31 -186 31 -180
rect -31 -220 -19 -186
rect 19 -220 31 -186
rect -31 -226 31 -220
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.75 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
