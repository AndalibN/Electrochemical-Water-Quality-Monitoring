magic
tech sky130A
magscale 1 2
timestamp 1665000004
<< checkpaint >>
rect 460 5580 4552 11338
rect 6355 -1349 9667 4409
<< error_s >>
rect 468 6497 503 6531
rect 469 6478 503 6497
rect 488 583 503 6478
rect 522 6444 557 6478
rect 522 583 556 6444
rect 4841 4526 4876 4560
rect 4842 4507 4876 4526
rect 1008 2825 1042 2879
rect 522 549 537 583
rect 1027 530 1042 2825
rect 1061 2791 1096 2825
rect 1061 530 1095 2791
rect 1061 496 1076 530
rect 4861 212 4876 4507
rect 4895 4473 4930 4507
rect 5580 4473 5615 4507
rect 4895 212 4929 4473
rect 5581 4454 5615 4473
rect 4895 178 4910 212
rect 5600 159 5615 4454
rect 5634 4420 5669 4454
rect 6319 4420 6354 4454
rect 5634 159 5668 4420
rect 6320 4401 6354 4420
rect 5634 125 5649 159
rect 6339 106 6354 4401
rect 6373 4367 6408 4401
rect 6373 106 6407 4367
rect 7059 2348 7093 2402
rect 6373 72 6388 106
rect 7078 53 7093 2348
rect 7112 2314 7147 2348
rect 7112 53 7146 2314
rect 7112 19 7127 53
use sky130_fd_pr__nfet_01v8_U7E5KL  XM1
timestamp 1664506894
transform 1 0 243 0 1 3557
box -296 -3010 296 3010
use sky130_fd_pr__nfet_01v8_U7E5KL  XM2
timestamp 1664506894
transform 1 0 782 0 1 3504
box -296 -3010 296 3010
use sky130_fd_pr__nfet_01v8_6WXQK8  XM3
timestamp 1664506894
transform 1 0 1321 0 1 1651
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_9QH3CS  XM4
timestamp 1664506894
transform 1 0 2116 0 1 8459
box -396 -1619 396 1619
use sky130_fd_pr__pfet_01v8_9QH3CS  XM5
timestamp 1664506894
transform 1 0 2896 0 1 8459
box -396 -1619 396 1619
use sky130_fd_pr__pfet_01v8_GGN3CJ  XM6
timestamp 1664506894
transform 1 0 3576 0 1 8459
box -296 -1619 296 1619
use sky130_fd_pr__pfet_01v8_GGN3CJ  XM7
timestamp 1664506894
transform 1 0 4156 0 1 8459
box -296 -1619 296 1619
use sky130_fd_pr__nfet_01v8_L9BG78  XM8
timestamp 1664506894
transform 1 0 4516 0 1 2386
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM9
timestamp 1664506894
transform 1 0 5255 0 1 2333
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM10
timestamp 1664506894
transform 1 0 5994 0 1 2280
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM11
timestamp 1664506894
transform 1 0 6733 0 1 2227
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_6WXQK8  XMB1
timestamp 1664506894
transform 1 0 7372 0 1 1174
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_9QH3CS  XMbias
timestamp 1664506894
transform 1 0 8011 0 1 1530
box -396 -1619 396 1619
<< end >>
