magic
tech sky130A
timestamp 1668017718
<< nmos >>
rect -15 -300 15 300
<< ndiff >>
rect -44 294 -15 300
rect -44 -294 -38 294
rect -21 -294 -15 294
rect -44 -300 -15 -294
rect 15 294 44 300
rect 15 -294 21 294
rect 38 -294 44 294
rect 15 -300 44 -294
<< ndiffc >>
rect -38 -294 -21 294
rect 21 -294 38 294
<< poly >>
rect -15 300 15 313
rect -15 -313 15 -300
<< locali >>
rect -38 294 -21 302
rect -38 -302 -21 -294
rect 21 294 38 302
rect 21 -302 38 -294
<< viali >>
rect -38 -294 -21 294
rect 21 -294 38 294
<< metal1 >>
rect -41 294 -18 300
rect -41 -294 -38 294
rect -21 -294 -18 294
rect -41 -300 -18 -294
rect 18 294 41 300
rect 18 -294 21 294
rect 38 -294 41 294
rect 18 -300 41 -294
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
