magic
tech sky130A
magscale 1 2
timestamp 1667324328
<< error_p >>
rect -95 1627 -33 1633
rect -95 1593 -83 1627
rect -95 1587 -33 1593
<< nmoslvt >>
rect -99 -1555 -29 1555
rect 29 -1555 99 1555
<< ndiff >>
rect -157 1543 -99 1555
rect -157 -1543 -145 1543
rect -111 -1543 -99 1543
rect -157 -1555 -99 -1543
rect -29 1543 29 1555
rect -29 -1543 -17 1543
rect 17 -1543 29 1543
rect -29 -1555 29 -1543
rect 99 1543 157 1555
rect 99 -1543 111 1543
rect 145 -1543 157 1543
rect 99 -1555 157 -1543
<< ndiffc >>
rect -145 -1543 -111 1543
rect -17 -1543 17 1543
rect 111 -1543 145 1543
<< poly >>
rect -99 1627 -29 1643
rect -99 1593 -83 1627
rect -45 1593 -29 1627
rect -99 1555 -29 1593
rect 29 1555 99 1585
rect -99 -1578 -29 -1555
rect 29 -1578 99 -1555
rect -99 -1648 99 -1578
<< polycont >>
rect -83 1593 -45 1627
<< locali >>
rect -99 1593 -83 1627
rect -45 1593 -29 1627
rect -145 1543 -111 1559
rect -145 -1559 -111 -1543
rect -17 1543 17 1559
rect -17 -1559 17 -1543
rect 111 1543 145 1559
rect 111 -1559 145 -1543
<< viali >>
rect -83 1593 -45 1627
rect -145 -1543 -111 1543
rect -17 -1543 17 1543
rect 111 -1543 145 1543
<< metal1 >>
rect -95 1627 -33 1633
rect -95 1593 -83 1627
rect -45 1593 -33 1627
rect -95 1587 -33 1593
rect -151 1543 -105 1555
rect -151 -1543 -145 1543
rect -111 -1543 -105 1543
rect -151 -1555 -105 -1543
rect -23 1543 23 1555
rect -23 -1543 -17 1543
rect 17 -1543 23 1543
rect -23 -1555 23 -1543
rect 105 1543 151 1555
rect 105 -1543 111 1543
rect 145 -1543 151 1543
rect 105 -1555 151 -1543
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 15.55 l 0.35 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
