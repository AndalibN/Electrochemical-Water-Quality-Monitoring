magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -1123 -298 1123 264
<< pmos >>
rect -1029 -236 -29 164
rect 29 -236 1029 164
<< pdiff >>
rect -1087 151 -1029 164
rect -1087 117 -1075 151
rect -1041 117 -1029 151
rect -1087 83 -1029 117
rect -1087 49 -1075 83
rect -1041 49 -1029 83
rect -1087 15 -1029 49
rect -1087 -19 -1075 15
rect -1041 -19 -1029 15
rect -1087 -53 -1029 -19
rect -1087 -87 -1075 -53
rect -1041 -87 -1029 -53
rect -1087 -121 -1029 -87
rect -1087 -155 -1075 -121
rect -1041 -155 -1029 -121
rect -1087 -189 -1029 -155
rect -1087 -223 -1075 -189
rect -1041 -223 -1029 -189
rect -1087 -236 -1029 -223
rect -29 151 29 164
rect -29 117 -17 151
rect 17 117 29 151
rect -29 83 29 117
rect -29 49 -17 83
rect 17 49 29 83
rect -29 15 29 49
rect -29 -19 -17 15
rect 17 -19 29 15
rect -29 -53 29 -19
rect -29 -87 -17 -53
rect 17 -87 29 -53
rect -29 -121 29 -87
rect -29 -155 -17 -121
rect 17 -155 29 -121
rect -29 -189 29 -155
rect -29 -223 -17 -189
rect 17 -223 29 -189
rect -29 -236 29 -223
rect 1029 151 1087 164
rect 1029 117 1041 151
rect 1075 117 1087 151
rect 1029 83 1087 117
rect 1029 49 1041 83
rect 1075 49 1087 83
rect 1029 15 1087 49
rect 1029 -19 1041 15
rect 1075 -19 1087 15
rect 1029 -53 1087 -19
rect 1029 -87 1041 -53
rect 1075 -87 1087 -53
rect 1029 -121 1087 -87
rect 1029 -155 1041 -121
rect 1075 -155 1087 -121
rect 1029 -189 1087 -155
rect 1029 -223 1041 -189
rect 1075 -223 1087 -189
rect 1029 -236 1087 -223
<< pdiffc >>
rect -1075 117 -1041 151
rect -1075 49 -1041 83
rect -1075 -19 -1041 15
rect -1075 -87 -1041 -53
rect -1075 -155 -1041 -121
rect -1075 -223 -1041 -189
rect -17 117 17 151
rect -17 49 17 83
rect -17 -19 17 15
rect -17 -87 17 -53
rect -17 -155 17 -121
rect -17 -223 17 -189
rect 1041 117 1075 151
rect 1041 49 1075 83
rect 1041 -19 1075 15
rect 1041 -87 1075 -53
rect 1041 -155 1075 -121
rect 1041 -223 1075 -189
<< poly >>
rect -1029 245 -29 261
rect -1029 211 -988 245
rect -954 211 -920 245
rect -886 211 -852 245
rect -818 211 -784 245
rect -750 211 -716 245
rect -682 211 -648 245
rect -614 211 -580 245
rect -546 211 -512 245
rect -478 211 -444 245
rect -410 211 -376 245
rect -342 211 -308 245
rect -274 211 -240 245
rect -206 211 -172 245
rect -138 211 -104 245
rect -70 211 -29 245
rect -1029 164 -29 211
rect 29 245 1029 261
rect 29 211 70 245
rect 104 211 138 245
rect 172 211 206 245
rect 240 211 274 245
rect 308 211 342 245
rect 376 211 410 245
rect 444 211 478 245
rect 512 211 546 245
rect 580 211 614 245
rect 648 211 682 245
rect 716 211 750 245
rect 784 211 818 245
rect 852 211 886 245
rect 920 211 954 245
rect 988 211 1029 245
rect 29 164 1029 211
rect -1029 -262 -29 -236
rect 29 -262 1029 -236
<< polycont >>
rect -988 211 -954 245
rect -920 211 -886 245
rect -852 211 -818 245
rect -784 211 -750 245
rect -716 211 -682 245
rect -648 211 -614 245
rect -580 211 -546 245
rect -512 211 -478 245
rect -444 211 -410 245
rect -376 211 -342 245
rect -308 211 -274 245
rect -240 211 -206 245
rect -172 211 -138 245
rect -104 211 -70 245
rect 70 211 104 245
rect 138 211 172 245
rect 206 211 240 245
rect 274 211 308 245
rect 342 211 376 245
rect 410 211 444 245
rect 478 211 512 245
rect 546 211 580 245
rect 614 211 648 245
rect 682 211 716 245
rect 750 211 784 245
rect 818 211 852 245
rect 886 211 920 245
rect 954 211 988 245
<< locali >>
rect -1029 211 -988 245
rect -944 211 -920 245
rect -872 211 -852 245
rect -800 211 -784 245
rect -728 211 -716 245
rect -656 211 -648 245
rect -584 211 -580 245
rect -478 211 -474 245
rect -410 211 -402 245
rect -342 211 -330 245
rect -274 211 -258 245
rect -206 211 -186 245
rect -138 211 -114 245
rect -70 211 -29 245
rect 29 211 70 245
rect 114 211 138 245
rect 186 211 206 245
rect 258 211 274 245
rect 330 211 342 245
rect 402 211 410 245
rect 474 211 478 245
rect 580 211 584 245
rect 648 211 656 245
rect 716 211 728 245
rect 784 211 800 245
rect 852 211 872 245
rect 920 211 944 245
rect 988 211 1029 245
rect -1075 151 -1041 168
rect -1075 83 -1041 91
rect -1075 15 -1041 19
rect -1075 -91 -1041 -87
rect -1075 -163 -1041 -155
rect -1075 -240 -1041 -223
rect -17 151 17 168
rect -17 83 17 91
rect -17 15 17 19
rect -17 -91 17 -87
rect -17 -163 17 -155
rect -17 -240 17 -223
rect 1041 151 1075 168
rect 1041 83 1075 91
rect 1041 15 1075 19
rect 1041 -91 1075 -87
rect 1041 -163 1075 -155
rect 1041 -240 1075 -223
<< viali >>
rect -978 211 -954 245
rect -954 211 -944 245
rect -906 211 -886 245
rect -886 211 -872 245
rect -834 211 -818 245
rect -818 211 -800 245
rect -762 211 -750 245
rect -750 211 -728 245
rect -690 211 -682 245
rect -682 211 -656 245
rect -618 211 -614 245
rect -614 211 -584 245
rect -546 211 -512 245
rect -474 211 -444 245
rect -444 211 -440 245
rect -402 211 -376 245
rect -376 211 -368 245
rect -330 211 -308 245
rect -308 211 -296 245
rect -258 211 -240 245
rect -240 211 -224 245
rect -186 211 -172 245
rect -172 211 -152 245
rect -114 211 -104 245
rect -104 211 -80 245
rect 80 211 104 245
rect 104 211 114 245
rect 152 211 172 245
rect 172 211 186 245
rect 224 211 240 245
rect 240 211 258 245
rect 296 211 308 245
rect 308 211 330 245
rect 368 211 376 245
rect 376 211 402 245
rect 440 211 444 245
rect 444 211 474 245
rect 512 211 546 245
rect 584 211 614 245
rect 614 211 618 245
rect 656 211 682 245
rect 682 211 690 245
rect 728 211 750 245
rect 750 211 762 245
rect 800 211 818 245
rect 818 211 834 245
rect 872 211 886 245
rect 886 211 906 245
rect 944 211 954 245
rect 954 211 978 245
rect -1075 117 -1041 125
rect -1075 91 -1041 117
rect -1075 49 -1041 53
rect -1075 19 -1041 49
rect -1075 -53 -1041 -19
rect -1075 -121 -1041 -91
rect -1075 -125 -1041 -121
rect -1075 -189 -1041 -163
rect -1075 -197 -1041 -189
rect -17 117 17 125
rect -17 91 17 117
rect -17 49 17 53
rect -17 19 17 49
rect -17 -53 17 -19
rect -17 -121 17 -91
rect -17 -125 17 -121
rect -17 -189 17 -163
rect -17 -197 17 -189
rect 1041 117 1075 125
rect 1041 91 1075 117
rect 1041 49 1075 53
rect 1041 19 1075 49
rect 1041 -53 1075 -19
rect 1041 -121 1075 -91
rect 1041 -125 1075 -121
rect 1041 -189 1075 -163
rect 1041 -197 1075 -189
<< metal1 >>
rect -1025 245 -33 251
rect -1025 211 -978 245
rect -944 211 -906 245
rect -872 211 -834 245
rect -800 211 -762 245
rect -728 211 -690 245
rect -656 211 -618 245
rect -584 211 -546 245
rect -512 211 -474 245
rect -440 211 -402 245
rect -368 211 -330 245
rect -296 211 -258 245
rect -224 211 -186 245
rect -152 211 -114 245
rect -80 211 -33 245
rect -1025 205 -33 211
rect 33 245 1025 251
rect 33 211 80 245
rect 114 211 152 245
rect 186 211 224 245
rect 258 211 296 245
rect 330 211 368 245
rect 402 211 440 245
rect 474 211 512 245
rect 546 211 584 245
rect 618 211 656 245
rect 690 211 728 245
rect 762 211 800 245
rect 834 211 872 245
rect 906 211 944 245
rect 978 211 1025 245
rect 33 205 1025 211
rect -1081 125 -1035 164
rect -1081 91 -1075 125
rect -1041 91 -1035 125
rect -1081 53 -1035 91
rect -1081 19 -1075 53
rect -1041 19 -1035 53
rect -1081 -19 -1035 19
rect -1081 -53 -1075 -19
rect -1041 -53 -1035 -19
rect -1081 -91 -1035 -53
rect -1081 -125 -1075 -91
rect -1041 -125 -1035 -91
rect -1081 -163 -1035 -125
rect -1081 -197 -1075 -163
rect -1041 -197 -1035 -163
rect -1081 -236 -1035 -197
rect -23 125 23 164
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -236 23 -197
rect 1035 125 1081 164
rect 1035 91 1041 125
rect 1075 91 1081 125
rect 1035 53 1081 91
rect 1035 19 1041 53
rect 1075 19 1081 53
rect 1035 -19 1081 19
rect 1035 -53 1041 -19
rect 1075 -53 1081 -19
rect 1035 -91 1081 -53
rect 1035 -125 1041 -91
rect 1075 -125 1081 -91
rect 1035 -163 1081 -125
rect 1035 -197 1041 -163
rect 1075 -197 1081 -163
rect 1035 -236 1081 -197
<< end >>
