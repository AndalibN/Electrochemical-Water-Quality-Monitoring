magic
tech sky130A
magscale 1 2
timestamp 1668221056
<< nwell >>
rect -2498 1724 1462 2367
rect -2498 -716 1465 1724
<< psubdiff >>
rect -2704 -3426 -2680 -2511
rect 2131 -3426 2155 -2511
<< nsubdiff >>
rect -2383 2156 1387 2229
rect -2383 2155 -985 2156
rect -2383 2154 -1423 2155
rect -1347 2154 -985 2155
rect -909 2154 1387 2156
rect -2383 1995 -2253 2154
rect 1292 1995 1387 2154
rect -2383 1895 1387 1995
<< psubdiffcont >>
rect -2680 -3426 2131 -2511
<< nsubdiffcont >>
rect -1423 2154 -1347 2155
rect -985 2154 -909 2156
rect -2253 1995 1292 2154
<< poly >>
rect -2633 1846 -2563 1880
rect -2633 1816 -982 1846
rect -2633 1814 -2563 1816
rect -2630 1742 -1304 1772
rect -2630 1701 -2560 1742
rect -1348 1640 -1304 1742
rect -1012 1549 -982 1816
rect -607 1742 -527 1746
rect -607 1729 731 1742
rect -607 1693 -587 1729
rect -545 1693 731 1729
rect -607 1685 731 1693
rect -607 1676 -527 1685
rect -250 1615 -170 1628
rect -250 1611 482 1615
rect -250 1608 -230 1611
rect -535 1575 -230 1608
rect -188 1575 482 1611
rect 670 1586 731 1685
rect -535 1566 482 1575
rect -535 1506 -475 1566
rect -417 1506 -357 1566
rect -250 1558 -170 1566
rect 422 1436 482 1566
rect -653 -508 -593 -460
rect -299 -508 -239 -460
rect 40 -508 364 -507
rect -653 -548 364 -508
rect 899 -597 1083 -550
rect -289 -1053 1169 -1023
rect -289 -1147 -250 -1053
rect 499 -1159 557 -1053
rect 1113 -1156 1169 -1053
rect -2462 -1300 -2285 -1253
rect -1358 -1863 -1065 -1807
rect -534 -1874 -472 -1813
rect 115 -1874 175 -1809
rect -534 -1922 175 -1874
rect 116 -1935 175 -1922
rect 883 -1886 926 -1820
rect 116 -1979 883 -1935
<< polycont >>
rect -587 1693 -545 1729
rect -230 1575 -188 1611
<< rmp >>
rect 883 -1979 926 -1886
<< locali >>
rect -2310 2156 1335 2190
rect -2310 2155 -985 2156
rect -2310 2154 -1423 2155
rect -1347 2154 -985 2155
rect -909 2154 1335 2156
rect -2310 1995 -2253 2154
rect 1292 1995 1335 2154
rect -2310 1948 1335 1995
rect -2630 1870 -2572 1878
rect -2630 1834 -2616 1870
rect -2582 1834 -2572 1870
rect -2630 1822 -2572 1834
rect -2626 1754 -2576 1762
rect -2626 1720 -2614 1754
rect -2580 1720 -2576 1754
rect -2626 1708 -2576 1720
rect -607 1729 -527 1746
rect -607 1693 -587 1729
rect -545 1693 -527 1729
rect -607 1676 -527 1693
rect -250 1611 -170 1628
rect -2186 1531 -1944 1585
rect -250 1575 -230 1611
rect -188 1575 -170 1611
rect -250 1558 -170 1575
rect -2002 -818 -1944 1531
rect -1342 -566 -1308 -483
rect 258 -566 292 1419
rect -1342 -600 292 -566
rect 258 -708 292 -600
rect 818 -514 888 44
rect 1092 -513 1163 29
rect 818 -610 864 -514
rect 812 -625 864 -610
rect 812 -626 872 -625
rect 812 -660 824 -626
rect 858 -660 872 -626
rect 812 -668 872 -660
rect 812 -673 864 -668
rect 915 -708 949 -557
rect 1117 -614 1163 -513
rect 1116 -628 1170 -614
rect 1116 -662 1124 -628
rect 1158 -662 1170 -628
rect 1116 -674 1170 -662
rect 258 -742 949 -708
rect -2003 -822 -1944 -818
rect -2003 -867 -1998 -822
rect -1949 -836 -1944 -822
rect -1949 -867 44 -836
rect -2003 -870 44 -867
rect -2003 -872 -1944 -870
rect 9 -988 44 -870
rect 9 -1018 427 -988
rect 10 -1022 427 -1018
rect 10 -1146 44 -1022
rect 393 -1153 427 -1022
rect -1171 -1894 -1137 -1197
rect -935 -1755 -901 -1165
rect -960 -1789 -901 -1755
rect -699 -1750 -665 -1181
rect 794 -1184 836 -742
rect 934 -823 992 -809
rect 934 -857 946 -823
rect 980 -857 992 -823
rect 934 -870 992 -857
rect -699 -1789 -640 -1750
rect -227 -1771 -193 -1195
rect 794 -1467 863 -1184
rect 940 -1329 986 -870
rect 1117 -914 1163 -674
rect 1117 -960 1378 -914
rect 1332 -1130 1378 -960
rect 1332 -1264 1414 -1130
rect -960 -1894 -926 -1789
rect -674 -1894 -640 -1789
rect -1171 -1928 -640 -1894
rect -2696 -3426 -2680 -2511
rect 2131 -3426 2147 -2511
<< viali >>
rect -1712 2065 -1667 2107
rect -1525 2094 -1480 2136
rect -1408 2101 -1363 2143
rect -970 2102 -925 2144
rect -468 2088 -423 2130
rect 123 2089 168 2131
rect 478 2091 523 2133
rect 598 2089 643 2131
rect 959 2089 1004 2131
rect 1224 2086 1269 2128
rect -1965 2016 -1920 2058
rect -2616 1834 -2582 1870
rect -2614 1720 -2580 1754
rect -587 1693 -545 1729
rect -230 1575 -188 1611
rect 824 -660 858 -626
rect 1124 -662 1158 -628
rect -1998 -867 -1949 -822
rect 946 -857 980 -823
rect -2397 -2835 -2352 -2793
rect -1866 -2834 -1821 -2792
rect -2524 -2880 -2479 -2838
rect -1424 -2840 -1379 -2798
rect -1058 -2840 -1013 -2798
rect -239 -2835 -194 -2793
rect 577 -2838 622 -2796
rect 1200 -2831 1245 -2789
rect 1608 -2826 1653 -2784
rect 1877 -2822 1922 -2780
rect -2321 -3103 -2276 -3061
<< metal1 >>
rect 2796 2247 2932 2257
rect 2796 2217 2808 2247
rect 2788 2167 2808 2217
rect -7116 2062 -6916 2141
rect -1539 2136 -1465 2145
rect -1726 2107 -1652 2116
rect -1970 2062 -1906 2072
rect -7116 2058 -1906 2062
rect -7116 2016 -1965 2058
rect -1920 2016 -1906 2058
rect -1726 2065 -1712 2107
rect -1667 2065 -1652 2107
rect -1539 2094 -1525 2136
rect -1480 2094 -1465 2136
rect -1539 2082 -1465 2094
rect -1422 2143 -1348 2152
rect -1422 2101 -1408 2143
rect -1363 2101 -1348 2143
rect -1422 2089 -1348 2101
rect -984 2144 -910 2153
rect -984 2102 -970 2144
rect -925 2102 -910 2144
rect 2796 2147 2808 2167
rect 2920 2222 2932 2247
rect 3877 2246 4005 2254
rect 3877 2222 3887 2246
rect 2920 2166 3887 2222
rect 2920 2147 2932 2166
rect -984 2090 -910 2102
rect -482 2130 -408 2139
rect -1726 2050 -1652 2065
rect -7116 2012 -1906 2016
rect -7116 1941 -6916 2012
rect -1970 2004 -1906 2012
rect -2632 1870 -2570 1880
rect -2632 1834 -2616 1870
rect -2582 1834 -2570 1870
rect -2632 1816 -2570 1834
rect -2632 1754 -2560 1772
rect -2632 1720 -2614 1754
rect -2580 1720 -2560 1754
rect -2632 1700 -2560 1720
rect -7118 1458 -6918 1658
rect -5586 1610 -5458 1618
rect -5586 1580 -5576 1610
rect -5638 1530 -5576 1580
rect -5586 1510 -5576 1530
rect -5464 1580 -5458 1610
rect -3928 1610 -3800 1618
rect -3928 1580 -3918 1610
rect -5464 1530 -3918 1580
rect -5464 1510 -5458 1530
rect -4630 1528 -4586 1530
rect -5586 1502 -5458 1510
rect -3928 1510 -3918 1530
rect -3806 1580 -3800 1610
rect -2190 1583 -2127 1584
rect -2309 1580 -2242 1581
rect -3806 1530 -2242 1580
rect -3806 1510 -3800 1530
rect -3066 1528 -2242 1530
rect -2190 1526 -2126 1583
rect -2189 1525 -2126 1526
rect -3928 1502 -3800 1510
rect -7116 1154 -6916 1354
rect -1702 1322 -1668 2050
rect -1517 1707 -1483 2082
rect -1530 1700 -1467 1707
rect -1530 1648 -1524 1700
rect -1472 1648 -1467 1700
rect -1530 1640 -1467 1648
rect -1401 1345 -1367 2089
rect -962 1493 -928 2090
rect -482 2088 -468 2130
rect -423 2088 -408 2130
rect -482 2076 -408 2088
rect 109 2131 183 2140
rect 109 2089 123 2131
rect 168 2089 183 2131
rect 109 2077 183 2089
rect 464 2133 538 2142
rect 464 2091 478 2133
rect 523 2091 538 2133
rect 464 2079 538 2091
rect 584 2131 658 2140
rect 584 2089 598 2131
rect 643 2089 658 2131
rect -599 1729 -533 1741
rect -599 1693 -587 1729
rect -545 1693 -533 1729
rect -599 1681 -533 1693
rect -888 1527 -665 1561
rect -962 1465 -913 1493
rect -947 1331 -913 1465
rect -5384 243 -5326 251
rect -4972 247 -4878 478
rect -5384 191 -5378 243
rect -5326 226 -5311 243
rect -5326 198 -5309 226
rect -5326 191 -5311 198
rect -5384 183 -5311 191
rect -4972 195 -4958 247
rect -4906 195 -4878 247
rect -5384 182 -5326 183
rect -7116 -573 -6916 -427
rect -7116 -609 -5621 -573
rect -7116 -627 -6916 -609
rect -5685 -616 -5621 -609
rect -5685 -668 -5678 -616
rect -5626 -668 -5621 -616
rect -5685 -677 -5621 -668
rect -5692 -809 -5628 -800
rect -7116 -831 -6916 -827
rect -5692 -831 -5685 -809
rect -7116 -861 -5685 -831
rect -5633 -831 -5628 -809
rect -5633 -861 -5616 -831
rect -7116 -867 -5616 -861
rect -7116 -1027 -6916 -867
rect -5692 -870 -5628 -867
rect -5690 -993 -5626 -984
rect -5887 -1045 -5683 -993
rect -5631 -1045 -5626 -993
rect -5887 -1047 -5626 -1045
rect -7116 -1299 -6916 -1227
rect -5887 -1299 -5839 -1047
rect -5690 -1054 -5626 -1047
rect -5711 -1104 -5615 -1094
rect -5711 -1156 -5684 -1104
rect -5632 -1156 -5615 -1104
rect -5711 -1165 -5615 -1156
rect -7116 -1348 -5839 -1299
rect -7116 -1427 -6916 -1348
rect -7116 -1736 -6916 -1629
rect -5683 -1736 -5643 -1165
rect -7116 -1772 -5643 -1736
rect -7116 -1829 -6916 -1772
rect -7116 -2154 -6916 -2059
rect -5714 -2150 -5650 -2141
rect -5714 -2154 -5707 -2150
rect -7116 -2190 -5707 -2154
rect -7116 -2259 -6916 -2190
rect -5714 -2202 -5707 -2190
rect -5655 -2154 -5650 -2150
rect -5655 -2190 -5637 -2154
rect -5655 -2202 -5650 -2190
rect -5714 -2211 -5650 -2202
rect -5378 -2848 -5326 182
rect -4972 171 -4878 195
rect -3314 261 -3220 573
rect -3314 209 -3292 261
rect -3240 209 -3220 261
rect -3314 182 -3220 209
rect -5268 66 -5140 74
rect -5268 36 -5258 66
rect -5282 -14 -5258 36
rect -5268 -34 -5258 -14
rect -5146 36 -5140 66
rect -3610 66 -3482 74
rect -4716 36 -4644 40
rect -3610 36 -3600 66
rect -5146 -14 -4644 36
rect -3624 -14 -3600 36
rect -5146 -34 -5140 -14
rect -5268 -42 -5140 -34
rect -4982 -876 -4925 -14
rect -3610 -34 -3600 -14
rect -3488 36 -3482 66
rect -3058 36 -2986 68
rect -3488 -14 -2986 36
rect -3488 -34 -3482 -14
rect -3610 -42 -3482 -34
rect -3216 -724 -3145 -14
rect -2369 -41 -2323 -40
rect -2369 -198 -2320 -41
rect -3218 -730 -3145 -724
rect -3218 -782 -3212 -730
rect -3160 -782 -3145 -730
rect -3218 -788 -3145 -782
rect -3215 -791 -3145 -788
rect -2368 -390 -2320 -198
rect -4986 -883 -4915 -876
rect -4988 -889 -4915 -883
rect -4988 -941 -4982 -889
rect -4930 -941 -4915 -889
rect -4988 -947 -4915 -941
rect -4985 -950 -4915 -947
rect -4982 -957 -4925 -950
rect -2519 -1250 -2473 -1249
rect -2519 -1303 -2400 -1250
rect -2368 -1253 -2333 -390
rect -2236 -484 -2202 -264
rect -2237 -491 -2174 -484
rect -2237 -544 -2232 -491
rect -2180 -544 -2174 -491
rect -2237 -550 -2174 -544
rect -2118 -1187 -2083 -130
rect -1866 -395 -1787 0
rect -1283 -377 -1249 -179
rect -1866 -491 -1802 -395
rect -1283 -406 -1236 -377
rect -1774 -483 -1711 -427
rect -1866 -544 -1859 -491
rect -1807 -544 -1802 -491
rect -1866 -550 -1802 -544
rect -1772 -601 -1716 -483
rect -1358 -496 -1292 -434
rect -1264 -524 -1236 -406
rect -1065 -474 -1031 612
rect -829 -474 -795 -145
rect -699 -428 -665 1527
rect -586 1449 -546 1681
rect -1065 -507 -783 -474
rect -1283 -550 -1236 -524
rect -1775 -611 -1711 -601
rect -1775 -664 -1768 -611
rect -1716 -664 -1711 -611
rect -1775 -670 -1711 -664
rect -1283 -729 -1249 -550
rect -1299 -735 -1235 -729
rect -1299 -787 -1293 -735
rect -1241 -787 -1235 -735
rect -1299 -793 -1235 -787
rect -2010 -810 -1938 -809
rect -2012 -813 -1938 -810
rect -2012 -870 -2003 -813
rect -1945 -870 -1938 -813
rect -2012 -879 -1938 -870
rect -2257 -1233 -1694 -1187
rect -2368 -1300 -2285 -1253
rect -2519 -1631 -2473 -1303
rect -2257 -1328 -2225 -1233
rect -2272 -1512 -2225 -1328
rect -2389 -2774 -2361 -1519
rect -1401 -1526 -1367 -1203
rect -1283 -1297 -1249 -793
rect -1053 -1482 -1019 -1197
rect -1861 -1864 -1822 -1526
rect -1861 -2773 -1833 -1864
rect -1668 -1868 -1632 -1678
rect -1664 -1961 -1632 -1868
rect -1414 -1789 -1367 -1526
rect -1665 -1970 -1596 -1961
rect -1665 -2022 -1654 -1970
rect -1602 -2022 -1596 -1970
rect -1665 -2029 -1596 -2022
rect -2413 -2793 -2334 -2774
rect -2540 -2838 -2462 -2819
rect -2540 -2848 -2524 -2838
rect -5378 -2876 -2524 -2848
rect -2540 -2880 -2524 -2876
rect -2479 -2880 -2462 -2838
rect -2413 -2835 -2397 -2793
rect -2352 -2835 -2334 -2793
rect -2413 -2855 -2334 -2835
rect -1882 -2792 -1803 -2773
rect -1414 -2779 -1386 -1789
rect -1283 -1817 -1249 -1643
rect -1358 -1857 -1249 -1817
rect -1358 -1863 -1292 -1857
rect -1054 -2186 -1019 -1482
rect -817 -1773 -783 -507
rect -581 -1771 -547 1449
rect -463 -428 -429 2076
rect -242 1611 -176 1623
rect -242 1575 -230 1611
rect -188 1575 -176 1611
rect -242 1563 -176 1575
rect -227 955 -193 1563
rect -228 -428 -193 955
rect -228 -939 -194 -428
rect -109 -492 -75 497
rect 129 -439 163 2077
rect 494 -477 528 2079
rect 584 2077 658 2089
rect 945 2131 1019 2140
rect 1242 2137 1276 2141
rect 2796 2137 2932 2147
rect 3877 2146 3887 2166
rect 3999 2216 4005 2246
rect 4987 2224 5051 2231
rect 5151 2224 5351 2301
rect 4987 2222 5351 2224
rect 3999 2166 4016 2216
rect 4987 2170 4992 2222
rect 5044 2170 5351 2222
rect 3999 2146 4005 2166
rect 4987 2161 5051 2170
rect 3877 2138 4005 2146
rect 945 2089 959 2131
rect 1004 2089 1019 2131
rect 945 2077 1019 2089
rect 1210 2128 1284 2137
rect 1210 2086 1224 2128
rect 1269 2086 1284 2128
rect 5151 2101 5351 2170
rect 606 -477 637 2077
rect 670 1584 733 1639
rect 974 1405 1008 2077
rect 1210 2074 1284 2086
rect 1242 1551 1276 2074
rect 1229 1544 1292 1551
rect 1229 1492 1235 1544
rect 1287 1492 1292 1544
rect 1229 1484 1292 1492
rect 3262 0 3408 14
rect 3262 -23 3278 0
rect 3261 -70 3278 -23
rect 3262 -100 3278 -70
rect 3390 -15 3408 0
rect 4351 5 4479 13
rect 4351 -15 4357 5
rect 3390 -71 4357 -15
rect 3390 -100 3408 -71
rect 3262 -116 3408 -100
rect 4351 -95 4357 -71
rect 4469 -15 4479 5
rect 4469 -65 4489 -15
rect 4469 -95 4479 -65
rect 4351 -103 4479 -95
rect 2906 -267 3042 -257
rect 2906 -279 2918 -267
rect -109 -538 113 -492
rect 69 -868 104 -538
rect 69 -904 353 -868
rect -228 -972 221 -939
rect -423 -996 -359 -990
rect -423 -1048 -417 -996
rect -365 -1048 -359 -996
rect -423 -1054 -359 -1048
rect 187 -1044 221 -972
rect -404 -1100 -370 -1054
rect 187 -1076 234 -1044
rect -302 -1097 -238 -1091
rect -421 -1155 -353 -1100
rect -302 -1149 -296 -1097
rect -244 -1101 -238 -1097
rect -244 -1111 -237 -1101
rect -244 -1145 -77 -1111
rect -244 -1149 -237 -1145
rect -302 -1154 -237 -1149
rect -6 -1154 59 -1100
rect 203 -1104 234 -1076
rect 114 -1152 234 -1104
rect -302 -1155 -238 -1154
rect 203 -1180 234 -1152
rect 187 -1223 234 -1180
rect 325 -1187 353 -904
rect 737 -974 783 -304
rect 1914 -347 2918 -279
rect 899 -597 965 -543
rect 1018 -597 1084 -543
rect 812 -625 872 -610
rect 1116 -625 1170 -614
rect 812 -626 1170 -625
rect 812 -660 824 -626
rect 858 -628 1170 -626
rect 858 -660 1124 -628
rect 812 -662 1124 -660
rect 1158 -662 1170 -628
rect 812 -668 1170 -662
rect 812 -673 872 -668
rect 1116 -674 1170 -668
rect 1179 -780 1811 -744
rect 934 -821 992 -809
rect 1179 -821 1209 -780
rect 934 -823 1209 -821
rect 934 -857 946 -823
rect 980 -857 1209 -823
rect 934 -870 992 -857
rect 1771 -938 1811 -780
rect 1914 -797 1968 -347
rect 2906 -367 2918 -347
rect 3030 -292 3042 -267
rect 3987 -268 4115 -260
rect 3987 -292 3997 -268
rect 3030 -348 3997 -292
rect 3030 -367 3042 -348
rect 2906 -377 3042 -367
rect 3987 -368 3997 -348
rect 4109 -298 4115 -268
rect 5006 -294 5070 -287
rect 5175 -294 5375 -200
rect 5006 -296 5375 -294
rect 4109 -348 4126 -298
rect 5006 -348 5011 -296
rect 5063 -348 5375 -296
rect 4109 -368 4115 -348
rect 5006 -357 5070 -348
rect 3987 -376 4115 -368
rect 5175 -400 5375 -348
rect 1911 -803 1975 -797
rect 1911 -855 1917 -803
rect 1969 -855 1975 -803
rect 1911 -861 1975 -855
rect 1771 -974 2421 -938
rect 737 -1016 1602 -974
rect 1421 -1050 1490 -1044
rect 1550 -1048 1602 -1016
rect 381 -1161 443 -1104
rect 499 -1161 561 -1104
rect 1112 -1158 1174 -1101
rect 1421 -1102 1430 -1050
rect 1482 -1102 1490 -1050
rect 1421 -1106 1490 -1102
rect 1540 -1104 1860 -1048
rect 1738 -1134 1768 -1104
rect 325 -1215 368 -1187
rect -469 -1725 -422 -1489
rect -469 -1782 -402 -1725
rect -892 -1865 -709 -1815
rect -818 -2038 -784 -1865
rect -538 -1870 -472 -1813
rect -831 -2045 -768 -2038
rect -831 -2097 -825 -2045
rect -773 -2097 -768 -2045
rect -831 -2105 -768 -2097
rect -1054 -2779 -1020 -2186
rect -442 -2389 -402 -1782
rect -452 -2395 -388 -2389
rect -452 -2447 -446 -2395
rect -394 -2447 -388 -2395
rect -452 -2453 -388 -2447
rect -227 -2774 -193 -1527
rect -52 -1964 -14 -1750
rect 187 -1771 221 -1223
rect 334 -1309 368 -1215
rect 570 -1791 620 -1400
rect 1738 -1418 1786 -1134
rect 1182 -1788 1236 -1513
rect 377 -1822 439 -1821
rect 377 -1878 443 -1822
rect 496 -1876 558 -1819
rect -60 -1971 5 -1964
rect -60 -2023 -54 -1971
rect -2 -2023 5 -1971
rect -60 -2030 5 -2023
rect -1882 -2834 -1866 -2792
rect -1821 -2834 -1803 -2792
rect -1882 -2854 -1803 -2834
rect -1440 -2798 -1361 -2779
rect -1440 -2840 -1424 -2798
rect -1379 -2840 -1361 -2798
rect -1440 -2860 -1361 -2840
rect -1074 -2798 -995 -2779
rect -1074 -2840 -1058 -2798
rect -1013 -2840 -995 -2798
rect -1074 -2860 -995 -2840
rect -255 -2793 -176 -2774
rect 586 -2777 620 -1791
rect 874 -1872 936 -1818
rect 992 -1872 1054 -1818
rect 1110 -1870 1172 -1816
rect 994 -2010 1052 -1872
rect 990 -2016 1054 -2010
rect 990 -2068 996 -2016
rect 1048 -2068 1054 -2016
rect 990 -2074 1054 -2068
rect 1202 -2770 1236 -1788
rect 1622 -2765 1656 -1511
rect 1876 -2761 1910 -1511
rect 2381 -2532 2421 -974
rect 3372 -2514 3518 -2498
rect 3372 -2532 3388 -2514
rect 2381 -2583 3388 -2532
rect 3371 -2584 3388 -2583
rect 3372 -2614 3388 -2584
rect 3500 -2529 3518 -2514
rect 4461 -2509 4589 -2501
rect 4461 -2529 4467 -2509
rect 3500 -2585 4467 -2529
rect 3500 -2614 3518 -2585
rect 3372 -2628 3518 -2614
rect 4461 -2609 4467 -2585
rect 4579 -2529 4589 -2509
rect 4579 -2579 4599 -2529
rect 4579 -2609 4589 -2579
rect 4461 -2617 4589 -2609
rect -255 -2835 -239 -2793
rect -194 -2835 -176 -2793
rect -255 -2855 -176 -2835
rect 561 -2796 640 -2777
rect 561 -2838 577 -2796
rect 622 -2838 640 -2796
rect 561 -2858 640 -2838
rect 1184 -2789 1263 -2770
rect 1184 -2831 1200 -2789
rect 1245 -2831 1263 -2789
rect 1184 -2851 1263 -2831
rect 1592 -2784 1671 -2765
rect 1592 -2826 1608 -2784
rect 1653 -2826 1671 -2784
rect 1592 -2846 1671 -2826
rect 1861 -2780 1940 -2761
rect 1861 -2822 1877 -2780
rect 1922 -2822 1940 -2780
rect 1861 -2842 1940 -2822
rect -2540 -2899 -2462 -2880
rect -7116 -3063 -6916 -2948
rect -2331 -3061 -2263 -3048
rect -2331 -3063 -2321 -3061
rect -7116 -3099 -2321 -3063
rect -7116 -3148 -6916 -3099
rect -2331 -3103 -2321 -3099
rect -2276 -3103 -2263 -3061
rect -2331 -3120 -2263 -3103
<< via1 >>
rect 2808 2147 2920 2247
rect -5576 1510 -5464 1610
rect -3918 1510 -3806 1610
rect -1524 1648 -1472 1700
rect -5378 191 -5326 243
rect -4958 195 -4906 247
rect -5678 -668 -5626 -616
rect -5685 -861 -5633 -809
rect -5683 -1045 -5631 -993
rect -5684 -1156 -5632 -1104
rect -5707 -2202 -5655 -2150
rect -3292 209 -3240 261
rect -5258 -34 -5146 66
rect -3600 -34 -3488 66
rect -3212 -782 -3160 -730
rect -4982 -941 -4930 -889
rect -2232 -544 -2180 -491
rect -1859 -544 -1807 -491
rect -1768 -664 -1716 -611
rect -1293 -787 -1241 -735
rect -2003 -822 -1945 -813
rect -2003 -867 -1998 -822
rect -1998 -867 -1949 -822
rect -1949 -867 -1945 -822
rect -2003 -870 -1945 -867
rect -1654 -2022 -1602 -1970
rect 3887 2146 3999 2246
rect 4992 2170 5044 2222
rect 1235 1492 1287 1544
rect 3278 -100 3390 0
rect 4357 -95 4469 5
rect -417 -1048 -365 -996
rect -296 -1149 -244 -1097
rect 2918 -367 3030 -267
rect 3997 -368 4109 -268
rect 5011 -348 5063 -296
rect 1917 -855 1969 -803
rect 1430 -1102 1482 -1050
rect -825 -2097 -773 -2045
rect -446 -2447 -394 -2395
rect -54 -2023 -2 -1971
rect 996 -2068 1048 -2016
rect 3388 -2614 3500 -2514
rect 4467 -2609 4579 -2509
<< metal2 >>
rect 2792 2251 2936 2263
rect 2792 2240 2802 2251
rect 1620 2177 2802 2240
rect -1537 1702 -1460 1715
rect -1537 1646 -1526 1702
rect -1470 1646 -1460 1702
rect -1537 1630 -1460 1646
rect -5592 1614 -5448 1626
rect -5592 1506 -5582 1614
rect -5460 1506 -5448 1614
rect -5592 1496 -5448 1506
rect -3934 1614 -3790 1626
rect -3934 1506 -3924 1614
rect -3802 1506 -3790 1614
rect -3934 1496 -3790 1506
rect 1222 1546 1299 1559
rect 1222 1490 1233 1546
rect 1289 1490 1299 1546
rect 1222 1474 1299 1490
rect -3302 261 -3230 284
rect -5384 243 -5309 255
rect -5384 191 -5378 243
rect -5326 232 -5309 243
rect -4964 247 -4900 253
rect -4964 232 -4958 247
rect -5326 202 -4958 232
rect -5326 191 -5309 202
rect -5384 182 -5309 191
rect -4964 195 -4958 202
rect -4906 232 -4900 247
rect -3302 232 -3292 261
rect -4906 209 -3292 232
rect -3240 209 -3230 261
rect -4906 202 -3230 209
rect -4906 195 -4900 202
rect -3302 197 -3230 202
rect -4964 189 -4900 195
rect -5274 70 -5130 82
rect -5274 -38 -5264 70
rect -5142 -38 -5130 70
rect -5274 -48 -5130 -38
rect -3616 70 -3472 82
rect -3616 -38 -3606 70
rect -3484 -38 -3472 70
rect -3616 -48 -3472 -38
rect -2237 -491 -2174 -484
rect -2237 -544 -2232 -491
rect -2180 -508 -2174 -491
rect -1866 -491 -1802 -481
rect -1866 -508 -1859 -491
rect -2180 -544 -1859 -508
rect -1807 -544 -1802 -491
rect -2237 -550 -1802 -544
rect -5685 -616 -5621 -607
rect -5685 -668 -5678 -616
rect -5626 -619 -5621 -616
rect -1775 -611 -1711 -601
rect -5626 -620 -2200 -619
rect -1775 -620 -1768 -611
rect -5626 -660 -1768 -620
rect -5626 -668 -5621 -660
rect -5397 -661 -1768 -660
rect -5685 -677 -5621 -668
rect -1775 -664 -1768 -661
rect -1716 -664 -1711 -611
rect -1775 -670 -1711 -664
rect 1620 -692 1659 2177
rect 2792 2143 2802 2177
rect 2924 2143 2936 2251
rect 2792 2133 2936 2143
rect 3871 2250 4015 2262
rect 3871 2142 3881 2250
rect 4003 2227 4015 2250
rect 4987 2227 5051 2231
rect 4003 2222 5051 2227
rect 4003 2170 4992 2222
rect 5044 2170 5051 2222
rect 4003 2165 5051 2170
rect 4003 2142 4015 2165
rect 4987 2161 5051 2165
rect 3871 2132 4015 2142
rect 3262 4 3408 14
rect 3262 -23 3274 4
rect 993 -722 1659 -692
rect 2297 -78 3274 -23
rect -3218 -730 -3154 -724
rect -3218 -782 -3212 -730
rect -3160 -745 -3154 -730
rect -1299 -735 -1235 -729
rect -1299 -745 -1293 -735
rect -3160 -775 -1293 -745
rect -3160 -782 -3154 -775
rect -3218 -788 -3154 -782
rect -1299 -787 -1293 -775
rect -1241 -748 -1235 -735
rect 993 -748 1027 -722
rect -1241 -778 1027 -748
rect -1241 -787 -1235 -778
rect -1299 -793 -1235 -787
rect -5692 -809 -5628 -800
rect 1911 -803 1975 -797
rect -5692 -861 -5685 -809
rect -5633 -822 -5628 -809
rect -2012 -813 -1939 -806
rect -5633 -823 -2435 -822
rect -2012 -823 -2003 -813
rect -5633 -853 -2003 -823
rect -5633 -861 -5628 -853
rect -5396 -854 -2003 -853
rect -5692 -870 -5628 -861
rect -2012 -870 -2003 -854
rect -1945 -870 -1939 -813
rect 1911 -815 1917 -803
rect -2012 -875 -1939 -870
rect 1306 -845 1917 -815
rect -4988 -889 -4924 -883
rect -4988 -941 -4982 -889
rect -4930 -904 -4924 -889
rect 1306 -904 1337 -845
rect 1911 -855 1917 -845
rect 1969 -855 1975 -803
rect 1911 -861 1975 -855
rect -4930 -934 1337 -904
rect 1421 -883 1494 -874
rect -4930 -941 -4924 -934
rect -4988 -947 -4924 -941
rect 1421 -939 1430 -883
rect 1486 -939 1494 -883
rect -5690 -993 -5626 -984
rect -5690 -1045 -5683 -993
rect -5631 -1002 -5626 -993
rect -423 -996 -359 -990
rect -5631 -1003 -849 -1002
rect -423 -1003 -417 -996
rect -5631 -1032 -417 -1003
rect -5631 -1045 -5626 -1032
rect -5264 -1033 -417 -1032
rect -5690 -1054 -5626 -1045
rect -423 -1048 -417 -1033
rect -365 -1048 -359 -996
rect -423 -1054 -359 -1048
rect 1421 -1050 1494 -939
rect -5711 -1104 -5615 -1094
rect -5711 -1156 -5684 -1104
rect -5632 -1110 -5615 -1104
rect -302 -1097 -238 -1091
rect -5632 -1111 -728 -1110
rect -302 -1111 -296 -1097
rect -5632 -1144 -296 -1111
rect -5632 -1156 -5615 -1144
rect -5244 -1145 -296 -1144
rect -302 -1149 -296 -1145
rect -244 -1101 -238 -1097
rect -244 -1149 -237 -1101
rect 1421 -1102 1430 -1050
rect 1482 -1102 1494 -1050
rect 1421 -1105 1494 -1102
rect 1421 -1106 1490 -1105
rect -302 -1154 -237 -1149
rect -302 -1155 -238 -1154
rect -5711 -1165 -5615 -1156
rect -1665 -1968 -1596 -1961
rect -60 -1968 5 -1964
rect -1665 -1970 5 -1968
rect -1665 -2022 -1654 -1970
rect -1602 -1971 5 -1970
rect -1602 -2002 -54 -1971
rect -1602 -2022 -1596 -2002
rect -61 -2006 -54 -2002
rect -1665 -2029 -1596 -2022
rect -60 -2023 -54 -2006
rect -2 -2023 5 -1971
rect -60 -2030 5 -2023
rect 990 -2016 1054 -2010
rect 990 -2026 996 -2016
rect -838 -2043 -761 -2030
rect -838 -2099 -827 -2043
rect -771 -2099 -761 -2043
rect 989 -2056 996 -2026
rect 990 -2068 996 -2056
rect 1048 -2068 1054 -2016
rect 990 -2074 1054 -2068
rect -838 -2115 -761 -2099
rect -5714 -2150 -5650 -2141
rect -5714 -2202 -5707 -2150
rect -5655 -2151 612 -2150
rect 999 -2151 1045 -2074
rect -5655 -2197 1044 -2151
rect -5655 -2202 -5650 -2197
rect -5246 -2198 1044 -2197
rect -5714 -2211 -5650 -2202
rect -452 -2395 -388 -2389
rect -452 -2447 -446 -2395
rect -394 -2412 -388 -2395
rect 2297 -2412 2331 -78
rect 3262 -104 3274 -78
rect 3396 -104 3408 4
rect 3262 -116 3408 -104
rect 4341 9 4485 19
rect 4341 -99 4353 9
rect 4475 -99 4485 9
rect 4341 -111 4485 -99
rect 2902 -263 3046 -251
rect 2902 -371 2912 -263
rect 3034 -371 3046 -263
rect 2902 -381 3046 -371
rect 3981 -264 4125 -252
rect 3981 -372 3991 -264
rect 4113 -287 4125 -264
rect 4113 -296 5070 -287
rect 4113 -348 5011 -296
rect 5063 -348 5070 -296
rect 4113 -355 5070 -348
rect 4113 -372 4125 -355
rect 5006 -357 5070 -355
rect 3981 -382 4125 -372
rect -394 -2446 2331 -2412
rect -394 -2447 -388 -2446
rect -452 -2453 -388 -2447
rect 3372 -2510 3518 -2498
rect 3372 -2618 3384 -2510
rect 3506 -2618 3518 -2510
rect 3372 -2628 3518 -2618
rect 4451 -2505 4595 -2495
rect 4451 -2613 4463 -2505
rect 4585 -2613 4595 -2505
rect 4451 -2625 4595 -2613
rect 3372 -2630 3516 -2628
<< via2 >>
rect 2802 2247 2924 2251
rect -1526 1700 -1470 1702
rect -1526 1648 -1524 1700
rect -1524 1648 -1472 1700
rect -1472 1648 -1470 1700
rect -1526 1646 -1470 1648
rect -5582 1610 -5460 1614
rect -5582 1510 -5576 1610
rect -5576 1510 -5464 1610
rect -5464 1510 -5460 1610
rect -5582 1506 -5460 1510
rect -3924 1610 -3802 1614
rect -3924 1510 -3918 1610
rect -3918 1510 -3806 1610
rect -3806 1510 -3802 1610
rect -3924 1506 -3802 1510
rect 1233 1544 1289 1546
rect 1233 1492 1235 1544
rect 1235 1492 1287 1544
rect 1287 1492 1289 1544
rect 1233 1490 1289 1492
rect -5264 66 -5142 70
rect -5264 -34 -5258 66
rect -5258 -34 -5146 66
rect -5146 -34 -5142 66
rect -5264 -38 -5142 -34
rect -3606 66 -3484 70
rect -3606 -34 -3600 66
rect -3600 -34 -3488 66
rect -3488 -34 -3484 66
rect -3606 -38 -3484 -34
rect 2802 2147 2808 2247
rect 2808 2147 2920 2247
rect 2920 2147 2924 2247
rect 2802 2143 2924 2147
rect 3881 2246 4003 2250
rect 3881 2146 3887 2246
rect 3887 2146 3999 2246
rect 3999 2146 4003 2246
rect 3881 2142 4003 2146
rect 3274 0 3396 4
rect 1430 -939 1486 -883
rect -827 -2045 -771 -2043
rect -827 -2097 -825 -2045
rect -825 -2097 -773 -2045
rect -773 -2097 -771 -2045
rect -827 -2099 -771 -2097
rect 3274 -100 3278 0
rect 3278 -100 3390 0
rect 3390 -100 3396 0
rect 3274 -104 3396 -100
rect 4353 5 4475 9
rect 4353 -95 4357 5
rect 4357 -95 4469 5
rect 4469 -95 4475 5
rect 4353 -99 4475 -95
rect 2912 -267 3034 -263
rect 2912 -367 2918 -267
rect 2918 -367 3030 -267
rect 3030 -367 3034 -267
rect 2912 -371 3034 -367
rect 3991 -268 4113 -264
rect 3991 -368 3997 -268
rect 3997 -368 4109 -268
rect 4109 -368 4113 -268
rect 3991 -372 4113 -368
rect 3384 -2514 3506 -2510
rect 3384 -2614 3388 -2514
rect 3388 -2614 3500 -2514
rect 3500 -2614 3506 -2514
rect 3384 -2618 3506 -2614
rect 4463 -2509 4585 -2505
rect 4463 -2609 4467 -2509
rect 4467 -2609 4579 -2509
rect 4579 -2609 4585 -2509
rect 4463 -2613 4585 -2609
<< metal3 >>
rect 2792 2255 2934 2261
rect 2792 2139 2798 2255
rect 2926 2139 2934 2255
rect 2792 2133 2934 2139
rect 3871 2254 4013 2260
rect 3871 2138 3877 2254
rect 4005 2138 4013 2254
rect 3871 2132 4013 2138
rect -1537 1702 -1460 1715
rect -1537 1646 -1526 1702
rect -1470 1646 -1460 1702
rect -1537 1630 -1460 1646
rect -5592 1618 -5450 1624
rect -5592 1502 -5586 1618
rect -5458 1502 -5450 1618
rect -5592 1496 -5450 1502
rect -3934 1618 -3792 1624
rect -3934 1502 -3928 1618
rect -3800 1502 -3792 1618
rect -3934 1496 -3792 1502
rect -5274 74 -5132 80
rect -5274 -42 -5268 74
rect -5140 -42 -5132 74
rect -5274 -48 -5132 -42
rect -3616 74 -3474 80
rect -3616 -42 -3610 74
rect -3482 -42 -3474 74
rect -3616 -48 -3474 -42
rect -1534 -2031 -1462 1630
rect 1222 1546 1299 1559
rect 1222 1490 1233 1546
rect 1289 1490 1299 1546
rect 1222 1474 1299 1490
rect 1230 -831 1293 1474
rect 3264 8 3406 14
rect 3264 -108 3272 8
rect 3400 -108 3406 8
rect 3264 -114 3406 -108
rect 4343 13 4485 19
rect 4343 -103 4351 13
rect 4479 -103 4485 13
rect 4343 -109 4485 -103
rect 2902 -259 3044 -253
rect 2902 -375 2908 -259
rect 3036 -375 3044 -259
rect 2902 -381 3044 -375
rect 3981 -260 4123 -254
rect 3981 -376 3987 -260
rect 4115 -376 4123 -260
rect 3981 -382 4123 -376
rect 1230 -883 1496 -831
rect 1230 -894 1430 -883
rect 1420 -939 1430 -894
rect 1486 -894 1496 -883
rect 1486 -939 1495 -894
rect 1420 -944 1495 -939
rect -838 -2031 -761 -2030
rect -1534 -2043 -761 -2031
rect -1534 -2099 -827 -2043
rect -771 -2099 -761 -2043
rect -1534 -2112 -761 -2099
rect -838 -2115 -761 -2112
rect 3374 -2506 3516 -2500
rect 3374 -2622 3382 -2506
rect 3510 -2622 3516 -2506
rect 3374 -2628 3516 -2622
rect 4453 -2501 4595 -2495
rect 4453 -2617 4461 -2501
rect 4589 -2617 4595 -2501
rect 4453 -2623 4595 -2617
<< via3 >>
rect 2798 2251 2926 2255
rect 2798 2143 2802 2251
rect 2802 2143 2924 2251
rect 2924 2143 2926 2251
rect 2798 2139 2926 2143
rect 3877 2250 4005 2254
rect 3877 2142 3881 2250
rect 3881 2142 4003 2250
rect 4003 2142 4005 2250
rect 3877 2138 4005 2142
rect -5586 1614 -5458 1618
rect -5586 1506 -5582 1614
rect -5582 1506 -5460 1614
rect -5460 1506 -5458 1614
rect -5586 1502 -5458 1506
rect -3928 1614 -3800 1618
rect -3928 1506 -3924 1614
rect -3924 1506 -3802 1614
rect -3802 1506 -3800 1614
rect -3928 1502 -3800 1506
rect -5268 70 -5140 74
rect -5268 -38 -5264 70
rect -5264 -38 -5142 70
rect -5142 -38 -5140 70
rect -5268 -42 -5140 -38
rect -3610 70 -3482 74
rect -3610 -38 -3606 70
rect -3606 -38 -3484 70
rect -3484 -38 -3482 70
rect -3610 -42 -3482 -38
rect 3272 4 3400 8
rect 3272 -104 3274 4
rect 3274 -104 3396 4
rect 3396 -104 3400 4
rect 3272 -108 3400 -104
rect 4351 9 4479 13
rect 4351 -99 4353 9
rect 4353 -99 4475 9
rect 4475 -99 4479 9
rect 4351 -103 4479 -99
rect 2908 -263 3036 -259
rect 2908 -371 2912 -263
rect 2912 -371 3034 -263
rect 3034 -371 3036 -263
rect 2908 -375 3036 -371
rect 3987 -264 4115 -260
rect 3987 -372 3991 -264
rect 3991 -372 4113 -264
rect 4113 -372 4115 -264
rect 3987 -376 4115 -372
rect 3382 -2510 3510 -2506
rect 3382 -2618 3384 -2510
rect 3384 -2618 3506 -2510
rect 3506 -2618 3510 -2510
rect 3382 -2622 3510 -2618
rect 4461 -2505 4589 -2501
rect 4461 -2613 4463 -2505
rect 4463 -2613 4585 -2505
rect 4585 -2613 4589 -2505
rect 4461 -2617 4589 -2613
<< metal4 >>
rect 2790 2255 2936 2263
rect 2790 2139 2798 2255
rect 2926 2139 2936 2255
rect 2790 2133 2936 2139
rect 3869 2254 4015 2262
rect 3869 2138 3877 2254
rect 4005 2138 4015 2254
rect 2812 2032 2916 2133
rect 3869 2132 4015 2138
rect 3891 2045 3995 2132
rect -5594 1618 -5448 1626
rect -5594 1502 -5586 1618
rect -5458 1502 -5448 1618
rect -5594 1496 -5448 1502
rect -3936 1618 -3790 1626
rect -3936 1502 -3928 1618
rect -3800 1502 -3790 1618
rect -3936 1496 -3790 1502
rect -5539 1240 -5476 1496
rect -3880 981 -3817 1496
rect -3878 932 -3817 981
rect -5234 82 -5174 456
rect -3576 82 -3516 626
rect -5276 74 -5130 82
rect -5276 -42 -5268 74
rect -5140 -42 -5130 74
rect -5276 -48 -5130 -42
rect -3618 74 -3472 82
rect -3618 -42 -3610 74
rect -3482 -42 -3472 74
rect 3282 14 3386 101
rect 4361 19 4465 107
rect -3618 -48 -3472 -42
rect 3262 8 3408 14
rect -5218 -60 -5158 -48
rect -3560 -60 -3500 -48
rect 3262 -108 3272 8
rect 3400 -108 3408 8
rect 3262 -116 3408 -108
rect 4341 13 4487 19
rect 4341 -103 4351 13
rect 4479 -103 4487 13
rect 4341 -111 4487 -103
rect 2900 -259 3046 -251
rect 2900 -375 2908 -259
rect 3036 -375 3046 -259
rect 2900 -381 3046 -375
rect 3979 -260 4125 -252
rect 3979 -376 3987 -260
rect 4115 -376 4125 -260
rect 2922 -406 3026 -381
rect 3979 -382 4125 -376
rect 4001 -406 4105 -382
rect 3392 -2498 3496 -2434
rect 4471 -2495 4575 -2434
rect 3372 -2506 3518 -2498
rect 3372 -2622 3382 -2506
rect 3510 -2622 3518 -2506
rect 3372 -2630 3518 -2622
rect 4451 -2501 4597 -2495
rect 4451 -2617 4461 -2501
rect 4589 -2617 4597 -2501
rect 4451 -2625 4597 -2617
<< labels >>
flabel metal1 -7116 -3148 -6916 -2948 0 FreeSans 256 0 0 0 GND
port 6 nsew
flabel metal1 -7116 1941 -6916 2141 0 FreeSans 256 0 0 0 VDD
port 7 nsew
flabel metal1 -7116 -2259 -6916 -2059 0 FreeSans 256 0 0 0 Vin
port 3 nsew
flabel metal1 -7116 -1829 -6916 -1629 0 FreeSans 256 0 0 0 Vbiasn
port 8 nsew
flabel metal1 -7116 -1427 -6916 -1227 0 FreeSans 256 0 0 0 Vip
port 2 nsew
flabel metal1 -7116 -1027 -6916 -827 0 FreeSans 256 0 0 0 Vcm
port 5 nsew
flabel metal1 -7116 -627 -6916 -427 0 FreeSans 256 0 0 0 Vbp
port 4 nsew
flabel metal1 5175 -400 5375 -200 0 FreeSans 256 0 0 0 Von
port 1 nsew
flabel metal1 5151 2101 5351 2301 0 FreeSans 256 0 0 0 Vop
port 0 nsew
rlabel metal1 -7096 1492 -6948 1632 1 Vabp
port 10 n
rlabel metal1 -7096 1180 -6938 1330 1 Vabn
port 11 n
<< end >>
