magic
tech sky130A
magscale 1 2
timestamp 1666663403
<< nmos >>
rect -45 -113 45 113
<< ndiff >>
rect -103 101 -45 113
rect -103 -101 -91 101
rect -57 -101 -45 101
rect -103 -113 -45 -101
rect 45 101 103 113
rect 45 -101 57 101
rect 91 -101 103 101
rect 45 -113 103 -101
<< ndiffc >>
rect -91 -101 -57 101
rect 57 -101 91 101
<< poly >>
rect -45 185 45 201
rect -45 151 -29 185
rect 29 151 45 185
rect -45 113 45 151
rect -45 -151 45 -113
rect -45 -185 -29 -151
rect 29 -185 45 -151
rect -45 -201 45 -185
<< polycont >>
rect -29 151 29 185
rect -29 -185 29 -151
<< locali >>
rect -45 151 -29 185
rect 29 151 45 185
rect -91 101 -57 117
rect -91 -117 -57 -101
rect 57 101 91 117
rect 57 -117 91 -101
rect -45 -185 -29 -151
rect 29 -185 45 -151
<< viali >>
rect -29 151 29 185
rect -91 -101 -57 101
rect 57 -101 91 101
rect -29 -185 29 -151
<< metal1 >>
rect -41 185 41 191
rect -41 151 -29 185
rect 29 151 41 185
rect -41 145 41 151
rect -97 101 -51 113
rect -97 -101 -91 101
rect -57 -101 -51 101
rect -97 -113 -51 -101
rect 51 101 97 113
rect 51 -101 57 101
rect 91 -101 97 101
rect 51 -113 97 -101
rect -41 -151 41 -145
rect -41 -185 -29 -151
rect 29 -185 41 -151
rect -41 -191 41 -185
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.13 l 0.45 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
