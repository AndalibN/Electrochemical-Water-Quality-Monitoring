magic
tech sky130A
timestamp 1662586819
<< nmos >>
rect -10 -25 10 25
<< ndiff >>
rect -39 19 -10 25
rect -39 -19 -33 19
rect -16 -19 -10 19
rect -39 -25 -10 -19
rect 10 19 39 25
rect 10 -19 16 19
rect 33 -19 39 19
rect 10 -25 39 -19
<< ndiffc >>
rect -33 -19 -16 19
rect 16 -19 33 19
<< poly >>
rect -10 25 10 38
rect -10 -38 10 -25
<< locali >>
rect -33 19 -16 27
rect -33 -27 -16 -19
rect 16 19 33 27
rect 16 -27 33 -19
<< viali >>
rect -33 -19 -16 19
rect 16 -19 33 19
<< metal1 >>
rect -36 19 -13 25
rect -36 -19 -33 19
rect -16 -19 -13 19
rect -36 -25 -13 -19
rect 13 19 36 25
rect 13 -19 16 19
rect 33 -19 36 19
rect 13 -25 36 -19
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
