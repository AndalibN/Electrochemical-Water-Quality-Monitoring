magic
tech sky130A
magscale 1 2
timestamp 1668714565
<< nmos >>
rect -861 -8300 -741 8300
rect -683 -8300 -563 8300
rect -505 -8300 -385 8300
rect -327 -8300 -207 8300
rect -149 -8300 -29 8300
rect 29 -8300 149 8300
rect 207 -8300 327 8300
rect 385 -8300 505 8300
rect 563 -8300 683 8300
rect 741 -8300 861 8300
<< ndiff >>
rect -919 8288 -861 8300
rect -919 -8288 -907 8288
rect -873 -8288 -861 8288
rect -919 -8300 -861 -8288
rect -741 8288 -683 8300
rect -741 -8288 -729 8288
rect -695 -8288 -683 8288
rect -741 -8300 -683 -8288
rect -563 8288 -505 8300
rect -563 -8288 -551 8288
rect -517 -8288 -505 8288
rect -563 -8300 -505 -8288
rect -385 8288 -327 8300
rect -385 -8288 -373 8288
rect -339 -8288 -327 8288
rect -385 -8300 -327 -8288
rect -207 8288 -149 8300
rect -207 -8288 -195 8288
rect -161 -8288 -149 8288
rect -207 -8300 -149 -8288
rect -29 8288 29 8300
rect -29 -8288 -17 8288
rect 17 -8288 29 8288
rect -29 -8300 29 -8288
rect 149 8288 207 8300
rect 149 -8288 161 8288
rect 195 -8288 207 8288
rect 149 -8300 207 -8288
rect 327 8288 385 8300
rect 327 -8288 339 8288
rect 373 -8288 385 8288
rect 327 -8300 385 -8288
rect 505 8288 563 8300
rect 505 -8288 517 8288
rect 551 -8288 563 8288
rect 505 -8300 563 -8288
rect 683 8288 741 8300
rect 683 -8288 695 8288
rect 729 -8288 741 8288
rect 683 -8300 741 -8288
rect 861 8288 919 8300
rect 861 -8288 873 8288
rect 907 -8288 919 8288
rect 861 -8300 919 -8288
<< ndiffc >>
rect -907 -8288 -873 8288
rect -729 -8288 -695 8288
rect -551 -8288 -517 8288
rect -373 -8288 -339 8288
rect -195 -8288 -161 8288
rect -17 -8288 17 8288
rect 161 -8288 195 8288
rect 339 -8288 373 8288
rect 517 -8288 551 8288
rect 695 -8288 729 8288
rect 873 -8288 907 8288
<< poly >>
rect -861 8372 -741 8388
rect -861 8338 -845 8372
rect -757 8338 -741 8372
rect -861 8300 -741 8338
rect -683 8372 -563 8388
rect -683 8338 -667 8372
rect -579 8338 -563 8372
rect -683 8300 -563 8338
rect -505 8372 -385 8388
rect -505 8338 -489 8372
rect -401 8338 -385 8372
rect -505 8300 -385 8338
rect -327 8372 -207 8388
rect -327 8338 -311 8372
rect -223 8338 -207 8372
rect -327 8300 -207 8338
rect -149 8372 -29 8388
rect -149 8338 -133 8372
rect -45 8338 -29 8372
rect -149 8300 -29 8338
rect 29 8372 149 8388
rect 29 8338 45 8372
rect 133 8338 149 8372
rect 29 8300 149 8338
rect 207 8372 327 8388
rect 207 8338 223 8372
rect 311 8338 327 8372
rect 207 8300 327 8338
rect 385 8372 505 8388
rect 385 8338 401 8372
rect 489 8338 505 8372
rect 385 8300 505 8338
rect 563 8372 683 8388
rect 563 8338 579 8372
rect 667 8338 683 8372
rect 563 8300 683 8338
rect 741 8372 861 8388
rect 741 8338 757 8372
rect 845 8338 861 8372
rect 741 8300 861 8338
rect -861 -8338 -741 -8300
rect -861 -8372 -845 -8338
rect -757 -8372 -741 -8338
rect -861 -8388 -741 -8372
rect -683 -8338 -563 -8300
rect -683 -8372 -667 -8338
rect -579 -8372 -563 -8338
rect -683 -8388 -563 -8372
rect -505 -8338 -385 -8300
rect -505 -8372 -489 -8338
rect -401 -8372 -385 -8338
rect -505 -8388 -385 -8372
rect -327 -8338 -207 -8300
rect -327 -8372 -311 -8338
rect -223 -8372 -207 -8338
rect -327 -8388 -207 -8372
rect -149 -8338 -29 -8300
rect -149 -8372 -133 -8338
rect -45 -8372 -29 -8338
rect -149 -8388 -29 -8372
rect 29 -8338 149 -8300
rect 29 -8372 45 -8338
rect 133 -8372 149 -8338
rect 29 -8388 149 -8372
rect 207 -8338 327 -8300
rect 207 -8372 223 -8338
rect 311 -8372 327 -8338
rect 207 -8388 327 -8372
rect 385 -8338 505 -8300
rect 385 -8372 401 -8338
rect 489 -8372 505 -8338
rect 385 -8388 505 -8372
rect 563 -8338 683 -8300
rect 563 -8372 579 -8338
rect 667 -8372 683 -8338
rect 563 -8388 683 -8372
rect 741 -8338 861 -8300
rect 741 -8372 757 -8338
rect 845 -8372 861 -8338
rect 741 -8388 861 -8372
<< polycont >>
rect -845 8338 -757 8372
rect -667 8338 -579 8372
rect -489 8338 -401 8372
rect -311 8338 -223 8372
rect -133 8338 -45 8372
rect 45 8338 133 8372
rect 223 8338 311 8372
rect 401 8338 489 8372
rect 579 8338 667 8372
rect 757 8338 845 8372
rect -845 -8372 -757 -8338
rect -667 -8372 -579 -8338
rect -489 -8372 -401 -8338
rect -311 -8372 -223 -8338
rect -133 -8372 -45 -8338
rect 45 -8372 133 -8338
rect 223 -8372 311 -8338
rect 401 -8372 489 -8338
rect 579 -8372 667 -8338
rect 757 -8372 845 -8338
<< locali >>
rect -861 8338 -845 8372
rect -757 8338 -741 8372
rect -683 8338 -667 8372
rect -579 8338 -563 8372
rect -505 8338 -489 8372
rect -401 8338 -385 8372
rect -327 8338 -311 8372
rect -223 8338 -207 8372
rect -149 8338 -133 8372
rect -45 8338 -29 8372
rect 29 8338 45 8372
rect 133 8338 149 8372
rect 207 8338 223 8372
rect 311 8338 327 8372
rect 385 8338 401 8372
rect 489 8338 505 8372
rect 563 8338 579 8372
rect 667 8338 683 8372
rect 741 8338 757 8372
rect 845 8338 861 8372
rect -907 8288 -873 8304
rect -907 -8304 -873 -8288
rect -729 8288 -695 8304
rect -729 -8304 -695 -8288
rect -551 8288 -517 8304
rect -551 -8304 -517 -8288
rect -373 8288 -339 8304
rect -373 -8304 -339 -8288
rect -195 8288 -161 8304
rect -195 -8304 -161 -8288
rect -17 8288 17 8304
rect -17 -8304 17 -8288
rect 161 8288 195 8304
rect 161 -8304 195 -8288
rect 339 8288 373 8304
rect 339 -8304 373 -8288
rect 517 8288 551 8304
rect 517 -8304 551 -8288
rect 695 8288 729 8304
rect 695 -8304 729 -8288
rect 873 8288 907 8304
rect 873 -8304 907 -8288
rect -861 -8372 -845 -8338
rect -757 -8372 -741 -8338
rect -683 -8372 -667 -8338
rect -579 -8372 -563 -8338
rect -505 -8372 -489 -8338
rect -401 -8372 -385 -8338
rect -327 -8372 -311 -8338
rect -223 -8372 -207 -8338
rect -149 -8372 -133 -8338
rect -45 -8372 -29 -8338
rect 29 -8372 45 -8338
rect 133 -8372 149 -8338
rect 207 -8372 223 -8338
rect 311 -8372 327 -8338
rect 385 -8372 401 -8338
rect 489 -8372 505 -8338
rect 563 -8372 579 -8338
rect 667 -8372 683 -8338
rect 741 -8372 757 -8338
rect 845 -8372 861 -8338
<< viali >>
rect -845 8338 -757 8372
rect -667 8338 -579 8372
rect -489 8338 -401 8372
rect -311 8338 -223 8372
rect -133 8338 -45 8372
rect 45 8338 133 8372
rect 223 8338 311 8372
rect 401 8338 489 8372
rect 579 8338 667 8372
rect 757 8338 845 8372
rect -907 -8288 -873 8288
rect -729 -8288 -695 8288
rect -551 -8288 -517 8288
rect -373 -8288 -339 8288
rect -195 -8288 -161 8288
rect -17 -8288 17 8288
rect 161 -8288 195 8288
rect 339 -8288 373 8288
rect 517 -8288 551 8288
rect 695 -8288 729 8288
rect 873 -8288 907 8288
rect -845 -8372 -757 -8338
rect -667 -8372 -579 -8338
rect -489 -8372 -401 -8338
rect -311 -8372 -223 -8338
rect -133 -8372 -45 -8338
rect 45 -8372 133 -8338
rect 223 -8372 311 -8338
rect 401 -8372 489 -8338
rect 579 -8372 667 -8338
rect 757 -8372 845 -8338
<< metal1 >>
rect -857 8372 -745 8378
rect -857 8338 -845 8372
rect -757 8338 -745 8372
rect -857 8332 -745 8338
rect -679 8372 -567 8378
rect -679 8338 -667 8372
rect -579 8338 -567 8372
rect -679 8332 -567 8338
rect -501 8372 -389 8378
rect -501 8338 -489 8372
rect -401 8338 -389 8372
rect -501 8332 -389 8338
rect -323 8372 -211 8378
rect -323 8338 -311 8372
rect -223 8338 -211 8372
rect -323 8332 -211 8338
rect -145 8372 -33 8378
rect -145 8338 -133 8372
rect -45 8338 -33 8372
rect -145 8332 -33 8338
rect 33 8372 145 8378
rect 33 8338 45 8372
rect 133 8338 145 8372
rect 33 8332 145 8338
rect 211 8372 323 8378
rect 211 8338 223 8372
rect 311 8338 323 8372
rect 211 8332 323 8338
rect 389 8372 501 8378
rect 389 8338 401 8372
rect 489 8338 501 8372
rect 389 8332 501 8338
rect 567 8372 679 8378
rect 567 8338 579 8372
rect 667 8338 679 8372
rect 567 8332 679 8338
rect 745 8372 857 8378
rect 745 8338 757 8372
rect 845 8338 857 8372
rect 745 8332 857 8338
rect -913 8288 -867 8300
rect -913 -8288 -907 8288
rect -873 -8288 -867 8288
rect -913 -8300 -867 -8288
rect -735 8288 -689 8300
rect -735 -8288 -729 8288
rect -695 -8288 -689 8288
rect -735 -8300 -689 -8288
rect -557 8288 -511 8300
rect -557 -8288 -551 8288
rect -517 -8288 -511 8288
rect -557 -8300 -511 -8288
rect -379 8288 -333 8300
rect -379 -8288 -373 8288
rect -339 -8288 -333 8288
rect -379 -8300 -333 -8288
rect -201 8288 -155 8300
rect -201 -8288 -195 8288
rect -161 -8288 -155 8288
rect -201 -8300 -155 -8288
rect -23 8288 23 8300
rect -23 -8288 -17 8288
rect 17 -8288 23 8288
rect -23 -8300 23 -8288
rect 155 8288 201 8300
rect 155 -8288 161 8288
rect 195 -8288 201 8288
rect 155 -8300 201 -8288
rect 333 8288 379 8300
rect 333 -8288 339 8288
rect 373 -8288 379 8288
rect 333 -8300 379 -8288
rect 511 8288 557 8300
rect 511 -8288 517 8288
rect 551 -8288 557 8288
rect 511 -8300 557 -8288
rect 689 8288 735 8300
rect 689 -8288 695 8288
rect 729 -8288 735 8288
rect 689 -8300 735 -8288
rect 867 8288 913 8300
rect 867 -8288 873 8288
rect 907 -8288 913 8288
rect 867 -8300 913 -8288
rect -857 -8338 -745 -8332
rect -857 -8372 -845 -8338
rect -757 -8372 -745 -8338
rect -857 -8378 -745 -8372
rect -679 -8338 -567 -8332
rect -679 -8372 -667 -8338
rect -579 -8372 -567 -8338
rect -679 -8378 -567 -8372
rect -501 -8338 -389 -8332
rect -501 -8372 -489 -8338
rect -401 -8372 -389 -8338
rect -501 -8378 -389 -8372
rect -323 -8338 -211 -8332
rect -323 -8372 -311 -8338
rect -223 -8372 -211 -8338
rect -323 -8378 -211 -8372
rect -145 -8338 -33 -8332
rect -145 -8372 -133 -8338
rect -45 -8372 -33 -8338
rect -145 -8378 -33 -8372
rect 33 -8338 145 -8332
rect 33 -8372 45 -8338
rect 133 -8372 145 -8338
rect 33 -8378 145 -8372
rect 211 -8338 323 -8332
rect 211 -8372 223 -8338
rect 311 -8372 323 -8338
rect 211 -8378 323 -8372
rect 389 -8338 501 -8332
rect 389 -8372 401 -8338
rect 489 -8372 501 -8338
rect 389 -8378 501 -8372
rect 567 -8338 679 -8332
rect 567 -8372 579 -8338
rect 667 -8372 679 -8338
rect 567 -8378 679 -8372
rect 745 -8338 857 -8332
rect 745 -8372 757 -8338
rect 845 -8372 857 -8338
rect 745 -8378 857 -8372
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 83 l 0.6 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
