magic
tech sky130A
magscale 1 2
timestamp 1669522289
<< error_p >>
rect 191917 524844 191918 524848
<< error_s >>
rect 471905 144063 471961 144076
rect 472107 144063 472375 144076
<< nwell >>
rect 76034 588188 76042 588306
rect 77982 588198 77992 588336
<< locali >>
rect 77982 588198 77992 588336
rect 79334 588224 79338 588244
rect 473947 144029 474002 144076
rect 471742 143976 471796 144019
rect 472156 143976 472210 144019
rect 472274 143976 472328 144020
rect 469811 143837 469866 143883
<< metal1 >>
rect 555848 644394 570748 646373
rect 11447 631068 16257 631627
rect 11447 627560 11934 631068
rect 15698 627560 16257 631068
rect 555848 630134 558070 644394
rect 568234 630134 570748 644394
rect 555848 628156 570748 630134
rect 11447 627028 16257 627560
rect 11524 602620 15728 627028
rect 127134 602620 209843 602887
rect 11524 599835 209843 602620
rect 11524 599642 128662 599835
rect 11524 599336 128666 599642
rect 11524 598416 113136 599336
rect 123468 598478 128666 599336
rect 108928 597880 113136 598416
rect 108932 597130 113128 597880
rect 99600 596241 101510 596540
rect 99600 595229 99968 596241
rect 101172 595760 101510 596241
rect 108932 596048 113130 597130
rect 101172 595530 108250 595760
rect 195468 595706 198174 599835
rect 101172 595229 101510 595530
rect 99600 594870 101510 595229
rect 105246 594999 109064 595176
rect 105246 594371 105428 594999
rect 105928 594998 109064 594999
rect 199624 595075 201786 595464
rect 105928 594371 106086 594998
rect 199624 594836 199918 595075
rect 105246 594176 106086 594371
rect 193894 594818 194254 594828
rect 193894 594768 195036 594818
rect 193894 594396 193984 594768
rect 194164 594396 195036 594768
rect 198410 594582 199918 594836
rect 193894 594336 195036 594396
rect 199624 594383 199918 594582
rect 201314 594383 201786 595075
rect 193894 594330 194254 594336
rect 105246 594174 106084 594176
rect 101706 593988 102292 594128
rect 101706 593552 101805 593988
rect 102177 593894 102292 593988
rect 118078 593977 119138 594148
rect 199624 593982 201786 594383
rect 102177 593666 109064 593894
rect 118078 593822 118287 593977
rect 102177 593552 102292 593666
rect 101706 593388 102292 593552
rect 113380 593410 118287 593822
rect 59644 593272 64808 593382
rect 118078 593285 118287 593410
rect 118979 593285 119138 593977
rect 59644 588280 85874 593272
rect 118078 593102 119138 593285
rect 195328 593438 198370 593568
rect 195328 593214 198366 593438
rect 109016 590868 113190 590870
rect 103178 590356 113190 590868
rect 195326 590356 198366 593214
rect 103178 588470 198366 590356
rect 59644 588264 77050 588280
rect 59644 567110 64808 588264
rect 76034 588188 76042 588264
rect 77982 588198 77992 588280
rect 79332 588198 79342 588280
rect 81855 582541 82253 582561
rect 81855 582489 82149 582541
rect 82201 582489 82253 582541
rect 81855 582471 82253 582489
rect 81855 582419 82149 582471
rect 82201 582419 82253 582471
rect 81855 582401 82253 582419
rect 81855 582349 82149 582401
rect 82201 582349 82253 582401
rect 81855 582331 82253 582349
rect 81855 582279 82149 582331
rect 82201 582279 82253 582331
rect 81855 582261 82253 582279
rect 81855 582209 82149 582261
rect 82201 582209 82253 582261
rect 81855 582140 82253 582209
rect 67536 576169 70924 576498
rect 67536 573493 68035 576169
rect 70583 575038 70924 576169
rect 103178 575038 109600 588470
rect 70583 573493 109600 575038
rect 67536 573188 109600 573493
rect 69072 573186 109600 573188
rect 59649 296487 64803 567110
rect 11848 291333 64803 296487
rect 76000 496004 79845 573186
rect 103178 573184 109600 573186
rect 206791 530472 209843 599835
rect 132927 527420 209843 530472
rect 132927 514865 135979 527420
rect 111402 513445 135979 514865
rect 102551 508083 112669 508299
rect 130965 500489 131015 501088
rect 119495 496004 127955 497268
rect 76000 494706 127955 496004
rect 11848 214140 17002 291333
rect 76000 285077 79845 494706
rect 119495 494704 127955 494706
rect 132927 461897 135979 513445
rect 45054 281232 79845 285077
rect 91209 458845 135979 461897
rect 11848 210248 12422 214140
rect 16570 210248 17002 214140
rect 11848 209892 17002 210248
rect 44859 142718 48899 281232
rect 91209 189279 94261 458845
rect 526360 231511 531111 231516
rect 531804 231511 537519 231516
rect 506865 231484 511616 231489
rect 512309 231484 518024 231489
rect 523210 231484 543816 231511
rect 486810 231452 491561 231457
rect 492254 231452 497969 231457
rect 503715 231452 543816 231484
rect 483655 231242 543816 231452
rect 483655 231178 517975 231242
rect 521803 231178 523479 231242
rect 524683 231178 537431 231242
rect 541323 231178 543816 231242
rect 483655 229028 483927 231178
rect 485131 231114 497879 231178
rect 501771 231114 503959 231178
rect 543499 229974 543816 231178
rect 440718 229020 483927 229028
rect 439606 227234 483927 229020
rect 439606 221804 440342 227234
rect 483655 224662 483927 227234
rect 485131 229657 487063 229974
rect 485131 227234 485451 229657
rect 485131 226062 485450 227234
rect 486810 226062 487063 229657
rect 485131 225802 487063 226062
rect 488267 229657 490135 229974
rect 488267 226062 488605 229657
rect 489766 226062 490135 229657
rect 488267 225802 490135 226062
rect 491275 229657 492503 229974
rect 491275 226062 491561 229657
rect 492254 226062 492503 229657
rect 491275 225802 492503 226062
rect 493707 229657 495447 229910
rect 493707 226062 494049 229657
rect 495075 226062 495447 229657
rect 493707 225802 495447 226062
rect 496587 229657 497879 229974
rect 496587 226062 496870 229657
rect 497638 226062 497879 229657
rect 496587 225802 497879 226062
rect 499083 229646 500567 229974
rect 499083 226062 499433 229646
rect 500230 226062 500567 229646
rect 499083 225802 500567 226062
rect 501771 229657 503959 229974
rect 501771 226062 502025 229657
rect 503715 226062 503959 229657
rect 501771 225802 503959 226062
rect 505227 229689 507095 229974
rect 505227 227266 505506 229689
rect 505227 226094 505505 227266
rect 506865 226094 507095 229689
rect 505227 225866 507095 226094
rect 508299 229689 510167 229974
rect 508299 226094 508660 229689
rect 509821 226094 510167 229689
rect 508299 225866 510167 226094
rect 511371 229689 512535 229974
rect 511371 226094 511616 229689
rect 512309 226094 512535 229689
rect 511371 225866 512535 226094
rect 513739 229689 515479 229974
rect 513739 226094 514104 229689
rect 515130 226094 515479 229689
rect 513739 225866 515479 226094
rect 516683 229689 517975 229974
rect 516683 226094 516925 229689
rect 517693 226094 517975 229689
rect 516683 225866 517975 226094
rect 519115 229678 520663 229974
rect 519115 226094 519488 229678
rect 520285 226094 520663 229678
rect 519115 225866 520663 226094
rect 521803 229689 523479 229974
rect 521803 226094 522080 229689
rect 523210 226094 523479 229689
rect 521803 225866 523479 226094
rect 524683 229716 526615 229974
rect 524683 227293 525001 229716
rect 524683 226121 525000 227293
rect 526360 226121 526615 229716
rect 524683 225866 526615 226121
rect 527819 229716 529687 229974
rect 527819 226121 528155 229716
rect 529316 226121 529687 229716
rect 527819 225866 529687 226121
rect 530827 229716 532055 229974
rect 530827 226121 531111 229716
rect 531804 226121 532055 229716
rect 530827 225866 532055 226121
rect 533259 229716 534999 229974
rect 533259 226121 533599 229716
rect 534625 226121 534999 229716
rect 533259 225866 534999 226121
rect 536139 229716 537431 229974
rect 536139 226121 536420 229716
rect 537188 226121 537431 229716
rect 536139 225866 537431 226121
rect 538635 229705 540119 229974
rect 538635 226121 538983 229705
rect 539780 226121 540119 229705
rect 538635 225866 540119 226121
rect 541323 229716 543816 229974
rect 541323 226121 541575 229716
rect 541323 225866 543793 226121
rect 543499 224726 543793 225866
rect 483655 224534 483991 224662
rect 488267 224534 490135 224662
rect 483655 224470 490135 224534
rect 493707 224470 495447 224662
rect 499083 224598 504023 224662
rect 508299 224598 510167 224662
rect 499083 224534 510167 224598
rect 513739 224534 515479 224662
rect 519115 224598 523543 224662
rect 527819 224598 529687 224726
rect 519115 224534 529687 224598
rect 533259 224534 534999 224726
rect 538635 224534 543793 224726
rect 499083 224470 543793 224534
rect 483655 224326 543793 224470
rect 483655 224299 524298 224326
rect 483655 224267 504243 224299
rect 489766 224233 494049 224267
rect 495075 224249 499433 224267
rect 509821 224265 514104 224299
rect 515130 224281 519488 224299
rect 529316 224292 533599 224326
rect 534625 224308 538983 224326
rect 439606 219622 455414 221804
rect 439606 212928 440342 219622
rect 450906 219346 455414 219622
rect 446975 217275 449725 217437
rect 446975 216711 447310 217275
rect 449474 216711 449725 217275
rect 446975 216630 449725 216711
rect 487570 209172 492321 209177
rect 493014 209172 498729 209177
rect 507395 209172 512146 209177
rect 512839 209172 518554 209177
rect 526906 209172 531657 209177
rect 532350 209172 538065 209177
rect 484415 208901 544362 209172
rect 484415 206748 484676 208901
rect 485880 208837 498692 208901
rect 502520 208837 504516 208901
rect 505720 208837 518468 208901
rect 522360 208837 524036 208901
rect 525176 208837 537988 208901
rect 541880 208837 544362 208901
rect 544056 207697 544362 208837
rect 477046 204954 484676 206748
rect 484415 202385 484676 204954
rect 485880 207377 487812 207697
rect 485880 204954 486211 207377
rect 485880 203782 486210 204954
rect 487570 203782 487812 207377
rect 485880 203525 487812 203782
rect 489016 207377 490884 207697
rect 489016 203782 489365 207377
rect 490526 203782 490884 207377
rect 489016 203525 490884 203782
rect 492088 207377 493252 207697
rect 492088 203782 492321 207377
rect 493014 203782 493252 207377
rect 492088 203525 493252 203782
rect 494456 207377 496196 207633
rect 494456 203782 494809 207377
rect 495835 203782 496196 207377
rect 494456 203525 496196 203782
rect 497336 207377 498692 207697
rect 497336 203782 497630 207377
rect 498398 203782 498692 207377
rect 497336 203525 498692 203782
rect 499832 207366 501380 207697
rect 499832 203782 500193 207366
rect 500990 203782 501380 207366
rect 499832 203525 501380 203782
rect 502520 207377 504516 207697
rect 502520 203782 502785 207377
rect 504240 206748 504516 207377
rect 504237 204954 504516 206748
rect 504240 203782 504516 204954
rect 502520 203525 504516 203782
rect 505720 207377 507652 207697
rect 505720 204954 506036 207377
rect 505720 203782 506035 204954
rect 507395 203782 507652 207377
rect 505720 203525 507652 203782
rect 508856 207377 510724 207697
rect 508856 203782 509190 207377
rect 510351 203782 510724 207377
rect 508856 203525 510724 203782
rect 511864 207377 513092 207697
rect 511864 203782 512146 207377
rect 512839 203782 513092 207377
rect 511864 203525 513092 203782
rect 514296 207377 516036 207633
rect 514296 203782 514634 207377
rect 515660 203782 516036 207377
rect 514296 203525 516036 203782
rect 517176 207377 518468 207697
rect 517176 203782 517455 207377
rect 518223 203782 518468 207377
rect 517176 203525 518468 203782
rect 519672 207366 521156 207697
rect 519672 203782 520018 207366
rect 520815 203782 521156 207366
rect 519672 203525 521156 203782
rect 522360 207377 524036 207697
rect 522360 203782 522610 207377
rect 523751 206748 524036 207377
rect 523748 204954 524036 206748
rect 523751 203782 524036 204954
rect 522360 203525 524036 203782
rect 525240 207377 527172 207697
rect 525240 204954 525547 207377
rect 525240 203782 525546 204954
rect 526906 203782 527172 207377
rect 525240 203525 527172 203782
rect 528312 207377 530244 207697
rect 528312 203782 528701 207377
rect 529862 203782 530244 207377
rect 528312 203525 530244 203782
rect 531384 207377 532612 207697
rect 531384 203782 531657 207377
rect 532350 203782 532612 207377
rect 531384 203525 532612 203782
rect 533752 207377 535492 207633
rect 533752 203782 534145 207377
rect 535171 203782 535492 207377
rect 533752 203525 535492 203782
rect 536696 207377 537988 207697
rect 536696 203782 536966 207377
rect 537734 203782 537988 207377
rect 536696 203525 537988 203782
rect 539192 207366 540676 207697
rect 539192 203782 539529 207366
rect 540326 203782 540676 207366
rect 539192 203525 540676 203782
rect 541880 207377 544362 207697
rect 541880 203782 542121 207377
rect 541880 203525 544339 203782
rect 543992 202385 544339 203525
rect 484415 202257 484740 202385
rect 489016 202257 490884 202385
rect 484415 202193 490884 202257
rect 494456 202193 496196 202385
rect 499832 202257 504580 202385
rect 508856 202257 510724 202385
rect 499832 202193 510724 202257
rect 514296 202193 516036 202385
rect 519672 202257 524100 202385
rect 528312 202257 530244 202385
rect 519672 202193 530244 202257
rect 533752 202193 535492 202385
rect 539192 202193 544339 202385
rect 484415 201987 544339 202193
rect 490526 201953 494809 201987
rect 495835 201969 500193 201987
rect 510351 201968 514634 201987
rect 515660 201969 520018 201987
rect 529862 201968 534145 201987
rect 535171 201969 539529 201987
rect 74531 189268 94261 189279
rect 74531 169255 109382 189268
rect 64648 167087 66472 167354
rect 64648 165691 64951 167087
rect 66155 167052 66472 167087
rect 66155 165730 70790 167052
rect 66155 165691 66472 165730
rect 64648 165362 66472 165691
rect 70546 165166 70790 165730
rect 74532 165494 88626 169255
rect 70546 164956 74109 165166
rect 67264 164704 74103 164914
rect 64846 163914 66490 164046
rect 67264 163914 67872 164704
rect 73858 164624 74110 164668
rect 64846 163893 67872 163914
rect 64846 162881 65091 163893
rect 66295 162881 67872 163893
rect 64846 162876 67872 162881
rect 68542 164464 74110 164624
rect 64846 162704 66490 162876
rect 65048 159194 66406 159346
rect 68542 159194 69524 164464
rect 65048 159173 69524 159194
rect 65048 158225 65247 159173
rect 66195 158225 69524 159173
rect 65048 158206 69524 158225
rect 65048 158030 66406 158206
rect 74617 142718 88744 158134
rect 44859 138967 88744 142718
rect 44859 41811 48952 138967
rect 106942 64678 109354 169255
rect 559502 168256 566449 628156
rect 559502 164498 566490 168256
rect 469924 161309 566490 164498
rect 469924 161301 565502 161309
rect 469924 150327 473121 161301
rect 469918 147935 473468 150327
rect 469924 147130 473468 147935
rect 473695 144071 473768 144142
rect 471847 143971 471940 144005
rect 471847 143962 471923 143971
rect 469535 142212 577709 142350
rect 469535 141095 575923 142212
rect 469523 140624 575923 141095
rect 577447 140624 577709 142212
rect 469523 140357 577709 140624
rect 106942 63026 107280 64678
rect 109060 63026 109354 64678
rect 106942 62650 109354 63026
rect 92276 61824 94497 61881
rect 102515 61486 106764 62038
rect 106323 58322 106764 61486
rect 106116 58204 107054 58322
rect 106116 57640 106287 58204
rect 106915 57640 107054 58204
rect 106116 57508 107054 57640
rect 81326 54740 81746 54887
rect 81326 54432 81406 54740
rect 81650 54432 81746 54740
rect 81326 54316 81746 54432
rect 99879 54864 100589 55041
rect 99879 54236 99937 54864
rect 100437 54236 100589 54864
rect 99879 54133 100589 54236
rect 99879 54132 100588 54133
rect 44859 39702 100481 41811
<< via1 >>
rect 11934 627560 15698 631068
rect 558070 630134 568234 644394
rect 99968 595229 101172 596241
rect 105428 594371 105928 594999
rect 193984 594396 194164 594768
rect 199918 594383 201314 595075
rect 101805 593552 102177 593988
rect 118287 593285 118979 593977
rect 82149 582489 82201 582541
rect 82149 582419 82201 582471
rect 82149 582349 82201 582401
rect 82149 582279 82201 582331
rect 82149 582209 82201 582261
rect 68035 573493 70583 576169
rect 124969 500569 125021 500621
rect 125129 500569 125181 500621
rect 125208 500569 125260 500621
rect 125288 500569 125340 500621
rect 124969 500499 125021 500551
rect 125048 500499 125100 500551
rect 125129 500499 125181 500551
rect 125208 500499 125260 500551
rect 125288 500499 125340 500551
rect 124969 500429 125021 500481
rect 125048 500429 125100 500481
rect 125129 500429 125181 500481
rect 125208 500429 125260 500481
rect 125288 500429 125340 500481
rect 12422 210248 16570 214140
rect 517975 231178 521803 231242
rect 523479 231178 524683 231242
rect 537431 231178 541323 231242
rect 483927 231114 485131 231178
rect 497879 231114 501771 231178
rect 503959 231114 543499 231178
rect 483927 229974 543499 231114
rect 483927 225802 485131 229974
rect 487063 225802 488267 229974
rect 490135 225802 491275 229974
rect 492503 229910 496587 229974
rect 492503 225802 493707 229910
rect 495447 225802 496587 229910
rect 497879 225802 499083 229974
rect 500567 225802 501771 229974
rect 503959 225866 505227 229974
rect 507095 225866 508299 229974
rect 510167 225866 511371 229974
rect 512535 225866 513739 229974
rect 515479 225866 516683 229974
rect 517975 225866 519115 229974
rect 520663 225866 521803 229974
rect 523479 225866 524683 229974
rect 526615 225866 527819 229974
rect 529687 225866 530827 229974
rect 532055 225866 533259 229974
rect 534999 225866 536139 229974
rect 537431 225866 538635 229974
rect 540119 225866 541323 229974
rect 503959 225802 543499 225866
rect 483927 224726 543499 225802
rect 483927 224662 527819 224726
rect 483991 224534 488267 224662
rect 490135 224470 493707 224662
rect 495447 224470 499083 224662
rect 504023 224598 508299 224662
rect 510167 224534 513739 224662
rect 515479 224534 519115 224662
rect 523543 224598 527819 224662
rect 529687 224534 533259 224726
rect 534999 224534 538635 224726
rect 447310 216711 449474 217275
rect 484676 208837 485880 208901
rect 498692 208837 502520 208901
rect 504516 208837 505720 208901
rect 518468 208837 522360 208901
rect 524036 208837 525176 208901
rect 537988 208837 541880 208901
rect 484676 207697 544056 208837
rect 484676 203525 485880 207697
rect 487812 203525 489016 207697
rect 490884 203525 492088 207697
rect 493252 207633 497336 207697
rect 493252 203525 494456 207633
rect 496196 203525 497336 207633
rect 498692 203525 499832 207697
rect 501380 203525 502520 207697
rect 504516 203525 505720 207697
rect 507652 203525 508856 207697
rect 510724 203525 511864 207697
rect 513092 207633 517176 207697
rect 513092 203525 514296 207633
rect 516036 203525 517176 207633
rect 518468 203525 519672 207697
rect 521156 203525 522360 207697
rect 524036 203525 525240 207697
rect 527172 203525 528312 207697
rect 530244 203525 531384 207697
rect 532612 207633 536696 207697
rect 532612 203525 533752 207633
rect 535492 203525 536696 207633
rect 537988 203525 539192 207697
rect 540676 203525 541880 207697
rect 484676 202385 543992 203525
rect 484740 202257 489016 202385
rect 490884 202193 494456 202385
rect 496196 202193 499832 202385
rect 504580 202257 508856 202385
rect 510724 202193 514296 202385
rect 516036 202193 519672 202385
rect 524100 202257 528312 202385
rect 530244 202193 533752 202385
rect 535492 202193 539192 202385
rect 64951 165691 66155 167087
rect 65091 162881 66295 163893
rect 65247 158225 66195 159173
rect 475328 142703 475380 142755
rect 475409 142704 475461 142756
rect 475490 142704 475542 142756
rect 475571 142704 475623 142756
rect 475652 142703 475704 142755
rect 475328 142622 475380 142674
rect 475409 142623 475461 142675
rect 475491 142621 475543 142673
rect 475571 142622 475623 142674
rect 475652 142622 475704 142674
rect 575923 140624 577447 142212
rect 107280 63026 109060 64678
rect 106287 57640 106915 58204
rect 81406 54432 81650 54740
rect 99937 54236 100437 54864
<< metal2 >>
rect 566589 690166 571598 690911
rect 566589 688210 567317 690166
rect 502484 686270 567317 688210
rect 570973 686270 571598 690166
rect 502484 685378 571598 686270
rect 11447 631068 16257 631627
rect 11447 627560 11934 631068
rect 15698 627560 16257 631068
rect 11447 627028 16257 627560
rect 67484 626039 73886 626978
rect 67484 621023 68344 626039
rect 72960 621023 73886 626039
rect 67484 620234 73886 621023
rect 69030 599046 72102 620234
rect 118068 614830 125192 616048
rect 118068 610214 119475 614830
rect 123611 610214 125192 614830
rect 118068 608944 125192 610214
rect 69004 599044 103712 599046
rect 69004 597710 103912 599044
rect 72244 597698 103912 597710
rect 99600 596248 101510 596540
rect 99600 595232 99947 596248
rect 101203 595232 101510 596248
rect 99600 595229 99968 595232
rect 101172 595229 101510 595232
rect 99600 594870 101510 595229
rect 103116 595178 103912 597698
rect 118072 595908 119138 608944
rect 120316 597866 120744 597870
rect 122238 597866 122710 598248
rect 120316 597272 122710 597866
rect 103116 594999 106088 595178
rect 103116 594812 105428 594999
rect 103108 594371 105428 594812
rect 105928 594371 106088 594999
rect 103108 594174 106088 594371
rect 118072 594858 119140 595908
rect 103116 594170 103912 594174
rect 33184 593988 102292 594128
rect 118072 594122 119142 594858
rect 33184 593711 101805 593988
rect 33184 591815 33649 593711
rect 36025 593552 101805 593711
rect 102177 593552 102292 593988
rect 36025 592948 102292 593552
rect 118078 593977 119138 594122
rect 118078 593285 118287 593977
rect 118979 593285 119138 593977
rect 118078 593102 119138 593285
rect 36025 591815 36516 592948
rect 33184 591326 36516 591815
rect 82132 582541 83318 582560
rect 82132 582489 82149 582541
rect 82201 582489 83318 582541
rect 82132 582471 83318 582489
rect 82132 582419 82149 582471
rect 82201 582419 83318 582471
rect 82132 582401 83318 582419
rect 82132 582349 82149 582401
rect 82201 582349 83318 582401
rect 82132 582331 83318 582349
rect 82132 582279 82149 582331
rect 82201 582279 83318 582331
rect 82132 582261 83318 582279
rect 82132 582209 82149 582261
rect 82201 582209 83318 582261
rect 82132 582008 83318 582209
rect 120316 581168 120744 597272
rect 122238 596856 122710 597272
rect 121470 595746 122642 596248
rect 121472 594390 121898 595746
rect 199624 595077 201786 595464
rect 199624 595075 199948 595077
rect 201284 595075 201786 595077
rect 193894 594770 194254 594828
rect 193894 594394 193966 594770
rect 194182 594394 194254 594770
rect 121472 591320 121900 594390
rect 193894 594330 194254 594394
rect 199624 594383 199918 595075
rect 201314 594383 201786 595075
rect 199624 594381 199948 594383
rect 201284 594381 201786 594383
rect 199624 593982 201786 594381
rect 131577 593730 131983 593788
rect 131577 593674 131739 593730
rect 131795 593674 131821 593730
rect 131877 593674 131983 593730
rect 131577 593623 131983 593674
rect 122284 592349 122656 592350
rect 122284 591973 122322 592349
rect 122618 591973 122656 592349
rect 122284 591972 122656 591973
rect 121472 590818 122708 591320
rect 121472 581525 121900 590818
rect 121472 581389 121530 581525
rect 121826 581389 121900 581525
rect 121472 581312 121900 581389
rect 11450 576169 70908 576520
rect 82502 576418 82576 581135
rect 120316 581032 120426 581168
rect 120642 581032 120744 581168
rect 120316 580976 120744 581032
rect 11450 574778 68035 576169
rect 11432 574314 68035 574778
rect 11432 571058 11957 574314
rect 15613 573493 68035 574314
rect 70583 573493 70908 576169
rect 15613 573187 70908 573493
rect 15613 571058 20780 573187
rect 45852 572555 47266 572810
rect 45852 571379 46120 572555
rect 47056 572554 47266 572555
rect 47056 572089 91288 572554
rect 47056 571873 90983 572089
rect 91199 571873 91288 572089
rect 47056 571706 91288 571873
rect 47056 571379 47266 571706
rect 45852 571140 47266 571379
rect 50732 571251 90778 571342
rect 11432 570648 20780 571058
rect 50732 571080 90491 571251
rect 11432 570604 16254 570648
rect 50732 569824 50950 571080
rect 51726 571035 90491 571080
rect 90707 571035 90778 571251
rect 51726 570550 90778 571035
rect 51726 569824 52016 570550
rect 50732 569574 52016 569824
rect 55500 569835 90162 569930
rect 55500 569619 89871 569835
rect 90087 569619 90162 569835
rect 55500 569523 90162 569619
rect 55500 568267 55842 569523
rect 56858 568866 90162 569523
rect 56858 568267 57226 568866
rect 55500 567942 57226 568267
rect 502484 243672 505316 685378
rect 566589 685375 571598 685378
rect 566486 682685 571541 682981
rect 438649 243249 505316 243672
rect 508167 682580 571541 682685
rect 508167 679853 567033 682580
rect 11848 214142 17002 215261
rect 11848 214140 12428 214142
rect 16564 214140 17002 214142
rect 11848 210248 12422 214140
rect 16570 210248 17002 214140
rect 438649 212496 438959 243249
rect 508167 242564 510999 679853
rect 566486 678444 567033 679853
rect 571009 678444 571541 682580
rect 566486 677985 571541 678444
rect 555848 644394 570748 646373
rect 555848 630134 558070 644394
rect 568234 630134 570748 644394
rect 555848 628156 570748 630134
rect 445402 241981 510999 242564
rect 513520 583422 515922 583674
rect 513520 582166 514045 583422
rect 515381 582166 515922 583422
rect 513520 242801 515922 582166
rect 542474 554928 548169 555589
rect 542474 541592 543521 554928
rect 546937 541592 548169 554928
rect 518813 494718 521215 494973
rect 518813 493302 519175 494718
rect 520831 493302 521215 494718
rect 445402 214771 445873 241981
rect 513520 241483 515923 242801
rect 456294 241076 515923 241483
rect 456294 240908 515922 241076
rect 446975 217275 449725 217437
rect 446975 216711 447310 217275
rect 449474 216711 449725 217275
rect 456294 216808 456848 240908
rect 513520 240904 515421 240908
rect 518813 239849 521215 493302
rect 446975 216630 449725 216711
rect 455064 216618 456848 216808
rect 458300 239152 521215 239849
rect 524067 450040 526469 450426
rect 524067 448464 524359 450040
rect 526095 448464 526469 450040
rect 458300 239151 519744 239152
rect 458300 216619 458937 239151
rect 524067 237885 526469 448464
rect 460198 237274 526469 237885
rect 460198 237273 525447 237274
rect 455064 216617 456485 216618
rect 458300 215580 458854 216619
rect 455857 215404 458854 215580
rect 445402 214300 446166 214771
rect 445695 213195 446166 214300
rect 438649 212376 441421 212496
rect 438649 212186 441422 212376
rect 455857 212185 456033 215404
rect 458300 215401 458854 215404
rect 460198 214833 460811 237273
rect 542474 233313 548169 541592
rect 553614 405600 556971 405945
rect 553614 403144 554301 405600
rect 556437 403144 556971 405600
rect 553614 402603 556971 403144
rect 553610 402563 556971 402603
rect 542475 233292 548167 233313
rect 542475 231511 542887 233292
rect 523241 231484 542887 231511
rect 503746 231452 542887 231484
rect 483691 231292 542887 231452
rect 483691 231242 523447 231292
rect 524623 231242 526647 231292
rect 483691 231212 517975 231242
rect 521803 231212 523447 231242
rect 524683 231212 526647 231242
rect 530703 231212 532007 231292
rect 536063 231242 542887 231292
rect 536063 231212 537431 231242
rect 541323 231212 542887 231242
rect 483691 224516 483927 231212
rect 485103 231178 487127 231212
rect 485131 231132 487127 231178
rect 491183 231132 492487 231212
rect 496543 231132 497847 231212
rect 501663 231178 504007 231212
rect 501771 231132 503959 231178
rect 547663 230116 548167 233292
rect 543503 230036 548167 230116
rect 485131 229657 487063 229956
rect 485131 226044 485486 229657
rect 486785 226044 487063 229657
rect 485131 225802 487063 226044
rect 488267 229657 490007 229956
rect 488267 226080 488580 229657
rect 489755 226080 490007 229657
rect 488267 225802 490007 226080
rect 491275 229640 492487 229956
rect 491275 226044 491550 229640
rect 492237 226044 492487 229640
rect 491275 225802 492487 226044
rect 493707 229657 495367 229910
rect 493707 226070 494032 229657
rect 495089 226070 495367 229657
rect 493707 225802 495367 226070
rect 496587 229648 497847 229956
rect 496587 226044 496884 229648
rect 497585 226044 497847 229648
rect 496587 225802 497847 226044
rect 499083 229657 500567 229956
rect 499083 226044 499380 229657
rect 500245 226044 500567 229657
rect 499083 225802 500567 226044
rect 501771 229657 503959 229956
rect 501771 226044 502040 229657
rect 502650 229652 503959 229657
rect 503746 226044 503959 229652
rect 501771 225852 503959 226044
rect 505227 229689 507095 229974
rect 505227 226076 505541 229689
rect 506840 226076 507095 229689
rect 505227 225866 507095 226076
rect 508303 229689 510087 229974
rect 508303 226112 508635 229689
rect 509810 226112 510087 229689
rect 508303 225866 510087 226112
rect 511371 229672 512535 229974
rect 511371 226076 511605 229672
rect 512292 226076 512535 229672
rect 511371 225866 512535 226076
rect 501771 225802 503927 225852
rect 513739 229689 515447 229974
rect 513739 226102 514087 229689
rect 515144 226102 515447 229689
rect 513739 225866 515447 226102
rect 516683 229680 517927 229974
rect 516683 226076 516939 229680
rect 517640 226076 517927 229680
rect 516683 225866 517927 226076
rect 519115 229689 520567 229974
rect 519115 226076 519435 229689
rect 520300 226076 520567 229689
rect 519115 225866 520567 226076
rect 521803 229689 523447 229974
rect 521803 226076 522095 229689
rect 522705 229684 523447 229689
rect 523241 226076 523447 229684
rect 521803 225866 523447 226076
rect 524683 229716 526615 229974
rect 524683 226103 525036 229716
rect 526335 226103 526615 229716
rect 524683 225866 526615 226103
rect 527823 229716 529527 229974
rect 527823 226139 528130 229716
rect 529305 226139 529527 229716
rect 527823 225866 529527 226139
rect 530827 229699 532007 229974
rect 530827 226103 531100 229699
rect 531787 226103 532007 229699
rect 530827 225866 532007 226103
rect 533259 229716 534887 229974
rect 533259 226129 533582 229716
rect 534639 226129 534887 229716
rect 533259 225866 534887 226129
rect 536139 229707 537431 229974
rect 536139 226103 536434 229707
rect 537135 226103 537431 229707
rect 536139 225866 537431 226103
rect 543499 229974 548167 230036
rect 538635 229716 540087 229974
rect 538635 226103 538930 229716
rect 539795 226103 540087 229716
rect 538635 225866 540087 226103
rect 541323 229716 548167 229974
rect 541323 226103 541590 229716
rect 542200 229711 548167 229716
rect 542475 229677 548167 229711
rect 541323 225866 543787 226103
rect 543499 225772 543787 225866
rect 543503 224596 543787 225772
rect 503903 224516 510087 224596
rect 513739 224534 515447 224596
rect 519115 224534 529527 224596
rect 533259 224534 534887 224596
rect 538635 224534 543787 224596
rect 513663 224516 515447 224534
rect 519103 224516 529527 224534
rect 533183 224516 534887 224534
rect 538543 224516 543787 224534
rect 483691 224436 490007 224516
rect 493707 224470 495447 224516
rect 499083 224470 543787 224516
rect 493663 224436 543787 224470
rect 483691 224308 543787 224436
rect 483691 224281 524292 224308
rect 483691 224249 504237 224281
rect 455440 212001 456033 212185
rect 456225 214659 460752 214833
rect 456225 214657 460630 214659
rect 456225 210940 456401 214657
rect 455408 210764 456401 210940
rect 11848 210246 12428 210248
rect 16564 210246 17002 210248
rect 11848 209892 17002 210246
rect 553610 210111 556967 402563
rect 559120 359429 562476 359447
rect 559120 359157 562477 359429
rect 559120 356701 559509 359157
rect 562125 356701 562477 359157
rect 553610 209215 556956 210111
rect 544141 209172 556956 209215
rect 484451 208941 556956 209172
rect 484451 202245 484661 208941
rect 485837 208901 487861 208941
rect 485880 208861 487861 208901
rect 491917 208861 493221 208941
rect 497277 208901 504501 208941
rect 505677 208901 507701 208941
rect 497277 208861 498692 208901
rect 502520 208861 504501 208901
rect 505720 208861 507701 208901
rect 511757 208861 513061 208941
rect 517117 208901 524021 208941
rect 517117 208861 518468 208901
rect 522360 208861 524021 208901
rect 525197 208861 527221 208941
rect 531277 208861 532581 208941
rect 536637 208901 556956 208941
rect 536637 208861 537988 208901
rect 541880 208861 556956 208901
rect 544077 207685 556956 208861
rect 485880 207377 487812 207685
rect 485880 203764 486246 207377
rect 487545 203764 487812 207377
rect 485880 203525 487812 203764
rect 489037 207377 490741 207685
rect 489037 203800 489340 207377
rect 490515 203800 490741 207377
rect 489037 203525 490741 203800
rect 492088 207360 493221 207685
rect 492088 203764 492310 207360
rect 492997 203764 493221 207360
rect 492088 203525 493221 203764
rect 494456 207377 496101 207633
rect 494456 203790 494792 207377
rect 495849 203790 496101 207377
rect 494456 203525 496101 203790
rect 497336 207368 498661 207685
rect 497336 203764 497644 207368
rect 498345 203764 498661 207368
rect 497336 203525 498661 203764
rect 499832 207377 501301 207685
rect 499832 203764 500140 207377
rect 501005 203764 501301 207377
rect 499832 203525 501301 203764
rect 502520 207377 504501 207685
rect 502520 203764 502800 207377
rect 503410 207372 504501 207377
rect 504276 203764 504501 207372
rect 502520 203525 504501 203764
rect 505720 207377 507652 207685
rect 505720 203764 506071 207377
rect 507370 203764 507652 207377
rect 505720 203525 507652 203764
rect 508877 207377 510581 207685
rect 508877 203800 509165 207377
rect 510340 203800 510581 207377
rect 508877 203525 510581 203800
rect 511864 207360 513061 207685
rect 511864 203764 512135 207360
rect 512822 203764 513061 207360
rect 511864 203525 513061 203764
rect 514296 207377 515941 207633
rect 514296 203790 514617 207377
rect 515674 203790 515941 207377
rect 514296 203525 515941 203790
rect 517176 207368 518421 207685
rect 517176 203764 517469 207368
rect 518170 203764 518421 207368
rect 517176 203525 518421 203764
rect 519672 207377 521141 207685
rect 519672 203764 519965 207377
rect 520830 203764 521141 207377
rect 519672 203525 521141 203764
rect 522360 207377 524021 207685
rect 522360 203764 522625 207377
rect 523235 207372 524021 207377
rect 523787 203764 524021 207372
rect 522360 203525 524021 203764
rect 525240 207377 527172 207685
rect 525240 203764 525582 207377
rect 526881 203764 527172 207377
rect 525240 203525 527172 203764
rect 528317 207377 530101 207685
rect 528317 203800 528676 207377
rect 529851 203800 530101 207377
rect 528317 203525 530101 203800
rect 531384 207360 532581 207685
rect 531384 203764 531646 207360
rect 532333 203764 532581 207360
rect 531384 203525 532581 203764
rect 533757 207377 535461 207633
rect 533757 203790 534128 207377
rect 535185 203790 535461 207377
rect 533757 203525 535461 203790
rect 536696 207368 537941 207685
rect 536696 203764 536980 207368
rect 537681 203764 537941 207368
rect 536696 203525 537941 203764
rect 539192 207377 540661 207685
rect 539192 203764 539476 207377
rect 540341 203764 540661 207377
rect 539192 203525 540661 203764
rect 541880 207398 556956 207685
rect 541880 207377 544362 207398
rect 541880 203764 542136 207377
rect 542746 207372 544362 207377
rect 559120 203796 562477 356701
rect 566807 316082 570323 316401
rect 566807 313226 567174 316082
rect 569870 313226 570323 316082
rect 544162 203764 562478 203796
rect 541880 203525 562478 203764
rect 543992 203421 562478 203525
rect 484451 202165 490741 202245
rect 494456 202193 496101 202245
rect 499832 202193 510581 202245
rect 514296 202193 515941 202245
rect 519672 202193 530101 202245
rect 543997 202245 562478 203421
rect 494397 202165 496101 202193
rect 499757 202165 510581 202193
rect 514237 202165 515941 202193
rect 519597 202165 530101 202193
rect 533757 202165 535461 202245
rect 539192 202193 562478 202245
rect 539117 202165 562478 202193
rect 484451 201979 562478 202165
rect 484451 201969 544333 201979
rect 64648 167097 66472 167354
rect 64648 167087 64965 167097
rect 66141 167087 66472 167097
rect 64648 165691 64951 167087
rect 66155 165691 66472 167087
rect 64648 165681 64965 165691
rect 66141 165681 66472 165691
rect 64648 165362 66472 165681
rect 89748 164941 92640 165382
rect 84545 164742 85468 164760
rect 89760 164578 90272 164808
rect 64846 163895 66490 164046
rect 64846 163893 65105 163895
rect 66281 163893 66490 163895
rect 64846 162881 65091 163893
rect 66295 162881 66490 163893
rect 64846 162879 65105 162881
rect 66281 162879 66490 162881
rect 64846 162704 66490 162879
rect 65048 159173 66406 159346
rect 65048 158225 65247 159173
rect 66195 158225 66406 159173
rect 65048 158030 66406 158225
rect 89783 151824 90078 164578
rect 48099 150415 90078 151824
rect 48099 72153 50125 150415
rect 92107 149214 92640 164941
rect 566807 160868 570323 313226
rect 52630 147519 92640 149214
rect 445889 157352 570323 160868
rect 572627 270712 577086 271155
rect 572627 268416 573278 270712
rect 576374 268416 577086 270712
rect 9453 70127 50125 72153
rect 9453 38985 11479 70127
rect 52634 66884 54574 147519
rect 9453 37569 9845 38985
rect 11021 37569 11479 38985
rect 9453 37223 11479 37569
rect 14472 64944 54574 66884
rect 14472 18084 16412 64944
rect 106942 64680 109354 64999
rect 106942 64678 107302 64680
rect 109038 64678 109354 64680
rect 106942 63026 107280 64678
rect 109060 63026 109354 64678
rect 106942 63024 107302 63026
rect 109038 63024 109354 63026
rect 106942 62650 109354 63024
rect 106116 58204 107054 58322
rect 106116 57640 106287 58204
rect 106915 57640 107054 58204
rect 106116 57508 107054 57640
rect 99879 54995 101295 55041
rect 7314 17702 16412 18084
rect 7314 16446 7605 17702
rect 8621 16446 16412 17702
rect 7314 16144 16412 16446
rect 78161 54740 81746 54887
rect 78161 54432 81406 54740
rect 81650 54432 81746 54740
rect 78161 54261 81746 54432
rect 99879 54864 103541 54995
rect 78161 17451 79781 54261
rect 99879 54236 99937 54864
rect 100437 54236 103541 54864
rect 99879 54137 103541 54236
rect 99879 54133 101295 54137
rect 102683 22578 103541 54137
rect 445889 22578 449405 157352
rect 572627 154868 577086 268416
rect 102683 19062 449405 22578
rect 451648 150409 577086 154868
rect 451648 17451 456107 150409
rect 475058 147348 476380 147408
rect 475058 147292 475421 147348
rect 475477 147292 475521 147348
rect 475577 147292 475621 147348
rect 475677 147292 475721 147348
rect 475777 147292 475821 147348
rect 475877 147292 475921 147348
rect 475977 147292 476021 147348
rect 476077 147292 476121 147348
rect 476177 147292 476380 147348
rect 475058 147249 476380 147292
rect 78161 12992 456107 17451
rect 457701 146941 465227 147119
rect 477118 147026 567690 147626
rect 457701 6399 458175 146941
rect 458720 146700 465235 146878
rect 458720 9716 459261 146700
rect 464944 145083 465322 145138
rect 464944 144867 465021 145083
rect 465237 144867 465322 145083
rect 464944 144822 465322 144867
rect 459942 144667 460412 144668
rect 459942 144489 465243 144667
rect 459942 13258 460412 144489
rect 476958 144337 564247 145086
rect 463628 143952 465233 144130
rect 463628 140866 464123 143952
rect 465010 143568 465248 143600
rect 465010 143432 465056 143568
rect 465192 143432 465248 143568
rect 465010 143402 465248 143432
rect 464874 143086 465390 143148
rect 464874 142790 464971 143086
rect 465267 142790 465390 143086
rect 464874 142712 465390 142790
rect 475247 142758 475823 142901
rect 475247 142702 475326 142758
rect 475382 142702 475407 142758
rect 475463 142702 475488 142758
rect 475544 142702 475569 142758
rect 475625 142702 475650 142758
rect 475706 142702 475823 142758
rect 475247 142676 475823 142702
rect 475247 142620 475326 142676
rect 475382 142620 475407 142676
rect 475463 142620 475488 142676
rect 475544 142620 475569 142676
rect 475625 142620 475650 142676
rect 475706 142620 475823 142676
rect 475247 142526 475823 142620
rect 463628 140864 464638 140866
rect 463628 140862 465038 140864
rect 465216 140862 466306 140864
rect 463628 140632 466306 140862
rect 463628 139388 464802 140632
rect 464550 139376 464802 139388
rect 466058 139376 466306 140632
rect 464550 139108 466306 139376
rect 563416 50018 564246 144337
rect 567040 94255 567690 147026
rect 575630 142212 577709 142436
rect 575630 142206 575923 142212
rect 577447 142206 577709 142212
rect 575630 140630 575897 142206
rect 577473 140630 577709 142206
rect 575630 140624 575923 140630
rect 577447 140624 577709 140630
rect 575630 140357 577709 140624
rect 567040 93799 567131 94255
rect 567587 93799 567690 94255
rect 567040 93708 567690 93799
rect 563194 49782 564398 50018
rect 563194 48766 563422 49782
rect 564118 48766 564398 49782
rect 563194 48556 564398 48766
rect 459942 12922 461676 13258
rect 459942 12226 460306 12922
rect 461322 12226 461676 12922
rect 459942 11886 461676 12226
rect 458720 9293 460749 9716
rect 458720 8037 459108 9293
rect 460364 8037 460749 9293
rect 458720 7710 460749 8037
rect 457696 5288 460059 6399
rect 457696 3792 458125 5288
rect 459461 3792 460059 5288
rect 457696 3274 460059 3792
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 567317 686270 570973 690166
rect 11948 627566 15684 631062
rect 68344 621023 72960 626039
rect 119475 610214 123611 614830
rect 99947 596241 101203 596248
rect 99947 595232 99968 596241
rect 99968 595232 101172 596241
rect 101172 595232 101203 596241
rect 33649 591815 36025 593711
rect 199948 595075 201284 595077
rect 131129 594412 131185 594468
rect 131210 594412 131266 594468
rect 131292 594412 131348 594468
rect 131373 594412 131429 594468
rect 131454 594412 131510 594468
rect 193966 594768 194182 594770
rect 193966 594396 193984 594768
rect 193984 594396 194164 594768
rect 194164 594396 194182 594768
rect 193966 594394 194182 594396
rect 131129 594330 131185 594386
rect 131210 594330 131266 594386
rect 131292 594330 131348 594386
rect 131373 594330 131429 594386
rect 131454 594330 131510 594386
rect 199948 594383 201284 595075
rect 199948 594381 201284 594383
rect 131739 593674 131795 593730
rect 131821 593674 131877 593730
rect 122322 591973 122618 592349
rect 121530 581389 121826 581525
rect 120426 581032 120642 581168
rect 11957 571058 15613 574314
rect 46120 571379 47056 572555
rect 90983 571873 91199 572089
rect 50950 569824 51726 571080
rect 90491 571035 90707 571251
rect 89871 569619 90087 569835
rect 55842 568267 56858 569523
rect 124952 499891 125008 499947
rect 125062 499892 125118 499948
rect 125282 499892 125338 499948
rect 12428 214140 16564 214142
rect 12428 210248 16564 214140
rect 567033 678444 571009 682580
rect 558084 630156 568220 644372
rect 514045 582166 515381 583422
rect 543521 541592 546937 554928
rect 519175 493302 520831 494718
rect 447324 216725 449460 217261
rect 524359 448464 526095 450040
rect 554301 403144 556437 405600
rect 523447 231242 524623 231292
rect 523447 231212 523479 231242
rect 523479 231212 524623 231242
rect 526647 231212 530703 231292
rect 532007 231212 536063 231292
rect 542887 231212 547663 233292
rect 483927 231178 485103 231212
rect 483927 231132 485103 231178
rect 487127 231132 491183 231212
rect 492487 231132 496543 231212
rect 497847 231178 501663 231212
rect 504007 231178 517975 231212
rect 517975 231178 521803 231212
rect 521803 231178 523479 231212
rect 523479 231178 524683 231212
rect 524683 231178 537431 231212
rect 537431 231178 541323 231212
rect 541323 231178 547663 231212
rect 497847 231132 497879 231178
rect 497879 231132 501663 231178
rect 504007 231132 543499 231178
rect 483927 231114 485131 231132
rect 485131 231114 497879 231132
rect 497879 231114 501771 231132
rect 501771 231114 503959 231132
rect 503959 231114 543499 231132
rect 483927 230036 543499 231114
rect 543499 230116 547663 231178
rect 543499 230036 543503 230116
rect 483927 229974 505183 230036
rect 507127 229974 508303 230036
rect 510087 229974 511183 230036
rect 483927 229956 485131 229974
rect 485131 229956 487063 229974
rect 487063 229956 488267 229974
rect 488267 229956 490135 229974
rect 490135 229956 491275 229974
rect 491275 229956 492503 229974
rect 492503 229956 496587 229974
rect 496587 229956 497879 229974
rect 497879 229956 499083 229974
rect 499083 229956 500567 229974
rect 500567 229956 501771 229974
rect 501771 229956 503959 229974
rect 503959 229956 505183 229974
rect 483927 225692 485103 229956
rect 487127 225692 488223 229956
rect 490007 225802 490135 229956
rect 490135 225802 491183 229956
rect 492487 225802 492503 229956
rect 492503 225802 493663 229956
rect 495367 229910 496543 229956
rect 495367 225802 495447 229910
rect 495447 225802 496543 229910
rect 497847 225802 497879 229956
rect 497879 225802 499023 229956
rect 490007 225692 491183 225802
rect 492487 225692 493663 225802
rect 495367 225692 496543 225802
rect 497847 225692 499023 225802
rect 500567 225692 501663 229956
rect 504007 225852 505183 229956
rect 507127 225866 508299 229974
rect 508299 225866 508303 229974
rect 510087 225866 510167 229974
rect 510167 225866 511183 229974
rect 503927 225802 503959 225852
rect 503959 225802 505183 225852
rect 503927 225772 505183 225802
rect 507127 225772 508303 225866
rect 510087 225772 511183 225866
rect 512567 225772 513663 230036
rect 515447 229974 516543 230036
rect 517927 229974 519103 230036
rect 520567 229974 521743 230036
rect 523447 229974 524623 230036
rect 526647 229974 527823 230036
rect 529527 229974 530703 230036
rect 532007 229974 533183 230036
rect 534887 229974 536063 230036
rect 515447 225866 515479 229974
rect 515479 225866 516543 229974
rect 517927 225866 517975 229974
rect 517975 225866 519103 229974
rect 520567 225866 520663 229974
rect 520663 225866 521743 229974
rect 523447 225866 523479 229974
rect 523479 225866 524623 229974
rect 526647 225866 527819 229974
rect 527819 225866 527823 229974
rect 529527 225866 529687 229974
rect 529687 225866 530703 229974
rect 532007 225866 532055 229974
rect 532055 225866 533183 229974
rect 534887 225866 534999 229974
rect 534999 225866 536063 229974
rect 515447 225772 516543 225866
rect 517927 225772 519103 225866
rect 520567 225772 521743 225866
rect 523447 225772 524623 225866
rect 526647 225772 527823 225866
rect 529527 225772 530703 225866
rect 532007 225772 533183 225866
rect 534887 225772 536063 225866
rect 537447 225772 538543 230036
rect 540087 229974 541263 230036
rect 540087 225866 540119 229974
rect 540119 225866 541263 229974
rect 540087 225772 541263 225866
rect 503927 225692 543499 225772
rect 483927 224726 543499 225692
rect 543499 224726 543503 225772
rect 483927 224662 527819 224726
rect 483927 224534 483991 224662
rect 483991 224534 488267 224662
rect 488267 224534 490135 224662
rect 483927 224516 490135 224534
rect 490135 224516 493707 224662
rect 493707 224516 495447 224662
rect 495447 224516 499083 224662
rect 499083 224598 504023 224662
rect 504023 224598 508299 224662
rect 508299 224598 510167 224662
rect 499083 224596 510167 224598
rect 510167 224596 513739 224662
rect 513739 224596 515479 224662
rect 515479 224596 519115 224662
rect 519115 224598 523543 224662
rect 523543 224598 527819 224662
rect 527819 224598 529687 224726
rect 519115 224596 529687 224598
rect 529687 224596 533259 224726
rect 533259 224596 534999 224726
rect 534999 224596 538635 224726
rect 538635 224596 543503 224726
rect 499083 224516 503903 224596
rect 510087 224534 510167 224596
rect 510167 224534 513663 224596
rect 515447 224534 515479 224596
rect 515479 224534 519103 224596
rect 529527 224534 529687 224596
rect 529687 224534 533183 224596
rect 534887 224534 534999 224596
rect 534999 224534 538543 224596
rect 510087 224516 513663 224534
rect 515447 224516 519103 224534
rect 529527 224516 533183 224534
rect 534887 224516 538543 224534
rect 490007 224470 490135 224516
rect 490135 224470 493663 224516
rect 490007 224436 493663 224470
rect 12428 210246 16564 210248
rect 559509 356701 562125 359157
rect 484661 208901 485837 208941
rect 484661 202385 484676 208901
rect 484676 208861 485837 208901
rect 487861 208861 491917 208941
rect 493221 208861 497277 208941
rect 504501 208901 505677 208941
rect 504501 208861 504516 208901
rect 504516 208861 505677 208901
rect 507701 208861 511757 208941
rect 513061 208861 517117 208941
rect 524021 208901 525197 208941
rect 524021 208861 524036 208901
rect 484676 208837 485880 208861
rect 485880 208837 498692 208861
rect 498692 208837 502520 208861
rect 502520 208837 504516 208861
rect 504516 208837 505720 208861
rect 505720 208837 518468 208861
rect 518468 208837 522360 208861
rect 522360 208837 524036 208861
rect 524036 208837 525176 208901
rect 525176 208861 525197 208901
rect 527221 208861 531277 208941
rect 532581 208861 536637 208941
rect 525176 208837 537988 208861
rect 537988 208837 541880 208861
rect 541880 208837 544077 208861
rect 484676 207697 544056 208837
rect 544056 207697 544077 208837
rect 484676 207685 485880 207697
rect 485880 207685 487812 207697
rect 487812 207685 489016 207697
rect 489016 207685 490884 207697
rect 490884 207685 492088 207697
rect 492088 207685 493252 207697
rect 493252 207685 497336 207697
rect 497336 207685 498692 207697
rect 498692 207685 499832 207697
rect 499832 207685 501380 207697
rect 501380 207685 502520 207697
rect 502520 207685 504516 207697
rect 504516 207685 505720 207697
rect 505720 207685 507652 207697
rect 507652 207685 508856 207697
rect 508856 207685 510724 207697
rect 510724 207685 511864 207697
rect 511864 207685 513092 207697
rect 513092 207685 517176 207697
rect 517176 207685 518468 207697
rect 518468 207685 519672 207697
rect 519672 207685 521156 207697
rect 521156 207685 522360 207697
rect 522360 207685 524036 207697
rect 524036 207685 525240 207697
rect 525240 207685 527172 207697
rect 527172 207685 528312 207697
rect 528312 207685 530244 207697
rect 530244 207685 531384 207697
rect 531384 207685 532612 207697
rect 532612 207685 536696 207697
rect 536696 207685 537988 207697
rect 537988 207685 539192 207697
rect 539192 207685 540676 207697
rect 540676 207685 541880 207697
rect 541880 207685 544077 207697
rect 484676 203421 485837 207685
rect 487861 203525 489016 207685
rect 489016 203525 489037 207685
rect 490741 203525 490884 207685
rect 490884 203525 491917 207685
rect 493221 203525 493252 207685
rect 493252 203525 494397 207685
rect 496101 207633 497277 207685
rect 496101 203525 496196 207633
rect 496196 203525 497277 207633
rect 498661 203525 498692 207685
rect 498692 203525 499757 207685
rect 501301 203525 501380 207685
rect 501380 203525 502477 207685
rect 504501 203525 504516 207685
rect 504516 203525 505677 207685
rect 507701 203525 508856 207685
rect 508856 203525 508877 207685
rect 510581 203525 510724 207685
rect 510724 203525 511757 207685
rect 513061 203525 513092 207685
rect 513092 203525 514237 207685
rect 515941 207633 517117 207685
rect 515941 203525 516036 207633
rect 516036 203525 517117 207633
rect 518421 203525 518468 207685
rect 518468 203525 519597 207685
rect 521141 203525 521156 207685
rect 521156 203525 522237 207685
rect 524021 203525 524036 207685
rect 524036 203525 525197 207685
rect 527221 203525 528312 207685
rect 528312 203525 528317 207685
rect 530101 203525 530244 207685
rect 530244 203525 531277 207685
rect 532581 203525 532612 207685
rect 532612 207633 533757 207685
rect 535461 207633 536637 207685
rect 532612 203525 533752 207633
rect 533752 203525 533757 207633
rect 535461 203525 535492 207633
rect 535492 203525 536637 207633
rect 537941 203525 537988 207685
rect 537988 203525 539117 207685
rect 540661 203525 540676 207685
rect 540676 203525 541757 207685
rect 567174 313226 569870 316082
rect 487861 203421 489037 203525
rect 490741 203421 491917 203525
rect 493221 203421 494397 203525
rect 496101 203421 497277 203525
rect 498661 203421 499757 203525
rect 501301 203421 502477 203525
rect 504501 203421 505677 203525
rect 507701 203421 508877 203525
rect 510581 203421 511757 203525
rect 513061 203421 514237 203525
rect 515941 203421 517117 203525
rect 518421 203421 519597 203525
rect 521141 203421 522237 203525
rect 524021 203421 525197 203525
rect 527221 203421 528317 203525
rect 530101 203421 531277 203525
rect 532581 203421 533757 203525
rect 535461 203421 536637 203525
rect 537941 203421 539117 203525
rect 540661 203421 541757 203525
rect 484676 202385 543992 203421
rect 543992 202385 543997 203421
rect 484661 202257 484740 202385
rect 484740 202257 489016 202385
rect 489016 202257 490884 202385
rect 484661 202245 490884 202257
rect 490884 202245 494456 202385
rect 494456 202245 496196 202385
rect 496196 202245 499832 202385
rect 499832 202257 504580 202385
rect 504580 202257 508856 202385
rect 508856 202257 510724 202385
rect 499832 202245 510724 202257
rect 510724 202245 514296 202385
rect 514296 202245 516036 202385
rect 516036 202245 519672 202385
rect 519672 202257 524100 202385
rect 524100 202257 528312 202385
rect 528312 202257 530244 202385
rect 519672 202245 530244 202257
rect 490741 202193 490884 202245
rect 490884 202193 494397 202245
rect 496101 202193 496196 202245
rect 496196 202193 499757 202245
rect 510581 202193 510724 202245
rect 510724 202193 514237 202245
rect 515941 202193 516036 202245
rect 516036 202193 519597 202245
rect 530101 202193 530244 202245
rect 530244 202193 533752 202385
rect 533752 202245 535492 202385
rect 535492 202245 539192 202385
rect 539192 202245 543997 202385
rect 533752 202193 533757 202245
rect 490741 202165 494397 202193
rect 496101 202165 499757 202193
rect 510581 202165 514237 202193
rect 515941 202165 519597 202193
rect 530101 202165 533757 202193
rect 535461 202193 535492 202245
rect 535492 202193 539117 202245
rect 535461 202165 539117 202193
rect 64965 167087 66141 167097
rect 64965 165691 66141 167087
rect 64965 165681 66141 165691
rect 84618 164673 84674 164729
rect 84698 164673 84754 164729
rect 84778 164673 84834 164729
rect 84858 164673 84914 164729
rect 84938 164673 84994 164729
rect 85018 164673 85074 164729
rect 85098 164673 85154 164729
rect 85178 164673 85234 164729
rect 85259 164672 85315 164728
rect 85351 164673 85407 164729
rect 79742 164215 79798 164271
rect 79742 164135 79798 164191
rect 79742 164055 79798 164111
rect 79742 163975 79798 164031
rect 79742 163895 79798 163951
rect 65105 163893 66281 163895
rect 65105 162881 66281 163893
rect 79742 163815 79798 163871
rect 79742 163735 79798 163791
rect 79742 163655 79798 163711
rect 79742 163575 79798 163631
rect 79742 163495 79798 163551
rect 65105 162879 66281 162881
rect 65253 158231 66189 159167
rect 573278 268416 576374 270712
rect 9845 37569 11021 38985
rect 107302 64678 109038 64680
rect 107302 63026 109038 64678
rect 107302 63024 109038 63026
rect 106293 57654 106909 58190
rect 7605 16446 8621 17702
rect 475421 147292 475477 147348
rect 475521 147292 475577 147348
rect 475621 147292 475677 147348
rect 475721 147292 475777 147348
rect 475821 147292 475877 147348
rect 475921 147292 475977 147348
rect 476021 147292 476077 147348
rect 476121 147292 476177 147348
rect 465021 144867 465237 145083
rect 465056 143432 465192 143568
rect 464971 142790 465267 143086
rect 475326 142755 475382 142758
rect 475326 142703 475328 142755
rect 475328 142703 475380 142755
rect 475380 142703 475382 142755
rect 475326 142702 475382 142703
rect 475407 142756 475463 142758
rect 475407 142704 475409 142756
rect 475409 142704 475461 142756
rect 475461 142704 475463 142756
rect 475407 142702 475463 142704
rect 475488 142756 475544 142758
rect 475488 142704 475490 142756
rect 475490 142704 475542 142756
rect 475542 142704 475544 142756
rect 475488 142702 475544 142704
rect 475569 142756 475625 142758
rect 475569 142704 475571 142756
rect 475571 142704 475623 142756
rect 475623 142704 475625 142756
rect 475569 142702 475625 142704
rect 475650 142755 475706 142758
rect 475650 142703 475652 142755
rect 475652 142703 475704 142755
rect 475704 142703 475706 142755
rect 475650 142702 475706 142703
rect 475326 142674 475382 142676
rect 475326 142622 475328 142674
rect 475328 142622 475380 142674
rect 475380 142622 475382 142674
rect 475326 142620 475382 142622
rect 475407 142675 475463 142676
rect 475407 142623 475409 142675
rect 475409 142623 475461 142675
rect 475461 142623 475463 142675
rect 475407 142620 475463 142623
rect 475488 142673 475544 142676
rect 475488 142621 475491 142673
rect 475491 142621 475543 142673
rect 475543 142621 475544 142673
rect 475488 142620 475544 142621
rect 475569 142674 475625 142676
rect 475569 142622 475571 142674
rect 475571 142622 475623 142674
rect 475623 142622 475625 142674
rect 475569 142620 475625 142622
rect 475650 142674 475706 142676
rect 475650 142622 475652 142674
rect 475652 142622 475704 142674
rect 475704 142622 475706 142674
rect 475650 142620 475706 142622
rect 464802 139376 466058 140632
rect 575897 140630 575923 142206
rect 575923 140630 577447 142206
rect 577447 140630 577473 142206
rect 567131 93799 567587 94255
rect 563422 48766 564118 49782
rect 460306 12226 461322 12922
rect 459108 8037 460364 9293
rect 458125 3792 459461 5288
<< metal3 >>
rect 16180 704800 21180 704810
rect 16180 702300 21194 704800
rect 16180 700290 21180 702300
rect 16160 696000 21180 700290
rect 44016 696000 48736 696008
rect 16150 690710 48736 696000
rect -800 685240 1700 685242
rect 18300 685240 36384 685250
rect -800 680260 36384 685240
rect -800 680250 18340 680260
rect -800 680242 1700 680250
rect -800 648619 1660 648642
rect -800 643842 16232 648619
rect -774 643805 16232 643842
rect -800 638635 1660 638642
rect 11444 638635 16232 643805
rect -800 633842 16232 638635
rect 11444 631627 16232 633842
rect 11444 631062 16257 631627
rect 11444 627566 11948 631062
rect 15684 627566 16257 631062
rect 11444 627037 16257 627566
rect 11447 627028 16257 627037
rect 31384 596448 36384 680260
rect 44016 606504 48736 690710
rect 68194 626978 73194 704800
rect 67484 626039 73886 626978
rect 67484 621023 68344 626039
rect 72960 621023 73886 626039
rect 67484 620234 73886 621023
rect 120194 616048 125194 704802
rect 566594 704800 571592 704801
rect 165594 702300 170598 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 703568 418394 704800
rect 413378 702300 418394 703568
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 175579 693838 324135 694407
rect 165594 691832 170594 692506
rect 165594 689288 166450 691832
rect 169714 689288 170594 691832
rect 175579 690814 320613 693838
rect 323557 690814 324135 693838
rect 175579 690389 324135 690814
rect 413378 692696 418390 702300
rect 175579 689880 179597 690389
rect 165594 684762 170594 689288
rect 118068 614830 125194 616048
rect 118068 610214 119475 614830
rect 123611 614492 125194 614830
rect 123611 610214 125192 614492
rect 118068 608944 125192 610214
rect 165596 606504 170594 684762
rect 44016 605004 120650 606504
rect 31380 596440 37860 596448
rect 67936 596440 72370 596444
rect 99600 596440 101510 596560
rect 31380 596248 101510 596440
rect 31380 595232 99947 596248
rect 101203 595232 101510 596248
rect 31380 594940 101510 595232
rect 31380 594936 41688 594940
rect 67936 594938 72370 594940
rect 99600 594870 101510 594940
rect 120042 594462 120650 605004
rect 33184 593711 36516 594128
rect 33184 591815 33649 593711
rect 36025 591815 36516 593711
rect 120040 592422 120650 594462
rect 121340 605006 170594 606504
rect 121340 605004 170592 605006
rect 121340 594744 121948 605004
rect 175576 603968 179600 689880
rect 413378 689500 418410 692696
rect 413398 681000 418410 689500
rect 200278 680996 418410 681000
rect 200076 678628 418410 680996
rect 200076 678502 418406 678628
rect 135464 602370 179600 603968
rect 200088 678500 418406 678502
rect 135464 597176 136816 602370
rect 200088 596078 201080 678500
rect 466186 677048 468686 702300
rect 566594 690911 571592 702300
rect 566589 690166 571598 690911
rect 566589 686270 567317 690166
rect 570973 686270 571598 690166
rect 566589 685375 571598 686270
rect 566501 682580 584800 682984
rect 566501 678444 567033 682580
rect 571009 678444 584800 682580
rect 566501 677984 584800 678444
rect 207091 674548 468686 677048
rect 199804 595464 201598 596078
rect 199624 595077 201786 595464
rect 193894 594774 194254 594828
rect 193894 594770 194002 594774
rect 194146 594770 194254 594774
rect 121340 594238 122734 594744
rect 193894 594394 193966 594770
rect 194182 594394 194254 594770
rect 193894 594390 194002 594394
rect 194146 594390 194254 594394
rect 193894 594330 194254 594390
rect 199624 594381 199948 595077
rect 201284 594381 201786 595077
rect 199624 593982 201786 594381
rect 131634 593734 131983 593788
rect 131634 593670 131735 593734
rect 131799 593670 131817 593734
rect 131881 593670 131983 593734
rect 131634 593623 131983 593670
rect 120040 592349 122714 592422
rect 120040 591973 122322 592349
rect 122618 591973 122714 592349
rect 120040 591902 122714 591973
rect 33184 591326 36516 591815
rect 11441 574778 20742 576490
rect 11432 574314 20742 574778
rect 11432 571058 11957 574314
rect 15613 571674 20742 574314
rect 15613 571058 16257 571674
rect 11432 570604 16257 571058
rect -800 564219 1660 564242
rect 11441 564219 16257 570604
rect -800 561763 16257 564219
rect -800 559442 16229 561763
rect -777 559405 16229 559442
rect -800 554235 1660 554242
rect 11441 554235 16229 559405
rect -803 551902 16229 554235
rect -803 549442 16246 551902
rect -803 549439 1663 549442
rect 33184 512822 36510 591326
rect 89790 581513 90096 581598
rect 89790 581289 89865 581513
rect 90009 581289 90096 581513
rect 121470 581529 121900 581596
rect 121470 581385 121526 581529
rect 121830 581385 121900 581529
rect 121470 581312 121900 581385
rect 89790 580396 90096 581289
rect 120316 581172 120744 581228
rect 45420 572555 47606 573056
rect 45420 571379 46120 572555
rect 47056 571379 47606 572555
rect 7142 511648 36510 512822
rect -800 511530 36510 511648
rect 7142 510896 36510 511530
rect 37928 551214 42430 551854
rect 37928 548430 38602 551214
rect 41546 548430 42430 551214
rect 37928 547750 42430 548430
rect 7142 510894 36502 510896
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 37928 472350 41254 547750
rect 36296 471852 41254 472350
rect 36296 469252 36953 471852
rect 6872 468420 36953 469252
rect -800 468308 36953 468420
rect 6872 467788 36953 468308
rect 40457 467788 41254 471852
rect 6872 467330 41254 467788
rect 6872 467324 41250 467330
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 45420 427328 47606 571379
rect 50730 571080 52020 571350
rect 50730 569824 50950 571080
rect 51726 569824 52020 571080
rect 50730 569576 52020 569824
rect 50724 569574 52020 569576
rect 50724 568512 52018 569574
rect 55500 569523 57212 569946
rect 89864 569926 90096 580396
rect 90482 581059 90714 581164
rect 90482 580995 90559 581059
rect 90623 580995 90714 581059
rect 90482 580979 90714 580995
rect 90482 580915 90559 580979
rect 90623 580915 90714 580979
rect 120316 581028 120422 581172
rect 120646 581028 120744 581172
rect 120316 580976 120744 581028
rect 90482 571342 90714 580915
rect 90974 580853 91212 580942
rect 90974 580789 91057 580853
rect 91121 580789 91212 580853
rect 90974 580773 91212 580789
rect 90974 580709 91057 580773
rect 91121 580709 91212 580773
rect 90974 572170 91212 580709
rect 207091 574172 209591 674548
rect 555848 644910 570748 646373
rect 555848 644571 570752 644910
rect 555848 644372 584800 644571
rect 555848 630156 558084 644372
rect 568220 639771 584800 644372
rect 568220 634584 570748 639771
rect 568220 630156 584800 634584
rect 555848 629784 584800 630156
rect 555848 628156 570748 629784
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 513520 583562 584800 583674
rect 513520 583422 577057 583562
rect 513520 582339 514045 583422
rect 513519 582166 514045 582339
rect 515381 582339 577057 583422
rect 515381 582166 515917 582339
rect 513519 581790 515917 582166
rect 90894 572089 91286 572170
rect 90894 571873 90983 572089
rect 91199 571873 91286 572089
rect 90894 571792 91286 571873
rect 114121 571672 209591 574172
rect 90420 571251 90776 571342
rect 90420 571035 90491 571251
rect 90707 571035 90776 571251
rect 90420 570954 90776 571035
rect 89806 569835 90162 569926
rect 89806 569619 89871 569835
rect 90087 569619 90162 569835
rect 89806 569538 90162 569619
rect 89864 569536 90096 569538
rect 43996 426927 47606 427328
rect 43996 426575 44638 426927
rect 6945 425198 44638 426575
rect -800 425086 44638 425198
rect 6945 424783 44638 425086
rect 47182 424783 47606 426927
rect 6945 424389 47606 424783
rect 43996 424388 47596 424389
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 50737 382224 52012 568512
rect 55500 568267 55842 569523
rect 56858 568267 57212 569523
rect 55500 566624 57212 568267
rect 5769 381976 52012 382224
rect -800 381864 52012 381976
rect 5769 380949 52012 381864
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 55571 340882 57201 566624
rect 114121 563122 116621 571672
rect 70303 560622 116621 563122
rect 70303 477270 72803 560622
rect 544585 555691 548067 555820
rect 542391 555469 548067 555691
rect 542295 555453 572140 555469
rect 542295 555345 572198 555453
rect 542295 554928 584800 555345
rect 542295 550669 543521 554928
rect 542391 541592 543521 550669
rect 546937 550669 584800 554928
rect 546937 545310 548067 550669
rect 554955 550545 584800 550669
rect 554955 545310 584800 545345
rect 546937 541592 584800 545310
rect 542391 540891 584800 541592
rect 542581 540545 584800 540891
rect 542581 540510 572426 540545
rect 186660 525028 191891 525562
rect 186660 523204 187358 525028
rect 191262 523204 191891 525028
rect 70303 475606 70706 477270
rect 72450 475606 72803 477270
rect 70303 475273 72803 475606
rect 186660 467969 191891 523204
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 518800 494973 521214 494977
rect 518800 494718 581097 494973
rect 518800 493302 519175 494718
rect 520831 494252 581097 494718
rect 520831 494140 584800 494252
rect 520831 493638 581097 494140
rect 520831 493302 521214 493638
rect 518800 492906 521214 493302
rect 82646 462738 191891 467969
rect 55571 340729 57204 340882
rect 55578 339542 57204 340729
rect 5790 338754 57204 339542
rect -800 338642 57204 338754
rect 5790 337912 57204 338642
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 2846 296492 8410 296865
rect 2844 296165 8410 296492
rect 2844 295532 3588 296165
rect -800 295420 3588 295532
rect -800 294238 480 294350
rect 2844 294078 3588 295420
rect -800 293056 480 293168
rect 2846 292101 3588 294078
rect 7732 292101 8410 296165
rect -800 291874 480 291986
rect 2846 291336 8410 292101
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 82646 254926 87877 462738
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 524071 450373 582463 450426
rect 524067 450040 582463 450373
rect 524067 448464 524359 450040
rect 526095 449830 582463 450040
rect 526095 449718 584800 449830
rect 526095 449085 582463 449718
rect 526095 448464 526461 449085
rect 524067 448044 526461 448464
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 553614 405600 580571 405945
rect 553614 403144 554301 405600
rect 556437 405408 580571 405600
rect 556437 405296 584800 405408
rect 556437 404815 580571 405296
rect 556437 403144 556971 404815
rect 553614 402563 556971 403144
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 562253 359447 582205 359472
rect 559120 359157 582205 359447
rect 559120 356701 559509 359157
rect 562125 358986 582205 359157
rect 562125 358874 584800 358986
rect 562125 358289 582205 358874
rect 562125 356701 562476 358289
rect 559120 356321 562476 356701
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 566803 316082 570308 316420
rect 566803 313226 567174 316082
rect 569870 314216 570308 316082
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 569870 313764 582518 314216
rect 569870 313652 584800 313764
rect 569870 313226 582518 313652
rect 566803 313212 582518 313226
rect 566803 312868 570308 313212
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 572605 270712 577066 271263
rect 572605 268416 573278 270712
rect 576374 270050 577066 270712
rect 583520 270412 584800 270524
rect 576374 269342 582479 270050
rect 576374 269230 584800 269342
rect 576374 268668 582479 269230
rect 576374 268416 577066 268668
rect 572605 267828 577066 268416
rect 6294 252510 87877 254926
rect -800 252398 87877 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect 6294 249695 87877 252398
rect 6294 249694 11528 249695
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect -800 214888 7711 219688
rect 2911 214679 7711 214888
rect 11848 214679 17002 215261
rect 2906 214142 17002 214679
rect 2906 210246 12428 214142
rect 16564 210246 17002 214142
rect 2906 209879 17002 210246
rect -800 209679 1660 209688
rect 2906 209679 7711 209879
rect -800 204888 7711 209679
rect -695 204879 7711 204888
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 28604 167390 31522 249695
rect 574844 235230 584800 240030
rect 542475 233292 548167 233663
rect 509823 231467 514086 231495
rect 529318 231494 533581 231522
rect 542475 231494 542887 233292
rect 547663 233289 548167 233292
rect 523229 231467 542887 231494
rect 489768 231435 494031 231463
rect 503734 231435 542887 231467
rect 483679 231292 542887 231435
rect 483679 231212 523447 231292
rect 524623 231289 526647 231292
rect 530703 231289 532007 231292
rect 536063 231289 542887 231292
rect 483679 231209 483927 231212
rect 485103 231209 487127 231212
rect 491183 231209 492487 231212
rect 496543 231209 497847 231212
rect 501663 231209 504007 231212
rect 483679 224505 483870 231209
rect 547694 230105 548167 233289
rect 485103 229640 487070 229956
rect 485103 226052 485474 229640
rect 486784 226052 487070 229640
rect 485103 225692 487070 226052
rect 488254 229640 490007 229956
rect 488254 226052 488579 229640
rect 489768 226052 490007 229640
rect 488254 225692 490007 226052
rect 491294 229640 492487 229956
rect 491294 226052 491563 229640
rect 492236 226052 492487 229640
rect 491294 225692 492487 226052
rect 493663 229640 495367 229956
rect 493663 226052 494031 229640
rect 495099 226052 495367 229640
rect 493663 225692 495367 226052
rect 496654 229640 497847 229956
rect 496654 226052 496894 229640
rect 497621 226052 497847 229640
rect 496654 225692 497847 226052
rect 499134 229640 500567 229956
rect 499134 226052 499416 229640
rect 500213 226052 500567 229640
rect 499134 225692 500567 226052
rect 501854 229640 503950 229956
rect 501854 226052 502008 229640
rect 503734 226052 503950 229640
rect 501854 225852 503950 226052
rect 501854 225692 503927 225852
rect 505183 229672 507127 230036
rect 505183 226084 505529 229672
rect 506839 226084 507127 229672
rect 505183 225772 507127 226084
rect 508303 229672 510087 230036
rect 508303 226084 508634 229672
rect 509823 226084 510087 229672
rect 508303 225772 510087 226084
rect 511294 229672 512510 230036
rect 511294 226084 511618 229672
rect 512291 226084 512510 229672
rect 511294 225772 512510 226084
rect 513694 229672 515447 230025
rect 513694 226084 514086 229672
rect 515154 226084 515447 229672
rect 513694 225772 515447 226084
rect 516734 229672 517927 230036
rect 516734 226084 516949 229672
rect 517676 226084 517927 229672
rect 516734 225772 517927 226084
rect 519134 229672 520567 230036
rect 519134 226084 519471 229672
rect 520268 226084 520567 229672
rect 519134 225772 520567 226084
rect 521934 229672 523447 230036
rect 521934 226084 522063 229672
rect 523229 226084 523447 229672
rect 521934 225772 523447 226084
rect 543503 230036 548167 230105
rect 524623 229699 526590 230036
rect 524623 226111 525024 229699
rect 526334 226111 526590 229699
rect 524623 225772 526590 226111
rect 527823 229699 529527 230036
rect 527823 226111 528129 229699
rect 529318 226111 529527 229699
rect 527823 225772 529527 226111
rect 530814 229699 532007 230036
rect 530814 226111 531113 229699
rect 531786 226111 532007 229699
rect 530814 225772 532007 226111
rect 533214 229699 534887 230036
rect 533214 226111 533581 229699
rect 534649 226111 534887 229699
rect 533214 225772 534887 226111
rect 536174 229699 537447 230036
rect 536174 226111 536444 229699
rect 537171 226111 537447 229699
rect 536174 225772 537447 226111
rect 538654 229699 540087 230036
rect 538654 226111 538966 229699
rect 539763 226111 540087 229699
rect 538654 225772 540087 226111
rect 541454 229699 548167 230036
rect 574844 230030 579544 235230
rect 541454 226111 541558 229699
rect 542475 229677 548167 229699
rect 551348 226126 584800 230030
rect 543501 226111 584800 226126
rect 541454 225772 584800 226111
rect 543503 225689 584800 225772
rect 543534 225275 584800 225689
rect 543534 224505 555659 225275
rect 582340 225230 584800 225275
rect 483679 224436 490007 224505
rect 493663 224436 495470 224505
rect 483679 224425 490110 224436
rect 493614 224425 495470 224436
rect 499134 224425 500670 224505
rect 501854 224425 555659 224505
rect 483679 224316 555659 224425
rect 483679 224289 524286 224316
rect 543501 224304 555659 224316
rect 483679 224257 504231 224289
rect 433033 218341 437788 218348
rect 433033 217437 449718 218341
rect 433033 217261 449725 217437
rect 433033 216725 447324 217261
rect 449460 216725 449725 217261
rect 433033 216662 449725 216725
rect 433033 173573 437788 216662
rect 446975 216630 449725 216662
rect 490528 209155 494791 209183
rect 510353 209155 514616 209183
rect 529864 209155 534127 209183
rect 484439 208941 544367 209155
rect 484439 208938 484661 208941
rect 485837 208938 487861 208941
rect 491917 208938 493221 208941
rect 497277 208938 504501 208941
rect 505677 208938 507701 208941
rect 511757 208938 513061 208941
rect 517117 208938 524021 208941
rect 525197 208938 527221 208941
rect 531277 208938 532581 208941
rect 536637 208938 544367 208941
rect 484439 202234 484625 208938
rect 544129 207754 544367 208938
rect 485837 207360 487825 207685
rect 485837 203772 486234 207360
rect 487544 203772 487825 207360
rect 485837 203421 487825 203772
rect 489037 207360 490741 207685
rect 489037 203772 489339 207360
rect 490528 203772 490741 207360
rect 489037 203421 490741 203772
rect 492049 207360 493221 207685
rect 492049 203772 492323 207360
rect 492996 203772 493221 207360
rect 492049 203421 493221 203772
rect 494397 207360 496101 207685
rect 494397 203772 494791 207360
rect 495859 203772 496101 207360
rect 494397 203421 496101 203772
rect 497409 207360 498661 207685
rect 497409 203772 497654 207360
rect 498381 203772 498661 207360
rect 497409 203421 498661 203772
rect 499889 207360 501301 207685
rect 499889 203772 500176 207360
rect 500973 203772 501301 207360
rect 499889 203421 501301 203772
rect 502609 207360 504465 207685
rect 502609 203772 502768 207360
rect 504264 203772 504465 207360
rect 502609 203421 504465 203772
rect 505677 207360 507665 207685
rect 505677 203772 506059 207360
rect 507369 203772 507665 207360
rect 505677 203421 507665 203772
rect 508877 207360 510581 207685
rect 508877 203772 509164 207360
rect 510353 203772 510581 207360
rect 508877 203421 510581 203772
rect 511809 207360 513061 207685
rect 511809 203772 512148 207360
rect 512821 203772 513061 207360
rect 511809 203421 513061 203772
rect 544077 207685 544367 207754
rect 514237 207360 515941 207685
rect 514237 203772 514616 207360
rect 515684 203772 515941 207360
rect 514237 203421 515941 203772
rect 517249 207360 518421 207685
rect 517249 203772 517479 207360
rect 518206 203772 518421 207360
rect 517249 203421 518421 203772
rect 519729 207360 521141 207685
rect 519729 203772 520001 207360
rect 520798 203772 521141 207360
rect 519729 203421 521141 203772
rect 522449 207360 523985 207685
rect 522449 203772 522593 207360
rect 523775 203772 523985 207360
rect 522449 203421 523985 203772
rect 525197 207360 527185 207685
rect 525197 203772 525570 207360
rect 526880 203772 527185 207360
rect 525197 203421 527185 203772
rect 528317 207360 530101 207685
rect 528317 203772 528675 207360
rect 529864 203772 530101 207360
rect 528317 203421 530101 203772
rect 531329 207360 532545 207685
rect 531329 203772 531659 207360
rect 532332 203772 532545 207360
rect 531329 203421 532545 203772
rect 533757 207360 535461 207685
rect 533757 203772 534127 207360
rect 535195 203772 535461 207360
rect 533757 203421 535461 203772
rect 536769 207360 537941 207685
rect 536769 203772 536990 207360
rect 537717 203772 537941 207360
rect 536769 203421 537941 203772
rect 539169 207360 540661 207685
rect 539169 203772 539512 207360
rect 540309 203772 540661 207360
rect 539169 203421 540661 203772
rect 541969 207360 544367 207685
rect 541969 203772 542104 207360
rect 541969 203421 544327 203772
rect 543997 203338 544327 203421
rect 544129 202234 544327 203338
rect 484439 202165 490741 202234
rect 494397 202165 496101 202234
rect 484439 202154 490865 202165
rect 494369 202154 496225 202165
rect 499889 202154 501505 202234
rect 502609 202165 510581 202234
rect 514237 202165 515941 202234
rect 502609 202154 510705 202165
rect 514209 202154 516065 202165
rect 519729 202154 521265 202234
rect 522449 202165 530101 202234
rect 533757 202165 535461 202234
rect 522449 202154 530225 202165
rect 533729 202154 535585 202165
rect 539169 202154 540785 202234
rect 541969 202154 544327 202234
rect 484439 201977 544327 202154
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 433033 173532 579709 173573
rect 433033 168774 580438 173532
rect 436258 168770 580438 168774
rect 28604 167097 66512 167390
rect 28604 165681 64965 167097
rect 66141 165681 66512 167097
rect 28604 165324 66512 165681
rect 28438 163895 66510 164066
rect 28438 162879 65105 163895
rect 66281 163548 66510 163895
rect 66281 162879 66506 163548
rect 28438 162680 66506 162879
rect 28438 162679 65133 162680
rect 28438 125256 31208 162679
rect 65048 159344 66406 159346
rect 5044 124888 31208 125256
rect -800 124776 31208 124888
rect 5044 124386 31208 124776
rect 41080 159167 66406 159344
rect 41080 158231 65253 159167
rect 66189 158231 66406 159167
rect 41080 158030 66406 158231
rect 41080 158027 65977 158030
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 41080 82054 43850 158027
rect 575676 151624 580438 168770
rect 582340 151624 584800 151630
rect 475058 147352 476380 147408
rect 475058 147288 475417 147352
rect 475481 147288 475517 147352
rect 475581 147288 475617 147352
rect 475681 147288 475717 147352
rect 475781 147288 475817 147352
rect 475881 147288 475917 147352
rect 475981 147288 476017 147352
rect 476081 147288 476117 147352
rect 476181 147288 476380 147352
rect 475058 147249 476380 147288
rect 575676 146862 584800 151624
rect 464944 145087 465322 145138
rect 464944 144863 465017 145087
rect 465241 144863 465322 145087
rect 464944 144822 465322 144863
rect 465010 143572 465248 143600
rect 465010 143428 465052 143572
rect 465196 143428 465248 143572
rect 465010 143402 465248 143428
rect 464766 143148 464934 143150
rect 464766 143086 465390 143148
rect 460984 143031 462372 143032
rect 464766 143031 464971 143086
rect 460984 143012 464971 143031
rect 4062 81666 43850 82054
rect -800 81554 43850 81666
rect 4062 81184 43850 81554
rect 460982 142857 464971 143012
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 106942 64684 109354 64999
rect 106942 63020 107298 64684
rect 109042 63020 109354 64684
rect 106942 62650 109354 63020
rect 106116 58190 107054 58322
rect 106116 57654 106293 58190
rect 106909 57654 107054 58190
rect 106116 57508 107054 57654
rect 9404 38985 11556 39232
rect 9404 38444 9845 38985
rect -800 38332 9845 38444
rect 9404 37569 9845 38332
rect 11021 37569 11556 38985
rect -800 37150 480 37262
rect 9404 37220 11556 37569
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect 106282 33569 106920 57508
rect 25257 32931 106920 33569
rect -800 32422 480 32534
rect 20849 20502 21484 20578
rect 20700 20434 21792 20502
rect 20700 20050 20977 20434
rect 21361 20050 21792 20434
rect 7312 17702 9026 18078
rect 7312 17022 7605 17702
rect -800 16910 7605 17022
rect 7312 16446 7605 16910
rect 8621 16446 9026 17702
rect 7312 16150 9026 16446
rect -800 15728 480 15840
rect -800 14546 480 14658
rect -800 13364 480 13476
rect -800 12182 480 12294
rect -800 11000 480 11112
rect -800 9818 480 9930
rect -800 8636 480 8748
rect 7534 8032 8626 8034
rect 20700 8032 21792 20050
rect 7534 7566 21792 8032
rect -800 7454 21792 7566
rect 7534 6940 21792 7454
rect 7534 6930 8626 6940
rect -800 6272 480 6384
rect -800 5090 480 5202
rect 25257 4748 25895 32931
rect 460982 17864 463239 142857
rect 464766 142790 464971 142857
rect 465267 142790 465390 143086
rect 464766 142712 465390 142790
rect 475246 142762 475823 142901
rect 475246 142698 475322 142762
rect 475386 142698 475403 142762
rect 475467 142698 475484 142762
rect 475548 142698 475565 142762
rect 475629 142698 475646 142762
rect 475710 142698 475823 142762
rect 475246 142680 475823 142698
rect 475246 142616 475322 142680
rect 475386 142616 475403 142680
rect 475467 142616 475484 142680
rect 475548 142616 475565 142680
rect 475629 142616 475646 142680
rect 475710 142616 475823 142680
rect 475246 142531 475823 142616
rect 575676 142436 578136 146862
rect 582340 146830 584800 146862
rect 575630 142206 578136 142436
rect 464550 140632 466306 140864
rect 464550 139376 464802 140632
rect 466058 139376 466306 140632
rect 575630 140630 575897 142206
rect 577473 141630 578136 142206
rect 577473 140630 584800 141630
rect 575630 140357 584800 140630
rect 464550 22714 466306 139376
rect 575658 139170 584800 140357
rect 575676 136830 584800 139170
rect 575676 136816 584762 136830
rect 583520 95118 584800 95230
rect 567040 94255 567690 94358
rect 567040 93799 567131 94255
rect 567587 94048 567690 94255
rect 567587 93936 584800 94048
rect 567587 93799 567690 93936
rect 567040 93708 567690 93799
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 563194 49782 564398 50018
rect 563194 48766 563422 49782
rect 564118 49390 564398 49782
rect 564118 49278 584800 49390
rect 564118 48766 564398 49278
rect 563194 48556 564398 48766
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 464550 22712 575192 22714
rect 464550 21750 576948 22712
rect 464538 21638 584800 21750
rect 464550 20962 576948 21638
rect 464550 20958 575134 20962
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 573544 17864 577376 17890
rect 460982 17022 577376 17864
rect 460982 16910 584800 17022
rect 460982 16124 577376 16910
rect 460982 16108 573780 16124
rect 575814 16108 577312 16124
rect 460982 16100 463239 16108
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect 583520 13364 584800 13476
rect 459942 13252 461676 13258
rect 459942 12922 577597 13252
rect 459942 12226 460306 12922
rect 461322 12294 577597 12922
rect 461322 12226 584800 12294
rect 459942 12182 584800 12226
rect 459942 11886 577597 12182
rect 461598 11884 462866 11886
rect 583520 11000 584800 11112
rect 583520 9818 584800 9930
rect 458720 9293 577522 9716
rect 458720 8037 459108 9293
rect 460364 8748 577522 9293
rect 460364 8636 584800 8748
rect 460364 8037 577522 8636
rect 458720 7731 577522 8037
rect 458720 7710 460749 7731
rect 583520 7454 584800 7566
rect 25254 4623 25895 4748
rect 457696 5649 460059 6399
rect 583520 6272 584800 6384
rect 457696 5288 577290 5649
rect 25254 4272 25894 4623
rect 7030 4020 25894 4272
rect -800 3908 25894 4020
rect 7030 3634 25894 3908
rect 25254 3632 25894 3634
rect 457696 3792 458125 5288
rect 459461 4020 577290 5288
rect 583520 5090 584800 5202
rect 459461 3908 584800 4020
rect 459461 3792 577290 3908
rect 457696 3274 577290 3792
rect 459443 3265 577290 3274
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 166450 689288 169714 691832
rect 320613 690814 323557 693838
rect 194002 594770 194146 594774
rect 131125 594468 131189 594472
rect 131125 594412 131129 594468
rect 131129 594412 131185 594468
rect 131185 594412 131189 594468
rect 131125 594408 131189 594412
rect 131206 594468 131270 594472
rect 131206 594412 131210 594468
rect 131210 594412 131266 594468
rect 131266 594412 131270 594468
rect 131206 594408 131270 594412
rect 131288 594468 131352 594472
rect 131288 594412 131292 594468
rect 131292 594412 131348 594468
rect 131348 594412 131352 594468
rect 131288 594408 131352 594412
rect 131369 594468 131433 594472
rect 131369 594412 131373 594468
rect 131373 594412 131429 594468
rect 131429 594412 131433 594468
rect 131369 594408 131433 594412
rect 131450 594468 131514 594472
rect 131450 594412 131454 594468
rect 131454 594412 131510 594468
rect 131510 594412 131514 594468
rect 131450 594408 131514 594412
rect 194002 594394 194146 594770
rect 194002 594390 194146 594394
rect 131125 594386 131189 594390
rect 131125 594330 131129 594386
rect 131129 594330 131185 594386
rect 131185 594330 131189 594386
rect 131125 594326 131189 594330
rect 131206 594386 131270 594390
rect 131206 594330 131210 594386
rect 131210 594330 131266 594386
rect 131266 594330 131270 594386
rect 131206 594326 131270 594330
rect 131288 594386 131352 594390
rect 131288 594330 131292 594386
rect 131292 594330 131348 594386
rect 131348 594330 131352 594386
rect 131288 594326 131352 594330
rect 131369 594386 131433 594390
rect 131369 594330 131373 594386
rect 131373 594330 131429 594386
rect 131429 594330 131433 594386
rect 131369 594326 131433 594330
rect 131450 594386 131514 594390
rect 131450 594330 131454 594386
rect 131454 594330 131510 594386
rect 131510 594330 131514 594386
rect 131450 594326 131514 594330
rect 131735 593730 131799 593734
rect 131735 593674 131739 593730
rect 131739 593674 131795 593730
rect 131795 593674 131799 593730
rect 131735 593670 131799 593674
rect 131817 593730 131881 593734
rect 131817 593674 131821 593730
rect 131821 593674 131877 593730
rect 131877 593674 131881 593730
rect 131817 593670 131881 593674
rect 89865 581289 90009 581513
rect 121526 581525 121830 581529
rect 121526 581389 121530 581525
rect 121530 581389 121826 581525
rect 121826 581389 121830 581525
rect 121526 581385 121830 581389
rect 38602 548430 41546 551214
rect 36953 467788 40457 471852
rect 90559 580995 90623 581059
rect 90559 580915 90623 580979
rect 120422 581168 120646 581172
rect 120422 581032 120426 581168
rect 120426 581032 120642 581168
rect 120642 581032 120646 581168
rect 120422 581028 120646 581032
rect 91057 580789 91121 580853
rect 91057 580709 91121 580773
rect 44638 424783 47182 426927
rect 187358 523204 191262 525028
rect 117469 515779 117693 515923
rect 117716 515779 117860 515923
rect 125070 499501 125134 499565
rect 125179 499501 125243 499565
rect 125294 499501 125358 499565
rect 70706 475606 72450 477270
rect 3588 292101 7732 296165
rect 542910 231289 547663 233289
rect 523470 231212 524623 231289
rect 524623 231212 526647 231289
rect 526647 231212 530703 231289
rect 530703 231212 532007 231289
rect 532007 231212 536063 231289
rect 536063 231212 542887 231289
rect 542887 231212 547663 231289
rect 523470 231209 547663 231212
rect 483870 224516 483927 231209
rect 483927 231132 485103 231209
rect 485103 231132 487127 231209
rect 487127 231132 491183 231209
rect 491183 231132 492487 231209
rect 492487 231132 496543 231209
rect 496543 231132 497847 231209
rect 497847 231132 501663 231209
rect 501663 231132 504007 231209
rect 504007 231132 547663 231209
rect 483927 230116 547663 231132
rect 547663 230116 547694 233289
rect 483927 230105 543503 230116
rect 543503 230105 547694 230116
rect 483927 230025 505134 230105
rect 483927 225609 485054 230025
rect 487070 229956 488254 230025
rect 490110 229956 491294 230025
rect 487070 225692 487127 229956
rect 487127 225692 488223 229956
rect 488223 225692 488254 229956
rect 490110 225692 491183 229956
rect 491183 225692 491294 229956
rect 487070 225609 488254 225692
rect 490110 225609 491294 225692
rect 492510 225609 493614 230025
rect 495470 229956 496654 230025
rect 497950 229956 499134 230025
rect 500670 229956 501854 230025
rect 503950 229956 505134 230025
rect 495470 225692 496543 229956
rect 496543 225692 496654 229956
rect 497950 225692 499023 229956
rect 499023 225692 499134 229956
rect 500670 225692 501663 229956
rect 501663 225692 501854 229956
rect 503950 225852 504007 229956
rect 504007 225852 505134 229956
rect 495470 225609 496654 225692
rect 497950 225609 499134 225692
rect 500670 225609 501854 225692
rect 503950 225689 505134 225852
rect 507150 225689 508254 230105
rect 510190 230036 511294 230105
rect 512510 230036 516734 230105
rect 518030 230036 519134 230105
rect 520750 230036 521934 230105
rect 510190 225772 511183 230036
rect 511183 225772 511294 230036
rect 512510 225772 512567 230036
rect 512567 225772 513663 230036
rect 513663 230025 515447 230036
rect 515447 230025 516543 230036
rect 513663 225772 513694 230025
rect 515550 225772 516543 230025
rect 516543 225772 516734 230036
rect 518030 225772 519103 230036
rect 519103 225772 519134 230036
rect 520750 225772 521743 230036
rect 521743 225772 521934 230036
rect 510190 225689 511294 225772
rect 512510 225689 513694 225772
rect 515550 225689 516734 225772
rect 518030 225689 519134 225772
rect 520750 225689 521934 225772
rect 523470 225689 524574 230105
rect 526590 230036 527774 230105
rect 529630 230036 530814 230105
rect 532030 230036 533214 230105
rect 535070 230036 536174 230105
rect 537470 230036 538654 230105
rect 540270 230036 541454 230105
rect 526590 225772 526647 230036
rect 526647 225772 527774 230036
rect 529630 225772 530703 230036
rect 530703 225772 530814 230036
rect 532030 225772 533183 230036
rect 533183 225772 533214 230036
rect 535070 225772 536063 230036
rect 536063 225772 536174 230036
rect 537470 225772 538543 230036
rect 538543 225772 538654 230036
rect 540270 225772 541263 230036
rect 541263 225772 541454 230036
rect 526590 225689 527774 225772
rect 529630 225689 530814 225772
rect 532030 225689 533214 225772
rect 535070 225689 536174 225772
rect 537470 225689 538654 225772
rect 540270 225689 541454 225772
rect 503950 225609 543503 225689
rect 483927 224596 543503 225609
rect 543503 224596 543534 225689
rect 483927 224516 503903 224596
rect 503903 224516 510087 224596
rect 510087 224516 513663 224596
rect 513663 224516 515447 224596
rect 515447 224516 519103 224596
rect 519103 224516 529527 224596
rect 529527 224516 533183 224596
rect 533183 224516 534887 224596
rect 534887 224516 538543 224596
rect 538543 224516 543534 224596
rect 483870 224505 490007 224516
rect 490007 224505 493663 224516
rect 493663 224505 543534 224516
rect 490110 224436 493614 224505
rect 490110 224425 493614 224436
rect 495470 224425 499134 224505
rect 500670 224425 501854 224505
rect 484625 202245 484661 208938
rect 484661 208861 485837 208938
rect 485837 208861 487861 208938
rect 487861 208861 491917 208938
rect 491917 208861 493221 208938
rect 493221 208861 497277 208938
rect 497277 208861 504501 208938
rect 504501 208861 505677 208938
rect 505677 208861 507701 208938
rect 507701 208861 511757 208938
rect 511757 208861 513061 208938
rect 513061 208861 517117 208938
rect 517117 208861 524021 208938
rect 524021 208861 525197 208938
rect 525197 208861 527221 208938
rect 527221 208861 531277 208938
rect 531277 208861 532581 208938
rect 532581 208861 536637 208938
rect 536637 208861 544129 208938
rect 484661 207754 544077 208861
rect 544077 207754 544129 208861
rect 484661 203338 485809 207754
rect 487825 207685 489009 207754
rect 490865 207685 492049 207754
rect 487825 203421 487861 207685
rect 487861 203421 489009 207685
rect 490865 203421 491917 207685
rect 491917 203421 492049 207685
rect 487825 203338 489009 203421
rect 490865 203338 492049 203421
rect 493265 203338 494369 207754
rect 496225 207685 497409 207754
rect 498705 207685 499889 207754
rect 501505 207685 502609 207754
rect 504465 207685 505649 207754
rect 507665 207685 508769 207754
rect 510705 207685 511809 207754
rect 496225 203421 497277 207685
rect 497277 203421 497409 207685
rect 498705 203421 499757 207685
rect 499757 203421 499889 207685
rect 501505 203421 502477 207685
rect 502477 203421 502609 207685
rect 504465 203421 504501 207685
rect 504501 203421 505649 207685
rect 507665 203421 507701 207685
rect 507701 203421 508769 207685
rect 510705 203421 511757 207685
rect 511757 203421 511809 207685
rect 496225 203338 497409 203421
rect 498705 203338 499889 203421
rect 501505 203338 502609 203421
rect 504465 203338 505649 203421
rect 507665 203338 508769 203421
rect 510705 203338 511809 203421
rect 513105 203338 514209 207754
rect 516065 207685 517249 207754
rect 518545 207685 519729 207754
rect 521265 207685 522449 207754
rect 523985 207685 525169 207754
rect 527185 207685 528289 207754
rect 530225 207685 531329 207754
rect 532545 207685 533729 207754
rect 535585 207685 536769 207754
rect 538065 207685 539169 207754
rect 540785 207685 541969 207754
rect 516065 203421 517117 207685
rect 517117 203421 517249 207685
rect 518545 203421 519597 207685
rect 519597 203421 519729 207685
rect 521265 203421 522237 207685
rect 522237 203421 522449 207685
rect 523985 203421 524021 207685
rect 524021 203421 525169 207685
rect 527185 203421 527221 207685
rect 527221 203421 528289 207685
rect 530225 203421 531277 207685
rect 531277 203421 531329 207685
rect 532545 203421 532581 207685
rect 532581 203421 533729 207685
rect 535585 203421 536637 207685
rect 536637 203421 536769 207685
rect 538065 203421 539117 207685
rect 539117 203421 539169 207685
rect 540785 203421 541757 207685
rect 541757 203421 541969 207685
rect 516065 203338 517249 203421
rect 518545 203338 519729 203421
rect 521265 203338 522449 203421
rect 523985 203338 525169 203421
rect 527185 203338 528289 203421
rect 530225 203338 531329 203421
rect 532545 203338 533729 203421
rect 535585 203338 536769 203421
rect 538065 203338 539169 203421
rect 540785 203338 541969 203421
rect 484661 202245 543997 203338
rect 543997 202245 544129 203338
rect 484625 202234 490741 202245
rect 490741 202234 494397 202245
rect 494397 202234 496101 202245
rect 496101 202234 499757 202245
rect 499757 202234 510581 202245
rect 510581 202234 514237 202245
rect 514237 202234 515941 202245
rect 515941 202234 519597 202245
rect 519597 202234 530101 202245
rect 530101 202234 533757 202245
rect 533757 202234 535461 202245
rect 535461 202234 539117 202245
rect 539117 202234 544129 202245
rect 490865 202165 494369 202234
rect 496225 202165 499757 202234
rect 499757 202165 499889 202234
rect 490865 202154 494369 202165
rect 496225 202154 499889 202165
rect 501505 202154 502609 202234
rect 510705 202165 514209 202234
rect 516065 202165 519597 202234
rect 519597 202165 519729 202234
rect 510705 202154 514209 202165
rect 516065 202154 519729 202165
rect 521265 202154 522449 202234
rect 530225 202165 533729 202234
rect 535585 202165 539117 202234
rect 539117 202165 539169 202234
rect 530225 202154 533729 202165
rect 535585 202154 539169 202165
rect 540785 202154 541969 202234
rect 84614 164729 84678 164733
rect 84614 164673 84618 164729
rect 84618 164673 84674 164729
rect 84674 164673 84678 164729
rect 84614 164669 84678 164673
rect 84694 164729 84758 164733
rect 84694 164673 84698 164729
rect 84698 164673 84754 164729
rect 84754 164673 84758 164729
rect 84694 164669 84758 164673
rect 84774 164729 84838 164733
rect 84774 164673 84778 164729
rect 84778 164673 84834 164729
rect 84834 164673 84838 164729
rect 84774 164669 84838 164673
rect 84854 164729 84918 164733
rect 84854 164673 84858 164729
rect 84858 164673 84914 164729
rect 84914 164673 84918 164729
rect 84854 164669 84918 164673
rect 84934 164729 84998 164733
rect 84934 164673 84938 164729
rect 84938 164673 84994 164729
rect 84994 164673 84998 164729
rect 84934 164669 84998 164673
rect 85014 164729 85078 164733
rect 85014 164673 85018 164729
rect 85018 164673 85074 164729
rect 85074 164673 85078 164729
rect 85014 164669 85078 164673
rect 85094 164729 85158 164733
rect 85094 164673 85098 164729
rect 85098 164673 85154 164729
rect 85154 164673 85158 164729
rect 85094 164669 85158 164673
rect 85174 164729 85238 164733
rect 85174 164673 85178 164729
rect 85178 164673 85234 164729
rect 85234 164673 85238 164729
rect 85174 164669 85238 164673
rect 85254 164728 85318 164733
rect 85254 164672 85259 164728
rect 85259 164672 85315 164728
rect 85315 164672 85318 164728
rect 85254 164669 85318 164672
rect 85347 164729 85411 164733
rect 85347 164673 85351 164729
rect 85351 164673 85407 164729
rect 85407 164673 85411 164729
rect 85347 164669 85411 164673
rect 79738 164271 79802 164275
rect 79738 164215 79742 164271
rect 79742 164215 79798 164271
rect 79798 164215 79802 164271
rect 79738 164211 79802 164215
rect 79738 164191 79802 164195
rect 79738 164135 79742 164191
rect 79742 164135 79798 164191
rect 79798 164135 79802 164191
rect 79738 164131 79802 164135
rect 79738 164111 79802 164115
rect 79738 164055 79742 164111
rect 79742 164055 79798 164111
rect 79798 164055 79802 164111
rect 79738 164051 79802 164055
rect 79738 164031 79802 164035
rect 79738 163975 79742 164031
rect 79742 163975 79798 164031
rect 79798 163975 79802 164031
rect 79738 163971 79802 163975
rect 79738 163951 79802 163955
rect 79738 163895 79742 163951
rect 79742 163895 79798 163951
rect 79798 163895 79802 163951
rect 79738 163891 79802 163895
rect 79738 163871 79802 163875
rect 79738 163815 79742 163871
rect 79742 163815 79798 163871
rect 79798 163815 79802 163871
rect 79738 163811 79802 163815
rect 79738 163791 79802 163795
rect 79738 163735 79742 163791
rect 79742 163735 79798 163791
rect 79798 163735 79802 163791
rect 79738 163731 79802 163735
rect 79738 163711 79802 163715
rect 79738 163655 79742 163711
rect 79742 163655 79798 163711
rect 79798 163655 79802 163711
rect 79738 163651 79802 163655
rect 79738 163631 79802 163635
rect 79738 163575 79742 163631
rect 79742 163575 79798 163631
rect 79798 163575 79802 163631
rect 79738 163571 79802 163575
rect 79738 163551 79802 163555
rect 79738 163495 79742 163551
rect 79742 163495 79798 163551
rect 79798 163495 79802 163551
rect 79738 163491 79802 163495
rect 475417 147348 475481 147352
rect 475417 147292 475421 147348
rect 475421 147292 475477 147348
rect 475477 147292 475481 147348
rect 475417 147288 475481 147292
rect 475517 147348 475581 147352
rect 475517 147292 475521 147348
rect 475521 147292 475577 147348
rect 475577 147292 475581 147348
rect 475517 147288 475581 147292
rect 475617 147348 475681 147352
rect 475617 147292 475621 147348
rect 475621 147292 475677 147348
rect 475677 147292 475681 147348
rect 475617 147288 475681 147292
rect 475717 147348 475781 147352
rect 475717 147292 475721 147348
rect 475721 147292 475777 147348
rect 475777 147292 475781 147348
rect 475717 147288 475781 147292
rect 475817 147348 475881 147352
rect 475817 147292 475821 147348
rect 475821 147292 475877 147348
rect 475877 147292 475881 147348
rect 475817 147288 475881 147292
rect 475917 147348 475981 147352
rect 475917 147292 475921 147348
rect 475921 147292 475977 147348
rect 475977 147292 475981 147348
rect 475917 147288 475981 147292
rect 476017 147348 476081 147352
rect 476017 147292 476021 147348
rect 476021 147292 476077 147348
rect 476077 147292 476081 147348
rect 476017 147288 476081 147292
rect 476117 147348 476181 147352
rect 476117 147292 476121 147348
rect 476121 147292 476177 147348
rect 476177 147292 476181 147348
rect 476117 147288 476181 147292
rect 465017 145083 465241 145087
rect 465017 144867 465021 145083
rect 465021 144867 465237 145083
rect 465237 144867 465241 145083
rect 465017 144863 465241 144867
rect 465052 143568 465196 143572
rect 465052 143432 465056 143568
rect 465056 143432 465192 143568
rect 465192 143432 465196 143568
rect 465052 143428 465196 143432
rect 107298 64680 109042 64684
rect 107298 63024 107302 64680
rect 107302 63024 109038 64680
rect 109038 63024 109042 64680
rect 107298 63020 109042 63024
rect 20977 20050 21361 20434
rect 475322 142758 475386 142762
rect 475322 142702 475326 142758
rect 475326 142702 475382 142758
rect 475382 142702 475386 142758
rect 475322 142698 475386 142702
rect 475403 142758 475467 142762
rect 475403 142702 475407 142758
rect 475407 142702 475463 142758
rect 475463 142702 475467 142758
rect 475403 142698 475467 142702
rect 475484 142758 475548 142762
rect 475484 142702 475488 142758
rect 475488 142702 475544 142758
rect 475544 142702 475548 142758
rect 475484 142698 475548 142702
rect 475565 142758 475629 142762
rect 475565 142702 475569 142758
rect 475569 142702 475625 142758
rect 475625 142702 475629 142758
rect 475565 142698 475629 142702
rect 475646 142758 475710 142762
rect 475646 142702 475650 142758
rect 475650 142702 475706 142758
rect 475706 142702 475710 142758
rect 475646 142698 475710 142702
rect 475322 142676 475386 142680
rect 475322 142620 475326 142676
rect 475326 142620 475382 142676
rect 475382 142620 475386 142676
rect 475322 142616 475386 142620
rect 475403 142676 475467 142680
rect 475403 142620 475407 142676
rect 475407 142620 475463 142676
rect 475463 142620 475467 142676
rect 475403 142616 475467 142620
rect 475484 142676 475548 142680
rect 475484 142620 475488 142676
rect 475488 142620 475544 142676
rect 475544 142620 475548 142676
rect 475484 142616 475548 142620
rect 475565 142676 475629 142680
rect 475565 142620 475569 142676
rect 475569 142620 475625 142676
rect 475625 142620 475629 142676
rect 475565 142616 475629 142620
rect 475646 142676 475710 142680
rect 475646 142620 475650 142676
rect 475650 142620 475706 142676
rect 475706 142620 475710 142676
rect 475646 142616 475710 142620
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 320117 693838 324135 694407
rect 165594 691832 170594 692506
rect 165594 689288 166450 691832
rect 169714 689288 170594 691832
rect 320117 690814 320613 693838
rect 323557 690814 324135 693838
rect 320117 690389 324135 690814
rect 165594 688526 170594 689288
rect 216844 687759 222114 688348
rect 216844 686724 217814 687759
rect 184756 684464 217814 686724
rect 184756 594827 186169 684464
rect 216844 684003 217814 684464
rect 221250 684003 222114 687759
rect 216844 683264 222114 684003
rect 184756 594774 194253 594827
rect 184756 594726 194002 594774
rect 141750 594390 194002 594726
rect 194146 594390 194253 594774
rect 141750 594208 194253 594390
rect 131630 593734 131748 593788
rect 131630 593670 131735 593734
rect 131630 593623 131748 593670
rect 41684 591932 89712 591934
rect 37928 590710 89712 591932
rect 37928 551854 41254 590710
rect 89483 581816 89712 590710
rect 89490 581782 89712 581816
rect 89792 581529 121900 581596
rect 89792 581513 121526 581529
rect 89792 581289 89865 581513
rect 90009 581385 121526 581513
rect 121830 581385 121900 581529
rect 90009 581312 121900 581385
rect 90009 581289 90096 581312
rect 89792 581200 90096 581289
rect 90482 581172 120744 581228
rect 90482 581059 120422 581172
rect 90482 580995 90559 581059
rect 90623 581028 120422 581059
rect 120646 581028 120744 581172
rect 90623 581020 120744 581028
rect 90623 580995 90732 581020
rect 90482 580979 90732 580995
rect 90482 580915 90559 580979
rect 90623 580915 90732 580979
rect 92254 580976 120744 581020
rect 90482 580844 90732 580915
rect 91026 580853 91152 580882
rect 91026 580789 91057 580853
rect 91121 580789 91152 580853
rect 91026 580773 91152 580789
rect 91026 580709 91057 580773
rect 91121 580709 91152 580773
rect 91026 580680 91152 580709
rect 37928 551214 42430 551854
rect 37928 548430 38602 551214
rect 41546 548430 42430 551214
rect 37928 547750 42430 548430
rect 101833 539626 103172 539836
rect 101833 539390 102055 539626
rect 102291 539390 102415 539626
rect 102651 539390 103172 539626
rect 101833 539277 103172 539390
rect 101833 539041 102053 539277
rect 102289 539041 102413 539277
rect 102649 539041 103172 539277
rect 101833 538834 103172 539041
rect 186640 525408 191917 525659
rect 128449 525028 191917 525408
rect 128449 524829 187358 525028
rect 186640 523204 187358 524829
rect 191262 524844 191917 525028
rect 191262 524788 191918 524844
rect 191262 523204 191917 524788
rect 186640 522626 191917 523204
rect 145661 502335 147444 502592
rect 144950 502074 147444 502335
rect 145661 501844 147444 502074
rect 110471 501470 110595 501772
rect 111463 501470 111598 501797
rect 112498 501470 112625 501783
rect 110131 501344 112625 501470
rect 104611 500923 106512 501019
rect 104611 500827 106896 500923
rect 104611 500683 107535 500827
rect 104611 500620 108845 500683
rect 110131 500620 110278 501344
rect 104611 500448 110279 500620
rect 104611 500385 108845 500448
rect 104611 500207 107535 500385
rect 104611 500106 106896 500207
rect 104611 500034 106512 500106
rect 95272 493461 110101 494394
rect 70254 477270 72893 477611
rect 70254 475606 70706 477270
rect 72450 475933 72893 477270
rect 117157 475933 117895 478544
rect 72450 475606 117895 475933
rect 70254 475195 117895 475606
rect 36296 471852 41254 472350
rect 36296 467788 36953 471852
rect 40457 470831 41254 471852
rect 40457 469993 76265 470831
rect 40457 467788 41254 469993
rect 36296 467330 41254 467788
rect 43996 427274 47596 427328
rect 43996 427272 70968 427274
rect 43996 426927 72262 427272
rect 43996 424783 44638 426927
rect 47182 424783 72262 426927
rect 43996 424388 72262 424783
rect 44002 424382 72262 424388
rect 70975 302419 72257 424382
rect 75427 307521 76265 469993
rect 75427 306683 132563 307521
rect 70975 301137 128187 302419
rect 2846 296171 8410 296865
rect 2846 296165 3622 296171
rect 7698 296165 8410 296171
rect 2846 292101 3588 296165
rect 7732 292101 8410 296165
rect 2846 292095 3622 292101
rect 7698 292095 8410 292101
rect 2846 291336 8410 292095
rect 97797 63408 98267 66513
rect 106942 64684 109354 64999
rect 106942 63418 107298 64684
rect 102603 63408 107298 63418
rect 95593 63142 107298 63408
rect 87866 63020 107298 63142
rect 109042 63020 109354 64684
rect 87866 62802 109354 63020
rect 95593 62637 109354 62802
rect 95593 62635 106989 62637
rect 95593 62632 103360 62635
rect 126905 29035 128187 301137
rect 131725 33127 132563 306683
rect 542475 233289 548167 233663
rect 542475 231494 542910 233289
rect 523210 231467 542910 231494
rect 503715 231435 542910 231467
rect 483653 231289 542910 231435
rect 483653 231209 523470 231289
rect 483653 224505 483870 231209
rect 485054 229640 487070 230025
rect 485054 226066 485448 229640
rect 486785 226066 487070 229640
rect 485054 225609 487070 226066
rect 488254 229640 490057 230025
rect 488254 226066 488580 229640
rect 489755 226066 490057 229640
rect 488254 225609 490057 226066
rect 491294 229640 492510 230025
rect 491294 226066 491550 229640
rect 492223 226066 492510 229640
rect 491294 225609 492510 226066
rect 493614 229640 495470 230025
rect 493614 226066 494018 229640
rect 495099 226066 495470 229640
rect 493614 225609 495470 226066
rect 496693 229640 497950 230025
rect 496693 226066 496894 229640
rect 497621 226066 497950 229640
rect 496693 225609 497950 226066
rect 499134 229640 500670 230025
rect 499134 226066 499416 229640
rect 500225 226066 500670 229640
rect 499134 225609 500670 226066
rect 501854 229640 503950 230025
rect 501854 226066 502020 229640
rect 503715 226066 503950 229640
rect 501854 225609 503950 226066
rect 505134 229672 507150 230105
rect 505134 226098 505503 229672
rect 506840 226098 507150 229672
rect 505134 225689 507150 226098
rect 508254 229672 510190 230105
rect 508254 226098 508635 229672
rect 509810 226098 510190 229672
rect 508254 225689 510190 226098
rect 511294 229672 512510 230105
rect 511294 226098 511605 229672
rect 512278 226098 512510 229672
rect 511294 225689 512510 226098
rect 513694 229672 515550 230025
rect 513694 226098 514073 229672
rect 515154 226098 515550 229672
rect 513694 225689 515550 226098
rect 516734 229672 518030 230105
rect 516734 226098 516949 229672
rect 517676 226098 518030 229672
rect 516734 225689 518030 226098
rect 519134 229672 520750 230105
rect 519134 226098 519471 229672
rect 520280 226098 520750 229672
rect 519134 225689 520750 226098
rect 521934 229672 523470 230105
rect 521934 226098 522075 229672
rect 523210 226098 523470 229672
rect 521934 225689 523470 226098
rect 524574 229699 526590 230105
rect 524574 226125 524998 229699
rect 526335 226125 526590 229699
rect 524574 225689 526590 226125
rect 527774 229699 529630 230105
rect 527774 226125 528130 229699
rect 529305 226125 529630 229699
rect 527774 225689 529630 226125
rect 530814 229699 532030 230105
rect 530814 226125 531100 229699
rect 531773 226125 532030 229699
rect 530814 225689 532030 226125
rect 533214 229699 535070 230105
rect 533214 226125 533568 229699
rect 534649 226125 535070 229699
rect 533214 225689 535070 226125
rect 536174 229699 537417 230105
rect 536174 226125 536444 229699
rect 537171 226125 537417 229699
rect 536174 225689 537417 226125
rect 538654 229699 540270 230105
rect 538654 226125 538966 229699
rect 539775 226125 540270 229699
rect 538654 225689 540270 226125
rect 547694 230105 548167 233289
rect 541454 229699 548167 230105
rect 541454 226125 541570 229699
rect 542475 229677 548167 229699
rect 541454 225689 543795 226125
rect 483653 224399 490057 224505
rect 543534 224505 543795 225689
rect 501854 224425 510217 224505
rect 496693 224399 498057 224425
rect 501813 224399 510217 224425
rect 516533 224399 543795 224505
rect 483653 224330 543795 224399
rect 483653 224303 524300 224330
rect 526335 224316 531100 224330
rect 531773 224316 536444 224330
rect 483653 224271 504245 224303
rect 506840 224289 511605 224303
rect 512278 224289 516949 224303
rect 486785 224257 491550 224271
rect 492223 224257 496894 224271
rect 484413 208938 544341 209155
rect 484413 202234 484625 208938
rect 485809 207360 487825 207754
rect 485809 203786 486208 207360
rect 487545 203786 487825 207360
rect 485809 203338 487825 203786
rect 489009 207360 490732 207754
rect 489009 203786 489340 207360
rect 490515 203786 490732 207360
rect 489009 203338 490732 203786
rect 492049 207360 493265 207754
rect 492049 203786 492310 207360
rect 492983 203786 493265 207360
rect 492049 203338 493265 203786
rect 494488 207360 496225 207754
rect 494488 203786 494778 207360
rect 495859 203786 496225 207360
rect 494488 203338 496225 203786
rect 497409 207360 498705 207754
rect 497409 203786 497654 207360
rect 498381 203786 498705 207360
rect 497409 203338 498705 203786
rect 499889 207360 501505 207754
rect 499889 203786 500176 207360
rect 500985 203786 501505 207360
rect 499889 203338 501505 203786
rect 502609 207360 504465 207754
rect 502609 203786 502780 207360
rect 504238 203786 504465 207360
rect 502609 203338 504465 203786
rect 505649 207360 507665 207754
rect 505649 203786 506033 207360
rect 507370 203786 507665 207360
rect 505649 203338 507665 203786
rect 508769 207360 510572 207754
rect 508769 203786 509165 207360
rect 510340 203786 510572 207360
rect 508769 203338 510572 203786
rect 511809 207360 513105 207754
rect 511809 203786 512135 207360
rect 512808 203786 513105 207360
rect 511809 203338 513105 203786
rect 514328 207360 516065 207754
rect 514328 203786 514603 207360
rect 515684 203786 516065 207360
rect 514328 203338 516065 203786
rect 517249 207360 518545 207754
rect 517249 203786 517479 207360
rect 518206 203786 518545 207360
rect 517249 203338 518545 203786
rect 519729 207360 521265 207754
rect 519729 203786 520001 207360
rect 520810 203786 521265 207360
rect 519729 203338 521265 203786
rect 522449 207360 523985 207754
rect 522449 203786 522605 207360
rect 523749 203786 523985 207360
rect 522449 203338 523985 203786
rect 525169 207360 527185 207754
rect 525169 203786 525544 207360
rect 526881 203786 527185 207360
rect 525169 203338 527185 203786
rect 528289 207360 530092 207754
rect 528289 203786 528676 207360
rect 529851 203786 530092 207360
rect 528289 203338 530092 203786
rect 531329 207360 532545 207754
rect 531329 203786 531646 207360
rect 532319 203786 532545 207360
rect 531329 203338 532545 203786
rect 533848 207360 535585 207754
rect 533848 203786 534114 207360
rect 535195 203786 535585 207360
rect 533848 203338 535585 203786
rect 536769 207360 538065 207754
rect 536769 203786 536990 207360
rect 537717 203786 538065 207360
rect 536769 203338 538065 203786
rect 539169 207360 540785 207754
rect 539169 203786 539512 207360
rect 540321 203786 540785 207360
rect 539169 203338 540785 203786
rect 544129 207754 544341 208938
rect 541969 207360 544341 207754
rect 541969 203786 542116 207360
rect 541969 203338 544341 203786
rect 544129 202234 544341 203338
rect 484413 202201 484652 202234
rect 544088 202201 544341 202234
rect 484413 202154 490865 202201
rect 494369 202154 496225 202201
rect 499889 202154 501505 202201
rect 502609 202154 510705 202201
rect 514209 202154 516065 202201
rect 519729 202154 521265 202201
rect 522449 202154 530225 202201
rect 533729 202154 535585 202201
rect 539169 202154 540785 202201
rect 541969 202154 544341 202201
rect 484413 201991 544341 202154
rect 487545 201977 492310 201991
rect 492983 201977 497654 201991
rect 507370 201977 512135 201991
rect 512808 201977 517479 201991
rect 526881 201977 531646 201991
rect 532319 201977 536990 201991
rect 475058 147352 476380 147408
rect 475058 147288 475417 147352
rect 475481 147288 475517 147352
rect 475581 147288 475617 147352
rect 475681 147288 475717 147352
rect 475781 147288 475817 147352
rect 475881 147288 475917 147352
rect 475981 147288 476017 147352
rect 476081 147288 476117 147352
rect 476181 147288 476380 147352
rect 475058 146749 476380 147288
rect 450922 145087 465322 145418
rect 450922 144863 465017 145087
rect 465241 144863 465322 145087
rect 450922 144822 465322 144863
rect 450922 33127 451760 144822
rect 453019 143598 461826 143781
rect 453019 143572 465248 143598
rect 453019 143428 465052 143572
rect 465196 143428 465248 143572
rect 453019 143409 465248 143428
rect 453019 142846 461826 143409
rect 131725 32289 451760 33127
rect 453021 142310 454308 142846
rect 453021 29035 454305 142310
rect 126905 27753 454305 29035
rect 127087 27693 453215 27753
rect 20849 20434 21484 20578
rect 20849 20050 20977 20434
rect 21361 20050 21484 20434
rect 20849 19943 21484 20050
<< via4 >>
rect 166524 689322 169640 691798
rect 320687 690928 323483 693724
rect 217814 684003 221250 687759
rect 102055 539390 102291 539626
rect 102415 539390 102651 539626
rect 102053 539041 102289 539277
rect 102413 539041 102649 539277
rect 3622 296165 7698 296171
rect 3622 292101 7698 296165
rect 3622 292095 7698 292101
rect 543177 231035 547573 233275
rect 483977 230159 547573 231035
rect 483977 225595 484853 230159
rect 487177 225595 488053 230159
rect 490057 230025 490933 230159
rect 490057 225609 490110 230025
rect 490110 225609 490933 230025
rect 490057 225595 490933 225609
rect 492617 225595 493493 230159
rect 495497 230025 496693 230159
rect 495497 225609 496654 230025
rect 496654 225609 496693 230025
rect 495497 225595 496693 225609
rect 498057 225595 498933 230159
rect 500937 225595 501813 230159
rect 504137 225595 505013 230159
rect 507337 225595 508213 230159
rect 510217 225595 511093 230159
rect 512777 225595 513653 230159
rect 515657 225595 516533 230159
rect 518217 225595 519093 230159
rect 520777 225595 521653 230159
rect 523657 225595 524533 230159
rect 526857 225595 527733 230159
rect 529737 225595 530613 230159
rect 532297 225595 533173 230159
rect 535177 225595 536053 230159
rect 537417 230105 538613 230159
rect 537417 225689 537470 230105
rect 537470 225689 538613 230105
rect 537417 225595 538613 225689
rect 540297 225595 541173 230159
rect 483977 224719 543413 225595
rect 490057 224505 496693 224719
rect 490057 224425 490110 224505
rect 490110 224425 493614 224505
rect 493614 224425 495470 224505
rect 495470 224425 496693 224505
rect 498057 224505 501813 224719
rect 510217 224505 516533 224719
rect 498057 224425 499134 224505
rect 499134 224425 500670 224505
rect 500670 224425 501813 224505
rect 490057 224399 496693 224425
rect 498057 224399 501813 224425
rect 510217 224399 516533 224505
rect 484652 207961 544088 208837
rect 484652 203077 485528 207961
rect 487852 203077 488728 207961
rect 490732 207754 491928 207961
rect 493612 207754 494488 207961
rect 490732 203338 490865 207754
rect 490865 203338 491928 207754
rect 493612 203338 494369 207754
rect 494369 203338 494488 207754
rect 490732 203077 491928 203338
rect 493612 203077 494488 203338
rect 496492 203077 497368 207961
rect 498732 203077 499608 207961
rect 501612 203077 502488 207961
rect 504492 203077 505368 207961
rect 507692 203077 508568 207961
rect 510572 207754 511768 207961
rect 513132 207754 514328 207961
rect 510572 203338 510705 207754
rect 510705 203338 511768 207754
rect 513132 203338 514209 207754
rect 514209 203338 514328 207754
rect 510572 203077 511768 203338
rect 513132 203077 514328 203338
rect 516332 203077 517208 207961
rect 518572 203077 519448 207961
rect 521452 203077 522328 207961
rect 524012 203077 524888 207961
rect 527212 203077 528088 207961
rect 530092 207754 531288 207961
rect 532652 207754 533848 207961
rect 530092 203338 530225 207754
rect 530225 203338 531288 207754
rect 532652 203338 533729 207754
rect 533729 203338 533848 207754
rect 530092 203077 531288 203338
rect 532652 203077 533848 203338
rect 535852 203077 536728 207961
rect 538092 203077 538968 207961
rect 540972 203077 541848 207961
rect 484652 202234 544088 203077
rect 484652 202201 490865 202234
rect 490865 202201 494369 202234
rect 494369 202201 496225 202234
rect 496225 202201 499889 202234
rect 499889 202201 501505 202234
rect 501505 202201 502609 202234
rect 502609 202201 510705 202234
rect 510705 202201 514209 202234
rect 514209 202201 516065 202234
rect 516065 202201 519729 202234
rect 519729 202201 521265 202234
rect 521265 202201 522449 202234
rect 522449 202201 530225 202234
rect 530225 202201 533729 202234
rect 533729 202201 535585 202234
rect 535585 202201 539169 202234
rect 539169 202201 540785 202234
rect 540785 202201 541969 202234
rect 541969 202201 544088 202234
rect 21051 20124 21287 20360
<< metal5 >>
rect 165594 702300 170598 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 165598 691852 170598 702300
rect 165594 691798 170594 691852
rect 165594 689322 166524 691798
rect 169640 689322 170594 691798
rect 165594 688526 170594 689322
rect 218600 688738 221100 702300
rect 320208 702291 323992 702300
rect 320208 694407 323930 702291
rect 320117 693724 324135 694407
rect 320117 690928 320687 693724
rect 323483 690928 324135 693724
rect 320117 690389 324135 690928
rect 216840 688292 222118 688738
rect 216844 687759 222114 688292
rect 216844 684003 217814 687759
rect 221250 684003 222114 687759
rect 216844 683264 222114 684003
rect 2846 296171 8410 296865
rect 2846 292095 3622 296171
rect 7698 292095 8410 296171
rect 2846 291336 8410 292095
rect 4640 86275 8279 291336
rect 542475 233275 548167 233663
rect 542475 231522 543177 233275
rect 523215 231495 543177 231522
rect 503720 231463 543177 231495
rect 483665 231035 543177 231463
rect 483665 224719 483977 231035
rect 547573 230159 548167 233275
rect 484853 229668 487177 230159
rect 484853 226052 485460 229668
rect 486785 226052 487177 229668
rect 484853 225595 487177 226052
rect 488053 229668 490057 230159
rect 488053 226052 488580 229668
rect 489755 226052 490057 229668
rect 488053 225595 490057 226052
rect 490933 229668 492617 230159
rect 490933 226052 491550 229668
rect 492237 226052 492617 229668
rect 490933 225595 492617 226052
rect 493493 229668 495497 230159
rect 493493 226052 494032 229668
rect 495099 226052 495497 229668
rect 493493 225595 495497 226052
rect 496693 229668 498057 230159
rect 496693 226052 496894 229668
rect 497595 226052 498057 229668
rect 496693 225595 498057 226052
rect 498933 229668 500937 230159
rect 498933 226052 499390 229668
rect 500225 226052 500937 229668
rect 498933 225595 500937 226052
rect 501813 229668 504137 230159
rect 501813 226052 502020 229668
rect 503720 226052 504137 229668
rect 501813 225595 504137 226052
rect 505013 229700 507337 230159
rect 505013 226084 505515 229700
rect 506840 226084 507337 229700
rect 505013 225595 507337 226084
rect 508213 229700 510217 230159
rect 508213 226084 508635 229700
rect 509810 226084 510217 229700
rect 508213 225595 510217 226084
rect 511093 229700 512777 230159
rect 511093 226084 511605 229700
rect 512292 226084 512777 229700
rect 511093 225595 512777 226084
rect 513653 229700 515657 230159
rect 513653 226084 514087 229700
rect 515154 226084 515657 229700
rect 513653 225595 515657 226084
rect 516533 229700 518217 230159
rect 516533 226084 516949 229700
rect 517650 226084 518217 229700
rect 516533 225595 518217 226084
rect 519093 229700 520777 230159
rect 519093 226084 519445 229700
rect 520280 226084 520777 229700
rect 519093 225595 520777 226084
rect 521653 229700 523657 230159
rect 521653 226084 522075 229700
rect 523215 226084 523657 229700
rect 521653 225595 523657 226084
rect 524533 229727 526857 230159
rect 524533 226111 525010 229727
rect 526335 226111 526857 229727
rect 524533 225595 526857 226111
rect 527733 229727 529737 230159
rect 527733 226111 528130 229727
rect 529305 226111 529737 229727
rect 527733 225595 529737 226111
rect 530613 229727 532297 230159
rect 530613 226111 531100 229727
rect 531787 226111 532297 229727
rect 530613 225595 532297 226111
rect 533173 229727 535177 230159
rect 533173 226111 533582 229727
rect 534649 226111 535177 229727
rect 533173 225595 535177 226111
rect 536053 229727 537417 230159
rect 536053 226111 536444 229727
rect 537145 226111 537417 229727
rect 536053 225595 537417 226111
rect 538613 229727 540297 230159
rect 538613 226111 538940 229727
rect 539775 226111 540297 229727
rect 538613 225595 540297 226111
rect 541173 229727 548167 230159
rect 541173 226111 541570 229727
rect 542475 229677 548167 229727
rect 541173 225595 543781 226111
rect 543413 224719 543781 225595
rect 483665 224399 490057 224719
rect 496693 224399 498057 224719
rect 501813 224399 510217 224719
rect 516533 224399 543781 224719
rect 483665 224316 543781 224399
rect 483665 224289 524286 224316
rect 529305 224302 533582 224316
rect 534649 224302 538940 224316
rect 483665 224257 504231 224289
rect 509810 224275 514087 224289
rect 515154 224275 519445 224289
rect 489755 224243 494032 224257
rect 495099 224243 499390 224257
rect 484425 208837 544341 209183
rect 484425 202201 484652 208837
rect 544088 207961 544341 208837
rect 485528 207388 487852 207961
rect 485528 203772 486220 207388
rect 487545 203772 487852 207388
rect 485528 203077 487852 203772
rect 488728 207388 490732 207961
rect 488728 203772 489340 207388
rect 490515 203772 490732 207388
rect 488728 203077 490732 203772
rect 491928 207388 493612 207961
rect 491928 203772 492310 207388
rect 492997 203772 493612 207388
rect 491928 203077 493612 203772
rect 494488 207388 496492 207961
rect 494488 203772 494792 207388
rect 495859 203772 496492 207388
rect 494488 203077 496492 203772
rect 497368 207388 498732 207961
rect 497368 203772 497654 207388
rect 498355 203772 498732 207388
rect 497368 203077 498732 203772
rect 499608 207388 501612 207961
rect 499608 203772 500150 207388
rect 500985 203772 501612 207388
rect 499608 203077 501612 203772
rect 502488 207388 504492 207961
rect 502488 203772 502780 207388
rect 504250 203772 504492 207388
rect 502488 203077 504492 203772
rect 505368 207388 507692 207961
rect 505368 203772 506045 207388
rect 507370 203772 507692 207388
rect 505368 203077 507692 203772
rect 508568 207388 510572 207961
rect 508568 203772 509165 207388
rect 510340 203772 510572 207388
rect 508568 203077 510572 203772
rect 511768 207388 513132 207961
rect 511768 203772 512135 207388
rect 512822 203772 513132 207388
rect 511768 203077 513132 203772
rect 514328 207388 516332 207961
rect 514328 203772 514617 207388
rect 515684 203772 516332 207388
rect 514328 203077 516332 203772
rect 517208 207388 518572 207961
rect 517208 203772 517479 207388
rect 518180 203772 518572 207388
rect 517208 203077 518572 203772
rect 519448 207388 521452 207961
rect 519448 203772 519975 207388
rect 520810 203772 521452 207388
rect 519448 203077 521452 203772
rect 522328 207388 524012 207961
rect 522328 203772 522605 207388
rect 523761 203772 524012 207388
rect 522328 203077 524012 203772
rect 524888 207388 527212 207961
rect 524888 203772 525556 207388
rect 526881 203772 527212 207388
rect 524888 203077 527212 203772
rect 528088 207388 530092 207961
rect 528088 203772 528676 207388
rect 529851 203772 530092 207388
rect 528088 203077 530092 203772
rect 531288 207388 532652 207961
rect 531288 203772 531646 207388
rect 532333 203772 532652 207388
rect 531288 203077 532652 203772
rect 533848 207388 535852 207961
rect 533848 203772 534128 207388
rect 535195 203772 535852 207388
rect 533848 203077 535852 203772
rect 536728 207388 538092 207961
rect 536728 203772 536990 207388
rect 537691 203772 538092 207388
rect 536728 203077 538092 203772
rect 538968 207388 540972 207961
rect 538968 203772 539486 207388
rect 540321 203772 540972 207388
rect 538968 203077 540972 203772
rect 541848 207388 544341 207961
rect 541848 203772 542116 207388
rect 541848 203077 544327 203772
rect 544088 202201 544327 203077
rect 484425 201977 544327 202201
rect 490515 201963 494792 201977
rect 495859 201963 500150 201977
rect 510340 201968 514617 201977
rect 515684 201968 519975 201977
rect 529851 201968 534128 201977
rect 535195 201968 539486 201977
rect 4640 85640 93103 86275
rect 75784 77252 89708 77715
rect 75784 77080 89709 77252
rect 75784 58994 76419 77080
rect 89074 66050 89709 77080
rect 88160 65020 89709 66050
rect 92468 66018 93103 85640
rect 88160 64992 89696 65020
rect 92464 64960 94000 66018
rect 70753 58992 74504 58993
rect 75153 58992 76419 58994
rect 20849 58358 76419 58992
rect 20849 58357 70780 58358
rect 71415 58357 76419 58358
rect 20849 20360 21484 58357
rect 20849 20124 21051 20360
rect 21287 20124 21484 20360
rect 20849 19943 21484 20124
use BGR1  BGR1_0
timestamp 1669522153
transform 1 0 75512 0 1 579984
box -2150 -5244 15700 8698
use PA_Lay_2  PA_Lay_2_0
timestamp 1669522153
transform 1 0 86952 0 1 41626
box -9932 -1382 18780 33188
use VCO  VCO_0
timestamp 1669522153
transform 1 0 195720 0 1 594808
box -808 -1396 2776 990
use biasAmp  biasAmp_0
timestamp 1669522153
transform 1 0 117256 0 1 587090
box -9186 2572 -2242 9318
use filter_op_amp  filter_op_amp_0
timestamp 1669522153
transform 1 0 472155 0 1 145116
box -7117 -3066 5267 2367
use lna_bk5  lna_bk5_0
timestamp 1669522153
transform 1 0 112389 0 1 501628
box -28856 -29561 65696 64408
use mixer_layout  mixer_layout_0
timestamp 1669522153
transform 1 0 76518 0 1 158348
box -2746 -924 13715 7860
use rldo_full  rldo_full_0
timestamp 1669522153
transform 1 0 435192 0 1 204384
box 4412 -1856 42026 15135
use tia  tia_0
timestamp 1669522153
transform 1 0 124008 0 1 590341
box -1768 -1627 18245 8897
<< labels >>
rlabel metal2 s 47804 -800 47916 480 4 wbs_adr_i[10]
port 1 nsew
rlabel metal2 s 41894 -800 42006 480 4 wbs_dat_i[8]
port 2 nsew
rlabel metal2 s 27710 -800 27822 480 4 wbs_dat_i[4]
port 3 nsew
rlabel metal2 s 52532 -800 52644 480 4 wbs_dat_i[11]
port 4 nsew
rlabel metal2 s 34802 -800 34914 480 4 wbs_dat_i[6]
port 5 nsew
rlabel metal2 s 70262 -800 70374 480 4 wbs_dat_i[16]
port 6 nsew
rlabel metal2 s 13526 -800 13638 480 4 wbs_dat_i[1]
port 7 nsew
rlabel metal2 s 20618 -800 20730 480 4 wbs_sel_i[2]
port 8 nsew
rlabel metal2 s 43076 -800 43188 480 4 wbs_dat_o[8]
port 9 nsew
rlabel metal2 s 60806 -800 60918 480 4 wbs_dat_o[13]
port 10 nsew
rlabel metal2 s 64352 -800 64464 480 4 wbs_dat_o[14]
port 11 nsew
rlabel metal2 s 22982 -800 23094 480 4 wbs_dat_i[3]
port 12 nsew
rlabel metal2 s 48986 -800 49098 480 4 wbs_dat_i[10]
port 13 nsew
rlabel metal2 s 18254 -800 18366 480 4 wbs_dat_i[2]
port 14 nsew
rlabel metal2 s 8798 -800 8910 480 4 wbs_dat_i[0]
port 15 nsew
rlabel metal2 s 56078 -800 56190 480 4 wbs_dat_i[12]
port 16 nsew
rlabel metal2 s 58442 -800 58554 480 4 wbs_adr_i[13]
port 17 nsew
rlabel metal2 s 45440 -800 45552 480 4 wbs_dat_i[9]
port 18 nsew
rlabel metal2 s 1706 -800 1818 480 4 wb_rst_i
port 19 nsew
rlabel metal2 s 54896 -800 55008 480 4 wbs_adr_i[12]
port 20 nsew
rlabel metal2 s 7616 -800 7728 480 4 wbs_adr_i[0]
port 21 nsew
rlabel metal2 s 39530 -800 39642 480 4 wbs_dat_o[7]
port 22 nsew
rlabel metal2 s 66716 -800 66828 480 4 wbs_dat_i[15]
port 23 nsew
rlabel metal2 s 2888 -800 3000 480 4 wbs_ack_o
port 24 nsew
rlabel metal2 s 26528 -800 26640 480 4 wbs_adr_i[4]
port 25 nsew
rlabel metal2 s 67898 -800 68010 480 4 wbs_dat_o[15]
port 26 nsew
rlabel metal2 s 63170 -800 63282 480 4 wbs_dat_i[14]
port 27 nsew
rlabel metal2 s 69080 -800 69192 480 4 wbs_adr_i[16]
port 28 nsew
rlabel metal2 s 5252 -800 5364 480 4 wbs_stb_i
port 29 nsew
rlabel metal2 s 9980 -800 10092 480 4 wbs_dat_o[0]
port 30 nsew
rlabel metal2 s 37166 -800 37278 480 4 wbs_adr_i[7]
port 31 nsew
rlabel metal2 s 12344 -800 12456 480 4 wbs_adr_i[1]
port 32 nsew
rlabel metal2 s 24164 -800 24276 480 4 wbs_dat_o[3]
port 33 nsew
rlabel metal2 s 72626 -800 72738 480 4 wbs_adr_i[17]
port 34 nsew
rlabel metal2 s 524 -800 636 480 4 wb_clk_i
port 35 nsew
rlabel metal2 s 4070 -800 4182 480 4 wbs_cyc_i
port 36 nsew
rlabel metal2 s 57260 -800 57372 480 4 wbs_dat_o[12]
port 37 nsew
rlabel metal2 s 40712 -800 40824 480 4 wbs_adr_i[8]
port 38 nsew
rlabel metal2 s 51350 -800 51462 480 4 wbs_adr_i[11]
port 39 nsew
rlabel metal2 s 38348 -800 38460 480 4 wbs_dat_i[7]
port 40 nsew
rlabel metal2 s 32438 -800 32550 480 4 wbs_dat_o[5]
port 41 nsew
rlabel metal2 s 46622 -800 46734 480 4 wbs_dat_o[9]
port 42 nsew
rlabel metal2 s 53714 -800 53826 480 4 wbs_dat_o[11]
port 43 nsew
rlabel metal2 s 31256 -800 31368 480 4 wbs_dat_i[5]
port 44 nsew
rlabel metal2 s 15890 -800 16002 480 4 wbs_sel_i[1]
port 45 nsew
rlabel metal2 s 25346 -800 25458 480 4 wbs_sel_i[3]
port 46 nsew
rlabel metal2 s 11162 -800 11274 480 4 wbs_sel_i[0]
port 47 nsew
rlabel metal2 s 44258 -800 44370 480 4 wbs_adr_i[9]
port 48 nsew
rlabel metal2 s 30074 -800 30186 480 4 wbs_adr_i[5]
port 49 nsew
rlabel metal2 s 65534 -800 65646 480 4 wbs_adr_i[15]
port 50 nsew
rlabel metal2 s 35984 -800 36096 480 4 wbs_dat_o[6]
port 51 nsew
rlabel metal2 s 21800 -800 21912 480 4 wbs_adr_i[3]
port 52 nsew
rlabel metal2 s 61988 -800 62100 480 4 wbs_adr_i[14]
port 53 nsew
rlabel metal2 s 59624 -800 59736 480 4 wbs_dat_i[13]
port 54 nsew
rlabel metal2 s 19436 -800 19548 480 4 wbs_dat_o[2]
port 55 nsew
rlabel metal2 s 28892 -800 29004 480 4 wbs_dat_o[4]
port 56 nsew
rlabel metal2 s 14708 -800 14820 480 4 wbs_dat_o[1]
port 57 nsew
rlabel metal2 s 50168 -800 50280 480 4 wbs_dat_o[10]
port 58 nsew
rlabel metal2 s 71444 -800 71556 480 4 wbs_dat_o[16]
port 59 nsew
rlabel metal2 s 17072 -800 17184 480 4 wbs_adr_i[2]
port 60 nsew
rlabel metal2 s 33620 -800 33732 480 4 wbs_adr_i[6]
port 61 nsew
rlabel metal2 s 6434 -800 6546 480 4 wbs_we_i
port 62 nsew
rlabel metal2 s 143546 -800 143658 480 4 la_data_in[5]
port 63 nsew
rlabel metal2 s 103358 -800 103470 480 4 wbs_dat_o[25]
port 64 nsew
rlabel metal2 s 83264 -800 83376 480 4 wbs_adr_i[20]
port 65 nsew
rlabel metal2 s 110450 -800 110562 480 4 wbs_dat_o[27]
port 66 nsew
rlabel metal2 s 124634 -800 124746 480 4 wbs_dat_o[31]
port 67 nsew
rlabel metal2 s 132908 -800 133020 480 4 la_data_in[2]
port 68 nsew
rlabel metal2 s 134090 -800 134202 480 4 la_data_out[2]
port 69 nsew
rlabel metal2 s 122270 -800 122382 480 4 wbs_adr_i[31]
port 70 nsew
rlabel metal2 s 76172 -800 76284 480 4 wbs_adr_i[18]
port 71 nsew
rlabel metal2 s 129362 -800 129474 480 4 la_data_in[1]
port 72 nsew
rlabel metal2 s 140000 -800 140112 480 4 la_data_in[4]
port 73 nsew
rlabel metal2 s 136454 -800 136566 480 4 la_data_in[3]
port 74 nsew
rlabel metal2 s 115178 -800 115290 480 4 wbs_adr_i[29]
port 75 nsew
rlabel metal2 s 128180 -800 128292 480 4 la_oenb[0]
port 76 nsew
rlabel metal2 s 85628 -800 85740 480 4 wbs_dat_o[20]
port 77 nsew
rlabel metal2 s 73808 -800 73920 480 4 wbs_dat_i[17]
port 78 nsew
rlabel metal2 s 123452 -800 123564 480 4 wbs_dat_i[31]
port 79 nsew
rlabel metal2 s 106904 -800 107016 480 4 wbs_dat_o[26]
port 80 nsew
rlabel metal2 s 80900 -800 81012 480 4 wbs_dat_i[19]
port 81 nsew
rlabel metal2 s 137636 -800 137748 480 4 la_data_out[3]
port 82 nsew
rlabel metal2 s 77354 -800 77466 480 4 wbs_dat_i[18]
port 83 nsew
rlabel metal2 s 131726 -800 131838 480 4 la_oenb[1]
port 84 nsew
rlabel metal2 s 145910 -800 146022 480 4 la_oenb[5]
port 85 nsew
rlabel metal2 s 104540 -800 104652 480 4 wbs_adr_i[26]
port 86 nsew
rlabel metal2 s 96266 -800 96378 480 4 wbs_dat_o[23]
port 87 nsew
rlabel metal2 s 98630 -800 98742 480 4 wbs_dat_i[24]
port 88 nsew
rlabel metal2 s 142364 -800 142476 480 4 la_oenb[4]
port 89 nsew
rlabel metal2 s 79718 -800 79830 480 4 wbs_adr_i[19]
port 90 nsew
rlabel metal2 s 119906 -800 120018 480 4 wbs_dat_i[30]
port 91 nsew
rlabel metal2 s 99812 -800 99924 480 4 wbs_dat_o[24]
port 92 nsew
rlabel metal2 s 86810 -800 86922 480 4 wbs_adr_i[21]
port 93 nsew
rlabel metal2 s 89174 -800 89286 480 4 wbs_dat_o[21]
port 94 nsew
rlabel metal2 s 109268 -800 109380 480 4 wbs_dat_i[27]
port 95 nsew
rlabel metal2 s 90356 -800 90468 480 4 wbs_adr_i[22]
port 96 nsew
rlabel metal2 s 93902 -800 94014 480 4 wbs_adr_i[23]
port 97 nsew
rlabel metal2 s 126998 -800 127110 480 4 la_data_out[0]
port 98 nsew
rlabel metal2 s 84446 -800 84558 480 4 wbs_dat_i[20]
port 99 nsew
rlabel metal2 s 74990 -800 75102 480 4 wbs_dat_o[17]
port 100 nsew
rlabel metal2 s 78536 -800 78648 480 4 wbs_dat_o[18]
port 101 nsew
rlabel metal2 s 82082 -800 82194 480 4 wbs_dat_o[19]
port 102 nsew
rlabel metal2 s 117542 -800 117654 480 4 wbs_dat_o[29]
port 103 nsew
rlabel metal2 s 91538 -800 91650 480 4 wbs_dat_i[22]
port 104 nsew
rlabel metal2 s 87992 -800 88104 480 4 wbs_dat_i[21]
port 105 nsew
rlabel metal2 s 138818 -800 138930 480 4 la_oenb[3]
port 106 nsew
rlabel metal2 s 118724 -800 118836 480 4 wbs_adr_i[30]
port 107 nsew
rlabel metal2 s 111632 -800 111744 480 4 wbs_adr_i[28]
port 108 nsew
rlabel metal2 s 144728 -800 144840 480 4 la_data_out[5]
port 109 nsew
rlabel metal2 s 121088 -800 121200 480 4 wbs_dat_o[30]
port 110 nsew
rlabel metal2 s 100994 -800 101106 480 4 wbs_adr_i[25]
port 111 nsew
rlabel metal2 s 112814 -800 112926 480 4 wbs_dat_i[28]
port 112 nsew
rlabel metal2 s 102176 -800 102288 480 4 wbs_dat_i[25]
port 113 nsew
rlabel metal2 s 92720 -800 92832 480 4 wbs_dat_o[22]
port 114 nsew
rlabel metal2 s 113996 -800 114108 480 4 wbs_dat_o[28]
port 115 nsew
rlabel metal2 s 95084 -800 95196 480 4 wbs_dat_i[23]
port 116 nsew
rlabel metal2 s 141182 -800 141294 480 4 la_data_out[4]
port 117 nsew
rlabel metal2 s 130544 -800 130656 480 4 la_data_out[1]
port 118 nsew
rlabel metal2 s 105722 -800 105834 480 4 wbs_dat_i[26]
port 119 nsew
rlabel metal2 s 116360 -800 116472 480 4 wbs_dat_i[29]
port 120 nsew
rlabel metal2 s 135272 -800 135384 480 4 la_oenb[2]
port 121 nsew
rlabel metal2 s 97448 -800 97560 480 4 wbs_adr_i[24]
port 122 nsew
rlabel metal2 s 125816 -800 125928 480 4 la_data_in[0]
port 123 nsew
rlabel metal2 s 108086 -800 108198 480 4 wbs_adr_i[27]
port 124 nsew
rlabel metal2 s 215648 -800 215760 480 4 la_data_out[25]
port 125 nsew
rlabel metal2 s 197918 -800 198030 480 4 la_data_out[20]
port 126 nsew
rlabel metal2 s 151820 -800 151932 480 4 la_data_out[7]
port 127 nsew
rlabel metal2 s 193190 -800 193302 480 4 la_data_in[19]
port 128 nsew
rlabel metal2 s 149456 -800 149568 480 4 la_oenb[6]
port 129 nsew
rlabel metal2 s 168368 -800 168480 480 4 la_data_in[12]
port 130 nsew
rlabel metal2 s 164822 -800 164934 480 4 la_data_in[11]
port 131 nsew
rlabel metal2 s 160094 -800 160206 480 4 la_oenb[9]
port 132 nsew
rlabel metal2 s 205010 -800 205122 480 4 la_data_out[22]
port 133 nsew
rlabel metal2 s 177824 -800 177936 480 4 la_oenb[14]
port 134 nsew
rlabel metal2 s 194372 -800 194484 480 4 la_data_out[19]
port 135 nsew
rlabel metal2 s 216830 -800 216942 480 4 la_oenb[25]
port 136 nsew
rlabel metal2 s 186098 -800 186210 480 4 la_data_in[17]
port 137 nsew
rlabel metal2 s 181370 -800 181482 480 4 la_oenb[15]
port 138 nsew
rlabel metal2 s 174278 -800 174390 480 4 la_oenb[13]
port 139 nsew
rlabel metal2 s 207374 -800 207486 480 4 la_data_in[23]
port 140 nsew
rlabel metal2 s 187280 -800 187392 480 4 la_data_out[17]
port 141 nsew
rlabel metal2 s 196736 -800 196848 480 4 la_data_in[20]
port 142 nsew
rlabel metal2 s 210920 -800 211032 480 4 la_data_in[24]
port 143 nsew
rlabel metal2 s 183734 -800 183846 480 4 la_data_out[16]
port 144 nsew
rlabel metal2 s 182552 -800 182664 480 4 la_data_in[16]
port 145 nsew
rlabel metal2 s 209738 -800 209850 480 4 la_oenb[23]
port 146 nsew
rlabel metal2 s 199100 -800 199212 480 4 la_oenb[20]
port 147 nsew
rlabel metal2 s 201464 -800 201576 480 4 la_data_out[21]
port 148 nsew
rlabel metal2 s 155366 -800 155478 480 4 la_data_out[8]
port 149 nsew
rlabel metal2 s 171914 -800 172026 480 4 la_data_in[13]
port 150 nsew
rlabel metal2 s 180188 -800 180300 480 4 la_data_out[15]
port 151 nsew
rlabel metal2 s 147092 -800 147204 480 4 la_data_in[6]
port 152 nsew
rlabel metal2 s 166004 -800 166116 480 4 la_data_out[11]
port 153 nsew
rlabel metal2 s 162458 -800 162570 480 4 la_data_out[10]
port 154 nsew
rlabel metal2 s 157730 -800 157842 480 4 la_data_in[9]
port 155 nsew
rlabel metal2 s 154184 -800 154296 480 4 la_data_in[8]
port 156 nsew
rlabel metal2 s 188462 -800 188574 480 4 la_oenb[17]
port 157 nsew
rlabel metal2 s 150638 -800 150750 480 4 la_data_in[7]
port 158 nsew
rlabel metal2 s 156548 -800 156660 480 4 la_oenb[8]
port 159 nsew
rlabel metal2 s 218012 -800 218124 480 4 la_data_in[26]
port 160 nsew
rlabel metal2 s 153002 -800 153114 480 4 la_oenb[7]
port 161 nsew
rlabel metal2 s 184916 -800 185028 480 4 la_oenb[16]
port 162 nsew
rlabel metal2 s 214466 -800 214578 480 4 la_data_in[25]
port 163 nsew
rlabel metal2 s 213284 -800 213396 480 4 la_oenb[24]
port 164 nsew
rlabel metal2 s 202646 -800 202758 480 4 la_oenb[21]
port 165 nsew
rlabel metal2 s 206192 -800 206304 480 4 la_oenb[22]
port 166 nsew
rlabel metal2 s 212102 -800 212214 480 4 la_data_out[24]
port 167 nsew
rlabel metal2 s 175460 -800 175572 480 4 la_data_in[14]
port 168 nsew
rlabel metal2 s 208556 -800 208668 480 4 la_data_out[23]
port 169 nsew
rlabel metal2 s 173096 -800 173208 480 4 la_data_out[13]
port 170 nsew
rlabel metal2 s 148274 -800 148386 480 4 la_data_out[6]
port 171 nsew
rlabel metal2 s 163640 -800 163752 480 4 la_oenb[10]
port 172 nsew
rlabel metal2 s 179006 -800 179118 480 4 la_data_in[15]
port 173 nsew
rlabel metal2 s 190826 -800 190938 480 4 la_data_out[18]
port 174 nsew
rlabel metal2 s 192008 -800 192120 480 4 la_oenb[18]
port 175 nsew
rlabel metal2 s 158912 -800 159024 480 4 la_data_out[9]
port 176 nsew
rlabel metal2 s 167186 -800 167298 480 4 la_oenb[11]
port 177 nsew
rlabel metal2 s 189644 -800 189756 480 4 la_data_in[18]
port 178 nsew
rlabel metal2 s 195554 -800 195666 480 4 la_oenb[19]
port 179 nsew
rlabel metal2 s 200282 -800 200394 480 4 la_data_in[21]
port 180 nsew
rlabel metal2 s 176642 -800 176754 480 4 la_data_out[14]
port 181 nsew
rlabel metal2 s 170732 -800 170844 480 4 la_oenb[12]
port 182 nsew
rlabel metal2 s 203828 -800 203940 480 4 la_data_in[22]
port 183 nsew
rlabel metal2 s 161276 -800 161388 480 4 la_data_in[10]
port 184 nsew
rlabel metal2 s 169550 -800 169662 480 4 la_data_out[12]
port 185 nsew
rlabel metal2 s 275930 -800 276042 480 4 la_data_out[42]
port 186 nsew
rlabel metal2 s 286568 -800 286680 480 4 la_data_out[45]
port 187 nsew
rlabel metal2 s 290114 -800 290226 480 4 la_data_out[46]
port 188 nsew
rlabel metal2 s 278294 -800 278406 480 4 la_data_in[43]
port 189 nsew
rlabel metal2 s 281840 -800 281952 480 4 la_data_in[44]
port 190 nsew
rlabel metal2 s 288932 -800 289044 480 4 la_data_in[46]
port 191 nsew
rlabel metal2 s 262928 -800 263040 480 4 la_oenb[38]
port 192 nsew
rlabel metal2 s 259382 -800 259494 480 4 la_oenb[37]
port 193 nsew
rlabel metal2 s 270020 -800 270132 480 4 la_oenb[40]
port 194 nsew
rlabel metal2 s 235742 -800 235854 480 4 la_data_in[31]
port 195 nsew
rlabel metal2 s 233378 -800 233490 480 4 la_data_out[30]
port 196 nsew
rlabel metal2 s 273566 -800 273678 480 4 la_oenb[41]
port 197 nsew
rlabel metal2 s 277112 -800 277224 480 4 la_oenb[42]
port 198 nsew
rlabel metal2 s 280658 -800 280770 480 4 la_oenb[43]
port 199 nsew
rlabel metal2 s 221558 -800 221670 480 4 la_data_in[27]
port 200 nsew
rlabel metal2 s 225104 -800 225216 480 4 la_data_in[28]
port 201 nsew
rlabel metal2 s 284204 -800 284316 480 4 la_oenb[44]
port 202 nsew
rlabel metal2 s 232196 -800 232308 480 4 la_data_in[30]
port 203 nsew
rlabel metal2 s 239288 -800 239400 480 4 la_data_in[32]
port 204 nsew
rlabel metal2 s 249926 -800 250038 480 4 la_data_in[35]
port 205 nsew
rlabel metal2 s 246380 -800 246492 480 4 la_data_in[34]
port 206 nsew
rlabel metal2 s 264110 -800 264222 480 4 la_data_in[39]
port 207 nsew
rlabel metal2 s 220376 -800 220488 480 4 la_oenb[26]
port 208 nsew
rlabel metal2 s 227468 -800 227580 480 4 la_oenb[28]
port 209 nsew
rlabel metal2 s 279476 -800 279588 480 4 la_data_out[43]
port 210 nsew
rlabel metal2 s 234560 -800 234672 480 4 la_oenb[30]
port 211 nsew
rlabel metal2 s 238106 -800 238218 480 4 la_oenb[31]
port 212 nsew
rlabel metal2 s 268838 -800 268950 480 4 la_data_out[40]
port 213 nsew
rlabel metal2 s 241652 -800 241764 480 4 la_oenb[32]
port 214 nsew
rlabel metal2 s 257018 -800 257130 480 4 la_data_in[37]
port 215 nsew
rlabel metal2 s 266474 -800 266586 480 4 la_oenb[39]
port 216 nsew
rlabel metal2 s 245198 -800 245310 480 4 la_oenb[33]
port 217 nsew
rlabel metal2 s 248744 -800 248856 480 4 la_oenb[34]
port 218 nsew
rlabel metal2 s 252290 -800 252402 480 4 la_oenb[35]
port 219 nsew
rlabel metal2 s 271202 -800 271314 480 4 la_data_in[41]
port 220 nsew
rlabel metal2 s 255836 -800 255948 480 4 la_oenb[36]
port 221 nsew
rlabel metal2 s 229832 -800 229944 480 4 la_data_out[29]
port 222 nsew
rlabel metal2 s 244016 -800 244128 480 4 la_data_out[33]
port 223 nsew
rlabel metal2 s 283022 -800 283134 480 4 la_data_out[44]
port 224 nsew
rlabel metal2 s 287750 -800 287862 480 4 la_oenb[45]
port 225 nsew
rlabel metal2 s 231014 -800 231126 480 4 la_oenb[29]
port 226 nsew
rlabel metal2 s 247562 -800 247674 480 4 la_data_out[34]
port 227 nsew
rlabel metal2 s 285386 -800 285498 480 4 la_data_in[45]
port 228 nsew
rlabel metal2 s 258200 -800 258312 480 4 la_data_out[37]
port 229 nsew
rlabel metal2 s 291296 -800 291408 480 4 la_oenb[46]
port 230 nsew
rlabel metal2 s 228650 -800 228762 480 4 la_data_in[29]
port 231 nsew
rlabel metal2 s 236924 -800 237036 480 4 la_data_out[31]
port 232 nsew
rlabel metal2 s 240470 -800 240582 480 4 la_data_out[32]
port 233 nsew
rlabel metal2 s 267656 -800 267768 480 4 la_data_in[40]
port 234 nsew
rlabel metal2 s 260564 -800 260676 480 4 la_data_in[38]
port 235 nsew
rlabel metal2 s 265292 -800 265404 480 4 la_data_out[39]
port 236 nsew
rlabel metal2 s 219194 -800 219306 480 4 la_data_out[26]
port 237 nsew
rlabel metal2 s 251108 -800 251220 480 4 la_data_out[35]
port 238 nsew
rlabel metal2 s 272384 -800 272496 480 4 la_data_out[41]
port 239 nsew
rlabel metal2 s 274748 -800 274860 480 4 la_data_in[42]
port 240 nsew
rlabel metal2 s 254654 -800 254766 480 4 la_data_out[36]
port 241 nsew
rlabel metal2 s 261746 -800 261858 480 4 la_data_out[38]
port 242 nsew
rlabel metal2 s 242834 -800 242946 480 4 la_data_in[33]
port 243 nsew
rlabel metal2 s 223922 -800 224034 480 4 la_oenb[27]
port 244 nsew
rlabel metal2 s 222740 -800 222852 480 4 la_data_out[27]
port 245 nsew
rlabel metal2 s 226286 -800 226398 480 4 la_data_out[28]
port 246 nsew
rlabel metal2 s 253472 -800 253584 480 4 la_data_in[36]
port 247 nsew
rlabel metal2 s 318482 -800 318594 480 4 la_data_out[54]
port 248 nsew
rlabel metal2 s 331484 -800 331596 480 4 la_data_in[58]
port 249 nsew
rlabel metal2 s 362216 -800 362328 480 4 la_oenb[66]
port 250 nsew
rlabel metal2 s 350396 -800 350508 480 4 la_data_out[63]
port 251 nsew
rlabel metal2 s 344486 -800 344598 480 4 la_oenb[61]
port 252 nsew
rlabel metal2 s 307844 -800 307956 480 4 la_data_out[51]
port 253 nsew
rlabel metal2 s 305480 -800 305592 480 4 la_oenb[50]
port 254 nsew
rlabel metal2 s 353942 -800 354054 480 4 la_data_out[64]
port 255 nsew
rlabel metal2 s 320846 -800 320958 480 4 la_data_in[55]
port 256 nsew
rlabel metal2 s 352760 -800 352872 480 4 la_data_in[64]
port 257 nsew
rlabel metal2 s 322028 -800 322140 480 4 la_data_out[55]
port 258 nsew
rlabel metal2 s 356306 -800 356418 480 4 la_data_in[65]
port 259 nsew
rlabel metal2 s 337394 -800 337506 480 4 la_oenb[59]
port 260 nsew
rlabel metal2 s 364580 -800 364692 480 4 la_data_out[67]
port 261 nsew
rlabel metal2 s 338576 -800 338688 480 4 la_data_in[60]
port 262 nsew
rlabel metal2 s 296024 -800 296136 480 4 la_data_in[48]
port 263 nsew
rlabel metal2 s 336212 -800 336324 480 4 la_data_out[59]
port 264 nsew
rlabel metal2 s 351578 -800 351690 480 4 la_oenb[63]
port 265 nsew
rlabel metal2 s 304298 -800 304410 480 4 la_data_out[50]
port 266 nsew
rlabel metal2 s 300752 -800 300864 480 4 la_data_out[49]
port 267 nsew
rlabel metal2 s 349214 -800 349326 480 4 la_data_in[63]
port 268 nsew
rlabel metal2 s 345668 -800 345780 480 4 la_data_in[62]
port 269 nsew
rlabel metal2 s 306662 -800 306774 480 4 la_data_in[51]
port 270 nsew
rlabel metal2 s 294842 -800 294954 480 4 la_oenb[47]
port 271 nsew
rlabel metal2 s 298388 -800 298500 480 4 la_oenb[48]
port 272 nsew
rlabel metal2 s 301934 -800 302046 480 4 la_oenb[49]
port 273 nsew
rlabel metal2 s 309026 -800 309138 480 4 la_oenb[51]
port 274 nsew
rlabel metal2 s 312572 -800 312684 480 4 la_oenb[52]
port 275 nsew
rlabel metal2 s 340940 -800 341052 480 4 la_oenb[60]
port 276 nsew
rlabel metal2 s 316118 -800 316230 480 4 la_oenb[53]
port 277 nsew
rlabel metal2 s 313754 -800 313866 480 4 la_data_in[53]
port 278 nsew
rlabel metal2 s 323210 -800 323322 480 4 la_oenb[55]
port 279 nsew
rlabel metal2 s 319664 -800 319776 480 4 la_oenb[54]
port 280 nsew
rlabel metal2 s 359852 -800 359964 480 4 la_data_in[66]
port 281 nsew
rlabel metal2 s 333848 -800 333960 480 4 la_oenb[58]
port 282 nsew
rlabel metal2 s 348032 -800 348144 480 4 la_oenb[62]
port 283 nsew
rlabel metal2 s 355124 -800 355236 480 4 la_oenb[64]
port 284 nsew
rlabel metal2 s 358670 -800 358782 480 4 la_oenb[65]
port 285 nsew
rlabel metal2 s 292478 -800 292590 480 4 la_data_in[47]
port 286 nsew
rlabel metal2 s 299570 -800 299682 480 4 la_data_in[49]
port 287 nsew
rlabel metal2 s 317300 -800 317412 480 4 la_data_in[54]
port 288 nsew
rlabel metal2 s 303116 -800 303228 480 4 la_data_in[50]
port 289 nsew
rlabel metal2 s 342122 -800 342234 480 4 la_data_in[61]
port 290 nsew
rlabel metal2 s 310208 -800 310320 480 4 la_data_in[52]
port 291 nsew
rlabel metal2 s 314936 -800 315048 480 4 la_data_out[53]
port 292 nsew
rlabel metal2 s 324392 -800 324504 480 4 la_data_in[56]
port 293 nsew
rlabel metal2 s 327938 -800 328050 480 4 la_data_in[57]
port 294 nsew
rlabel metal2 s 335030 -800 335142 480 4 la_data_in[59]
port 295 nsew
rlabel metal2 s 293660 -800 293772 480 4 la_data_out[47]
port 296 nsew
rlabel metal2 s 325574 -800 325686 480 4 la_data_out[56]
port 297 nsew
rlabel metal2 s 326756 -800 326868 480 4 la_oenb[56]
port 298 nsew
rlabel metal2 s 329120 -800 329232 480 4 la_data_out[57]
port 299 nsew
rlabel metal2 s 311390 -800 311502 480 4 la_data_out[52]
port 300 nsew
rlabel metal2 s 332666 -800 332778 480 4 la_data_out[58]
port 301 nsew
rlabel metal2 s 339758 -800 339870 480 4 la_data_out[60]
port 302 nsew
rlabel metal2 s 343304 -800 343416 480 4 la_data_out[61]
port 303 nsew
rlabel metal2 s 346850 -800 346962 480 4 la_data_out[62]
port 304 nsew
rlabel metal2 s 357488 -800 357600 480 4 la_data_out[65]
port 305 nsew
rlabel metal2 s 297206 -800 297318 480 4 la_data_out[48]
port 306 nsew
rlabel metal2 s 361034 -800 361146 480 4 la_data_out[66]
port 307 nsew
rlabel metal2 s 363398 -800 363510 480 4 la_data_in[67]
port 308 nsew
rlabel metal2 s 330302 -800 330414 480 4 la_oenb[57]
port 309 nsew
rlabel metal2 s 424862 -800 424974 480 4 la_data_out[84]
port 310 nsew
rlabel metal2 s 416588 -800 416700 480 4 la_data_in[82]
port 311 nsew
rlabel metal2 s 403586 -800 403698 480 4 la_data_out[78]
port 312 nsew
rlabel metal2 s 366944 -800 367056 480 4 la_data_in[68]
port 313 nsew
rlabel metal2 s 376400 -800 376512 480 4 la_oenb[70]
port 314 nsew
rlabel metal2 s 404768 -800 404880 480 4 la_oenb[78]
port 315 nsew
rlabel metal2 s 368126 -800 368238 480 4 la_data_out[68]
port 316 nsew
rlabel metal2 s 422498 -800 422610 480 4 la_oenb[83]
port 317 nsew
rlabel metal2 s 415406 -800 415518 480 4 la_oenb[81]
port 318 nsew
rlabel metal2 s 383492 -800 383604 480 4 la_oenb[72]
port 319 nsew
rlabel metal2 s 375218 -800 375330 480 4 la_data_out[70]
port 320 nsew
rlabel metal2 s 371672 -800 371784 480 4 la_data_out[69]
port 321 nsew
rlabel metal2 s 420134 -800 420246 480 4 la_data_in[83]
port 322 nsew
rlabel metal2 s 411860 -800 411972 480 4 la_oenb[80]
port 323 nsew
rlabel metal2 s 428408 -800 428520 480 4 la_data_out[85]
port 324 nsew
rlabel metal2 s 431954 -800 432066 480 4 la_data_out[86]
port 325 nsew
rlabel metal2 s 417770 -800 417882 480 4 la_data_out[82]
port 326 nsew
rlabel metal2 s 436682 -800 436794 480 4 la_oenb[87]
port 327 nsew
rlabel metal2 s 397676 -800 397788 480 4 la_oenb[76]
port 328 nsew
rlabel metal2 s 365762 -800 365874 480 4 la_oenb[67]
port 329 nsew
rlabel metal2 s 381128 -800 381240 480 4 la_data_in[72]
port 330 nsew
rlabel metal2 s 407132 -800 407244 480 4 la_data_out[79]
port 331 nsew
rlabel metal2 s 421316 -800 421428 480 4 la_data_out[83]
port 332 nsew
rlabel metal2 s 389402 -800 389514 480 4 la_data_out[74]
port 333 nsew
rlabel metal2 s 377582 -800 377694 480 4 la_data_in[71]
port 334 nsew
rlabel metal2 s 387038 -800 387150 480 4 la_oenb[73]
port 335 nsew
rlabel metal2 s 435500 -800 435612 480 4 la_data_out[87]
port 336 nsew
rlabel metal2 s 384674 -800 384786 480 4 la_data_in[73]
port 337 nsew
rlabel metal2 s 391766 -800 391878 480 4 la_data_in[75]
port 338 nsew
rlabel metal2 s 410678 -800 410790 480 4 la_data_out[80]
port 339 nsew
rlabel metal2 s 372854 -800 372966 480 4 la_oenb[69]
port 340 nsew
rlabel metal2 s 398858 -800 398970 480 4 la_data_in[77]
port 341 nsew
rlabel metal2 s 388220 -800 388332 480 4 la_data_in[74]
port 342 nsew
rlabel metal2 s 402404 -800 402516 480 4 la_data_in[78]
port 343 nsew
rlabel metal2 s 405950 -800 406062 480 4 la_data_in[79]
port 344 nsew
rlabel metal2 s 413042 -800 413154 480 4 la_data_in[81]
port 345 nsew
rlabel metal2 s 423680 -800 423792 480 4 la_data_in[84]
port 346 nsew
rlabel metal2 s 427226 -800 427338 480 4 la_data_in[85]
port 347 nsew
rlabel metal2 s 430772 -800 430884 480 4 la_data_in[86]
port 348 nsew
rlabel metal2 s 434318 -800 434430 480 4 la_data_in[87]
port 349 nsew
rlabel metal2 s 370490 -800 370602 480 4 la_data_in[69]
port 350 nsew
rlabel metal2 s 369308 -800 369420 480 4 la_oenb[68]
port 351 nsew
rlabel metal2 s 379946 -800 380058 480 4 la_oenb[71]
port 352 nsew
rlabel metal2 s 390584 -800 390696 480 4 la_oenb[74]
port 353 nsew
rlabel metal2 s 394130 -800 394242 480 4 la_oenb[75]
port 354 nsew
rlabel metal2 s 401222 -800 401334 480 4 la_oenb[77]
port 355 nsew
rlabel metal2 s 426044 -800 426156 480 4 la_oenb[84]
port 356 nsew
rlabel metal2 s 429590 -800 429702 480 4 la_oenb[85]
port 357 nsew
rlabel metal2 s 433136 -800 433248 480 4 la_oenb[86]
port 358 nsew
rlabel metal2 s 374036 -800 374148 480 4 la_data_in[70]
port 359 nsew
rlabel metal2 s 378764 -800 378876 480 4 la_data_out[71]
port 360 nsew
rlabel metal2 s 382310 -800 382422 480 4 la_data_out[72]
port 361 nsew
rlabel metal2 s 385856 -800 385968 480 4 la_data_out[73]
port 362 nsew
rlabel metal2 s 392948 -800 393060 480 4 la_data_out[75]
port 363 nsew
rlabel metal2 s 418952 -800 419064 480 4 la_oenb[82]
port 364 nsew
rlabel metal2 s 396494 -800 396606 480 4 la_data_out[76]
port 365 nsew
rlabel metal2 s 400040 -800 400152 480 4 la_data_out[77]
port 366 nsew
rlabel metal2 s 414224 -800 414336 480 4 la_data_out[81]
port 367 nsew
rlabel metal2 s 395312 -800 395424 480 4 la_data_in[76]
port 368 nsew
rlabel metal2 s 408314 -800 408426 480 4 la_oenb[79]
port 369 nsew
rlabel metal2 s 409496 -800 409608 480 4 la_data_in[80]
port 370 nsew
rlabel metal2 s 465050 -800 465162 480 4 la_oenb[95]
port 371 nsew
rlabel metal2 s 498146 -800 498258 480 4 la_data_in[105]
port 372 nsew
rlabel metal2 s 467414 -800 467526 480 4 la_data_out[96]
port 373 nsew
rlabel metal2 s 453230 -800 453342 480 4 la_data_out[92]
port 374 nsew
rlabel metal2 s 469778 -800 469890 480 4 la_data_in[97]
port 375 nsew
rlabel metal2 s 486326 -800 486438 480 4 la_oenb[101]
port 376 nsew
rlabel metal2 s 448502 -800 448614 480 4 la_data_in[91]
port 377 nsew
rlabel metal2 s 437864 -800 437976 480 4 la_data_in[88]
port 378 nsew
rlabel metal2 s 483962 -800 484074 480 4 la_data_in[101]
port 379 nsew
rlabel metal2 s 463868 -800 463980 480 4 la_data_out[95]
port 380 nsew
rlabel metal2 s 443774 -800 443886 480 4 la_oenb[89]
port 381 nsew
rlabel metal2 s 450866 -800 450978 480 4 la_oenb[91]
port 382 nsew
rlabel metal2 s 449684 -800 449796 480 4 la_data_out[91]
port 383 nsew
rlabel metal2 s 442592 -800 442704 480 4 la_data_out[89]
port 384 nsew
rlabel metal2 s 499328 -800 499440 480 4 la_data_out[105]
port 385 nsew
rlabel metal2 s 439046 -800 439158 480 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 440228 -800 440340 480 4 la_oenb[88]
port 387 nsew
rlabel metal2 s 500510 -800 500622 480 4 la_oenb[105]
port 388 nsew
rlabel metal2 s 441410 -800 441522 480 4 la_data_in[89]
port 389 nsew
rlabel metal2 s 457958 -800 458070 480 4 la_oenb[93]
port 390 nsew
rlabel metal2 s 507602 -800 507714 480 4 la_oenb[107]
port 391 nsew
rlabel metal2 s 493418 -800 493530 480 4 la_oenb[103]
port 392 nsew
rlabel metal2 s 474506 -800 474618 480 4 la_data_out[98]
port 393 nsew
rlabel metal2 s 504056 -800 504168 480 4 la_oenb[106]
port 394 nsew
rlabel metal2 s 446138 -800 446250 480 4 la_data_out[90]
port 395 nsew
rlabel metal2 s 496964 -800 497076 480 4 la_oenb[104]
port 396 nsew
rlabel metal2 s 489872 -800 489984 480 4 la_oenb[102]
port 397 nsew
rlabel metal2 s 491054 -800 491166 480 4 la_data_in[103]
port 398 nsew
rlabel metal2 s 462686 -800 462798 480 4 la_data_in[95]
port 399 nsew
rlabel metal2 s 479234 -800 479346 480 4 la_oenb[99]
port 400 nsew
rlabel metal2 s 470960 -800 471072 480 4 la_data_out[97]
port 401 nsew
rlabel metal2 s 509966 -800 510078 480 4 la_data_out[108]
port 402 nsew
rlabel metal2 s 506420 -800 506532 480 4 la_data_out[107]
port 403 nsew
rlabel metal2 s 494600 -800 494712 480 4 la_data_in[104]
port 404 nsew
rlabel metal2 s 505238 -800 505350 480 4 la_data_in[107]
port 405 nsew
rlabel metal2 s 481598 -800 481710 480 4 la_data_out[100]
port 406 nsew
rlabel metal2 s 460322 -800 460434 480 4 la_data_out[94]
port 407 nsew
rlabel metal2 s 482780 -800 482892 480 4 la_oenb[100]
port 408 nsew
rlabel metal2 s 452048 -800 452160 480 4 la_data_in[92]
port 409 nsew
rlabel metal2 s 478052 -800 478164 480 4 la_data_out[99]
port 410 nsew
rlabel metal2 s 502874 -800 502986 480 4 la_data_out[106]
port 411 nsew
rlabel metal2 s 447320 -800 447432 480 4 la_oenb[90]
port 412 nsew
rlabel metal2 s 454412 -800 454524 480 4 la_oenb[92]
port 413 nsew
rlabel metal2 s 461504 -800 461616 480 4 la_oenb[94]
port 414 nsew
rlabel metal2 s 468596 -800 468708 480 4 la_oenb[96]
port 415 nsew
rlabel metal2 s 472142 -800 472254 480 4 la_oenb[97]
port 416 nsew
rlabel metal2 s 475688 -800 475800 480 4 la_oenb[98]
port 417 nsew
rlabel metal2 s 487508 -800 487620 480 4 la_data_in[102]
port 418 nsew
rlabel metal2 s 501692 -800 501804 480 4 la_data_in[106]
port 419 nsew
rlabel metal2 s 508784 -800 508896 480 4 la_data_in[108]
port 420 nsew
rlabel metal2 s 480416 -800 480528 480 4 la_data_in[100]
port 421 nsew
rlabel metal2 s 444956 -800 445068 480 4 la_data_in[90]
port 422 nsew
rlabel metal2 s 455594 -800 455706 480 4 la_data_in[93]
port 423 nsew
rlabel metal2 s 459140 -800 459252 480 4 la_data_in[94]
port 424 nsew
rlabel metal2 s 466232 -800 466344 480 4 la_data_in[96]
port 425 nsew
rlabel metal2 s 473324 -800 473436 480 4 la_data_in[98]
port 426 nsew
rlabel metal2 s 476870 -800 476982 480 4 la_data_in[99]
port 427 nsew
rlabel metal2 s 488690 -800 488802 480 4 la_data_out[102]
port 428 nsew
rlabel metal2 s 485144 -800 485256 480 4 la_data_out[101]
port 429 nsew
rlabel metal2 s 492236 -800 492348 480 4 la_data_out[103]
port 430 nsew
rlabel metal2 s 495782 -800 495894 480 4 la_data_out[104]
port 431 nsew
rlabel metal2 s 456776 -800 456888 480 4 la_data_out[93]
port 432 nsew
rlabel metal2 s 548972 -800 549084 480 4 la_data_out[119]
port 433 nsew
rlabel metal2 s 570248 -800 570360 480 4 la_data_out[125]
port 434 nsew
rlabel metal2 s 579704 -800 579816 480 4 user_clock2
port 435 nsew
rlabel metal2 s 533606 -800 533718 480 4 la_data_in[115]
port 436 nsew
rlabel metal2 s 583250 -800 583362 480 4 user_irq[2]
port 437 nsew
rlabel metal2 s 541880 -800 541992 480 4 la_data_out[117]
port 438 nsew
rlabel metal2 s 561974 -800 562086 480 4 la_data_in[123]
port 439 nsew
rlabel metal2 s 566702 -800 566814 480 4 la_data_out[124]
port 440 nsew
rlabel metal2 s 534788 -800 534900 480 4 la_data_out[115]
port 441 nsew
rlabel metal2 s 574976 -800 575088 480 4 la_oenb[126]
port 442 nsew
rlabel metal2 s 552518 -800 552630 480 4 la_data_out[120]
port 443 nsew
rlabel metal2 s 531242 -800 531354 480 4 la_data_out[114]
port 444 nsew
rlabel metal2 s 572612 -800 572724 480 4 la_data_in[126]
port 445 nsew
rlabel metal2 s 520604 -800 520716 480 4 la_data_out[111]
port 446 nsew
rlabel metal2 s 582068 -800 582180 480 4 user_irq[1]
port 447 nsew
rlabel metal2 s 564338 -800 564450 480 4 la_oenb[123]
port 448 nsew
rlabel metal2 s 563156 -800 563268 480 4 la_data_out[123]
port 449 nsew
rlabel metal2 s 537152 -800 537264 480 4 la_data_in[116]
port 450 nsew
rlabel metal2 s 538334 -800 538446 480 4 la_data_out[116]
port 451 nsew
rlabel metal2 s 559610 -800 559722 480 4 la_data_out[122]
port 452 nsew
rlabel metal2 s 573794 -800 573906 480 4 la_data_out[126]
port 453 nsew
rlabel metal2 s 577340 -800 577452 480 4 la_data_out[127]
port 454 nsew
rlabel metal2 s 513512 -800 513624 480 4 la_data_out[109]
port 455 nsew
rlabel metal2 s 532424 -800 532536 480 4 la_oenb[114]
port 456 nsew
rlabel metal2 s 518240 -800 518352 480 4 la_oenb[110]
port 457 nsew
rlabel metal2 s 519422 -800 519534 480 4 la_data_in[111]
port 458 nsew
rlabel metal2 s 546608 -800 546720 480 4 la_oenb[118]
port 459 nsew
rlabel metal2 s 543062 -800 543174 480 4 la_oenb[117]
port 460 nsew
rlabel metal2 s 556064 -800 556176 480 4 la_data_out[121]
port 461 nsew
rlabel metal2 s 545426 -800 545538 480 4 la_data_out[118]
port 462 nsew
rlabel metal2 s 576158 -800 576270 480 4 la_data_in[127]
port 463 nsew
rlabel metal2 s 580886 -800 580998 480 4 user_irq[0]
port 464 nsew
rlabel metal2 s 569066 -800 569178 480 4 la_data_in[125]
port 465 nsew
rlabel metal2 s 578522 -800 578634 480 4 la_oenb[127]
port 466 nsew
rlabel metal2 s 547790 -800 547902 480 4 la_data_in[119]
port 467 nsew
rlabel metal2 s 522968 -800 523080 480 4 la_data_in[112]
port 468 nsew
rlabel metal2 s 521786 -800 521898 480 4 la_oenb[111]
port 469 nsew
rlabel metal2 s 554882 -800 554994 480 4 la_data_in[121]
port 470 nsew
rlabel metal2 s 527696 -800 527808 480 4 la_data_out[113]
port 471 nsew
rlabel metal2 s 551336 -800 551448 480 4 la_data_in[120]
port 472 nsew
rlabel metal2 s 558428 -800 558540 480 4 la_data_in[122]
port 473 nsew
rlabel metal2 s 515876 -800 515988 480 4 la_data_in[110]
port 474 nsew
rlabel metal2 s 517058 -800 517170 480 4 la_data_out[110]
port 475 nsew
rlabel metal2 s 567884 -800 567996 480 4 la_oenb[124]
port 476 nsew
rlabel metal2 s 528878 -800 528990 480 4 la_oenb[113]
port 477 nsew
rlabel metal2 s 539516 -800 539628 480 4 la_oenb[116]
port 478 nsew
rlabel metal2 s 553700 -800 553812 480 4 la_oenb[120]
port 479 nsew
rlabel metal2 s 525332 -800 525444 480 4 la_oenb[112]
port 480 nsew
rlabel metal2 s 512330 -800 512442 480 4 la_data_in[109]
port 481 nsew
rlabel metal2 s 560792 -800 560904 480 4 la_oenb[122]
port 482 nsew
rlabel metal2 s 526514 -800 526626 480 4 la_data_in[113]
port 483 nsew
rlabel metal2 s 524150 -800 524262 480 4 la_data_out[112]
port 484 nsew
rlabel metal2 s 571430 -800 571542 480 4 la_oenb[125]
port 485 nsew
rlabel metal2 s 530060 -800 530172 480 4 la_data_in[114]
port 486 nsew
rlabel metal2 s 565520 -800 565632 480 4 la_data_in[124]
port 487 nsew
rlabel metal2 s 535970 -800 536082 480 4 la_oenb[115]
port 488 nsew
rlabel metal2 s 514694 -800 514806 480 4 la_oenb[109]
port 489 nsew
rlabel metal2 s 544244 -800 544356 480 4 la_data_in[118]
port 490 nsew
rlabel metal2 s 557246 -800 557358 480 4 la_oenb[121]
port 491 nsew
rlabel metal2 s 511148 -800 511260 480 4 la_oenb[108]
port 492 nsew
rlabel metal2 s 540698 -800 540810 480 4 la_data_in[117]
port 493 nsew
rlabel metal2 s 550154 -800 550266 480 4 la_oenb[119]
port 494 nsew
rlabel metal4 s 175894 702300 180894 704800 4 io_analog[6]
port 495 nsew
rlabel metal4 s 217294 702300 222294 704800 4 io_analog[5]
port 496 nsew
rlabel metal4 s 227594 702300 232594 704800 4 io_analog[5]
port 496 nsew
rlabel metal4 s 318994 702300 323994 704800 4 io_analog[4]
port 497 nsew
rlabel metal4 s 329294 702300 334294 704800 4 io_analog[4]
port 497 nsew
rlabel metal3 s 583520 495322 584800 495434 4 gpio_noesd[5]
port 498 nsew
rlabel metal3 s 566594 702300 571594 704800 4 io_analog[1]
port 499 nsew
rlabel metal3 s 583520 358874 584800 358986 4 gpio_analog[2]
port 500 nsew
rlabel metal3 s 582340 540545 584800 545345 4 vdda1
port 501 nsew
rlabel metal3 s 582340 550545 584800 555345 4 vdda1
port 501 nsew
rlabel metal3 s 583520 588290 584800 588402 4 io_out[13]
port 502 nsew
rlabel metal3 s 583520 498868 584800 498980 4 io_out[12]
port 503 nsew
rlabel metal3 s 583520 589472 584800 589584 4 io_oeb[13]
port 504 nsew
rlabel metal3 s 583520 364784 584800 364896 4 io_oeb[9]
port 505 nsew
rlabel metal3 s 583520 410024 584800 410136 4 io_out[10]
port 506 nsew
rlabel metal3 s 583520 361238 584800 361350 4 io_in_3v3[9]
port 507 nsew
rlabel metal3 s 583520 407660 584800 407772 4 io_in_3v3[10]
port 508 nsew
rlabel metal3 s 582340 629784 584800 634584 4 vccd1
port 509 nsew
rlabel metal3 s 582340 639771 584800 644571 4 vccd1
port 509 nsew
rlabel metal3 s 583520 411206 584800 411318 4 io_oeb[10]
port 510 nsew
rlabel metal3 s 583520 496504 584800 496616 4 io_in_3v3[12]
port 511 nsew
rlabel metal3 s 318994 702300 323994 704800 4 io_analog[4]
port 497 nsew
rlabel metal3 s 329294 702300 334294 704800 4 io_analog[4]
port 497 nsew
rlabel metal3 s 583520 450900 584800 451012 4 gpio_noesd[4]
port 512 nsew
rlabel metal3 s 583520 452082 584800 452194 4 io_in_3v3[11]
port 513 nsew
rlabel metal3 s 465394 702300 470394 704800 4 io_analog[2]
port 514 nsew
rlabel metal3 s 583520 363602 584800 363714 4 io_out[9]
port 515 nsew
rlabel metal3 s 583520 583562 584800 583674 4 gpio_analog[6]
port 516 nsew
rlabel metal3 s 510594 702340 515394 704800 4 vssa1
port 517 nsew
rlabel metal3 s 520594 702340 525394 704800 4 vssa1
port 517 nsew
rlabel metal3 s 583520 587108 584800 587220 4 io_in[13]
port 518 nsew
rlabel metal3 s 413394 702300 418394 704800 4 io_analog[3]
port 519 nsew
rlabel metal3 s 583520 449718 584800 449830 4 gpio_analog[4]
port 520 nsew
rlabel metal3 s 583520 360056 584800 360168 4 gpio_noesd[2]
port 521 nsew
rlabel metal3 s 583520 584744 584800 584856 4 gpio_noesd[6]
port 522 nsew
rlabel metal3 s 583520 455628 584800 455740 4 io_oeb[11]
port 523 nsew
rlabel metal3 s 326794 702300 328994 704800 4 io_clamp_high[0]
port 524 nsew
rlabel metal3 s 583520 494140 584800 494252 4 gpio_analog[5]
port 525 nsew
rlabel metal3 s 583520 408842 584800 408954 4 io_in[10]
port 526 nsew
rlabel metal3 s 583520 405296 584800 405408 4 gpio_analog[3]
port 527 nsew
rlabel metal3 s 583520 585926 584800 586038 4 io_in_3v3[13]
port 528 nsew
rlabel metal3 s 582300 677984 584800 682984 4 io_analog[0]
port 529 nsew
rlabel metal3 s 324294 702300 326494 704800 4 io_clamp_low[0]
port 530 nsew
rlabel metal3 s 583520 362420 584800 362532 4 io_in[9]
port 531 nsew
rlabel metal3 s 583520 454446 584800 454558 4 io_out[11]
port 532 nsew
rlabel metal3 s 583520 453264 584800 453376 4 io_in[11]
port 533 nsew
rlabel metal3 s 583520 497686 584800 497798 4 io_in[12]
port 534 nsew
rlabel metal3 s 583520 406478 584800 406590 4 gpio_noesd[3]
port 535 nsew
rlabel metal3 s 583520 500050 584800 500162 4 io_oeb[12]
port 536 nsew
rlabel metal3 s -800 423904 480 424016 4 gpio_noesd[9]
port 537 nsew
rlabel metal3 s 175894 702300 180894 704800 4 io_analog[6]
port 495 nsew
rlabel metal3 s 68194 702300 73194 704800 4 io_analog[8]
port 538 nsew
rlabel metal3 s -800 465944 480 466056 4 io_in_3v3[15]
port 539 nsew
rlabel metal3 s -800 506802 480 506914 4 io_out[14]
port 540 nsew
rlabel metal3 s -800 381864 480 381976 4 gpio_analog[10]
port 541 nsew
rlabel metal3 s -800 505620 480 505732 4 io_oeb[14]
port 542 nsew
rlabel metal3 s 16194 702300 21194 704800 4 io_analog[9]
port 543 nsew
rlabel metal3 s -800 378318 480 378430 4 io_in[17]
port 544 nsew
rlabel metal3 s -800 425086 480 425198 4 gpio_analog[9]
port 545 nsew
rlabel metal3 s 225094 702300 227294 704800 4 io_clamp_high[1]
port 546 nsew
rlabel metal3 s 0 680242 1700 685242 4 io_analog[10]
port 547 nsew
rlabel metal3 s 120194 702300 125194 704800 4 io_analog[7]
port 548 nsew
rlabel metal3 s 173394 702300 175594 704800 4 io_clamp_high[2]
port 549 nsew
rlabel metal3 s -800 421540 480 421652 4 io_in[16]
port 550 nsew
rlabel metal3 s 217294 702300 222294 704800 4 io_analog[5]
port 496 nsew
rlabel metal3 s 227594 702300 232594 704800 4 io_analog[5]
port 496 nsew
rlabel metal3 s -800 422722 480 422834 4 io_in_3v3[16]
port 551 nsew
rlabel metal3 s -800 462398 480 462510 4 io_oeb[15]
port 552 nsew
rlabel metal3 s -800 419176 480 419288 4 io_oeb[16]
port 553 nsew
rlabel metal3 s -800 375954 480 376066 4 io_oeb[17]
port 554 nsew
rlabel metal3 s -800 467126 480 467238 4 gpio_noesd[8]
port 555 nsew
rlabel metal3 s 222594 702300 224794 704800 4 io_clamp_low[1]
port 556 nsew
rlabel metal3 s -800 420358 480 420470 4 io_out[16]
port 557 nsew
rlabel metal3 s 170894 702300 173094 704800 4 io_clamp_low[2]
port 558 nsew
rlabel metal3 s -800 379500 480 379612 4 io_in_3v3[17]
port 559 nsew
rlabel metal3 s 0 633842 1660 638642 4 vccd2
port 560 nsew
rlabel metal3 s 0 643842 1660 648642 4 vccd2
port 560 nsew
rlabel metal3 s -800 509166 480 509278 4 io_in_3v3[14]
port 561 nsew
rlabel metal3 s -800 511530 480 511642 4 gpio_analog[7]
port 562 nsew
rlabel metal3 s -800 377136 480 377248 4 io_out[17]
port 563 nsew
rlabel metal3 s -800 468308 480 468420 4 gpio_analog[8]
port 564 nsew
rlabel metal3 s -800 464762 480 464874 4 io_in[15]
port 565 nsew
rlabel metal3 s 0 549442 1660 554242 4 vssa2
port 566 nsew
rlabel metal3 s 0 559442 1660 564242 4 vssa2
port 566 nsew
rlabel metal3 s -800 380682 480 380794 4 gpio_noesd[10]
port 567 nsew
rlabel metal3 s -800 507984 480 508096 4 io_in[14]
port 568 nsew
rlabel metal3 s -800 510348 480 510460 4 gpio_noesd[7]
port 569 nsew
rlabel metal3 s 165598 702300 170598 704800 4 io_analog[6]
port 495 nsew
rlabel metal3 s -800 463580 480 463692 4 io_out[15]
port 570 nsew
rlabel metal3 s -800 333914 480 334026 4 io_out[18]
port 571 nsew
rlabel metal3 s -800 80372 480 80484 4 gpio_noesd[15]
port 572 nsew
rlabel metal3 s -800 251216 480 251328 4 gpio_noesd[13]
port 573 nsew
rlabel metal3 s -800 3908 480 4020 4 io_in[26]
port 574 nsew
rlabel metal3 s -800 16910 480 17022 4 gpio_analog[17]
port 575 nsew
rlabel metal3 s -800 13364 480 13476 4 io_in[24]
port 576 nsew
rlabel metal3 s -800 34786 480 34898 4 io_in[23]
port 577 nsew
rlabel metal3 s -800 35968 480 36080 4 io_in_3v3[23]
port 578 nsew
rlabel metal3 s -800 124776 480 124888 4 gpio_analog[14]
port 579 nsew
rlabel metal3 s -800 78008 480 78120 4 io_in[22]
port 580 nsew
rlabel metal3 s -800 1544 480 1656 4 io_oeb[26]
port 581 nsew
rlabel metal3 s -800 335096 480 335208 4 io_in[18]
port 582 nsew
rlabel metal3 s -800 76826 480 76938 4 io_out[22]
port 583 nsew
rlabel metal3 s 0 162888 1660 167688 4 vssd2
port 584 nsew
rlabel metal3 s 0 172888 1660 177688 4 vssd2
port 584 nsew
rlabel metal3 s -800 122412 480 122524 4 io_in_3v3[21]
port 585 nsew
rlabel metal3 s -800 32422 480 32534 4 io_oeb[23]
port 586 nsew
rlabel metal3 s -800 118866 480 118978 4 io_oeb[21]
port 587 nsew
rlabel metal3 s -800 11000 480 11112 4 io_oeb[24]
port 588 nsew
rlabel metal3 s -800 9818 480 9930 4 io_in_3v3[25]
port 589 nsew
rlabel metal3 s 0 204888 1660 209688 4 vdda2
port 590 nsew
rlabel metal3 s 0 214888 1660 219688 4 vdda2
port 590 nsew
rlabel metal3 s -800 252398 480 252510 4 gpio_analog[13]
port 591 nsew
rlabel metal3 s -800 5090 480 5202 4 io_in_3v3[26]
port 592 nsew
rlabel metal3 s -800 293056 480 293168 4 io_in_3v3[19]
port 593 nsew
rlabel metal3 s -800 246488 480 246600 4 io_oeb[20]
port 594 nsew
rlabel metal3 s -800 336278 480 336390 4 io_in_3v3[18]
port 595 nsew
rlabel metal3 s -800 15728 480 15840 4 gpio_noesd[17]
port 596 nsew
rlabel metal3 s -800 250034 480 250146 4 io_in_3v3[20]
port 597 nsew
rlabel metal3 s -800 294238 480 294350 4 gpio_noesd[12]
port 598 nsew
rlabel metal3 s -800 37150 480 37262 4 gpio_noesd[16]
port 599 nsew
rlabel metal3 s -800 2726 480 2838 4 io_out[26]
port 600 nsew
rlabel metal3 s -800 81554 480 81666 4 gpio_analog[15]
port 601 nsew
rlabel metal3 s -800 295420 480 295532 4 gpio_analog[12]
port 602 nsew
rlabel metal3 s -800 7454 480 7566 4 io_out[25]
port 603 nsew
rlabel metal3 s -800 12182 480 12294 4 io_out[24]
port 604 nsew
rlabel metal3 s -800 248852 480 248964 4 io_in[20]
port 605 nsew
rlabel metal3 s -800 337460 480 337572 4 gpio_noesd[11]
port 606 nsew
rlabel metal3 s -800 33604 480 33716 4 io_out[23]
port 607 nsew
rlabel metal3 s -800 8636 480 8748 4 io_in[25]
port 608 nsew
rlabel metal3 s -800 14546 480 14658 4 io_in_3v3[24]
port 609 nsew
rlabel metal3 s -800 38332 480 38444 4 gpio_analog[16]
port 610 nsew
rlabel metal3 s -800 338642 480 338754 4 gpio_analog[11]
port 611 nsew
rlabel metal3 s -800 123594 480 123706 4 gpio_noesd[14]
port 612 nsew
rlabel metal3 s -800 120048 480 120160 4 io_out[21]
port 613 nsew
rlabel metal3 s -800 332732 480 332844 4 io_oeb[18]
port 614 nsew
rlabel metal3 s -800 291874 480 291986 4 io_in[19]
port 615 nsew
rlabel metal3 s -800 247670 480 247782 4 io_out[20]
port 616 nsew
rlabel metal3 s -800 121230 480 121342 4 io_in[21]
port 617 nsew
rlabel metal3 s -800 290692 480 290804 4 io_out[19]
port 618 nsew
rlabel metal3 s -800 289510 480 289622 4 io_oeb[19]
port 619 nsew
rlabel metal3 s -800 79190 480 79302 4 io_in_3v3[22]
port 620 nsew
rlabel metal3 s -800 75644 480 75756 4 io_oeb[22]
port 621 nsew
rlabel metal3 s -800 6272 480 6384 4 io_oeb[25]
port 622 nsew
rlabel metal3 s 583520 93936 584800 94048 4 io_out[6]
port 623 nsew
rlabel metal3 s 583520 49278 584800 49390 4 io_out[5]
port 624 nsew
rlabel metal3 s 583520 1544 584800 1656 4 io_in_3v3[0]
port 625 nsew
rlabel metal3 s 583520 9818 584800 9930 4 io_oeb[1]
port 626 nsew
rlabel metal3 s 583520 272776 584800 272888 4 io_in[7]
port 627 nsew
rlabel metal3 s 583520 7454 584800 7566 4 io_in[1]
port 628 nsew
rlabel metal3 s 583520 19274 584800 19386 4 io_oeb[3]
port 629 nsew
rlabel metal3 s 583520 6272 584800 6384 4 io_in_3v3[1]
port 630 nsew
rlabel metal3 s 583520 275140 584800 275252 4 io_oeb[7]
port 631 nsew
rlabel metal3 s 583520 48096 584800 48208 4 io_in[5]
port 632 nsew
rlabel metal3 s 583520 95118 584800 95230 4 io_oeb[6]
port 633 nsew
rlabel metal3 s 583520 16910 584800 17022 4 io_in[3]
port 634 nsew
rlabel metal3 s 583520 318380 584800 318492 4 io_out[8]
port 635 nsew
rlabel metal3 s 583520 314834 584800 314946 4 gpio_noesd[1]
port 636 nsew
rlabel metal3 s 583520 12182 584800 12294 4 io_in[2]
port 637 nsew
rlabel metal3 s 583520 91572 584800 91684 4 io_in_3v3[6]
port 638 nsew
rlabel metal3 s 583520 5090 584800 5202 4 io_oeb[0]
port 639 nsew
rlabel metal3 s 583520 2726 584800 2838 4 io_in[0]
port 640 nsew
rlabel metal3 s 583520 92754 584800 92866 4 io_in[6]
port 641 nsew
rlabel metal3 s 583520 316016 584800 316128 4 io_in_3v3[8]
port 642 nsew
rlabel metal3 s 583520 13364 584800 13476 4 io_out[2]
port 643 nsew
rlabel metal3 s 583520 46914 584800 47026 4 io_in_3v3[5]
port 644 nsew
rlabel metal3 s 582340 181430 584800 186230 4 vssd1
port 645 nsew
rlabel metal3 s 583520 317198 584800 317310 4 io_in[8]
port 646 nsew
rlabel metal3 s 583520 18092 584800 18204 4 io_out[3]
port 647 nsew
rlabel metal3 s 582340 191430 584800 196230 4 vssd1
port 645 nsew
rlabel metal3 s 583520 22820 584800 22932 4 io_out[4]
port 648 nsew
rlabel metal3 s 583520 8636 584800 8748 4 io_out[1]
port 649 nsew
rlabel metal3 s 583520 273958 584800 274070 4 io_out[7]
port 650 nsew
rlabel metal3 s 583520 271594 584800 271706 4 io_in_3v3[7]
port 651 nsew
rlabel metal3 s 582340 136830 584800 141630 4 vssa1
port 517 nsew
rlabel metal3 s 583520 270412 584800 270524 4 gpio_noesd[0]
port 652 nsew
rlabel metal3 s 583520 319562 584800 319674 4 io_oeb[8]
port 653 nsew
rlabel metal3 s 583520 11000 584800 11112 4 io_in_3v3[2]
port 654 nsew
rlabel metal3 s 582340 146830 584800 151630 4 vssa1
port 517 nsew
rlabel metal3 s 583520 15728 584800 15840 4 io_in_3v3[3]
port 655 nsew
rlabel metal3 s 583520 24002 584800 24114 4 io_oeb[4]
port 656 nsew
rlabel metal3 s 582340 225230 584800 230030 4 vdda1
port 501 nsew
rlabel metal3 s 583520 269230 584800 269342 4 gpio_analog[0]
port 657 nsew
rlabel metal3 s 583520 21638 584800 21750 4 io_in[4]
port 658 nsew
rlabel metal3 s 582340 235230 584800 240030 4 vdda1
port 501 nsew
rlabel metal3 s 583520 50460 584800 50572 4 io_oeb[5]
port 659 nsew
rlabel metal3 s 583520 3908 584800 4020 4 io_out[0]
port 660 nsew
rlabel metal3 s 583520 14546 584800 14658 4 io_oeb[2]
port 661 nsew
rlabel metal3 s 583520 20456 584800 20568 4 io_in_3v3[4]
port 662 nsew
rlabel metal3 s 583520 313652 584800 313764 4 gpio_analog[1]
port 663 nsew
rlabel metal5 s 165594 702300 170594 704800 4 io_analog[6]
port 495 nsew
rlabel metal5 s 175894 702300 180894 704800 4 io_analog[6]
port 495 nsew
rlabel metal5 s 217294 702300 222294 704800 4 io_analog[5]
port 496 nsew
rlabel metal5 s 227594 702300 232594 704800 4 io_analog[5]
port 496 nsew
rlabel metal5 s 318994 702300 323994 704800 4 io_analog[4]
port 497 nsew
rlabel metal5 s 329294 702300 334294 704800 4 io_analog[4]
port 497 nsew
<< end >>
