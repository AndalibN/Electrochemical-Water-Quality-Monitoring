magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_s >>
rect 5009 13166 5015 13172
rect 5247 13166 5253 13172
rect 5003 13160 5009 13166
rect 5253 13160 5259 13166
rect 5003 12922 5009 12928
rect 5253 12922 5259 12928
rect 5009 12916 5015 12922
rect 5247 12916 5253 12922
rect -2235 -197 -2171 -196
rect -2235 -259 -2234 -197
rect -2172 -259 -2171 -197
rect -2235 -260 -2171 -259
rect 18576 -962 18626 -947
rect 18548 -990 18626 -975
<< pwell >>
rect -10861 6165 -10652 6170
rect -9402 6165 -9193 6170
rect -10867 5928 -9170 6165
rect -10861 5 -10652 5928
rect -9402 5 -9193 5928
rect -3642 5326 -3488 5356
rect -4828 5208 -3474 5326
rect -10885 -167 -9150 5
rect -10861 -191 -10652 -167
rect -9402 -191 -9193 -167
rect -4796 -392 -4686 5208
rect -3642 -392 -3488 5208
rect -4844 -510 -3450 -392
rect -4796 -526 -4686 -510
rect -3642 -550 -3488 -510
rect 12300 -772 12464 422
rect 12179 -920 12298 -902
rect 11558 -1021 12298 -920
rect 18840 -990 19220 950
rect 11576 -2722 11666 -1021
rect 12179 -2722 12283 -1021
rect 11558 -2823 12298 -2722
rect 11576 -2838 11666 -2823
rect 12179 -2832 12283 -2823
rect 10720 -5240 11544 -4534
<< psubdiff >>
rect -10835 6139 -10678 6144
rect -9376 6139 -9219 6144
rect -10841 6110 -9196 6139
rect -10841 5954 -10817 6110
rect -10835 -21 -10817 5954
rect -10859 -112 -10817 -21
rect -10715 5954 -9321 6008
rect -10715 -21 -10678 5954
rect -9376 -21 -9321 5954
rect -10715 -78 -9321 -21
rect -10715 -112 -10681 -78
rect -10647 -112 -10613 -78
rect -10579 -112 -10545 -78
rect -10511 -112 -10477 -78
rect -10443 -112 -10409 -78
rect -10375 -112 -10341 -78
rect -10307 -112 -10273 -78
rect -10239 -112 -10205 -78
rect -10171 -112 -10137 -78
rect -10103 -112 -10069 -78
rect -10035 -112 -10001 -78
rect -9967 -112 -9933 -78
rect -9899 -112 -9865 -78
rect -9831 -112 -9797 -78
rect -9763 -112 -9729 -78
rect -9695 -112 -9661 -78
rect -9627 -112 -9593 -78
rect -9559 -112 -9525 -78
rect -9491 -112 -9457 -78
rect -9423 -112 -9389 -78
rect -9355 -112 -9321 -78
rect -9219 5954 -9196 6110
rect -3616 5300 -3514 5330
rect -4802 5284 -3500 5300
rect -4802 5250 -4758 5284
rect -4724 5250 -4657 5284
rect -4623 5250 -4589 5284
rect -4555 5250 -4521 5284
rect -4487 5250 -4453 5284
rect -4419 5250 -4385 5284
rect -4351 5250 -4317 5284
rect -4283 5250 -4249 5284
rect -4215 5250 -4181 5284
rect -4147 5250 -4113 5284
rect -4079 5250 -4045 5284
rect -4011 5250 -3977 5284
rect -3943 5250 -3909 5284
rect -3875 5250 -3841 5284
rect -3807 5250 -3773 5284
rect -3739 5250 -3705 5284
rect -3671 5276 -3500 5284
rect -3671 5250 -3616 5276
rect -4802 5234 -3616 5250
rect -4770 5179 -4712 5234
rect -4770 5145 -4758 5179
rect -4724 5145 -4712 5179
rect -4770 5111 -4712 5145
rect -4770 5077 -4758 5111
rect -4724 5077 -4712 5111
rect -4770 5043 -4712 5077
rect -4770 5009 -4758 5043
rect -4724 5009 -4712 5043
rect -4770 4975 -4712 5009
rect -4770 4941 -4758 4975
rect -4724 4941 -4712 4975
rect -4770 4907 -4712 4941
rect -4770 4873 -4758 4907
rect -4724 4873 -4712 4907
rect -4770 4839 -4712 4873
rect -4770 4805 -4758 4839
rect -4724 4805 -4712 4839
rect -4770 4771 -4712 4805
rect -4770 4737 -4758 4771
rect -4724 4737 -4712 4771
rect -4770 4703 -4712 4737
rect -4770 4669 -4758 4703
rect -4724 4669 -4712 4703
rect -4770 4635 -4712 4669
rect -4770 4601 -4758 4635
rect -4724 4601 -4712 4635
rect -4770 4567 -4712 4601
rect -4770 4533 -4758 4567
rect -4724 4533 -4712 4567
rect -4770 4499 -4712 4533
rect -4770 4465 -4758 4499
rect -4724 4465 -4712 4499
rect -4770 4431 -4712 4465
rect -4770 4397 -4758 4431
rect -4724 4397 -4712 4431
rect -4770 4363 -4712 4397
rect -4770 4329 -4758 4363
rect -4724 4329 -4712 4363
rect -4770 4295 -4712 4329
rect -4770 4261 -4758 4295
rect -4724 4261 -4712 4295
rect -4770 4227 -4712 4261
rect -4770 4193 -4758 4227
rect -4724 4193 -4712 4227
rect -4770 4159 -4712 4193
rect -4770 4125 -4758 4159
rect -4724 4125 -4712 4159
rect -4770 4091 -4712 4125
rect -4770 4057 -4758 4091
rect -4724 4057 -4712 4091
rect -4770 4023 -4712 4057
rect -4770 3989 -4758 4023
rect -4724 3989 -4712 4023
rect -4770 3955 -4712 3989
rect -4770 3921 -4758 3955
rect -4724 3921 -4712 3955
rect -4770 3887 -4712 3921
rect -4770 3853 -4758 3887
rect -4724 3853 -4712 3887
rect -4770 3819 -4712 3853
rect -4770 3785 -4758 3819
rect -4724 3785 -4712 3819
rect -4770 3751 -4712 3785
rect -4770 3717 -4758 3751
rect -4724 3717 -4712 3751
rect -4770 3683 -4712 3717
rect -4770 3649 -4758 3683
rect -4724 3649 -4712 3683
rect -4770 3615 -4712 3649
rect -4770 3581 -4758 3615
rect -4724 3581 -4712 3615
rect -4770 3547 -4712 3581
rect -4770 3513 -4758 3547
rect -4724 3513 -4712 3547
rect -4770 3479 -4712 3513
rect -4770 3445 -4758 3479
rect -4724 3445 -4712 3479
rect -4770 3411 -4712 3445
rect -4770 3377 -4758 3411
rect -4724 3377 -4712 3411
rect -4770 3343 -4712 3377
rect -4770 3309 -4758 3343
rect -4724 3309 -4712 3343
rect -4770 3275 -4712 3309
rect -4770 3241 -4758 3275
rect -4724 3241 -4712 3275
rect -4770 3207 -4712 3241
rect -4770 3173 -4758 3207
rect -4724 3173 -4712 3207
rect -4770 3139 -4712 3173
rect -4770 3105 -4758 3139
rect -4724 3105 -4712 3139
rect -4770 3071 -4712 3105
rect -4770 3037 -4758 3071
rect -4724 3037 -4712 3071
rect -4770 3003 -4712 3037
rect -4770 2969 -4758 3003
rect -4724 2969 -4712 3003
rect -4770 2935 -4712 2969
rect -4770 2901 -4758 2935
rect -4724 2901 -4712 2935
rect -4770 2867 -4712 2901
rect -4770 2833 -4758 2867
rect -4724 2833 -4712 2867
rect -4770 2799 -4712 2833
rect -4770 2765 -4758 2799
rect -4724 2765 -4712 2799
rect -4770 2731 -4712 2765
rect -4770 2697 -4758 2731
rect -4724 2697 -4712 2731
rect -4770 2663 -4712 2697
rect -4770 2629 -4758 2663
rect -4724 2629 -4712 2663
rect -4770 2595 -4712 2629
rect -4770 2561 -4758 2595
rect -4724 2561 -4712 2595
rect -4770 2527 -4712 2561
rect -4770 2493 -4758 2527
rect -4724 2493 -4712 2527
rect -4770 2459 -4712 2493
rect -4770 2425 -4758 2459
rect -4724 2425 -4712 2459
rect -4770 2391 -4712 2425
rect -4770 2357 -4758 2391
rect -4724 2357 -4712 2391
rect -4770 2323 -4712 2357
rect -4770 2289 -4758 2323
rect -4724 2289 -4712 2323
rect -4770 2255 -4712 2289
rect -4770 2221 -4758 2255
rect -4724 2221 -4712 2255
rect -4770 2187 -4712 2221
rect -4770 2153 -4758 2187
rect -4724 2153 -4712 2187
rect -4770 2119 -4712 2153
rect -4770 2085 -4758 2119
rect -4724 2085 -4712 2119
rect -4770 2051 -4712 2085
rect -4770 2017 -4758 2051
rect -4724 2017 -4712 2051
rect -4770 1983 -4712 2017
rect -4770 1949 -4758 1983
rect -4724 1949 -4712 1983
rect -4770 1915 -4712 1949
rect -4770 1881 -4758 1915
rect -4724 1881 -4712 1915
rect -4770 1847 -4712 1881
rect -4770 1813 -4758 1847
rect -4724 1813 -4712 1847
rect -4770 1779 -4712 1813
rect -4770 1745 -4758 1779
rect -4724 1745 -4712 1779
rect -4770 1711 -4712 1745
rect -4770 1677 -4758 1711
rect -4724 1677 -4712 1711
rect -4770 1643 -4712 1677
rect -4770 1609 -4758 1643
rect -4724 1609 -4712 1643
rect -4770 1575 -4712 1609
rect -4770 1541 -4758 1575
rect -4724 1541 -4712 1575
rect -4770 1507 -4712 1541
rect -4770 1473 -4758 1507
rect -4724 1473 -4712 1507
rect -4770 1439 -4712 1473
rect -4770 1405 -4758 1439
rect -4724 1405 -4712 1439
rect -4770 1371 -4712 1405
rect -4770 1337 -4758 1371
rect -4724 1337 -4712 1371
rect -4770 1303 -4712 1337
rect -4770 1269 -4758 1303
rect -4724 1269 -4712 1303
rect -4770 1235 -4712 1269
rect -4770 1201 -4758 1235
rect -4724 1201 -4712 1235
rect -4770 1167 -4712 1201
rect -4770 1133 -4758 1167
rect -4724 1133 -4712 1167
rect -4770 1099 -4712 1133
rect -4770 1065 -4758 1099
rect -4724 1065 -4712 1099
rect -4770 1031 -4712 1065
rect -4770 997 -4758 1031
rect -4724 997 -4712 1031
rect -4770 963 -4712 997
rect -4770 929 -4758 963
rect -4724 929 -4712 963
rect -4770 895 -4712 929
rect -4770 861 -4758 895
rect -4724 861 -4712 895
rect -4770 827 -4712 861
rect -4770 793 -4758 827
rect -4724 793 -4712 827
rect -4770 759 -4712 793
rect -4770 725 -4758 759
rect -4724 725 -4712 759
rect -4770 691 -4712 725
rect -4770 657 -4758 691
rect -4724 657 -4712 691
rect -4770 623 -4712 657
rect -4770 589 -4758 623
rect -4724 589 -4712 623
rect -4770 555 -4712 589
rect -4770 521 -4758 555
rect -4724 521 -4712 555
rect -4770 487 -4712 521
rect -4770 453 -4758 487
rect -4724 453 -4712 487
rect -4770 419 -4712 453
rect -4770 385 -4758 419
rect -4724 385 -4712 419
rect -4770 351 -4712 385
rect -4770 317 -4758 351
rect -4724 317 -4712 351
rect -4770 283 -4712 317
rect -4770 249 -4758 283
rect -4724 249 -4712 283
rect -4770 215 -4712 249
rect -4770 181 -4758 215
rect -4724 181 -4712 215
rect -4770 147 -4712 181
rect -4770 113 -4758 147
rect -4724 113 -4712 147
rect -4770 79 -4712 113
rect -4770 45 -4758 79
rect -4724 45 -4712 79
rect -4770 11 -4712 45
rect -9219 -112 -9176 -21
rect -10859 -141 -9176 -112
rect -4770 -23 -4758 11
rect -4724 -23 -4712 11
rect -4770 -57 -4712 -23
rect -4770 -91 -4758 -57
rect -4724 -91 -4712 -57
rect -4770 -125 -4712 -91
rect -10835 -165 -10678 -141
rect -9376 -165 -9219 -141
rect -4770 -159 -4758 -125
rect -4724 -159 -4712 -125
rect -4770 -193 -4712 -159
rect -4770 -227 -4758 -193
rect -4724 -227 -4712 -193
rect -4770 -261 -4712 -227
rect -4770 -295 -4758 -261
rect -4724 -295 -4712 -261
rect -4770 -329 -4712 -295
rect -4770 -363 -4758 -329
rect -4724 -363 -4712 -329
rect -4770 -418 -4712 -363
rect -4818 -434 -3616 -418
rect -4818 -468 -4758 -434
rect -4724 -468 -4657 -434
rect -4623 -468 -4589 -434
rect -4555 -468 -4521 -434
rect -4487 -468 -4453 -434
rect -4419 -468 -4385 -434
rect -4351 -468 -4317 -434
rect -4283 -468 -4249 -434
rect -4215 -468 -4181 -434
rect -4147 -468 -4113 -434
rect -4079 -468 -4045 -434
rect -4011 -468 -3977 -434
rect -3943 -468 -3909 -434
rect -3875 -468 -3841 -434
rect -3807 -468 -3773 -434
rect -3739 -468 -3705 -434
rect -3671 -468 -3616 -434
rect -4818 -470 -3616 -468
rect -3514 5234 -3500 5276
rect 18866 881 19194 924
rect 12326 352 12438 396
rect -3514 -470 -3476 -418
rect -4818 -484 -3476 -470
rect -4770 -500 -4712 -484
rect -3616 -524 -3514 -484
rect 12326 -702 12331 352
rect 12433 -702 12438 352
rect 12326 -746 12438 -702
rect 18866 -921 18877 881
rect 19183 -921 19194 881
rect 12205 -946 12257 -928
rect 11584 -954 12272 -946
rect 11584 -988 11674 -954
rect 11708 -988 11742 -954
rect 11776 -988 11810 -954
rect 11844 -988 11878 -954
rect 11912 -988 11946 -954
rect 11980 -988 12014 -954
rect 12048 -988 12082 -954
rect 12116 -988 12150 -954
rect 12184 -988 12218 -954
rect 12252 -988 12272 -954
rect 18866 -964 19194 -921
rect 11584 -995 12272 -988
rect 11602 -1039 11640 -995
rect 11602 -1073 11604 -1039
rect 11638 -1073 11640 -1039
rect 11602 -1107 11640 -1073
rect 11602 -1141 11604 -1107
rect 11638 -1141 11640 -1107
rect 11602 -1175 11640 -1141
rect 11602 -1209 11604 -1175
rect 11638 -1209 11640 -1175
rect 11602 -1243 11640 -1209
rect 11602 -1277 11604 -1243
rect 11638 -1277 11640 -1243
rect 11602 -1311 11640 -1277
rect 11602 -1345 11604 -1311
rect 11638 -1345 11640 -1311
rect 11602 -1379 11640 -1345
rect 11602 -1413 11604 -1379
rect 11638 -1413 11640 -1379
rect 11602 -1447 11640 -1413
rect 11602 -1481 11604 -1447
rect 11638 -1481 11640 -1447
rect 11602 -1515 11640 -1481
rect 11602 -1549 11604 -1515
rect 11638 -1549 11640 -1515
rect 11602 -1583 11640 -1549
rect 11602 -1617 11604 -1583
rect 11638 -1617 11640 -1583
rect 11602 -1651 11640 -1617
rect 11602 -1685 11604 -1651
rect 11638 -1685 11640 -1651
rect 11602 -1719 11640 -1685
rect 11602 -1753 11604 -1719
rect 11638 -1753 11640 -1719
rect 11602 -1787 11640 -1753
rect 11602 -1821 11604 -1787
rect 11638 -1821 11640 -1787
rect 11602 -1855 11640 -1821
rect 11602 -1889 11604 -1855
rect 11638 -1889 11640 -1855
rect 11602 -1923 11640 -1889
rect 11602 -1957 11604 -1923
rect 11638 -1957 11640 -1923
rect 11602 -1991 11640 -1957
rect 11602 -2025 11604 -1991
rect 11638 -2025 11640 -1991
rect 11602 -2059 11640 -2025
rect 11602 -2093 11604 -2059
rect 11638 -2093 11640 -2059
rect 11602 -2127 11640 -2093
rect 11602 -2161 11604 -2127
rect 11638 -2161 11640 -2127
rect 11602 -2195 11640 -2161
rect 11602 -2229 11604 -2195
rect 11638 -2229 11640 -2195
rect 11602 -2263 11640 -2229
rect 11602 -2297 11604 -2263
rect 11638 -2297 11640 -2263
rect 11602 -2331 11640 -2297
rect 11602 -2365 11604 -2331
rect 11638 -2365 11640 -2331
rect 11602 -2399 11640 -2365
rect 11602 -2433 11604 -2399
rect 11638 -2433 11640 -2399
rect 11602 -2467 11640 -2433
rect 11602 -2501 11604 -2467
rect 11638 -2501 11640 -2467
rect 11602 -2535 11640 -2501
rect 11602 -2569 11604 -2535
rect 11638 -2569 11640 -2535
rect 11602 -2603 11640 -2569
rect 11602 -2637 11604 -2603
rect 11638 -2637 11640 -2603
rect 11602 -2671 11640 -2637
rect 11602 -2705 11604 -2671
rect 11638 -2705 11640 -2671
rect 11602 -2748 11640 -2705
rect 12205 -1039 12257 -995
rect 12205 -1073 12214 -1039
rect 12248 -1073 12257 -1039
rect 12205 -1107 12257 -1073
rect 12205 -1141 12214 -1107
rect 12248 -1141 12257 -1107
rect 12205 -1175 12257 -1141
rect 12205 -1209 12214 -1175
rect 12248 -1209 12257 -1175
rect 12205 -1243 12257 -1209
rect 12205 -1277 12214 -1243
rect 12248 -1277 12257 -1243
rect 12205 -1311 12257 -1277
rect 12205 -1345 12214 -1311
rect 12248 -1345 12257 -1311
rect 12205 -1379 12257 -1345
rect 12205 -1413 12214 -1379
rect 12248 -1413 12257 -1379
rect 12205 -1447 12257 -1413
rect 12205 -1481 12214 -1447
rect 12248 -1481 12257 -1447
rect 12205 -1515 12257 -1481
rect 12205 -1549 12214 -1515
rect 12248 -1549 12257 -1515
rect 12205 -1583 12257 -1549
rect 12205 -1617 12214 -1583
rect 12248 -1617 12257 -1583
rect 12205 -1651 12257 -1617
rect 12205 -1685 12214 -1651
rect 12248 -1685 12257 -1651
rect 12205 -1719 12257 -1685
rect 12205 -1753 12214 -1719
rect 12248 -1753 12257 -1719
rect 12205 -1787 12257 -1753
rect 12205 -1821 12214 -1787
rect 12248 -1821 12257 -1787
rect 12205 -1855 12257 -1821
rect 12205 -1889 12214 -1855
rect 12248 -1889 12257 -1855
rect 12205 -1923 12257 -1889
rect 12205 -1957 12214 -1923
rect 12248 -1957 12257 -1923
rect 12205 -1991 12257 -1957
rect 12205 -2025 12214 -1991
rect 12248 -2025 12257 -1991
rect 12205 -2059 12257 -2025
rect 12205 -2093 12214 -2059
rect 12248 -2093 12257 -2059
rect 12205 -2127 12257 -2093
rect 12205 -2161 12214 -2127
rect 12248 -2161 12257 -2127
rect 12205 -2195 12257 -2161
rect 12205 -2229 12214 -2195
rect 12248 -2229 12257 -2195
rect 12205 -2263 12257 -2229
rect 12205 -2297 12214 -2263
rect 12248 -2297 12257 -2263
rect 12205 -2331 12257 -2297
rect 12205 -2365 12214 -2331
rect 12248 -2365 12257 -2331
rect 12205 -2399 12257 -2365
rect 12205 -2433 12214 -2399
rect 12248 -2433 12257 -2399
rect 12205 -2467 12257 -2433
rect 12205 -2501 12214 -2467
rect 12248 -2501 12257 -2467
rect 12205 -2535 12257 -2501
rect 12205 -2569 12214 -2535
rect 12248 -2569 12257 -2535
rect 12205 -2603 12257 -2569
rect 12205 -2637 12214 -2603
rect 12248 -2637 12257 -2603
rect 12205 -2671 12257 -2637
rect 12205 -2705 12214 -2671
rect 12248 -2705 12257 -2671
rect 12205 -2748 12257 -2705
rect 11584 -2756 12272 -2748
rect 11584 -2790 11674 -2756
rect 11708 -2790 11742 -2756
rect 11776 -2790 11810 -2756
rect 11844 -2790 11878 -2756
rect 11912 -2790 11946 -2756
rect 11980 -2790 12014 -2756
rect 12048 -2790 12082 -2756
rect 12116 -2790 12150 -2756
rect 12184 -2790 12272 -2756
rect 11584 -2797 12272 -2790
rect 11602 -2812 11640 -2797
rect 12205 -2806 12257 -2797
rect 10746 -4564 11518 -4560
rect 10746 -5210 10775 -4564
rect 11489 -5210 11518 -4564
rect 10746 -5214 11518 -5210
<< psubdiffcont >>
rect -10817 6008 -9219 6110
rect -10817 -112 -10715 6008
rect -10681 -112 -10647 -78
rect -10613 -112 -10579 -78
rect -10545 -112 -10511 -78
rect -10477 -112 -10443 -78
rect -10409 -112 -10375 -78
rect -10341 -112 -10307 -78
rect -10273 -112 -10239 -78
rect -10205 -112 -10171 -78
rect -10137 -112 -10103 -78
rect -10069 -112 -10035 -78
rect -10001 -112 -9967 -78
rect -9933 -112 -9899 -78
rect -9865 -112 -9831 -78
rect -9797 -112 -9763 -78
rect -9729 -112 -9695 -78
rect -9661 -112 -9627 -78
rect -9593 -112 -9559 -78
rect -9525 -112 -9491 -78
rect -9457 -112 -9423 -78
rect -9389 -112 -9355 -78
rect -9321 -112 -9219 6008
rect -4758 5250 -4724 5284
rect -4657 5250 -4623 5284
rect -4589 5250 -4555 5284
rect -4521 5250 -4487 5284
rect -4453 5250 -4419 5284
rect -4385 5250 -4351 5284
rect -4317 5250 -4283 5284
rect -4249 5250 -4215 5284
rect -4181 5250 -4147 5284
rect -4113 5250 -4079 5284
rect -4045 5250 -4011 5284
rect -3977 5250 -3943 5284
rect -3909 5250 -3875 5284
rect -3841 5250 -3807 5284
rect -3773 5250 -3739 5284
rect -3705 5250 -3671 5284
rect -4758 5145 -4724 5179
rect -4758 5077 -4724 5111
rect -4758 5009 -4724 5043
rect -4758 4941 -4724 4975
rect -4758 4873 -4724 4907
rect -4758 4805 -4724 4839
rect -4758 4737 -4724 4771
rect -4758 4669 -4724 4703
rect -4758 4601 -4724 4635
rect -4758 4533 -4724 4567
rect -4758 4465 -4724 4499
rect -4758 4397 -4724 4431
rect -4758 4329 -4724 4363
rect -4758 4261 -4724 4295
rect -4758 4193 -4724 4227
rect -4758 4125 -4724 4159
rect -4758 4057 -4724 4091
rect -4758 3989 -4724 4023
rect -4758 3921 -4724 3955
rect -4758 3853 -4724 3887
rect -4758 3785 -4724 3819
rect -4758 3717 -4724 3751
rect -4758 3649 -4724 3683
rect -4758 3581 -4724 3615
rect -4758 3513 -4724 3547
rect -4758 3445 -4724 3479
rect -4758 3377 -4724 3411
rect -4758 3309 -4724 3343
rect -4758 3241 -4724 3275
rect -4758 3173 -4724 3207
rect -4758 3105 -4724 3139
rect -4758 3037 -4724 3071
rect -4758 2969 -4724 3003
rect -4758 2901 -4724 2935
rect -4758 2833 -4724 2867
rect -4758 2765 -4724 2799
rect -4758 2697 -4724 2731
rect -4758 2629 -4724 2663
rect -4758 2561 -4724 2595
rect -4758 2493 -4724 2527
rect -4758 2425 -4724 2459
rect -4758 2357 -4724 2391
rect -4758 2289 -4724 2323
rect -4758 2221 -4724 2255
rect -4758 2153 -4724 2187
rect -4758 2085 -4724 2119
rect -4758 2017 -4724 2051
rect -4758 1949 -4724 1983
rect -4758 1881 -4724 1915
rect -4758 1813 -4724 1847
rect -4758 1745 -4724 1779
rect -4758 1677 -4724 1711
rect -4758 1609 -4724 1643
rect -4758 1541 -4724 1575
rect -4758 1473 -4724 1507
rect -4758 1405 -4724 1439
rect -4758 1337 -4724 1371
rect -4758 1269 -4724 1303
rect -4758 1201 -4724 1235
rect -4758 1133 -4724 1167
rect -4758 1065 -4724 1099
rect -4758 997 -4724 1031
rect -4758 929 -4724 963
rect -4758 861 -4724 895
rect -4758 793 -4724 827
rect -4758 725 -4724 759
rect -4758 657 -4724 691
rect -4758 589 -4724 623
rect -4758 521 -4724 555
rect -4758 453 -4724 487
rect -4758 385 -4724 419
rect -4758 317 -4724 351
rect -4758 249 -4724 283
rect -4758 181 -4724 215
rect -4758 113 -4724 147
rect -4758 45 -4724 79
rect -4758 -23 -4724 11
rect -4758 -91 -4724 -57
rect -4758 -159 -4724 -125
rect -4758 -227 -4724 -193
rect -4758 -295 -4724 -261
rect -4758 -363 -4724 -329
rect -4758 -468 -4724 -434
rect -4657 -468 -4623 -434
rect -4589 -468 -4555 -434
rect -4521 -468 -4487 -434
rect -4453 -468 -4419 -434
rect -4385 -468 -4351 -434
rect -4317 -468 -4283 -434
rect -4249 -468 -4215 -434
rect -4181 -468 -4147 -434
rect -4113 -468 -4079 -434
rect -4045 -468 -4011 -434
rect -3977 -468 -3943 -434
rect -3909 -468 -3875 -434
rect -3841 -468 -3807 -434
rect -3773 -468 -3739 -434
rect -3705 -468 -3671 -434
rect -3616 -470 -3514 5276
rect 12331 -702 12433 352
rect 18877 -921 19183 881
rect 11674 -988 11708 -954
rect 11742 -988 11776 -954
rect 11810 -988 11844 -954
rect 11878 -988 11912 -954
rect 11946 -988 11980 -954
rect 12014 -988 12048 -954
rect 12082 -988 12116 -954
rect 12150 -988 12184 -954
rect 12218 -988 12252 -954
rect 11604 -1073 11638 -1039
rect 11604 -1141 11638 -1107
rect 11604 -1209 11638 -1175
rect 11604 -1277 11638 -1243
rect 11604 -1345 11638 -1311
rect 11604 -1413 11638 -1379
rect 11604 -1481 11638 -1447
rect 11604 -1549 11638 -1515
rect 11604 -1617 11638 -1583
rect 11604 -1685 11638 -1651
rect 11604 -1753 11638 -1719
rect 11604 -1821 11638 -1787
rect 11604 -1889 11638 -1855
rect 11604 -1957 11638 -1923
rect 11604 -2025 11638 -1991
rect 11604 -2093 11638 -2059
rect 11604 -2161 11638 -2127
rect 11604 -2229 11638 -2195
rect 11604 -2297 11638 -2263
rect 11604 -2365 11638 -2331
rect 11604 -2433 11638 -2399
rect 11604 -2501 11638 -2467
rect 11604 -2569 11638 -2535
rect 11604 -2637 11638 -2603
rect 11604 -2705 11638 -2671
rect 12214 -1073 12248 -1039
rect 12214 -1141 12248 -1107
rect 12214 -1209 12248 -1175
rect 12214 -1277 12248 -1243
rect 12214 -1345 12248 -1311
rect 12214 -1413 12248 -1379
rect 12214 -1481 12248 -1447
rect 12214 -1549 12248 -1515
rect 12214 -1617 12248 -1583
rect 12214 -1685 12248 -1651
rect 12214 -1753 12248 -1719
rect 12214 -1821 12248 -1787
rect 12214 -1889 12248 -1855
rect 12214 -1957 12248 -1923
rect 12214 -2025 12248 -1991
rect 12214 -2093 12248 -2059
rect 12214 -2161 12248 -2127
rect 12214 -2229 12248 -2195
rect 12214 -2297 12248 -2263
rect 12214 -2365 12248 -2331
rect 12214 -2433 12248 -2399
rect 12214 -2501 12248 -2467
rect 12214 -2569 12248 -2535
rect 12214 -2637 12248 -2603
rect 12214 -2705 12248 -2671
rect 11674 -2790 11708 -2756
rect 11742 -2790 11776 -2756
rect 11810 -2790 11844 -2756
rect 11878 -2790 11912 -2756
rect 11946 -2790 11980 -2756
rect 12014 -2790 12048 -2756
rect 12082 -2790 12116 -2756
rect 12150 -2790 12184 -2756
rect 10775 -5210 11489 -4564
<< locali >>
rect -10833 6136 -9204 6139
rect -10835 6110 -9204 6136
rect -10835 -21 -10817 6110
rect -10851 -112 -10817 -21
rect -10715 5954 -9321 6008
rect -10715 -21 -10678 5954
rect -9376 5240 -9321 5954
rect -9380 5178 -9321 5240
rect -10128 352 -10094 668
rect -9900 382 -9866 676
rect -9901 352 -9866 382
rect -10129 348 -9866 352
rect -10129 306 -9867 348
rect -9376 -21 -9321 5178
rect -10715 -78 -9321 -21
rect -10715 -112 -10681 -78
rect -10647 -112 -10613 -78
rect -10579 -112 -10545 -78
rect -10511 -112 -10477 -78
rect -10443 -112 -10409 -78
rect -10375 -112 -10341 -78
rect -10307 -112 -10273 -78
rect -10239 -112 -10205 -78
rect -10171 -112 -10137 -78
rect -10103 -112 -10069 -78
rect -10035 -112 -10001 -78
rect -9967 -112 -9933 -78
rect -9899 -112 -9865 -78
rect -9831 -112 -9797 -78
rect -9763 -112 -9729 -78
rect -9695 -112 -9661 -78
rect -9627 -112 -9593 -78
rect -9559 -112 -9525 -78
rect -9491 -112 -9457 -78
rect -9423 -112 -9389 -78
rect -9355 -112 -9321 -78
rect -9219 5954 -9204 6110
rect -3616 5300 -3514 5322
rect -4794 5284 -3508 5300
rect -4794 5250 -4758 5284
rect -4724 5250 -4657 5284
rect -4623 5250 -4589 5284
rect -4555 5250 -4521 5284
rect -4487 5250 -4453 5284
rect -4419 5250 -4385 5284
rect -4351 5250 -4317 5284
rect -4283 5250 -4249 5284
rect -4215 5250 -4181 5284
rect -4147 5250 -4113 5284
rect -4079 5250 -4045 5284
rect -4011 5250 -3977 5284
rect -3943 5250 -3909 5284
rect -3875 5250 -3841 5284
rect -3807 5250 -3773 5284
rect -3739 5250 -3705 5284
rect -3671 5276 -3508 5284
rect -3671 5250 -3616 5276
rect -4794 5240 -3616 5250
rect -9219 5234 -3616 5240
rect -9219 5179 -4712 5234
rect -9219 5178 -4758 5179
rect -4770 5145 -4758 5178
rect -4724 5145 -4712 5179
rect -4770 5111 -4712 5145
rect -4770 5077 -4758 5111
rect -4724 5077 -4712 5111
rect -4770 5043 -4712 5077
rect -4770 5009 -4758 5043
rect -4724 5009 -4712 5043
rect -4770 4975 -4712 5009
rect -4770 4941 -4758 4975
rect -4724 4941 -4712 4975
rect -4770 4907 -4712 4941
rect -4770 4873 -4758 4907
rect -4724 4873 -4712 4907
rect -4770 4839 -4712 4873
rect -4770 4805 -4758 4839
rect -4724 4805 -4712 4839
rect -4770 4771 -4712 4805
rect -4770 4737 -4758 4771
rect -4724 4737 -4712 4771
rect -4770 4703 -4712 4737
rect -4770 4669 -4758 4703
rect -4724 4669 -4712 4703
rect -4770 4635 -4712 4669
rect -4770 4601 -4758 4635
rect -4724 4601 -4712 4635
rect -4770 4567 -4712 4601
rect -4770 4533 -4758 4567
rect -4724 4533 -4712 4567
rect -4770 4499 -4712 4533
rect -4770 4465 -4758 4499
rect -4724 4465 -4712 4499
rect -4770 4431 -4712 4465
rect -4770 4397 -4758 4431
rect -4724 4397 -4712 4431
rect -4770 4363 -4712 4397
rect -4770 4329 -4758 4363
rect -4724 4329 -4712 4363
rect -4770 4295 -4712 4329
rect -4770 4261 -4758 4295
rect -4724 4261 -4712 4295
rect -4770 4227 -4712 4261
rect -4770 4193 -4758 4227
rect -4724 4193 -4712 4227
rect -4770 4159 -4712 4193
rect -4770 4125 -4758 4159
rect -4724 4125 -4712 4159
rect -4770 4091 -4712 4125
rect -4770 4057 -4758 4091
rect -4724 4057 -4712 4091
rect -4770 4023 -4712 4057
rect -4770 3989 -4758 4023
rect -4724 3989 -4712 4023
rect -4770 3955 -4712 3989
rect -4770 3921 -4758 3955
rect -4724 3921 -4712 3955
rect -4770 3887 -4712 3921
rect -4770 3853 -4758 3887
rect -4724 3853 -4712 3887
rect -4770 3819 -4712 3853
rect -4770 3785 -4758 3819
rect -4724 3785 -4712 3819
rect -4770 3751 -4712 3785
rect -4770 3717 -4758 3751
rect -4724 3717 -4712 3751
rect -4770 3683 -4712 3717
rect -4770 3649 -4758 3683
rect -4724 3649 -4712 3683
rect -4770 3615 -4712 3649
rect -4770 3581 -4758 3615
rect -4724 3581 -4712 3615
rect -4770 3547 -4712 3581
rect -4770 3513 -4758 3547
rect -4724 3513 -4712 3547
rect -4770 3479 -4712 3513
rect -4770 3445 -4758 3479
rect -4724 3445 -4712 3479
rect -4770 3411 -4712 3445
rect -4770 3377 -4758 3411
rect -4724 3377 -4712 3411
rect -4770 3343 -4712 3377
rect -4770 3309 -4758 3343
rect -4724 3309 -4712 3343
rect -4770 3275 -4712 3309
rect -4770 3241 -4758 3275
rect -4724 3241 -4712 3275
rect -4770 3207 -4712 3241
rect -4770 3173 -4758 3207
rect -4724 3173 -4712 3207
rect -4770 3139 -4712 3173
rect -4770 3105 -4758 3139
rect -4724 3105 -4712 3139
rect -4770 3071 -4712 3105
rect -4770 3037 -4758 3071
rect -4724 3037 -4712 3071
rect -4770 3003 -4712 3037
rect -4770 2969 -4758 3003
rect -4724 2969 -4712 3003
rect -4770 2935 -4712 2969
rect -4770 2901 -4758 2935
rect -4724 2901 -4712 2935
rect -4770 2867 -4712 2901
rect -4770 2833 -4758 2867
rect -4724 2833 -4712 2867
rect -4770 2799 -4712 2833
rect -4770 2765 -4758 2799
rect -4724 2765 -4712 2799
rect -4770 2731 -4712 2765
rect -4770 2697 -4758 2731
rect -4724 2697 -4712 2731
rect -4770 2663 -4712 2697
rect -4770 2629 -4758 2663
rect -4724 2629 -4712 2663
rect -4770 2595 -4712 2629
rect -4770 2561 -4758 2595
rect -4724 2561 -4712 2595
rect -4770 2527 -4712 2561
rect -4770 2493 -4758 2527
rect -4724 2493 -4712 2527
rect -4770 2459 -4712 2493
rect -4770 2425 -4758 2459
rect -4724 2425 -4712 2459
rect -4770 2391 -4712 2425
rect -4770 2357 -4758 2391
rect -4724 2357 -4712 2391
rect -4770 2323 -4712 2357
rect -4770 2289 -4758 2323
rect -4724 2289 -4712 2323
rect -4770 2255 -4712 2289
rect -4770 2221 -4758 2255
rect -4724 2221 -4712 2255
rect -4770 2187 -4712 2221
rect -4770 2153 -4758 2187
rect -4724 2153 -4712 2187
rect -4770 2119 -4712 2153
rect -4770 2085 -4758 2119
rect -4724 2085 -4712 2119
rect -4770 2051 -4712 2085
rect -4770 2017 -4758 2051
rect -4724 2017 -4712 2051
rect -4770 1983 -4712 2017
rect -4770 1949 -4758 1983
rect -4724 1949 -4712 1983
rect -4770 1915 -4712 1949
rect -4770 1881 -4758 1915
rect -4724 1881 -4712 1915
rect -4770 1847 -4712 1881
rect -4770 1813 -4758 1847
rect -4724 1813 -4712 1847
rect -4770 1779 -4712 1813
rect -4770 1745 -4758 1779
rect -4724 1745 -4712 1779
rect -4770 1711 -4712 1745
rect -4770 1677 -4758 1711
rect -4724 1677 -4712 1711
rect -4770 1643 -4712 1677
rect -4770 1609 -4758 1643
rect -4724 1609 -4712 1643
rect -4770 1575 -4712 1609
rect -4770 1541 -4758 1575
rect -4724 1541 -4712 1575
rect -4770 1507 -4712 1541
rect -4770 1473 -4758 1507
rect -4724 1473 -4712 1507
rect -4770 1439 -4712 1473
rect -4770 1405 -4758 1439
rect -4724 1405 -4712 1439
rect -4770 1371 -4712 1405
rect -4770 1337 -4758 1371
rect -4724 1337 -4712 1371
rect -4770 1303 -4712 1337
rect -4770 1269 -4758 1303
rect -4724 1269 -4712 1303
rect -4770 1235 -4712 1269
rect -4770 1201 -4758 1235
rect -4724 1201 -4712 1235
rect -4770 1167 -4712 1201
rect -4770 1133 -4758 1167
rect -4724 1133 -4712 1167
rect -4770 1099 -4712 1133
rect -4770 1065 -4758 1099
rect -4724 1065 -4712 1099
rect -4770 1031 -4712 1065
rect -4770 997 -4758 1031
rect -4724 997 -4712 1031
rect -4770 963 -4712 997
rect -4770 929 -4758 963
rect -4724 929 -4712 963
rect -4770 895 -4712 929
rect -4770 861 -4758 895
rect -4724 861 -4712 895
rect -4770 827 -4712 861
rect -4770 793 -4758 827
rect -4724 793 -4712 827
rect -4770 759 -4712 793
rect -4770 725 -4758 759
rect -4724 725 -4712 759
rect -4770 691 -4712 725
rect -4770 657 -4758 691
rect -4724 657 -4712 691
rect -4770 623 -4712 657
rect -4770 589 -4758 623
rect -4724 589 -4712 623
rect -4770 555 -4712 589
rect -4770 521 -4758 555
rect -4724 521 -4712 555
rect -4770 487 -4712 521
rect -4770 453 -4758 487
rect -4724 453 -4712 487
rect -4770 419 -4712 453
rect -4770 385 -4758 419
rect -4724 385 -4712 419
rect -4770 351 -4712 385
rect -4770 317 -4758 351
rect -4724 317 -4712 351
rect -4770 283 -4712 317
rect -4770 249 -4758 283
rect -4724 249 -4712 283
rect -4770 215 -4712 249
rect -4770 181 -4758 215
rect -4724 181 -4712 215
rect -4770 147 -4712 181
rect -4770 113 -4758 147
rect -4724 113 -4712 147
rect -4770 79 -4712 113
rect -4770 45 -4758 79
rect -4724 45 -4712 79
rect -4770 11 -4712 45
rect -9219 -112 -9184 -21
rect -10851 -141 -9184 -112
rect -4770 -23 -4758 11
rect -4724 -23 -4712 11
rect -4770 -57 -4712 -23
rect -4770 -91 -4758 -57
rect -4724 -91 -4712 -57
rect -4770 -125 -4712 -91
rect -10835 -157 -10678 -141
rect -9376 -157 -9219 -141
rect -4770 -159 -4758 -125
rect -4724 -159 -4712 -125
rect -4770 -193 -4712 -159
rect -4770 -227 -4758 -193
rect -4724 -227 -4712 -193
rect -4770 -261 -4712 -227
rect -4770 -295 -4758 -261
rect -4724 -295 -4712 -261
rect -4770 -329 -4712 -295
rect -4770 -363 -4758 -329
rect -4724 -363 -4712 -329
rect -4770 -418 -4712 -363
rect -4286 -326 -4252 -88
rect -4058 -326 -4024 -80
rect -4286 -364 -4024 -326
rect -4810 -434 -3616 -418
rect -4810 -468 -4758 -434
rect -4724 -468 -4657 -434
rect -4623 -468 -4589 -434
rect -4555 -468 -4521 -434
rect -4487 -468 -4453 -434
rect -4419 -468 -4385 -434
rect -4351 -468 -4317 -434
rect -4283 -468 -4249 -434
rect -4215 -468 -4181 -434
rect -4147 -468 -4113 -434
rect -4079 -468 -4045 -434
rect -4011 -468 -3977 -434
rect -3943 -468 -3909 -434
rect -3875 -468 -3841 -434
rect -3807 -468 -3773 -434
rect -3739 -468 -3705 -434
rect -3671 -468 -3616 -434
rect -4810 -470 -3616 -468
rect -3514 5234 -3508 5276
rect 4920 5196 5102 5197
rect -3514 5074 5102 5196
rect -3514 -470 -3484 -418
rect -4810 -484 -3484 -470
rect -4770 -492 -4712 -484
rect -3616 -516 -3514 -484
rect 2318 -4938 2814 5074
rect 4920 -1358 5102 5074
rect 12366 1476 12436 1485
rect 16600 1476 16646 1546
rect 12366 1444 16646 1476
rect 12366 1386 25368 1444
rect 10890 780 10944 792
rect 12366 780 12436 1386
rect 16598 1228 25368 1386
rect 16600 1168 16646 1228
rect 19008 916 19052 1228
rect 10890 716 12436 780
rect 10890 -1358 10944 716
rect 12366 388 12436 716
rect 18866 881 19194 916
rect 12326 352 12438 388
rect 12326 -702 12331 352
rect 12433 -702 12438 352
rect 12326 -738 12438 -702
rect 18866 -921 18877 881
rect 19183 -921 19194 881
rect 12205 -946 12257 -936
rect 11592 -954 12264 -946
rect 11592 -988 11674 -954
rect 11708 -988 11742 -954
rect 11776 -988 11810 -954
rect 11844 -988 11878 -954
rect 11912 -988 11946 -954
rect 11980 -988 12014 -954
rect 12048 -988 12082 -954
rect 12116 -988 12150 -954
rect 12184 -988 12218 -954
rect 12252 -988 12264 -954
rect 18866 -956 19194 -921
rect 11592 -995 12264 -988
rect 11602 -1039 11640 -995
rect 11602 -1073 11604 -1039
rect 11638 -1073 11640 -1039
rect 11602 -1107 11640 -1073
rect 11602 -1141 11604 -1107
rect 11638 -1141 11640 -1107
rect 11602 -1175 11640 -1141
rect 11602 -1209 11604 -1175
rect 11638 -1209 11640 -1175
rect 11602 -1243 11640 -1209
rect 11602 -1277 11604 -1243
rect 11638 -1277 11640 -1243
rect 11602 -1311 11640 -1277
rect 11602 -1345 11604 -1311
rect 11638 -1345 11640 -1311
rect 11602 -1350 11640 -1345
rect 11562 -1358 11640 -1350
rect 4920 -1379 11640 -1358
rect 4920 -1413 11604 -1379
rect 11638 -1413 11640 -1379
rect 4920 -1447 11640 -1413
rect 4920 -1460 11604 -1447
rect 11562 -1466 11604 -1460
rect 11602 -1481 11604 -1466
rect 11638 -1481 11640 -1447
rect 11602 -1515 11640 -1481
rect 11602 -1549 11604 -1515
rect 11638 -1549 11640 -1515
rect 11602 -1583 11640 -1549
rect 11602 -1617 11604 -1583
rect 11638 -1617 11640 -1583
rect 11602 -1651 11640 -1617
rect 11602 -1685 11604 -1651
rect 11638 -1685 11640 -1651
rect 11602 -1719 11640 -1685
rect 11602 -1753 11604 -1719
rect 11638 -1753 11640 -1719
rect 11602 -1787 11640 -1753
rect 11602 -1821 11604 -1787
rect 11638 -1821 11640 -1787
rect 11602 -1855 11640 -1821
rect 11602 -1889 11604 -1855
rect 11638 -1889 11640 -1855
rect 11602 -1923 11640 -1889
rect 11602 -1957 11604 -1923
rect 11638 -1957 11640 -1923
rect 11602 -1991 11640 -1957
rect 11602 -2025 11604 -1991
rect 11638 -2025 11640 -1991
rect 11602 -2059 11640 -2025
rect 11602 -2093 11604 -2059
rect 11638 -2093 11640 -2059
rect 11602 -2127 11640 -2093
rect 11602 -2161 11604 -2127
rect 11638 -2161 11640 -2127
rect 11602 -2195 11640 -2161
rect 11602 -2229 11604 -2195
rect 11638 -2229 11640 -2195
rect 11602 -2263 11640 -2229
rect 11602 -2297 11604 -2263
rect 11638 -2297 11640 -2263
rect 11602 -2331 11640 -2297
rect 11602 -2365 11604 -2331
rect 11638 -2365 11640 -2331
rect 11602 -2399 11640 -2365
rect 11602 -2433 11604 -2399
rect 11638 -2433 11640 -2399
rect 11602 -2467 11640 -2433
rect 11602 -2501 11604 -2467
rect 11638 -2501 11640 -2467
rect 11602 -2535 11640 -2501
rect 11602 -2569 11604 -2535
rect 11638 -2569 11640 -2535
rect 11602 -2603 11640 -2569
rect 11602 -2637 11604 -2603
rect 11638 -2637 11640 -2603
rect 11602 -2671 11640 -2637
rect 11602 -2705 11604 -2671
rect 11638 -2705 11640 -2671
rect 11602 -2748 11640 -2705
rect 12205 -1039 12257 -995
rect 12205 -1073 12214 -1039
rect 12248 -1073 12257 -1039
rect 12205 -1107 12257 -1073
rect 12205 -1141 12214 -1107
rect 12248 -1141 12257 -1107
rect 12205 -1175 12257 -1141
rect 12205 -1209 12214 -1175
rect 12248 -1209 12257 -1175
rect 12205 -1243 12257 -1209
rect 12205 -1277 12214 -1243
rect 12248 -1277 12257 -1243
rect 12205 -1311 12257 -1277
rect 12205 -1345 12214 -1311
rect 12248 -1345 12257 -1311
rect 12205 -1379 12257 -1345
rect 12205 -1413 12214 -1379
rect 12248 -1413 12257 -1379
rect 12205 -1447 12257 -1413
rect 12205 -1481 12214 -1447
rect 12248 -1481 12257 -1447
rect 12205 -1515 12257 -1481
rect 12205 -1549 12214 -1515
rect 12248 -1549 12257 -1515
rect 12205 -1583 12257 -1549
rect 12205 -1617 12214 -1583
rect 12248 -1617 12257 -1583
rect 12205 -1651 12257 -1617
rect 12205 -1685 12214 -1651
rect 12248 -1685 12257 -1651
rect 12205 -1719 12257 -1685
rect 12205 -1753 12214 -1719
rect 12248 -1753 12257 -1719
rect 12205 -1787 12257 -1753
rect 12205 -1821 12214 -1787
rect 12248 -1821 12257 -1787
rect 12205 -1855 12257 -1821
rect 12205 -1889 12214 -1855
rect 12248 -1889 12257 -1855
rect 12205 -1923 12257 -1889
rect 12205 -1957 12214 -1923
rect 12248 -1957 12257 -1923
rect 12205 -1991 12257 -1957
rect 12205 -2025 12214 -1991
rect 12248 -2025 12257 -1991
rect 12205 -2059 12257 -2025
rect 12205 -2093 12214 -2059
rect 12248 -2093 12257 -2059
rect 12205 -2127 12257 -2093
rect 12205 -2161 12214 -2127
rect 12248 -2161 12257 -2127
rect 12205 -2195 12257 -2161
rect 12205 -2229 12214 -2195
rect 12248 -2229 12257 -2195
rect 12205 -2263 12257 -2229
rect 12205 -2297 12214 -2263
rect 12248 -2297 12257 -2263
rect 12205 -2331 12257 -2297
rect 12205 -2365 12214 -2331
rect 12248 -2365 12257 -2331
rect 12205 -2399 12257 -2365
rect 12205 -2433 12214 -2399
rect 12248 -2433 12257 -2399
rect 12205 -2467 12257 -2433
rect 12205 -2501 12214 -2467
rect 12248 -2501 12257 -2467
rect 12205 -2535 12257 -2501
rect 12205 -2569 12214 -2535
rect 12248 -2569 12257 -2535
rect 12205 -2603 12257 -2569
rect 12205 -2637 12214 -2603
rect 12248 -2637 12257 -2603
rect 12205 -2671 12257 -2637
rect 12205 -2705 12214 -2671
rect 12248 -2705 12257 -2671
rect 12205 -2748 12257 -2705
rect 11592 -2756 12264 -2748
rect 11592 -2790 11674 -2756
rect 11708 -2790 11742 -2756
rect 11776 -2790 11810 -2756
rect 11844 -2790 11878 -2756
rect 11912 -2790 11946 -2756
rect 11980 -2790 12014 -2756
rect 12048 -2790 12082 -2756
rect 12116 -2790 12150 -2756
rect 12184 -2790 12264 -2756
rect 11592 -2797 12264 -2790
rect 11602 -2804 11640 -2797
rect 11302 -3408 11376 -3388
rect 11302 -3442 11323 -3408
rect 11357 -3442 11376 -3408
rect 11302 -4560 11376 -3442
rect 11854 -4453 11996 -4436
rect 11854 -4559 11870 -4453
rect 11976 -4559 11996 -4453
rect -1936 -5096 2814 -4938
rect 10754 -4564 11510 -4560
rect -1936 -5112 2424 -5096
rect 10754 -5210 10775 -4564
rect 11489 -4632 11510 -4564
rect 11854 -4632 11996 -4559
rect 11489 -4696 11996 -4632
rect 11489 -5067 11510 -4696
rect 12088 -5067 12164 -2797
rect 12205 -2798 12257 -2797
rect 11489 -5108 12164 -5067
rect 11489 -5116 12098 -5108
rect 11489 -5210 11510 -5116
rect 10754 -5214 11510 -5210
<< viali >>
rect 11323 -3442 11357 -3408
rect 11870 -4559 11976 -4453
<< metal1 >>
rect -1558 19046 280 19160
rect -1558 18098 -1307 19046
rect -39 18098 280 19046
rect -10172 6957 -10054 6990
rect -10172 6905 -10134 6957
rect -10082 6905 -10054 6957
rect -10172 5576 -10054 6905
rect -10242 148 -10208 5424
rect -10128 488 -10094 5576
rect -9856 5470 -9798 6671
rect -1558 6530 280 18098
rect -10014 148 -9980 5424
rect -9900 488 -9866 5424
rect -9786 148 -9752 5424
rect -5242 5076 -4606 5078
rect -7498 5074 -6336 5076
rect -5242 5074 -4600 5076
rect -8648 5070 -4600 5074
rect -8852 5068 -4600 5070
rect -9060 5032 -4600 5068
rect -9060 5030 -5216 5032
rect -9060 5028 -8848 5030
rect -8648 5028 -7486 5030
rect -6378 5028 -5216 5030
rect -9060 2670 -9030 5028
rect -4636 4984 -4600 5032
rect -4288 4984 -4058 4986
rect -4636 4956 -4058 4984
rect -4636 4954 -4252 4956
rect -4636 4738 -4600 4954
rect -9060 2644 -9028 2670
rect -9058 148 -9028 2644
rect -10420 120 -9028 148
rect -10420 114 -9032 120
rect -10420 112 -9702 114
rect -4400 -242 -4366 4828
rect -4286 -108 -4252 4954
rect -4018 4876 -3678 4922
rect -3708 4830 -3680 4876
rect -2972 4832 -2706 4834
rect -2972 4830 -2518 4832
rect -3730 4828 -2518 4830
rect -4172 -242 -4138 4828
rect -4058 -108 -4024 4828
rect -3944 3240 -3910 4828
rect -3730 4780 -2498 4828
rect -3730 4776 -2962 4780
rect -2856 4778 -2590 4780
rect -3944 3168 -2642 3240
rect -3944 3133 -2636 3168
rect -3944 3081 -2717 3133
rect -2665 3081 -2636 3133
rect -3944 3052 -2636 3081
rect -3944 3038 -2642 3052
rect -3944 -242 -3910 3038
rect -2556 2962 -2498 4780
rect 12586 3027 23592 6964
rect -2556 2956 -2496 2962
rect -2554 810 -2496 2956
rect 12585 2664 23592 3027
rect 12585 1308 12808 2664
rect 12674 1166 12712 1308
rect 12668 1164 12712 1166
rect 12668 852 12706 1164
rect 15940 1002 16178 1012
rect 16458 1002 16486 1004
rect 15940 996 16486 1002
rect 15940 982 18620 996
rect 15188 950 15338 980
rect 15938 950 15968 982
rect 16140 952 18620 982
rect 15188 900 15966 950
rect 16140 928 16486 952
rect 16140 922 16302 928
rect 16140 920 16178 922
rect -3294 790 -2496 810
rect -3302 674 -2496 790
rect -3302 664 -2504 674
rect -3302 -150 -3240 664
rect 15188 338 15338 900
rect 18582 892 18620 952
rect -3328 -193 -3088 -150
rect -4408 -286 -3896 -242
rect -3328 -245 -3169 -193
rect -3117 -245 -3088 -193
rect -3328 -286 -3088 -245
rect -4408 -288 -4126 -286
rect 12668 -498 12706 -94
rect 15188 -413 15379 338
rect 12674 -744 12712 -498
rect 13001 -509 15379 -413
rect 13001 -575 15306 -509
rect 12971 -707 15306 -575
rect 12971 -744 13037 -707
rect 12540 -770 13037 -744
rect 12015 -780 13037 -770
rect 12015 -818 13008 -780
rect 11831 -822 13008 -818
rect 11831 -869 12089 -822
rect 12540 -824 13008 -822
rect 12540 -825 12611 -824
rect 11942 -1060 12008 -1059
rect 12044 -1060 12089 -869
rect 12529 -1007 18626 -975
rect 12529 -1059 12659 -1007
rect 12711 -1059 18626 -1007
rect 11942 -1092 12121 -1060
rect 11942 -1093 12008 -1092
rect 11883 -2912 11917 -1127
rect 12001 -1176 12035 -1127
rect 12090 -1176 12121 -1092
rect 12001 -1214 12121 -1176
rect 12529 -1214 18626 -1059
rect 12001 -2469 12035 -1214
rect 12090 -1215 12121 -1214
rect 11169 -3033 11380 -3004
rect 11169 -3085 11198 -3033
rect 11250 -3085 11380 -3033
rect 11169 -3120 11380 -3085
rect 11300 -3408 11380 -3120
rect 11300 -3442 11323 -3408
rect 11357 -3442 11380 -3408
rect 11300 -3466 11380 -3442
rect 11846 -4453 11998 -2912
rect 11846 -4559 11870 -4453
rect 11976 -4559 11998 -4453
rect 11846 -4590 11998 -4559
<< via1 >>
rect -1307 18098 -39 19046
rect -10134 6905 -10082 6957
rect 5009 12922 5253 13166
rect -2717 3081 -2665 3133
rect -3169 -245 -3117 -193
rect 12659 -1059 12711 -1007
rect 11198 -3085 11250 -3033
<< metal2 >>
rect -1548 22376 300 22466
rect -1548 21520 -1214 22376
rect 122 21520 300 22376
rect -1548 19046 300 21520
rect -1548 18098 -1307 19046
rect -39 18098 300 19046
rect -1548 17946 300 18098
rect 4941 13769 5315 13832
rect 4941 13553 5028 13769
rect 5244 13553 5315 13769
rect 4941 13166 5315 13553
rect 4941 12922 5009 13166
rect 5253 12922 5315 13166
rect 4941 12842 5315 12922
rect -10172 7428 -10054 7442
rect -10172 7372 -10138 7428
rect -10082 7372 -10054 7428
rect -10172 6957 -10054 7372
rect -10172 6905 -10134 6957
rect -10082 6905 -10054 6957
rect -10172 6866 -10054 6905
rect -2752 3134 -2080 3176
rect -2752 3133 -2159 3134
rect -2752 3081 -2717 3133
rect -2665 3081 -2159 3133
rect -2752 3078 -2159 3081
rect -2103 3078 -2080 3134
rect -2752 3042 -2080 3078
rect -3204 -192 -2532 -150
rect -3204 -193 -2611 -192
rect -3204 -245 -3169 -193
rect -3117 -245 -2611 -193
rect -3204 -248 -2611 -245
rect -2555 -248 -2532 -192
rect -3204 -284 -2532 -248
rect 12529 -1007 12997 -975
rect 12529 -1059 12659 -1007
rect 12711 -1059 12997 -1007
rect 12529 -1680 12997 -1059
rect 12529 -1736 12783 -1680
rect 12839 -1736 12997 -1680
rect 12529 -1770 12997 -1736
rect 10613 -3030 11285 -2994
rect 10613 -3086 10636 -3030
rect 10692 -3033 11285 -3030
rect 10692 -3085 11198 -3033
rect 11250 -3085 11285 -3033
rect 10692 -3086 11285 -3085
rect 10613 -3128 11285 -3086
<< via2 >>
rect -1214 21520 122 22376
rect 5028 13553 5244 13769
rect -10138 7372 -10082 7428
rect -2159 3078 -2103 3134
rect -2611 -248 -2555 -192
rect 12783 -1736 12839 -1680
rect 10636 -3086 10692 -3030
<< metal3 >>
rect -1942 33938 924 34392
rect -1942 32114 -1564 33938
rect 580 32114 924 33938
rect -1942 29400 924 32114
rect -1942 29264 934 29400
rect -1932 26332 934 29264
rect -1936 24272 934 26332
rect -1936 22376 930 24272
rect -1936 21520 -1214 22376
rect 122 21520 930 22376
rect -1936 21204 930 21520
rect 4706 14295 5576 14370
rect 4706 14151 4833 14295
rect 5057 14151 5576 14295
rect 4706 13769 5576 14151
rect 4706 13553 5028 13769
rect 5244 13553 5576 13769
rect 4706 13500 5576 13553
rect -10168 7804 -10044 7816
rect -10168 7740 -10138 7804
rect -10074 7740 -10044 7804
rect -10168 7428 -10044 7740
rect -10168 7372 -10138 7428
rect -10082 7372 -10044 7428
rect -10168 7352 -10044 7372
rect -2188 3134 -1704 3170
rect -2188 3078 -2159 3134
rect -2103 3130 -1704 3134
rect -2103 3078 -1783 3130
rect -2188 3066 -1783 3078
rect -1719 3066 -1704 3130
rect -2188 3042 -1704 3066
rect -2640 -192 -2156 -156
rect -2640 -248 -2611 -192
rect -2555 -196 -2156 -192
rect -2555 -248 -2235 -196
rect -2640 -260 -2235 -248
rect -2171 -260 -2156 -196
rect -2640 -284 -2156 -260
rect 12529 -1680 12999 -1662
rect 12529 -1736 12783 -1680
rect 12839 -1736 12999 -1680
rect 12529 -2063 12999 -1736
rect 12529 -2127 12563 -2063
rect 12627 -2127 12999 -2063
rect 12529 -2146 12999 -2127
rect 10237 -3018 10721 -2994
rect 10237 -3082 10252 -3018
rect 10316 -3030 10721 -3018
rect 10316 -3082 10636 -3030
rect 10237 -3086 10636 -3082
rect 10692 -3086 10721 -3030
rect 10237 -3122 10721 -3086
<< via3 >>
rect -1564 32114 580 33938
rect 4833 14151 5057 14295
rect -10138 7740 -10074 7804
rect -1783 3066 -1719 3130
rect -2235 -260 -2171 -196
rect 12563 -2127 12627 -2063
rect 10252 -3082 10316 -3018
<< metal4 >>
rect -10554 25749 -9882 38208
rect -2884 35122 16204 36162
rect -2874 33938 1832 35122
rect -2874 32114 -1564 33938
rect 580 32114 1832 33938
rect -2874 31566 1832 32114
rect -10554 25238 9090 25749
rect -10554 7804 -9882 25238
rect 8960 23173 9090 25238
rect 16060 23428 16738 23780
rect 13764 23201 16738 23428
rect 8960 23036 12534 23173
rect 12051 19559 12534 23036
rect 4708 18678 11195 19484
rect 12051 18887 15999 19559
rect 4708 14295 5576 18678
rect 4708 14151 4833 14295
rect 5057 14151 5576 14295
rect 4708 14050 5576 14151
rect -10554 7740 -10138 7804
rect -10074 7740 -9882 7804
rect -10554 7704 -9882 7740
rect -1804 3130 -1355 3158
rect -1804 3066 -1783 3130
rect -1719 3066 -1355 3130
rect -1804 3038 -1355 3066
rect -1482 2849 1416 3026
rect 1017 -3515 1416 2849
rect 12529 -2063 12999 -2046
rect 12529 -2127 12563 -2063
rect 12627 -2127 12999 -2063
rect 3171 -2978 5778 -2970
rect 3171 -2990 10134 -2978
rect 3171 -3018 10337 -2990
rect 3171 -3082 10252 -3018
rect 10316 -3082 10337 -3018
rect 3171 -3110 10337 -3082
rect 3171 -3123 10134 -3110
rect 3171 -3359 3284 -3123
rect 3520 -3165 10134 -3123
rect 3520 -3359 5778 -3165
rect 3171 -3483 5778 -3359
rect -3005 -4109 1416 -3515
rect -3006 -8167 -2284 -4109
rect 12529 -11434 12999 -2127
rect 12529 -11670 12644 -11434
rect 12880 -11670 12999 -11434
rect 12529 -11768 12999 -11670
rect 32562 -14989 32762 708
rect 4270 -15106 32762 -14989
rect 2821 -22907 9680 -22284
rect 4768 -23822 5588 -22907
<< via4 >>
rect -7596 -1378 -6720 -822
rect 3284 -3359 3520 -3123
rect 12644 -11670 12880 -11434
<< metal5 >>
rect -10557 37208 7296 38208
rect -28744 -611 -27675 -400
rect -28856 -822 -6516 -611
rect -28856 -1378 -7596 -822
rect -6720 -1378 -6516 -822
rect -28856 -1590 -6516 -1378
rect -28744 -28336 -27675 -1590
rect 3192 -3123 3605 -2971
rect 3192 -3359 3284 -3123
rect 3520 -3359 3605 -3123
rect 3192 -5356 3605 -3359
rect 3238 -8176 3586 -5356
rect 3192 -8829 3605 -8176
rect 973 -8830 3605 -8829
rect -24150 -9304 -19438 -8856
rect -54 -8860 3605 -8830
rect -24974 -9992 -19438 -9304
rect -76 -9405 3605 -8860
rect -76 -9696 1186 -9405
rect 3192 -9407 3605 -9405
rect -24974 -12022 -23048 -9992
rect -25010 -21310 -23048 -12022
rect -76 -13282 720 -9696
rect 1748 -11383 12999 -11213
rect 1662 -11434 12999 -11383
rect 1662 -11670 12644 -11434
rect 12880 -11670 12999 -11434
rect 1662 -11769 12999 -11670
rect -25010 -23304 -23084 -21310
rect -68 -23132 690 -13282
rect -7532 -23304 690 -23132
rect -25010 -23340 690 -23304
rect -25010 -23958 482 -23340
rect -25010 -24028 -6536 -23958
rect -23462 -24096 -6536 -24028
rect 1662 -28336 2090 -11769
rect -28744 -28362 32796 -28336
rect 35266 -28362 36120 -9204
rect -28744 -29312 36120 -28362
rect -28744 -29561 32796 -29312
rect 35266 -29406 36120 -29312
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC1
timestamp 1669522153
transform 1 0 9723 0 1 21290
box -1711 -1972 1710 1995
use sky130_fd_pr__cap_mim_m3_1_FLZ2GZ  XC3
timestamp 1669522153
transform 1 0 6250 0 1 -18718
box -3568 -3814 3668 3729
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC4
timestamp 1669522153
transform 1 0 14527 0 1 21308
box -1711 -1972 1710 1995
use sky130_fd_pr__nfet_01v8_TAQE79  XM2
timestamp 1669522153
transform 1 0 -9997 0 1 2956
box -283 -2568 283 2568
use sky130_fd_pr__nfet_01v8_PAV6Y8  XM3
timestamp 1669522153
transform 1 0 11959 0 1 -1798
box -114 -755 114 755
use sky130_fd_pr__cap_mim_m3_1_LJH8TW  sky130_fd_pr__cap_mim_m3_1_LJH8TW_0
timestamp 1669522153
transform 1 0 -801 0 1 1362
box -1489 -1360 1488 1796
use sky130_fd_pr__nfet_01v8_TAQE79  sky130_fd_pr__nfet_01v8_TAQE79_0
timestamp 1669522153
transform 1 0 -4155 0 1 2360
box -283 -2568 283 2568
use sky130_fd_pr__res_xhigh_po_0p35_8U82AX  sky130_fd_pr__res_xhigh_po_0p35_8U82AX_0
timestamp 1669522153
transform 1 0 12687 0 1 376
box -35 -502 35 502
use sky130_fd_pr__res_xhigh_po_0p35_957LLN  sky130_fd_pr__res_xhigh_po_0p35_957LLN_0
timestamp 1669522153
transform 1 0 18601 0 1 -26
box -35 -942 35 942
use sq_ind_6p5n_f  sq_ind_6p5n_f_0
timestamp 1669522153
transform 1 0 9808 0 -1 39808
box -3200 -24600 24600 6756
use sq_ind_13n_f  sq_ind_13n_f_0
timestamp 1669522153
transform 0 -1 39496 1 0 -5372
box -4800 -26200 26200 4717
use sqr_ind_0p502n  sqr_ind_0p502n_0
timestamp 1669522153
transform 1 0 -20518 0 1 -8350
box 200 -13600 13200 1099
<< labels >>
rlabel locali s 10770 -5214 11494 -4560 4 GND
port 1 nsew
rlabel metal1 s 20408 4420 23150 6956 4 VDD
port 2 nsew
rlabel metal4 s 4768 -23822 5588 -23084 4 RFIN
port 3 nsew
rlabel metal4 s 16310 23440 16548 23660 4 RFOUT
port 4 nsew
<< end >>
