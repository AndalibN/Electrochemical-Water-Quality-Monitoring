magic
tech sky130A
magscale 1 2
timestamp 1668715771
<< psubdiff >>
rect -10835 6139 -10678 6144
rect -9376 6139 -9219 6144
rect -10841 6120 -10817 6139
rect -9220 6120 -9196 6139
rect -10841 5954 -10835 6120
rect -9219 5954 -9196 6120
rect -3616 5306 -3514 5330
rect -4802 5234 -4778 5300
rect -3514 5234 -3500 5300
rect -10859 -141 -10835 -21
rect -9200 -141 -9176 -21
rect -10835 -165 -10678 -141
rect -9376 -165 -9219 -141
rect 16371 409 16762 433
rect 12326 372 12438 396
rect -4818 -484 -4794 -418
rect -3500 -484 -3476 -418
rect -4770 -500 -4712 -484
rect -3616 -524 -3514 -500
rect 16371 -550 16762 -526
rect 12326 -746 12438 -722
rect 12205 -946 12257 -928
rect 11584 -974 11608 -946
rect 12248 -952 12272 -946
rect 11584 -995 11602 -974
rect 12257 -995 12272 -952
rect 11584 -2788 11602 -2748
rect 12257 -2782 12272 -2748
rect 11584 -2797 11608 -2788
rect 12248 -2797 12272 -2782
rect 11602 -2812 11640 -2797
rect 12205 -2806 12257 -2797
rect 10746 -5214 10770 -4560
rect 11494 -5214 11518 -4560
<< psubdiffcont >>
rect -10817 6120 -9220 6139
rect -10835 5954 -9219 6120
rect -10835 -21 -10678 5954
rect -9376 -21 -9219 5954
rect -3616 5300 -3514 5306
rect -4778 5234 -3514 5300
rect -10835 -141 -9200 -21
rect -4770 -418 -4712 5234
rect -3616 -418 -3514 5234
rect -4794 -484 -3500 -418
rect -3616 -500 -3514 -484
rect 12326 -722 12438 372
rect 16371 -526 16762 409
rect 11608 -952 12248 -946
rect 11608 -974 12257 -952
rect 11602 -995 12257 -974
rect 11602 -2748 11640 -995
rect 12205 -2748 12257 -995
rect 11602 -2782 12257 -2748
rect 11602 -2788 12248 -2782
rect 11608 -2797 12248 -2788
rect 10770 -5214 11494 -4560
<< locali >>
rect -10833 6136 -10817 6139
rect -10835 6120 -10817 6136
rect -9220 6120 -9204 6139
rect -9219 5954 -9204 6120
rect -9380 5178 -9376 5240
rect -10128 352 -10094 668
rect -9900 382 -9866 676
rect -9901 352 -9866 382
rect -10129 348 -9866 352
rect -10129 306 -9867 348
rect -3616 5306 -3514 5322
rect -4794 5240 -4778 5300
rect -9219 5234 -4778 5240
rect -3514 5234 -3508 5300
rect -9219 5178 -4770 5234
rect -10851 -141 -10835 -21
rect -9200 -141 -9184 -21
rect -10835 -157 -10678 -141
rect -9376 -157 -9219 -141
rect -4286 -326 -4252 -88
rect -4058 -326 -4024 -80
rect -4286 -364 -4024 -326
rect 4920 5196 5102 5197
rect -3514 5074 5102 5196
rect -4810 -484 -4794 -418
rect -3500 -484 -3484 -418
rect -4770 -492 -4712 -484
rect -3616 -516 -3514 -500
rect 2318 -4938 2814 5074
rect 4920 -1358 5102 5074
rect 12366 1476 12436 1485
rect 16600 1476 16646 1546
rect 12366 1444 16646 1476
rect 12366 1386 25368 1444
rect 10890 780 10944 792
rect 12366 780 12436 1386
rect 16598 1228 25368 1386
rect 10890 716 12436 780
rect 10890 -1358 10944 716
rect 12366 388 12436 716
rect 16600 534 16646 1228
rect 16600 425 16670 534
rect 16371 409 16762 425
rect 12326 372 12438 388
rect 16371 -542 16762 -526
rect 12326 -738 12438 -722
rect 12205 -946 12257 -936
rect 11592 -974 11608 -946
rect 12248 -952 12264 -946
rect 11592 -995 11602 -974
rect 12257 -995 12264 -952
rect 11562 -1358 11602 -1350
rect 4920 -1460 11602 -1358
rect 11562 -1466 11602 -1460
rect 11592 -2788 11602 -2748
rect 12257 -2782 12264 -2748
rect 11592 -2797 11608 -2788
rect 12248 -2797 12264 -2782
rect 11602 -2804 11640 -2797
rect 11302 -3404 11376 -3388
rect 11302 -3446 11310 -3404
rect 11370 -3446 11376 -3404
rect 11302 -4560 11376 -3446
rect 11854 -4448 11996 -4436
rect -1936 -5096 2814 -4938
rect -1936 -5112 2424 -5096
rect 10754 -5214 10770 -4560
rect 11494 -4632 11510 -4560
rect 11854 -4564 11866 -4448
rect 11980 -4564 11996 -4448
rect 11854 -4632 11996 -4564
rect 11494 -4696 11996 -4632
rect 11494 -5067 11510 -4696
rect 12088 -5067 12164 -2797
rect 12205 -2798 12257 -2797
rect 11494 -5108 12164 -5067
rect 11494 -5116 12098 -5108
rect 11494 -5214 11510 -5116
<< viali >>
rect 11310 -3446 11370 -3404
rect 11866 -4564 11980 -4448
<< metal1 >>
rect -1748 19058 280 19160
rect -1748 18086 -1320 19058
rect -26 18086 280 19058
rect -1748 15844 280 18086
rect 11960 15844 12210 16334
rect -1748 15080 12210 15844
rect -1748 15012 280 15080
rect -1772 14346 280 15012
rect 11960 14432 12210 15080
rect 11948 14390 12210 14432
rect 11948 14294 12204 14390
rect 4618 13200 5094 13234
rect 4618 12912 4738 13200
rect 5000 12912 5094 13200
rect 4618 11938 5094 12912
rect 11994 12484 12194 14294
rect 13030 12484 13166 12504
rect 11994 12446 13166 12484
rect 12002 12294 13166 12446
rect 12960 12112 13166 12294
rect 4786 9450 4984 11938
rect 12960 9664 13122 12112
rect 12964 9572 13116 9664
rect 12006 9530 13116 9572
rect 11994 9450 13116 9530
rect 4786 9382 13078 9450
rect 4786 9250 12382 9382
rect 11994 8234 12194 9250
rect 11756 7654 12194 8234
rect 11994 7232 12194 7654
rect 20136 7232 23624 7236
rect -10172 6974 -10054 6990
rect -10172 6888 -10146 6974
rect -10070 6888 -10054 6974
rect -10172 6586 -10054 6888
rect 11994 6964 23624 7232
rect -10156 6500 -10070 6586
rect -10128 5716 -10094 6500
rect 11994 5860 12194 6964
rect 11994 5842 12190 5860
rect 11266 5836 12190 5842
rect 9442 5832 12190 5836
rect 5786 5828 12190 5832
rect 3948 5824 12190 5828
rect 318 5822 12190 5824
rect -3232 5820 12190 5822
rect -5082 5818 12190 5820
rect -8278 5814 -7116 5816
rect -6022 5814 12190 5818
rect -9428 5810 12190 5814
rect -9632 5808 12190 5810
rect -9840 5792 12190 5808
rect -9840 5786 11310 5792
rect -9840 5782 9472 5786
rect -9840 5778 5816 5782
rect -9840 5774 3996 5778
rect -9840 5772 454 5774
rect -9840 5770 -5996 5772
rect -5082 5770 -3214 5772
rect -9840 5768 -9628 5770
rect -9428 5768 -8266 5770
rect -7158 5768 -5996 5770
rect -10128 5594 -10082 5716
rect -9840 5706 -9810 5768
rect -9856 5678 -9798 5706
rect -9836 5598 -9806 5678
rect -10242 148 -10208 5424
rect -10128 488 -10094 5594
rect -9856 5470 -9798 5598
rect 19960 5486 23624 6964
rect -10014 148 -9980 5424
rect -9900 488 -9866 5424
rect -9786 148 -9752 5424
rect 18778 5419 23624 5486
rect -5242 5076 -4606 5078
rect -7498 5074 -6336 5076
rect -5242 5074 -4600 5076
rect -8648 5070 -4600 5074
rect -8852 5068 -4600 5070
rect -9060 5032 -4600 5068
rect -9060 5030 -5216 5032
rect -9060 5028 -8848 5030
rect -8648 5028 -7486 5030
rect -6378 5028 -5216 5030
rect -9060 2670 -9030 5028
rect -4636 4984 -4600 5032
rect -4288 4984 -4058 4986
rect -4636 4956 -4058 4984
rect -4636 4954 -4252 4956
rect -4636 4738 -4600 4954
rect -9060 2644 -9028 2670
rect -9058 148 -9028 2644
rect -10420 120 -9028 148
rect -10420 114 -9032 120
rect -10420 112 -9702 114
rect -4400 -242 -4366 4828
rect -4286 -108 -4252 4954
rect -4018 4876 -3678 4922
rect -3708 4830 -3680 4876
rect -2972 4832 -2706 4834
rect -2972 4830 -2518 4832
rect -3730 4828 -2518 4830
rect -4172 -242 -4138 4828
rect -4058 -108 -4024 4828
rect -3944 3240 -3910 4828
rect -3730 4780 -2498 4828
rect -3730 4776 -2962 4780
rect -2856 4778 -2590 4780
rect -3944 3168 -2642 3240
rect -3944 3160 -2636 3168
rect -3944 3054 -2736 3160
rect -2646 3054 -2636 3160
rect -3944 3052 -2636 3054
rect -3944 3038 -2642 3052
rect -3944 -242 -3910 3038
rect -2556 2962 -2498 4780
rect 19960 4184 23624 5419
rect 19960 3693 20376 4184
rect 12622 3413 20376 3693
rect 12585 3064 20376 3413
rect 12585 3027 20196 3064
rect -2556 2956 -2496 2962
rect -2554 810 -2496 2956
rect -3294 790 -2496 810
rect -3302 674 -2496 790
rect -3302 664 -2504 674
rect -3302 -150 -3240 664
rect 12585 383 12808 3027
rect 12541 322 12808 383
rect 15188 950 15338 980
rect 15188 900 15944 950
rect 15188 338 15338 900
rect 12541 318 12711 322
rect 12541 171 12612 318
rect -3328 -166 -3088 -150
rect -4408 -286 -3896 -242
rect -3328 -272 -3188 -166
rect -3098 -272 -3088 -166
rect -3328 -286 -3088 -272
rect -4408 -288 -4126 -286
rect 15188 -413 15379 338
rect 13001 -509 15379 -413
rect 13001 -575 15306 -509
rect 12540 -744 12611 -637
rect 12971 -707 15306 -575
rect 12971 -744 13037 -707
rect 12540 -770 13037 -744
rect 12015 -780 13037 -770
rect 12015 -818 13008 -780
rect 11831 -822 13008 -818
rect 11831 -869 12089 -822
rect 12540 -824 13008 -822
rect 12540 -825 12611 -824
rect 11942 -1060 12008 -1059
rect 12044 -1060 12089 -869
rect 15890 -888 15956 -450
rect 15560 -895 15956 -888
rect 12778 -974 15956 -895
rect 12778 -975 15952 -974
rect 11942 -1092 12121 -1060
rect 11942 -1093 12008 -1092
rect 11883 -2912 11917 -1127
rect 12001 -1176 12035 -1127
rect 12090 -1176 12121 -1092
rect 12001 -1214 12121 -1176
rect 12778 -1114 12894 -975
rect 15560 -976 15952 -975
rect 12778 -1204 12780 -1114
rect 12886 -1204 12894 -1114
rect 12778 -1214 12894 -1204
rect 12001 -2469 12035 -1214
rect 12090 -1215 12121 -1214
rect 11169 -3006 11380 -3004
rect 11169 -3112 11179 -3006
rect 11269 -3112 11380 -3006
rect 11169 -3120 11380 -3112
rect 11300 -3404 11380 -3120
rect 11300 -3446 11310 -3404
rect 11370 -3446 11380 -3404
rect 11300 -3466 11380 -3446
rect 11846 -4448 11998 -2912
rect 11846 -4564 11866 -4448
rect 11980 -4564 11998 -4448
rect 11846 -4590 11998 -4564
<< via1 >>
rect -1320 18086 -26 19058
rect 4738 12912 5000 13200
rect -10146 6888 -10070 6974
rect -2736 3054 -2646 3160
rect -3188 -272 -3098 -166
rect 12780 -1204 12886 -1114
rect 11179 -3112 11269 -3006
<< metal2 >>
rect -1548 22396 300 22466
rect -1548 21500 -1250 22396
rect 158 21500 300 22396
rect -1548 19058 300 21500
rect -1548 18086 -1320 19058
rect -26 18086 300 19058
rect -1548 17946 300 18086
rect 4680 13790 5054 13830
rect 4680 13564 4738 13790
rect 4994 13564 5054 13790
rect 4680 13200 5054 13564
rect 4680 12912 4738 13200
rect 5000 12912 5054 13200
rect 4680 12840 5054 12912
rect -10172 7430 -10054 7442
rect -10172 7370 -10150 7430
rect -10070 7370 -10054 7430
rect -10172 6974 -10054 7370
rect -10172 6888 -10146 6974
rect -10070 6888 -10054 6974
rect -10172 6866 -10054 6888
rect -2752 3160 -2080 3176
rect -2752 3054 -2736 3160
rect -2646 3156 -2080 3160
rect -2646 3056 -2172 3156
rect -2090 3056 -2080 3156
rect -2646 3054 -2080 3056
rect -2752 3042 -2080 3054
rect -3204 -166 -2532 -150
rect -3204 -272 -3188 -166
rect -3098 -170 -2532 -166
rect -3098 -270 -2624 -170
rect -2542 -270 -2532 -170
rect -3098 -272 -2532 -270
rect -3204 -284 -2532 -272
rect 12768 -1114 12902 -1098
rect 12768 -1204 12780 -1114
rect 12886 -1204 12902 -1114
rect 12768 -1678 12902 -1204
rect 12768 -1760 12782 -1678
rect 12882 -1760 12902 -1678
rect 12768 -1770 12902 -1760
rect 10613 -3006 11285 -2994
rect 10613 -3008 11179 -3006
rect 10613 -3108 10623 -3008
rect 10705 -3108 11179 -3008
rect 10613 -3112 11179 -3108
rect 11269 -3112 11285 -3006
rect 10613 -3128 11285 -3112
<< via2 >>
rect -1250 21500 158 22396
rect 4738 13564 4994 13790
rect -10150 7370 -10070 7430
rect -2172 3056 -2090 3156
rect -2624 -270 -2542 -170
rect 12782 -1760 12882 -1678
rect 10623 -3108 10705 -3008
<< metal3 >>
rect -1942 33954 924 34392
rect -1942 32098 -1572 33954
rect 588 32098 924 33954
rect -1942 29400 924 32098
rect -1942 29264 934 29400
rect -1932 26332 934 29264
rect -1936 24272 934 26332
rect -1936 22396 930 24272
rect -1936 21500 -1250 22396
rect 158 21500 930 22396
rect -1936 21204 930 21500
rect 4682 14332 5048 14370
rect 4682 14114 4748 14332
rect 4982 14114 5048 14332
rect 4682 13790 5048 14114
rect 4682 13564 4738 13790
rect 4994 13564 5048 13790
rect 4682 13500 5048 13564
rect -10168 7804 -10044 7816
rect -10168 7740 -10146 7804
rect -10066 7740 -10044 7804
rect -10168 7430 -10044 7740
rect -10168 7370 -10150 7430
rect -10070 7370 -10044 7430
rect -10168 7352 -10044 7370
rect -2188 3156 -1704 3170
rect -2188 3056 -2172 3156
rect -2090 3148 -1704 3156
rect -2090 3056 -1792 3148
rect -2188 3048 -1792 3056
rect -1710 3048 -1704 3148
rect -2188 3042 -1704 3048
rect -2640 -170 -2156 -156
rect -2640 -270 -2624 -170
rect -2542 -178 -2156 -170
rect -2542 -270 -2244 -178
rect -2640 -278 -2244 -270
rect -2162 -278 -2156 -178
rect -2640 -284 -2156 -278
rect 12768 -1678 12896 -1662
rect 12768 -1760 12782 -1678
rect 12882 -1760 12896 -1678
rect 12768 -2058 12896 -1760
rect 12768 -2140 12774 -2058
rect 12874 -2140 12896 -2058
rect 12768 -2146 12896 -2140
rect 10237 -3000 10721 -2994
rect 10237 -3100 10243 -3000
rect 10325 -3008 10721 -3000
rect 10325 -3100 10623 -3008
rect 10237 -3108 10623 -3100
rect 10705 -3108 10721 -3008
rect 10237 -3122 10721 -3108
<< via3 >>
rect -1572 32098 588 33954
rect 4748 14114 4982 14332
rect -10146 7740 -10066 7804
rect -1792 3048 -1710 3148
rect -2244 -278 -2162 -178
rect 12774 -2140 12874 -2058
rect 10243 -3100 10325 -3000
<< metal4 >>
rect -13282 38314 -11178 38468
rect -13282 36108 -13128 38314
rect -11436 36108 -11178 38314
rect -13282 31672 -11178 36108
rect -2884 35122 16204 36162
rect -13406 31534 -11178 31672
rect -2874 33954 1832 35122
rect -2874 32098 -1572 33954
rect 588 32098 1832 33954
rect -2874 31566 1832 32098
rect -13406 30770 -11230 31534
rect -13386 26930 -11282 30770
rect 9000 26950 9318 26958
rect 4024 26946 9318 26950
rect 1880 26930 9318 26946
rect -13386 26352 9318 26930
rect -13386 26286 4644 26352
rect -13386 25482 1978 26286
rect -13386 15040 -11282 25482
rect 9000 23118 9318 26352
rect 16060 23290 16738 23780
rect 16030 23286 16738 23290
rect 13764 23162 16738 23286
rect 13764 23160 16210 23162
rect 8958 23036 12366 23118
rect 8958 22928 9068 23036
rect 10130 22892 10234 23036
rect 11300 22920 11402 23036
rect 12192 23034 12366 23036
rect 4708 19556 5026 19562
rect 8448 19556 8558 19696
rect 4708 19482 8558 19556
rect 9622 19482 9732 19704
rect 10790 19482 10900 19698
rect 4708 19396 10900 19482
rect 12224 19462 12366 23034
rect 13764 22928 13868 23160
rect 14936 22928 15038 23160
rect 16106 22928 16210 23160
rect 13332 19718 13358 19722
rect 13252 19462 13362 19716
rect 14422 19462 14532 19704
rect 15596 19462 15700 19708
rect 12224 19458 15700 19462
rect 4708 19018 5026 19396
rect 8448 19392 10900 19396
rect 12222 19336 15700 19458
rect 12222 19334 13246 19336
rect 12222 19240 12376 19334
rect 4708 18678 11736 19018
rect 4708 15760 5026 18678
rect 4708 15750 5036 15760
rect -13386 14642 -10034 15040
rect 4698 14658 5036 15750
rect -13386 14624 -11282 14642
rect -10164 7966 -10070 14642
rect 4688 14332 5036 14658
rect 4688 14114 4748 14332
rect 4982 14114 5036 14332
rect 4688 14026 5036 14114
rect 4688 14004 5010 14026
rect -10164 7804 -10040 7966
rect -10164 7740 -10146 7804
rect -10066 7740 -10040 7804
rect -10164 7726 -10040 7740
rect -1804 3148 -1643 3158
rect -1804 3048 -1792 3148
rect -1710 3048 -1643 3148
rect -1804 3038 -1643 3048
rect -1803 2938 -1647 3038
rect 1404 2982 1685 3201
rect 598 2940 1685 2982
rect 596 2938 1685 2940
rect -2053 2911 1685 2938
rect -2053 2849 659 2911
rect -1482 2770 -1378 2849
rect -464 2771 -360 2849
rect 544 2771 659 2849
rect -1923 -168 -1813 -44
rect -2256 -172 -1813 -168
rect -903 -172 -799 -47
rect 116 -172 220 -47
rect -2256 -178 686 -172
rect -2256 -278 -2244 -178
rect -2162 -278 686 -178
rect -2256 -288 686 -278
rect -1840 -608 -1503 -288
rect -7700 -769 -1503 -608
rect -7700 -1431 -7640 -769
rect -6676 -1431 -1503 -769
rect -7700 -1552 -1503 -1431
rect -1840 -1553 -1503 -1552
rect 1404 -3215 1685 2911
rect 12764 -2058 12884 -2046
rect 12764 -2140 12774 -2058
rect 12874 -2140 12884 -2058
rect 12764 -2249 12884 -2140
rect 12752 -2519 12939 -2249
rect 12698 -2665 12939 -2519
rect 3171 -2978 5778 -2970
rect 3171 -2990 10134 -2978
rect 3171 -3000 10337 -2990
rect 3171 -3057 10243 -3000
rect -3094 -3510 1711 -3215
rect 3171 -3425 3243 -3057
rect 3561 -3100 10243 -3057
rect 10325 -3100 10337 -3000
rect 3561 -3110 10337 -3100
rect 3561 -3165 10134 -3110
rect 12698 -3127 12914 -2665
rect 3561 -3425 5778 -3165
rect 3171 -3483 5778 -3425
rect -3362 -4109 1711 -3510
rect -16890 -7376 -5572 -7136
rect -17028 -7584 -5572 -7376
rect -17028 -7756 -5504 -7584
rect -17028 -8718 -16444 -7756
rect -5848 -10920 -5504 -7756
rect -3362 -8694 -2906 -4109
rect -3340 -8832 -3128 -8694
rect -3594 -9656 -3128 -8832
rect -4016 -10920 -3126 -9656
rect -5848 -11126 -3126 -10920
rect -5778 -11470 -3126 -11126
rect -4016 -11684 -3126 -11470
rect -3608 -11702 -3126 -11684
rect -3606 -11707 -3126 -11702
rect 12347 -11292 12982 -3127
rect 12347 -11697 12401 -11292
rect 12941 -11697 12982 -11292
rect 12347 -11751 12982 -11697
rect 3806 -12852 4130 -12825
rect 32562 -12852 33294 1062
rect 3755 -13160 33294 -12852
rect 3755 -13290 32796 -13160
rect 3806 -14863 4130 -13290
rect 3806 -14876 9858 -14863
rect 3433 -14978 9858 -14876
rect 3433 -14990 9891 -14978
rect 4266 -15282 4369 -14990
rect 6109 -15281 6213 -14990
rect 7947 -15280 8051 -14990
rect 9787 -15281 9891 -14990
rect 3447 -22395 3538 -22151
rect 3440 -22399 3897 -22395
rect 5291 -22399 5382 -22151
rect 7127 -22399 7218 -22152
rect 8960 -22399 9051 -22152
rect 3440 -22533 9924 -22399
rect 5005 -23084 5301 -22533
rect 4768 -23822 5588 -23084
<< via4 >>
rect -13128 36108 -11436 38314
rect -7640 -1431 -6676 -769
rect 3243 -3425 3561 -3057
rect 12401 -11697 12941 -11292
<< metal5 >>
rect -13306 46350 -5208 46454
rect -13306 45284 -4756 46350
rect -13302 38314 -11298 45284
rect -13302 36108 -13128 38314
rect -11436 36108 -11298 38314
rect -5428 38140 -4756 45284
rect -5572 37276 7296 38140
rect -13302 35788 -11298 36108
rect -28744 -611 -27675 -400
rect -28856 -769 -6516 -611
rect -28856 -1431 -7640 -769
rect -6676 -1431 -6516 -769
rect -28856 -1590 -6516 -1431
rect -28744 -28336 -27675 -1590
rect 3192 -3057 3605 -2971
rect 3192 -3425 3243 -3057
rect 3561 -3425 3605 -3057
rect 3192 -5356 3605 -3425
rect 3238 -8176 3586 -5356
rect 3192 -8829 3605 -8176
rect 973 -8830 3605 -8829
rect -24150 -9304 -19438 -8856
rect -54 -8860 3605 -8830
rect -24974 -9992 -19438 -9304
rect -76 -9405 3605 -8860
rect -76 -9696 1186 -9405
rect 3192 -9407 3605 -9405
rect -24974 -12022 -23048 -9992
rect -25010 -21310 -23048 -12022
rect -76 -13282 720 -9696
rect 1748 -11292 12999 -11213
rect 1748 -11383 12401 -11292
rect 1662 -11697 12401 -11383
rect 12941 -11697 12999 -11292
rect 1662 -11769 12999 -11697
rect -25010 -23304 -23084 -21310
rect -68 -23132 690 -13282
rect -7532 -23304 690 -23132
rect -25010 -23340 690 -23304
rect -25010 -23958 482 -23340
rect -25010 -24028 -6536 -23958
rect -23462 -24096 -6536 -24028
rect 1662 -28336 2090 -11769
rect -28744 -28362 32796 -28336
rect 35266 -28362 36120 -9204
rect -28744 -29312 36120 -28362
rect -28744 -29561 32796 -29312
rect 35266 -29406 36120 -29312
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC1
timestamp 1667951165
transform 1 0 9723 0 1 21290
box -1711 -1620 1710 1640
use sky130_fd_pr__cap_mim_m3_1_FLZ2GZ  XC3
timestamp 1667951165
transform 1 0 6250 0 1 -18718
box -3568 -3440 3668 3440
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC4
timestamp 1667951165
transform 1 0 14527 0 1 21308
box -1711 -1620 1710 1640
use sky130_fd_pr__nfet_01v8_TAQE79  XM2
timestamp 1668019001
transform 1 0 -9997 0 1 2956
box -257 -2568 257 2568
use sky130_fd_pr__nfet_01v8_PAV6Y8  XM3
timestamp 1668017392
transform 1 0 11959 0 1 -1798
box -88 -755 88 755
use sky130_fd_pr__cap_mim_m3_1_LJH8TW  sky130_fd_pr__cap_mim_m3_1_LJH8TW_1
timestamp 1667951165
transform 1 0 -801 0 1 1362
box -1489 -1410 1488 1410
use sky130_fd_pr__nfet_01v8_TAQE79  sky130_fd_pr__nfet_01v8_TAQE79_0
timestamp 1668019001
transform 1 0 -4155 0 1 2360
box -257 -2568 257 2568
use sky130_fd_pr__res_xhigh_po_0p35_BELDZV  sky130_fd_pr__res_xhigh_po_0p35_BELDZV_0
timestamp 1668226266
transform -1 0 12576 0 1 -217
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_Y9Q9SK  sky130_fd_pr__res_xhigh_po_0p35_Y9Q9SK_0
timestamp 1668226266
transform -1 0 15923 0 -1 56
box -37 -932 37 932
use sq_ind_6p5n_f  sq_ind_6p5n_f_0
timestamp 1668222614
transform 1 0 9808 0 -1 39808
box -3200 -24600 24600 6756
use sq_ind_13n_f  sq_ind_13n_f_0
timestamp 1668222539
transform 0 -1 39496 1 0 -5372
box -4800 -26200 26200 6756
use sqr_ind_0p502n  sqr_ind_0p502n_0
timestamp 1668384124
transform 1 0 -20518 0 1 -8350
box 1200 -12000 11600 -300
<< labels >>
rlabel metal4 16310 23440 16548 23660 1 RFOUT
port 1 n
rlabel metal4 4768 -23822 5588 -23084 1 RFIN
port 2 n
rlabel metal1 20408 4420 23150 6956 1 VDD
port 4 n
rlabel psubdiffcont 10770 -5214 11494 -4560 1 GND
port 3 n
<< end >>
