magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -1098 -740 948 742
<< pmos >>
rect -754 -624 -714 626
rect -656 -624 -616 626
rect -558 -624 -518 626
rect -460 -624 -420 626
rect -362 -624 -322 626
rect -264 -624 -224 626
rect -166 -624 -126 626
rect -68 -624 -28 626
rect 30 -624 70 626
rect 128 -624 168 626
rect 226 -624 266 626
rect 324 -624 364 626
rect 422 -624 462 626
rect 520 -624 560 626
rect 618 -624 658 626
rect 716 -624 756 626
<< pdiff >>
rect -812 596 -754 626
rect -812 562 -800 596
rect -766 562 -754 596
rect -812 528 -754 562
rect -812 494 -800 528
rect -766 494 -754 528
rect -812 460 -754 494
rect -812 426 -800 460
rect -766 426 -754 460
rect -812 392 -754 426
rect -812 358 -800 392
rect -766 358 -754 392
rect -812 324 -754 358
rect -812 290 -800 324
rect -766 290 -754 324
rect -812 256 -754 290
rect -812 222 -800 256
rect -766 222 -754 256
rect -812 188 -754 222
rect -812 154 -800 188
rect -766 154 -754 188
rect -812 120 -754 154
rect -812 86 -800 120
rect -766 86 -754 120
rect -812 52 -754 86
rect -812 18 -800 52
rect -766 18 -754 52
rect -812 -16 -754 18
rect -812 -50 -800 -16
rect -766 -50 -754 -16
rect -812 -84 -754 -50
rect -812 -118 -800 -84
rect -766 -118 -754 -84
rect -812 -152 -754 -118
rect -812 -186 -800 -152
rect -766 -186 -754 -152
rect -812 -220 -754 -186
rect -812 -254 -800 -220
rect -766 -254 -754 -220
rect -812 -288 -754 -254
rect -812 -322 -800 -288
rect -766 -322 -754 -288
rect -812 -356 -754 -322
rect -812 -390 -800 -356
rect -766 -390 -754 -356
rect -812 -424 -754 -390
rect -812 -458 -800 -424
rect -766 -458 -754 -424
rect -812 -492 -754 -458
rect -812 -526 -800 -492
rect -766 -526 -754 -492
rect -812 -560 -754 -526
rect -812 -594 -800 -560
rect -766 -594 -754 -560
rect -812 -624 -754 -594
rect -714 596 -656 626
rect -714 562 -702 596
rect -668 562 -656 596
rect -714 528 -656 562
rect -714 494 -702 528
rect -668 494 -656 528
rect -714 460 -656 494
rect -714 426 -702 460
rect -668 426 -656 460
rect -714 392 -656 426
rect -714 358 -702 392
rect -668 358 -656 392
rect -714 324 -656 358
rect -714 290 -702 324
rect -668 290 -656 324
rect -714 256 -656 290
rect -714 222 -702 256
rect -668 222 -656 256
rect -714 188 -656 222
rect -714 154 -702 188
rect -668 154 -656 188
rect -714 120 -656 154
rect -714 86 -702 120
rect -668 86 -656 120
rect -714 52 -656 86
rect -714 18 -702 52
rect -668 18 -656 52
rect -714 -16 -656 18
rect -714 -50 -702 -16
rect -668 -50 -656 -16
rect -714 -84 -656 -50
rect -714 -118 -702 -84
rect -668 -118 -656 -84
rect -714 -152 -656 -118
rect -714 -186 -702 -152
rect -668 -186 -656 -152
rect -714 -220 -656 -186
rect -714 -254 -702 -220
rect -668 -254 -656 -220
rect -714 -288 -656 -254
rect -714 -322 -702 -288
rect -668 -322 -656 -288
rect -714 -356 -656 -322
rect -714 -390 -702 -356
rect -668 -390 -656 -356
rect -714 -424 -656 -390
rect -714 -458 -702 -424
rect -668 -458 -656 -424
rect -714 -492 -656 -458
rect -714 -526 -702 -492
rect -668 -526 -656 -492
rect -714 -560 -656 -526
rect -714 -594 -702 -560
rect -668 -594 -656 -560
rect -714 -624 -656 -594
rect -616 596 -558 626
rect -616 562 -604 596
rect -570 562 -558 596
rect -616 528 -558 562
rect -616 494 -604 528
rect -570 494 -558 528
rect -616 460 -558 494
rect -616 426 -604 460
rect -570 426 -558 460
rect -616 392 -558 426
rect -616 358 -604 392
rect -570 358 -558 392
rect -616 324 -558 358
rect -616 290 -604 324
rect -570 290 -558 324
rect -616 256 -558 290
rect -616 222 -604 256
rect -570 222 -558 256
rect -616 188 -558 222
rect -616 154 -604 188
rect -570 154 -558 188
rect -616 120 -558 154
rect -616 86 -604 120
rect -570 86 -558 120
rect -616 52 -558 86
rect -616 18 -604 52
rect -570 18 -558 52
rect -616 -16 -558 18
rect -616 -50 -604 -16
rect -570 -50 -558 -16
rect -616 -84 -558 -50
rect -616 -118 -604 -84
rect -570 -118 -558 -84
rect -616 -152 -558 -118
rect -616 -186 -604 -152
rect -570 -186 -558 -152
rect -616 -220 -558 -186
rect -616 -254 -604 -220
rect -570 -254 -558 -220
rect -616 -288 -558 -254
rect -616 -322 -604 -288
rect -570 -322 -558 -288
rect -616 -356 -558 -322
rect -616 -390 -604 -356
rect -570 -390 -558 -356
rect -616 -424 -558 -390
rect -616 -458 -604 -424
rect -570 -458 -558 -424
rect -616 -492 -558 -458
rect -616 -526 -604 -492
rect -570 -526 -558 -492
rect -616 -560 -558 -526
rect -616 -594 -604 -560
rect -570 -594 -558 -560
rect -616 -624 -558 -594
rect -518 596 -460 626
rect -518 562 -506 596
rect -472 562 -460 596
rect -518 528 -460 562
rect -518 494 -506 528
rect -472 494 -460 528
rect -518 460 -460 494
rect -518 426 -506 460
rect -472 426 -460 460
rect -518 392 -460 426
rect -518 358 -506 392
rect -472 358 -460 392
rect -518 324 -460 358
rect -518 290 -506 324
rect -472 290 -460 324
rect -518 256 -460 290
rect -518 222 -506 256
rect -472 222 -460 256
rect -518 188 -460 222
rect -518 154 -506 188
rect -472 154 -460 188
rect -518 120 -460 154
rect -518 86 -506 120
rect -472 86 -460 120
rect -518 52 -460 86
rect -518 18 -506 52
rect -472 18 -460 52
rect -518 -16 -460 18
rect -518 -50 -506 -16
rect -472 -50 -460 -16
rect -518 -84 -460 -50
rect -518 -118 -506 -84
rect -472 -118 -460 -84
rect -518 -152 -460 -118
rect -518 -186 -506 -152
rect -472 -186 -460 -152
rect -518 -220 -460 -186
rect -518 -254 -506 -220
rect -472 -254 -460 -220
rect -518 -288 -460 -254
rect -518 -322 -506 -288
rect -472 -322 -460 -288
rect -518 -356 -460 -322
rect -518 -390 -506 -356
rect -472 -390 -460 -356
rect -518 -424 -460 -390
rect -518 -458 -506 -424
rect -472 -458 -460 -424
rect -518 -492 -460 -458
rect -518 -526 -506 -492
rect -472 -526 -460 -492
rect -518 -560 -460 -526
rect -518 -594 -506 -560
rect -472 -594 -460 -560
rect -518 -624 -460 -594
rect -420 596 -362 626
rect -420 562 -408 596
rect -374 562 -362 596
rect -420 528 -362 562
rect -420 494 -408 528
rect -374 494 -362 528
rect -420 460 -362 494
rect -420 426 -408 460
rect -374 426 -362 460
rect -420 392 -362 426
rect -420 358 -408 392
rect -374 358 -362 392
rect -420 324 -362 358
rect -420 290 -408 324
rect -374 290 -362 324
rect -420 256 -362 290
rect -420 222 -408 256
rect -374 222 -362 256
rect -420 188 -362 222
rect -420 154 -408 188
rect -374 154 -362 188
rect -420 120 -362 154
rect -420 86 -408 120
rect -374 86 -362 120
rect -420 52 -362 86
rect -420 18 -408 52
rect -374 18 -362 52
rect -420 -16 -362 18
rect -420 -50 -408 -16
rect -374 -50 -362 -16
rect -420 -84 -362 -50
rect -420 -118 -408 -84
rect -374 -118 -362 -84
rect -420 -152 -362 -118
rect -420 -186 -408 -152
rect -374 -186 -362 -152
rect -420 -220 -362 -186
rect -420 -254 -408 -220
rect -374 -254 -362 -220
rect -420 -288 -362 -254
rect -420 -322 -408 -288
rect -374 -322 -362 -288
rect -420 -356 -362 -322
rect -420 -390 -408 -356
rect -374 -390 -362 -356
rect -420 -424 -362 -390
rect -420 -458 -408 -424
rect -374 -458 -362 -424
rect -420 -492 -362 -458
rect -420 -526 -408 -492
rect -374 -526 -362 -492
rect -420 -560 -362 -526
rect -420 -594 -408 -560
rect -374 -594 -362 -560
rect -420 -624 -362 -594
rect -322 596 -264 626
rect -322 562 -310 596
rect -276 562 -264 596
rect -322 528 -264 562
rect -322 494 -310 528
rect -276 494 -264 528
rect -322 460 -264 494
rect -322 426 -310 460
rect -276 426 -264 460
rect -322 392 -264 426
rect -322 358 -310 392
rect -276 358 -264 392
rect -322 324 -264 358
rect -322 290 -310 324
rect -276 290 -264 324
rect -322 256 -264 290
rect -322 222 -310 256
rect -276 222 -264 256
rect -322 188 -264 222
rect -322 154 -310 188
rect -276 154 -264 188
rect -322 120 -264 154
rect -322 86 -310 120
rect -276 86 -264 120
rect -322 52 -264 86
rect -322 18 -310 52
rect -276 18 -264 52
rect -322 -16 -264 18
rect -322 -50 -310 -16
rect -276 -50 -264 -16
rect -322 -84 -264 -50
rect -322 -118 -310 -84
rect -276 -118 -264 -84
rect -322 -152 -264 -118
rect -322 -186 -310 -152
rect -276 -186 -264 -152
rect -322 -220 -264 -186
rect -322 -254 -310 -220
rect -276 -254 -264 -220
rect -322 -288 -264 -254
rect -322 -322 -310 -288
rect -276 -322 -264 -288
rect -322 -356 -264 -322
rect -322 -390 -310 -356
rect -276 -390 -264 -356
rect -322 -424 -264 -390
rect -322 -458 -310 -424
rect -276 -458 -264 -424
rect -322 -492 -264 -458
rect -322 -526 -310 -492
rect -276 -526 -264 -492
rect -322 -560 -264 -526
rect -322 -594 -310 -560
rect -276 -594 -264 -560
rect -322 -624 -264 -594
rect -224 596 -166 626
rect -224 562 -212 596
rect -178 562 -166 596
rect -224 528 -166 562
rect -224 494 -212 528
rect -178 494 -166 528
rect -224 460 -166 494
rect -224 426 -212 460
rect -178 426 -166 460
rect -224 392 -166 426
rect -224 358 -212 392
rect -178 358 -166 392
rect -224 324 -166 358
rect -224 290 -212 324
rect -178 290 -166 324
rect -224 256 -166 290
rect -224 222 -212 256
rect -178 222 -166 256
rect -224 188 -166 222
rect -224 154 -212 188
rect -178 154 -166 188
rect -224 120 -166 154
rect -224 86 -212 120
rect -178 86 -166 120
rect -224 52 -166 86
rect -224 18 -212 52
rect -178 18 -166 52
rect -224 -16 -166 18
rect -224 -50 -212 -16
rect -178 -50 -166 -16
rect -224 -84 -166 -50
rect -224 -118 -212 -84
rect -178 -118 -166 -84
rect -224 -152 -166 -118
rect -224 -186 -212 -152
rect -178 -186 -166 -152
rect -224 -220 -166 -186
rect -224 -254 -212 -220
rect -178 -254 -166 -220
rect -224 -288 -166 -254
rect -224 -322 -212 -288
rect -178 -322 -166 -288
rect -224 -356 -166 -322
rect -224 -390 -212 -356
rect -178 -390 -166 -356
rect -224 -424 -166 -390
rect -224 -458 -212 -424
rect -178 -458 -166 -424
rect -224 -492 -166 -458
rect -224 -526 -212 -492
rect -178 -526 -166 -492
rect -224 -560 -166 -526
rect -224 -594 -212 -560
rect -178 -594 -166 -560
rect -224 -624 -166 -594
rect -126 596 -68 626
rect -126 562 -114 596
rect -80 562 -68 596
rect -126 528 -68 562
rect -126 494 -114 528
rect -80 494 -68 528
rect -126 460 -68 494
rect -126 426 -114 460
rect -80 426 -68 460
rect -126 392 -68 426
rect -126 358 -114 392
rect -80 358 -68 392
rect -126 324 -68 358
rect -126 290 -114 324
rect -80 290 -68 324
rect -126 256 -68 290
rect -126 222 -114 256
rect -80 222 -68 256
rect -126 188 -68 222
rect -126 154 -114 188
rect -80 154 -68 188
rect -126 120 -68 154
rect -126 86 -114 120
rect -80 86 -68 120
rect -126 52 -68 86
rect -126 18 -114 52
rect -80 18 -68 52
rect -126 -16 -68 18
rect -126 -50 -114 -16
rect -80 -50 -68 -16
rect -126 -84 -68 -50
rect -126 -118 -114 -84
rect -80 -118 -68 -84
rect -126 -152 -68 -118
rect -126 -186 -114 -152
rect -80 -186 -68 -152
rect -126 -220 -68 -186
rect -126 -254 -114 -220
rect -80 -254 -68 -220
rect -126 -288 -68 -254
rect -126 -322 -114 -288
rect -80 -322 -68 -288
rect -126 -356 -68 -322
rect -126 -390 -114 -356
rect -80 -390 -68 -356
rect -126 -424 -68 -390
rect -126 -458 -114 -424
rect -80 -458 -68 -424
rect -126 -492 -68 -458
rect -126 -526 -114 -492
rect -80 -526 -68 -492
rect -126 -560 -68 -526
rect -126 -594 -114 -560
rect -80 -594 -68 -560
rect -126 -624 -68 -594
rect -28 596 30 626
rect -28 562 -16 596
rect 18 562 30 596
rect -28 528 30 562
rect -28 494 -16 528
rect 18 494 30 528
rect -28 460 30 494
rect -28 426 -16 460
rect 18 426 30 460
rect -28 392 30 426
rect -28 358 -16 392
rect 18 358 30 392
rect -28 324 30 358
rect -28 290 -16 324
rect 18 290 30 324
rect -28 256 30 290
rect -28 222 -16 256
rect 18 222 30 256
rect -28 188 30 222
rect -28 154 -16 188
rect 18 154 30 188
rect -28 120 30 154
rect -28 86 -16 120
rect 18 86 30 120
rect -28 52 30 86
rect -28 18 -16 52
rect 18 18 30 52
rect -28 -16 30 18
rect -28 -50 -16 -16
rect 18 -50 30 -16
rect -28 -84 30 -50
rect -28 -118 -16 -84
rect 18 -118 30 -84
rect -28 -152 30 -118
rect -28 -186 -16 -152
rect 18 -186 30 -152
rect -28 -220 30 -186
rect -28 -254 -16 -220
rect 18 -254 30 -220
rect -28 -288 30 -254
rect -28 -322 -16 -288
rect 18 -322 30 -288
rect -28 -356 30 -322
rect -28 -390 -16 -356
rect 18 -390 30 -356
rect -28 -424 30 -390
rect -28 -458 -16 -424
rect 18 -458 30 -424
rect -28 -492 30 -458
rect -28 -526 -16 -492
rect 18 -526 30 -492
rect -28 -560 30 -526
rect -28 -594 -16 -560
rect 18 -594 30 -560
rect -28 -624 30 -594
rect 70 596 128 626
rect 70 562 82 596
rect 116 562 128 596
rect 70 528 128 562
rect 70 494 82 528
rect 116 494 128 528
rect 70 460 128 494
rect 70 426 82 460
rect 116 426 128 460
rect 70 392 128 426
rect 70 358 82 392
rect 116 358 128 392
rect 70 324 128 358
rect 70 290 82 324
rect 116 290 128 324
rect 70 256 128 290
rect 70 222 82 256
rect 116 222 128 256
rect 70 188 128 222
rect 70 154 82 188
rect 116 154 128 188
rect 70 120 128 154
rect 70 86 82 120
rect 116 86 128 120
rect 70 52 128 86
rect 70 18 82 52
rect 116 18 128 52
rect 70 -16 128 18
rect 70 -50 82 -16
rect 116 -50 128 -16
rect 70 -84 128 -50
rect 70 -118 82 -84
rect 116 -118 128 -84
rect 70 -152 128 -118
rect 70 -186 82 -152
rect 116 -186 128 -152
rect 70 -220 128 -186
rect 70 -254 82 -220
rect 116 -254 128 -220
rect 70 -288 128 -254
rect 70 -322 82 -288
rect 116 -322 128 -288
rect 70 -356 128 -322
rect 70 -390 82 -356
rect 116 -390 128 -356
rect 70 -424 128 -390
rect 70 -458 82 -424
rect 116 -458 128 -424
rect 70 -492 128 -458
rect 70 -526 82 -492
rect 116 -526 128 -492
rect 70 -560 128 -526
rect 70 -594 82 -560
rect 116 -594 128 -560
rect 70 -624 128 -594
rect 168 596 226 626
rect 168 562 180 596
rect 214 562 226 596
rect 168 528 226 562
rect 168 494 180 528
rect 214 494 226 528
rect 168 460 226 494
rect 168 426 180 460
rect 214 426 226 460
rect 168 392 226 426
rect 168 358 180 392
rect 214 358 226 392
rect 168 324 226 358
rect 168 290 180 324
rect 214 290 226 324
rect 168 256 226 290
rect 168 222 180 256
rect 214 222 226 256
rect 168 188 226 222
rect 168 154 180 188
rect 214 154 226 188
rect 168 120 226 154
rect 168 86 180 120
rect 214 86 226 120
rect 168 52 226 86
rect 168 18 180 52
rect 214 18 226 52
rect 168 -16 226 18
rect 168 -50 180 -16
rect 214 -50 226 -16
rect 168 -84 226 -50
rect 168 -118 180 -84
rect 214 -118 226 -84
rect 168 -152 226 -118
rect 168 -186 180 -152
rect 214 -186 226 -152
rect 168 -220 226 -186
rect 168 -254 180 -220
rect 214 -254 226 -220
rect 168 -288 226 -254
rect 168 -322 180 -288
rect 214 -322 226 -288
rect 168 -356 226 -322
rect 168 -390 180 -356
rect 214 -390 226 -356
rect 168 -424 226 -390
rect 168 -458 180 -424
rect 214 -458 226 -424
rect 168 -492 226 -458
rect 168 -526 180 -492
rect 214 -526 226 -492
rect 168 -560 226 -526
rect 168 -594 180 -560
rect 214 -594 226 -560
rect 168 -624 226 -594
rect 266 596 324 626
rect 266 562 278 596
rect 312 562 324 596
rect 266 528 324 562
rect 266 494 278 528
rect 312 494 324 528
rect 266 460 324 494
rect 266 426 278 460
rect 312 426 324 460
rect 266 392 324 426
rect 266 358 278 392
rect 312 358 324 392
rect 266 324 324 358
rect 266 290 278 324
rect 312 290 324 324
rect 266 256 324 290
rect 266 222 278 256
rect 312 222 324 256
rect 266 188 324 222
rect 266 154 278 188
rect 312 154 324 188
rect 266 120 324 154
rect 266 86 278 120
rect 312 86 324 120
rect 266 52 324 86
rect 266 18 278 52
rect 312 18 324 52
rect 266 -16 324 18
rect 266 -50 278 -16
rect 312 -50 324 -16
rect 266 -84 324 -50
rect 266 -118 278 -84
rect 312 -118 324 -84
rect 266 -152 324 -118
rect 266 -186 278 -152
rect 312 -186 324 -152
rect 266 -220 324 -186
rect 266 -254 278 -220
rect 312 -254 324 -220
rect 266 -288 324 -254
rect 266 -322 278 -288
rect 312 -322 324 -288
rect 266 -356 324 -322
rect 266 -390 278 -356
rect 312 -390 324 -356
rect 266 -424 324 -390
rect 266 -458 278 -424
rect 312 -458 324 -424
rect 266 -492 324 -458
rect 266 -526 278 -492
rect 312 -526 324 -492
rect 266 -560 324 -526
rect 266 -594 278 -560
rect 312 -594 324 -560
rect 266 -624 324 -594
rect 364 596 422 626
rect 364 562 376 596
rect 410 562 422 596
rect 364 528 422 562
rect 364 494 376 528
rect 410 494 422 528
rect 364 460 422 494
rect 364 426 376 460
rect 410 426 422 460
rect 364 392 422 426
rect 364 358 376 392
rect 410 358 422 392
rect 364 324 422 358
rect 364 290 376 324
rect 410 290 422 324
rect 364 256 422 290
rect 364 222 376 256
rect 410 222 422 256
rect 364 188 422 222
rect 364 154 376 188
rect 410 154 422 188
rect 364 120 422 154
rect 364 86 376 120
rect 410 86 422 120
rect 364 52 422 86
rect 364 18 376 52
rect 410 18 422 52
rect 364 -16 422 18
rect 364 -50 376 -16
rect 410 -50 422 -16
rect 364 -84 422 -50
rect 364 -118 376 -84
rect 410 -118 422 -84
rect 364 -152 422 -118
rect 364 -186 376 -152
rect 410 -186 422 -152
rect 364 -220 422 -186
rect 364 -254 376 -220
rect 410 -254 422 -220
rect 364 -288 422 -254
rect 364 -322 376 -288
rect 410 -322 422 -288
rect 364 -356 422 -322
rect 364 -390 376 -356
rect 410 -390 422 -356
rect 364 -424 422 -390
rect 364 -458 376 -424
rect 410 -458 422 -424
rect 364 -492 422 -458
rect 364 -526 376 -492
rect 410 -526 422 -492
rect 364 -560 422 -526
rect 364 -594 376 -560
rect 410 -594 422 -560
rect 364 -624 422 -594
rect 462 596 520 626
rect 462 562 474 596
rect 508 562 520 596
rect 462 528 520 562
rect 462 494 474 528
rect 508 494 520 528
rect 462 460 520 494
rect 462 426 474 460
rect 508 426 520 460
rect 462 392 520 426
rect 462 358 474 392
rect 508 358 520 392
rect 462 324 520 358
rect 462 290 474 324
rect 508 290 520 324
rect 462 256 520 290
rect 462 222 474 256
rect 508 222 520 256
rect 462 188 520 222
rect 462 154 474 188
rect 508 154 520 188
rect 462 120 520 154
rect 462 86 474 120
rect 508 86 520 120
rect 462 52 520 86
rect 462 18 474 52
rect 508 18 520 52
rect 462 -16 520 18
rect 462 -50 474 -16
rect 508 -50 520 -16
rect 462 -84 520 -50
rect 462 -118 474 -84
rect 508 -118 520 -84
rect 462 -152 520 -118
rect 462 -186 474 -152
rect 508 -186 520 -152
rect 462 -220 520 -186
rect 462 -254 474 -220
rect 508 -254 520 -220
rect 462 -288 520 -254
rect 462 -322 474 -288
rect 508 -322 520 -288
rect 462 -356 520 -322
rect 462 -390 474 -356
rect 508 -390 520 -356
rect 462 -424 520 -390
rect 462 -458 474 -424
rect 508 -458 520 -424
rect 462 -492 520 -458
rect 462 -526 474 -492
rect 508 -526 520 -492
rect 462 -560 520 -526
rect 462 -594 474 -560
rect 508 -594 520 -560
rect 462 -624 520 -594
rect 560 596 618 626
rect 560 562 572 596
rect 606 562 618 596
rect 560 528 618 562
rect 560 494 572 528
rect 606 494 618 528
rect 560 460 618 494
rect 560 426 572 460
rect 606 426 618 460
rect 560 392 618 426
rect 560 358 572 392
rect 606 358 618 392
rect 560 324 618 358
rect 560 290 572 324
rect 606 290 618 324
rect 560 256 618 290
rect 560 222 572 256
rect 606 222 618 256
rect 560 188 618 222
rect 560 154 572 188
rect 606 154 618 188
rect 560 120 618 154
rect 560 86 572 120
rect 606 86 618 120
rect 560 52 618 86
rect 560 18 572 52
rect 606 18 618 52
rect 560 -16 618 18
rect 560 -50 572 -16
rect 606 -50 618 -16
rect 560 -84 618 -50
rect 560 -118 572 -84
rect 606 -118 618 -84
rect 560 -152 618 -118
rect 560 -186 572 -152
rect 606 -186 618 -152
rect 560 -220 618 -186
rect 560 -254 572 -220
rect 606 -254 618 -220
rect 560 -288 618 -254
rect 560 -322 572 -288
rect 606 -322 618 -288
rect 560 -356 618 -322
rect 560 -390 572 -356
rect 606 -390 618 -356
rect 560 -424 618 -390
rect 560 -458 572 -424
rect 606 -458 618 -424
rect 560 -492 618 -458
rect 560 -526 572 -492
rect 606 -526 618 -492
rect 560 -560 618 -526
rect 560 -594 572 -560
rect 606 -594 618 -560
rect 560 -624 618 -594
rect 658 596 716 626
rect 658 562 670 596
rect 704 562 716 596
rect 658 528 716 562
rect 658 494 670 528
rect 704 494 716 528
rect 658 460 716 494
rect 658 426 670 460
rect 704 426 716 460
rect 658 392 716 426
rect 658 358 670 392
rect 704 358 716 392
rect 658 324 716 358
rect 658 290 670 324
rect 704 290 716 324
rect 658 256 716 290
rect 658 222 670 256
rect 704 222 716 256
rect 658 188 716 222
rect 658 154 670 188
rect 704 154 716 188
rect 658 120 716 154
rect 658 86 670 120
rect 704 86 716 120
rect 658 52 716 86
rect 658 18 670 52
rect 704 18 716 52
rect 658 -16 716 18
rect 658 -50 670 -16
rect 704 -50 716 -16
rect 658 -84 716 -50
rect 658 -118 670 -84
rect 704 -118 716 -84
rect 658 -152 716 -118
rect 658 -186 670 -152
rect 704 -186 716 -152
rect 658 -220 716 -186
rect 658 -254 670 -220
rect 704 -254 716 -220
rect 658 -288 716 -254
rect 658 -322 670 -288
rect 704 -322 716 -288
rect 658 -356 716 -322
rect 658 -390 670 -356
rect 704 -390 716 -356
rect 658 -424 716 -390
rect 658 -458 670 -424
rect 704 -458 716 -424
rect 658 -492 716 -458
rect 658 -526 670 -492
rect 704 -526 716 -492
rect 658 -560 716 -526
rect 658 -594 670 -560
rect 704 -594 716 -560
rect 658 -624 716 -594
rect 756 596 814 626
rect 756 562 768 596
rect 802 562 814 596
rect 756 528 814 562
rect 756 494 768 528
rect 802 494 814 528
rect 756 460 814 494
rect 756 426 768 460
rect 802 426 814 460
rect 756 392 814 426
rect 756 358 768 392
rect 802 358 814 392
rect 756 324 814 358
rect 756 290 768 324
rect 802 290 814 324
rect 756 256 814 290
rect 756 222 768 256
rect 802 222 814 256
rect 756 188 814 222
rect 756 154 768 188
rect 802 154 814 188
rect 756 120 814 154
rect 756 86 768 120
rect 802 86 814 120
rect 756 52 814 86
rect 756 18 768 52
rect 802 18 814 52
rect 756 -16 814 18
rect 756 -50 768 -16
rect 802 -50 814 -16
rect 756 -84 814 -50
rect 756 -118 768 -84
rect 802 -118 814 -84
rect 756 -152 814 -118
rect 756 -186 768 -152
rect 802 -186 814 -152
rect 756 -220 814 -186
rect 756 -254 768 -220
rect 802 -254 814 -220
rect 756 -288 814 -254
rect 756 -322 768 -288
rect 802 -322 814 -288
rect 756 -356 814 -322
rect 756 -390 768 -356
rect 802 -390 814 -356
rect 756 -424 814 -390
rect 756 -458 768 -424
rect 802 -458 814 -424
rect 756 -492 814 -458
rect 756 -526 768 -492
rect 802 -526 814 -492
rect 756 -560 814 -526
rect 756 -594 768 -560
rect 802 -594 814 -560
rect 756 -624 814 -594
<< pdiffc >>
rect -800 562 -766 596
rect -800 494 -766 528
rect -800 426 -766 460
rect -800 358 -766 392
rect -800 290 -766 324
rect -800 222 -766 256
rect -800 154 -766 188
rect -800 86 -766 120
rect -800 18 -766 52
rect -800 -50 -766 -16
rect -800 -118 -766 -84
rect -800 -186 -766 -152
rect -800 -254 -766 -220
rect -800 -322 -766 -288
rect -800 -390 -766 -356
rect -800 -458 -766 -424
rect -800 -526 -766 -492
rect -800 -594 -766 -560
rect -702 562 -668 596
rect -702 494 -668 528
rect -702 426 -668 460
rect -702 358 -668 392
rect -702 290 -668 324
rect -702 222 -668 256
rect -702 154 -668 188
rect -702 86 -668 120
rect -702 18 -668 52
rect -702 -50 -668 -16
rect -702 -118 -668 -84
rect -702 -186 -668 -152
rect -702 -254 -668 -220
rect -702 -322 -668 -288
rect -702 -390 -668 -356
rect -702 -458 -668 -424
rect -702 -526 -668 -492
rect -702 -594 -668 -560
rect -604 562 -570 596
rect -604 494 -570 528
rect -604 426 -570 460
rect -604 358 -570 392
rect -604 290 -570 324
rect -604 222 -570 256
rect -604 154 -570 188
rect -604 86 -570 120
rect -604 18 -570 52
rect -604 -50 -570 -16
rect -604 -118 -570 -84
rect -604 -186 -570 -152
rect -604 -254 -570 -220
rect -604 -322 -570 -288
rect -604 -390 -570 -356
rect -604 -458 -570 -424
rect -604 -526 -570 -492
rect -604 -594 -570 -560
rect -506 562 -472 596
rect -506 494 -472 528
rect -506 426 -472 460
rect -506 358 -472 392
rect -506 290 -472 324
rect -506 222 -472 256
rect -506 154 -472 188
rect -506 86 -472 120
rect -506 18 -472 52
rect -506 -50 -472 -16
rect -506 -118 -472 -84
rect -506 -186 -472 -152
rect -506 -254 -472 -220
rect -506 -322 -472 -288
rect -506 -390 -472 -356
rect -506 -458 -472 -424
rect -506 -526 -472 -492
rect -506 -594 -472 -560
rect -408 562 -374 596
rect -408 494 -374 528
rect -408 426 -374 460
rect -408 358 -374 392
rect -408 290 -374 324
rect -408 222 -374 256
rect -408 154 -374 188
rect -408 86 -374 120
rect -408 18 -374 52
rect -408 -50 -374 -16
rect -408 -118 -374 -84
rect -408 -186 -374 -152
rect -408 -254 -374 -220
rect -408 -322 -374 -288
rect -408 -390 -374 -356
rect -408 -458 -374 -424
rect -408 -526 -374 -492
rect -408 -594 -374 -560
rect -310 562 -276 596
rect -310 494 -276 528
rect -310 426 -276 460
rect -310 358 -276 392
rect -310 290 -276 324
rect -310 222 -276 256
rect -310 154 -276 188
rect -310 86 -276 120
rect -310 18 -276 52
rect -310 -50 -276 -16
rect -310 -118 -276 -84
rect -310 -186 -276 -152
rect -310 -254 -276 -220
rect -310 -322 -276 -288
rect -310 -390 -276 -356
rect -310 -458 -276 -424
rect -310 -526 -276 -492
rect -310 -594 -276 -560
rect -212 562 -178 596
rect -212 494 -178 528
rect -212 426 -178 460
rect -212 358 -178 392
rect -212 290 -178 324
rect -212 222 -178 256
rect -212 154 -178 188
rect -212 86 -178 120
rect -212 18 -178 52
rect -212 -50 -178 -16
rect -212 -118 -178 -84
rect -212 -186 -178 -152
rect -212 -254 -178 -220
rect -212 -322 -178 -288
rect -212 -390 -178 -356
rect -212 -458 -178 -424
rect -212 -526 -178 -492
rect -212 -594 -178 -560
rect -114 562 -80 596
rect -114 494 -80 528
rect -114 426 -80 460
rect -114 358 -80 392
rect -114 290 -80 324
rect -114 222 -80 256
rect -114 154 -80 188
rect -114 86 -80 120
rect -114 18 -80 52
rect -114 -50 -80 -16
rect -114 -118 -80 -84
rect -114 -186 -80 -152
rect -114 -254 -80 -220
rect -114 -322 -80 -288
rect -114 -390 -80 -356
rect -114 -458 -80 -424
rect -114 -526 -80 -492
rect -114 -594 -80 -560
rect -16 562 18 596
rect -16 494 18 528
rect -16 426 18 460
rect -16 358 18 392
rect -16 290 18 324
rect -16 222 18 256
rect -16 154 18 188
rect -16 86 18 120
rect -16 18 18 52
rect -16 -50 18 -16
rect -16 -118 18 -84
rect -16 -186 18 -152
rect -16 -254 18 -220
rect -16 -322 18 -288
rect -16 -390 18 -356
rect -16 -458 18 -424
rect -16 -526 18 -492
rect -16 -594 18 -560
rect 82 562 116 596
rect 82 494 116 528
rect 82 426 116 460
rect 82 358 116 392
rect 82 290 116 324
rect 82 222 116 256
rect 82 154 116 188
rect 82 86 116 120
rect 82 18 116 52
rect 82 -50 116 -16
rect 82 -118 116 -84
rect 82 -186 116 -152
rect 82 -254 116 -220
rect 82 -322 116 -288
rect 82 -390 116 -356
rect 82 -458 116 -424
rect 82 -526 116 -492
rect 82 -594 116 -560
rect 180 562 214 596
rect 180 494 214 528
rect 180 426 214 460
rect 180 358 214 392
rect 180 290 214 324
rect 180 222 214 256
rect 180 154 214 188
rect 180 86 214 120
rect 180 18 214 52
rect 180 -50 214 -16
rect 180 -118 214 -84
rect 180 -186 214 -152
rect 180 -254 214 -220
rect 180 -322 214 -288
rect 180 -390 214 -356
rect 180 -458 214 -424
rect 180 -526 214 -492
rect 180 -594 214 -560
rect 278 562 312 596
rect 278 494 312 528
rect 278 426 312 460
rect 278 358 312 392
rect 278 290 312 324
rect 278 222 312 256
rect 278 154 312 188
rect 278 86 312 120
rect 278 18 312 52
rect 278 -50 312 -16
rect 278 -118 312 -84
rect 278 -186 312 -152
rect 278 -254 312 -220
rect 278 -322 312 -288
rect 278 -390 312 -356
rect 278 -458 312 -424
rect 278 -526 312 -492
rect 278 -594 312 -560
rect 376 562 410 596
rect 376 494 410 528
rect 376 426 410 460
rect 376 358 410 392
rect 376 290 410 324
rect 376 222 410 256
rect 376 154 410 188
rect 376 86 410 120
rect 376 18 410 52
rect 376 -50 410 -16
rect 376 -118 410 -84
rect 376 -186 410 -152
rect 376 -254 410 -220
rect 376 -322 410 -288
rect 376 -390 410 -356
rect 376 -458 410 -424
rect 376 -526 410 -492
rect 376 -594 410 -560
rect 474 562 508 596
rect 474 494 508 528
rect 474 426 508 460
rect 474 358 508 392
rect 474 290 508 324
rect 474 222 508 256
rect 474 154 508 188
rect 474 86 508 120
rect 474 18 508 52
rect 474 -50 508 -16
rect 474 -118 508 -84
rect 474 -186 508 -152
rect 474 -254 508 -220
rect 474 -322 508 -288
rect 474 -390 508 -356
rect 474 -458 508 -424
rect 474 -526 508 -492
rect 474 -594 508 -560
rect 572 562 606 596
rect 572 494 606 528
rect 572 426 606 460
rect 572 358 606 392
rect 572 290 606 324
rect 572 222 606 256
rect 572 154 606 188
rect 572 86 606 120
rect 572 18 606 52
rect 572 -50 606 -16
rect 572 -118 606 -84
rect 572 -186 606 -152
rect 572 -254 606 -220
rect 572 -322 606 -288
rect 572 -390 606 -356
rect 572 -458 606 -424
rect 572 -526 606 -492
rect 572 -594 606 -560
rect 670 562 704 596
rect 670 494 704 528
rect 670 426 704 460
rect 670 358 704 392
rect 670 290 704 324
rect 670 222 704 256
rect 670 154 704 188
rect 670 86 704 120
rect 670 18 704 52
rect 670 -50 704 -16
rect 670 -118 704 -84
rect 670 -186 704 -152
rect 670 -254 704 -220
rect 670 -322 704 -288
rect 670 -390 704 -356
rect 670 -458 704 -424
rect 670 -526 704 -492
rect 670 -594 704 -560
rect 768 562 802 596
rect 768 494 802 528
rect 768 426 802 460
rect 768 358 802 392
rect 768 290 802 324
rect 768 222 802 256
rect 768 154 802 188
rect 768 86 802 120
rect 768 18 802 52
rect 768 -50 802 -16
rect 768 -118 802 -84
rect 768 -186 802 -152
rect 768 -254 802 -220
rect 768 -322 802 -288
rect 768 -390 802 -356
rect 768 -458 802 -424
rect 768 -526 802 -492
rect 768 -594 802 -560
<< poly >>
rect -1088 695 658 732
rect -1088 593 -1049 695
rect -947 694 658 695
rect -947 593 -910 694
rect -1088 556 -910 593
rect -1088 -591 -910 -554
rect -1088 -693 -1049 -591
rect -947 -692 -910 -591
rect -868 -650 -828 652
rect -754 626 -714 652
rect -656 626 -616 694
rect -558 626 -518 694
rect -460 626 -420 652
rect -362 626 -322 652
rect -264 626 -224 694
rect -166 626 -126 694
rect -68 626 -28 652
rect 30 626 70 652
rect 128 626 168 694
rect 226 626 266 694
rect 324 626 364 652
rect 422 626 462 652
rect 520 626 560 694
rect 618 626 658 694
rect 716 626 756 652
rect -754 -692 -714 -624
rect -656 -650 -616 -624
rect -558 -650 -518 -624
rect -460 -692 -420 -624
rect -362 -692 -322 -624
rect -264 -650 -224 -624
rect -166 -650 -126 -624
rect -68 -692 -28 -624
rect 30 -692 70 -624
rect 128 -650 168 -624
rect 226 -650 266 -624
rect 324 -692 364 -624
rect 422 -692 462 -624
rect 520 -650 560 -624
rect 618 -650 658 -624
rect 716 -692 756 -624
rect 830 -650 870 652
rect -947 -693 756 -692
rect -1088 -730 756 -693
<< polycont >>
rect -1049 593 -947 695
rect -1049 -693 -947 -591
<< locali >>
rect -1088 697 -910 732
rect -1088 591 -1051 697
rect -945 591 -910 697
rect -1088 556 -910 591
rect -800 596 -766 630
rect -800 528 -766 560
rect -800 460 -766 488
rect -800 392 -766 416
rect -800 324 -766 344
rect -800 256 -766 272
rect -800 188 -766 200
rect -800 120 -766 128
rect -800 52 -766 56
rect -800 -54 -766 -50
rect -800 -126 -766 -118
rect -800 -198 -766 -186
rect -800 -270 -766 -254
rect -800 -342 -766 -322
rect -800 -414 -766 -390
rect -800 -486 -766 -458
rect -1088 -589 -910 -554
rect -1088 -695 -1051 -589
rect -945 -695 -910 -589
rect -800 -558 -766 -526
rect -800 -628 -766 -594
rect -702 596 -668 630
rect -702 528 -668 560
rect -702 460 -668 488
rect -702 392 -668 416
rect -702 324 -668 344
rect -702 256 -668 272
rect -702 188 -668 200
rect -702 120 -668 128
rect -702 52 -668 56
rect -702 -54 -668 -50
rect -702 -126 -668 -118
rect -702 -198 -668 -186
rect -702 -270 -668 -254
rect -702 -342 -668 -322
rect -702 -414 -668 -390
rect -702 -486 -668 -458
rect -702 -558 -668 -526
rect -702 -628 -668 -594
rect -604 596 -570 630
rect -604 528 -570 560
rect -604 460 -570 488
rect -604 392 -570 416
rect -604 324 -570 344
rect -604 256 -570 272
rect -604 188 -570 200
rect -604 120 -570 128
rect -604 52 -570 56
rect -604 -54 -570 -50
rect -604 -126 -570 -118
rect -604 -198 -570 -186
rect -604 -270 -570 -254
rect -604 -342 -570 -322
rect -604 -414 -570 -390
rect -604 -486 -570 -458
rect -604 -558 -570 -526
rect -604 -628 -570 -594
rect -506 596 -472 630
rect -506 528 -472 560
rect -506 460 -472 488
rect -506 392 -472 416
rect -506 324 -472 344
rect -506 256 -472 272
rect -506 188 -472 200
rect -506 120 -472 128
rect -506 52 -472 56
rect -506 -54 -472 -50
rect -506 -126 -472 -118
rect -506 -198 -472 -186
rect -506 -270 -472 -254
rect -506 -342 -472 -322
rect -506 -414 -472 -390
rect -506 -486 -472 -458
rect -506 -558 -472 -526
rect -506 -628 -472 -594
rect -408 596 -374 630
rect -408 528 -374 560
rect -408 460 -374 488
rect -408 392 -374 416
rect -408 324 -374 344
rect -408 256 -374 272
rect -408 188 -374 200
rect -408 120 -374 128
rect -408 52 -374 56
rect -408 -54 -374 -50
rect -408 -126 -374 -118
rect -408 -198 -374 -186
rect -408 -270 -374 -254
rect -408 -342 -374 -322
rect -408 -414 -374 -390
rect -408 -486 -374 -458
rect -408 -558 -374 -526
rect -408 -628 -374 -594
rect -310 596 -276 630
rect -310 528 -276 560
rect -310 460 -276 488
rect -310 392 -276 416
rect -310 324 -276 344
rect -310 256 -276 272
rect -310 188 -276 200
rect -310 120 -276 128
rect -310 52 -276 56
rect -310 -54 -276 -50
rect -310 -126 -276 -118
rect -310 -198 -276 -186
rect -310 -270 -276 -254
rect -310 -342 -276 -322
rect -310 -414 -276 -390
rect -310 -486 -276 -458
rect -310 -558 -276 -526
rect -310 -628 -276 -594
rect -212 596 -178 630
rect -212 528 -178 560
rect -212 460 -178 488
rect -212 392 -178 416
rect -212 324 -178 344
rect -212 256 -178 272
rect -212 188 -178 200
rect -212 120 -178 128
rect -212 52 -178 56
rect -212 -54 -178 -50
rect -212 -126 -178 -118
rect -212 -198 -178 -186
rect -212 -270 -178 -254
rect -212 -342 -178 -322
rect -212 -414 -178 -390
rect -212 -486 -178 -458
rect -212 -558 -178 -526
rect -212 -628 -178 -594
rect -114 596 -80 630
rect -114 528 -80 560
rect -114 460 -80 488
rect -114 392 -80 416
rect -114 324 -80 344
rect -114 256 -80 272
rect -114 188 -80 200
rect -114 120 -80 128
rect -114 52 -80 56
rect -114 -54 -80 -50
rect -114 -126 -80 -118
rect -114 -198 -80 -186
rect -114 -270 -80 -254
rect -114 -342 -80 -322
rect -114 -414 -80 -390
rect -114 -486 -80 -458
rect -114 -558 -80 -526
rect -114 -628 -80 -594
rect -16 596 18 630
rect -16 528 18 560
rect -16 460 18 488
rect -16 392 18 416
rect -16 324 18 344
rect -16 256 18 272
rect -16 188 18 200
rect -16 120 18 128
rect -16 52 18 56
rect -16 -54 18 -50
rect -16 -126 18 -118
rect -16 -198 18 -186
rect -16 -270 18 -254
rect -16 -342 18 -322
rect -16 -414 18 -390
rect -16 -486 18 -458
rect -16 -558 18 -526
rect -16 -628 18 -594
rect 82 596 116 630
rect 82 528 116 560
rect 82 460 116 488
rect 82 392 116 416
rect 82 324 116 344
rect 82 256 116 272
rect 82 188 116 200
rect 82 120 116 128
rect 82 52 116 56
rect 82 -54 116 -50
rect 82 -126 116 -118
rect 82 -198 116 -186
rect 82 -270 116 -254
rect 82 -342 116 -322
rect 82 -414 116 -390
rect 82 -486 116 -458
rect 82 -558 116 -526
rect 82 -628 116 -594
rect 180 596 214 630
rect 180 528 214 560
rect 180 460 214 488
rect 180 392 214 416
rect 180 324 214 344
rect 180 256 214 272
rect 180 188 214 200
rect 180 120 214 128
rect 180 52 214 56
rect 180 -54 214 -50
rect 180 -126 214 -118
rect 180 -198 214 -186
rect 180 -270 214 -254
rect 180 -342 214 -322
rect 180 -414 214 -390
rect 180 -486 214 -458
rect 180 -558 214 -526
rect 180 -628 214 -594
rect 278 596 312 630
rect 278 528 312 560
rect 278 460 312 488
rect 278 392 312 416
rect 278 324 312 344
rect 278 256 312 272
rect 278 188 312 200
rect 278 120 312 128
rect 278 52 312 56
rect 278 -54 312 -50
rect 278 -126 312 -118
rect 278 -198 312 -186
rect 278 -270 312 -254
rect 278 -342 312 -322
rect 278 -414 312 -390
rect 278 -486 312 -458
rect 278 -558 312 -526
rect 278 -628 312 -594
rect 376 596 410 630
rect 376 528 410 560
rect 376 460 410 488
rect 376 392 410 416
rect 376 324 410 344
rect 376 256 410 272
rect 376 188 410 200
rect 376 120 410 128
rect 376 52 410 56
rect 376 -54 410 -50
rect 376 -126 410 -118
rect 376 -198 410 -186
rect 376 -270 410 -254
rect 376 -342 410 -322
rect 376 -414 410 -390
rect 376 -486 410 -458
rect 376 -558 410 -526
rect 376 -628 410 -594
rect 474 596 508 630
rect 474 528 508 560
rect 474 460 508 488
rect 474 392 508 416
rect 474 324 508 344
rect 474 256 508 272
rect 474 188 508 200
rect 474 120 508 128
rect 474 52 508 56
rect 474 -54 508 -50
rect 474 -126 508 -118
rect 474 -198 508 -186
rect 474 -270 508 -254
rect 474 -342 508 -322
rect 474 -414 508 -390
rect 474 -486 508 -458
rect 474 -558 508 -526
rect 474 -628 508 -594
rect 572 596 606 630
rect 572 528 606 560
rect 572 460 606 488
rect 572 392 606 416
rect 572 324 606 344
rect 572 256 606 272
rect 572 188 606 200
rect 572 120 606 128
rect 572 52 606 56
rect 572 -54 606 -50
rect 572 -126 606 -118
rect 572 -198 606 -186
rect 572 -270 606 -254
rect 572 -342 606 -322
rect 572 -414 606 -390
rect 572 -486 606 -458
rect 572 -558 606 -526
rect 572 -628 606 -594
rect 670 596 704 630
rect 670 528 704 560
rect 670 460 704 488
rect 670 392 704 416
rect 670 324 704 344
rect 670 256 704 272
rect 670 188 704 200
rect 670 120 704 128
rect 670 52 704 56
rect 670 -54 704 -50
rect 670 -126 704 -118
rect 670 -198 704 -186
rect 670 -270 704 -254
rect 670 -342 704 -322
rect 670 -414 704 -390
rect 670 -486 704 -458
rect 670 -558 704 -526
rect 670 -628 704 -594
rect 768 596 802 630
rect 768 528 802 560
rect 768 460 802 488
rect 768 392 802 416
rect 768 324 802 344
rect 768 256 802 272
rect 768 188 802 200
rect 768 120 802 128
rect 768 52 802 56
rect 768 -54 802 -50
rect 768 -126 802 -118
rect 768 -198 802 -186
rect 768 -270 802 -254
rect 768 -342 802 -322
rect 768 -414 802 -390
rect 768 -486 802 -458
rect 768 -558 802 -526
rect 768 -628 802 -594
rect -1088 -730 -910 -695
<< viali >>
rect -1051 695 -945 697
rect -1051 593 -1049 695
rect -1049 593 -947 695
rect -947 593 -945 695
rect -1051 591 -945 593
rect -800 562 -766 594
rect -800 560 -766 562
rect -800 494 -766 522
rect -800 488 -766 494
rect -800 426 -766 450
rect -800 416 -766 426
rect -800 358 -766 378
rect -800 344 -766 358
rect -800 290 -766 306
rect -800 272 -766 290
rect -800 222 -766 234
rect -800 200 -766 222
rect -800 154 -766 162
rect -800 128 -766 154
rect -800 86 -766 90
rect -800 56 -766 86
rect -800 -16 -766 18
rect -800 -84 -766 -54
rect -800 -88 -766 -84
rect -800 -152 -766 -126
rect -800 -160 -766 -152
rect -800 -220 -766 -198
rect -800 -232 -766 -220
rect -800 -288 -766 -270
rect -800 -304 -766 -288
rect -800 -356 -766 -342
rect -800 -376 -766 -356
rect -800 -424 -766 -414
rect -800 -448 -766 -424
rect -800 -492 -766 -486
rect -800 -520 -766 -492
rect -1051 -591 -945 -589
rect -1051 -693 -1049 -591
rect -1049 -693 -947 -591
rect -947 -693 -945 -591
rect -1051 -695 -945 -693
rect -800 -560 -766 -558
rect -800 -592 -766 -560
rect -702 562 -668 594
rect -702 560 -668 562
rect -702 494 -668 522
rect -702 488 -668 494
rect -702 426 -668 450
rect -702 416 -668 426
rect -702 358 -668 378
rect -702 344 -668 358
rect -702 290 -668 306
rect -702 272 -668 290
rect -702 222 -668 234
rect -702 200 -668 222
rect -702 154 -668 162
rect -702 128 -668 154
rect -702 86 -668 90
rect -702 56 -668 86
rect -702 -16 -668 18
rect -702 -84 -668 -54
rect -702 -88 -668 -84
rect -702 -152 -668 -126
rect -702 -160 -668 -152
rect -702 -220 -668 -198
rect -702 -232 -668 -220
rect -702 -288 -668 -270
rect -702 -304 -668 -288
rect -702 -356 -668 -342
rect -702 -376 -668 -356
rect -702 -424 -668 -414
rect -702 -448 -668 -424
rect -702 -492 -668 -486
rect -702 -520 -668 -492
rect -702 -560 -668 -558
rect -702 -592 -668 -560
rect -604 562 -570 594
rect -604 560 -570 562
rect -604 494 -570 522
rect -604 488 -570 494
rect -604 426 -570 450
rect -604 416 -570 426
rect -604 358 -570 378
rect -604 344 -570 358
rect -604 290 -570 306
rect -604 272 -570 290
rect -604 222 -570 234
rect -604 200 -570 222
rect -604 154 -570 162
rect -604 128 -570 154
rect -604 86 -570 90
rect -604 56 -570 86
rect -604 -16 -570 18
rect -604 -84 -570 -54
rect -604 -88 -570 -84
rect -604 -152 -570 -126
rect -604 -160 -570 -152
rect -604 -220 -570 -198
rect -604 -232 -570 -220
rect -604 -288 -570 -270
rect -604 -304 -570 -288
rect -604 -356 -570 -342
rect -604 -376 -570 -356
rect -604 -424 -570 -414
rect -604 -448 -570 -424
rect -604 -492 -570 -486
rect -604 -520 -570 -492
rect -604 -560 -570 -558
rect -604 -592 -570 -560
rect -506 562 -472 594
rect -506 560 -472 562
rect -506 494 -472 522
rect -506 488 -472 494
rect -506 426 -472 450
rect -506 416 -472 426
rect -506 358 -472 378
rect -506 344 -472 358
rect -506 290 -472 306
rect -506 272 -472 290
rect -506 222 -472 234
rect -506 200 -472 222
rect -506 154 -472 162
rect -506 128 -472 154
rect -506 86 -472 90
rect -506 56 -472 86
rect -506 -16 -472 18
rect -506 -84 -472 -54
rect -506 -88 -472 -84
rect -506 -152 -472 -126
rect -506 -160 -472 -152
rect -506 -220 -472 -198
rect -506 -232 -472 -220
rect -506 -288 -472 -270
rect -506 -304 -472 -288
rect -506 -356 -472 -342
rect -506 -376 -472 -356
rect -506 -424 -472 -414
rect -506 -448 -472 -424
rect -506 -492 -472 -486
rect -506 -520 -472 -492
rect -506 -560 -472 -558
rect -506 -592 -472 -560
rect -408 562 -374 594
rect -408 560 -374 562
rect -408 494 -374 522
rect -408 488 -374 494
rect -408 426 -374 450
rect -408 416 -374 426
rect -408 358 -374 378
rect -408 344 -374 358
rect -408 290 -374 306
rect -408 272 -374 290
rect -408 222 -374 234
rect -408 200 -374 222
rect -408 154 -374 162
rect -408 128 -374 154
rect -408 86 -374 90
rect -408 56 -374 86
rect -408 -16 -374 18
rect -408 -84 -374 -54
rect -408 -88 -374 -84
rect -408 -152 -374 -126
rect -408 -160 -374 -152
rect -408 -220 -374 -198
rect -408 -232 -374 -220
rect -408 -288 -374 -270
rect -408 -304 -374 -288
rect -408 -356 -374 -342
rect -408 -376 -374 -356
rect -408 -424 -374 -414
rect -408 -448 -374 -424
rect -408 -492 -374 -486
rect -408 -520 -374 -492
rect -408 -560 -374 -558
rect -408 -592 -374 -560
rect -310 562 -276 594
rect -310 560 -276 562
rect -310 494 -276 522
rect -310 488 -276 494
rect -310 426 -276 450
rect -310 416 -276 426
rect -310 358 -276 378
rect -310 344 -276 358
rect -310 290 -276 306
rect -310 272 -276 290
rect -310 222 -276 234
rect -310 200 -276 222
rect -310 154 -276 162
rect -310 128 -276 154
rect -310 86 -276 90
rect -310 56 -276 86
rect -310 -16 -276 18
rect -310 -84 -276 -54
rect -310 -88 -276 -84
rect -310 -152 -276 -126
rect -310 -160 -276 -152
rect -310 -220 -276 -198
rect -310 -232 -276 -220
rect -310 -288 -276 -270
rect -310 -304 -276 -288
rect -310 -356 -276 -342
rect -310 -376 -276 -356
rect -310 -424 -276 -414
rect -310 -448 -276 -424
rect -310 -492 -276 -486
rect -310 -520 -276 -492
rect -310 -560 -276 -558
rect -310 -592 -276 -560
rect -212 562 -178 594
rect -212 560 -178 562
rect -212 494 -178 522
rect -212 488 -178 494
rect -212 426 -178 450
rect -212 416 -178 426
rect -212 358 -178 378
rect -212 344 -178 358
rect -212 290 -178 306
rect -212 272 -178 290
rect -212 222 -178 234
rect -212 200 -178 222
rect -212 154 -178 162
rect -212 128 -178 154
rect -212 86 -178 90
rect -212 56 -178 86
rect -212 -16 -178 18
rect -212 -84 -178 -54
rect -212 -88 -178 -84
rect -212 -152 -178 -126
rect -212 -160 -178 -152
rect -212 -220 -178 -198
rect -212 -232 -178 -220
rect -212 -288 -178 -270
rect -212 -304 -178 -288
rect -212 -356 -178 -342
rect -212 -376 -178 -356
rect -212 -424 -178 -414
rect -212 -448 -178 -424
rect -212 -492 -178 -486
rect -212 -520 -178 -492
rect -212 -560 -178 -558
rect -212 -592 -178 -560
rect -114 562 -80 594
rect -114 560 -80 562
rect -114 494 -80 522
rect -114 488 -80 494
rect -114 426 -80 450
rect -114 416 -80 426
rect -114 358 -80 378
rect -114 344 -80 358
rect -114 290 -80 306
rect -114 272 -80 290
rect -114 222 -80 234
rect -114 200 -80 222
rect -114 154 -80 162
rect -114 128 -80 154
rect -114 86 -80 90
rect -114 56 -80 86
rect -114 -16 -80 18
rect -114 -84 -80 -54
rect -114 -88 -80 -84
rect -114 -152 -80 -126
rect -114 -160 -80 -152
rect -114 -220 -80 -198
rect -114 -232 -80 -220
rect -114 -288 -80 -270
rect -114 -304 -80 -288
rect -114 -356 -80 -342
rect -114 -376 -80 -356
rect -114 -424 -80 -414
rect -114 -448 -80 -424
rect -114 -492 -80 -486
rect -114 -520 -80 -492
rect -114 -560 -80 -558
rect -114 -592 -80 -560
rect -16 562 18 594
rect -16 560 18 562
rect -16 494 18 522
rect -16 488 18 494
rect -16 426 18 450
rect -16 416 18 426
rect -16 358 18 378
rect -16 344 18 358
rect -16 290 18 306
rect -16 272 18 290
rect -16 222 18 234
rect -16 200 18 222
rect -16 154 18 162
rect -16 128 18 154
rect -16 86 18 90
rect -16 56 18 86
rect -16 -16 18 18
rect -16 -84 18 -54
rect -16 -88 18 -84
rect -16 -152 18 -126
rect -16 -160 18 -152
rect -16 -220 18 -198
rect -16 -232 18 -220
rect -16 -288 18 -270
rect -16 -304 18 -288
rect -16 -356 18 -342
rect -16 -376 18 -356
rect -16 -424 18 -414
rect -16 -448 18 -424
rect -16 -492 18 -486
rect -16 -520 18 -492
rect -16 -560 18 -558
rect -16 -592 18 -560
rect 82 562 116 594
rect 82 560 116 562
rect 82 494 116 522
rect 82 488 116 494
rect 82 426 116 450
rect 82 416 116 426
rect 82 358 116 378
rect 82 344 116 358
rect 82 290 116 306
rect 82 272 116 290
rect 82 222 116 234
rect 82 200 116 222
rect 82 154 116 162
rect 82 128 116 154
rect 82 86 116 90
rect 82 56 116 86
rect 82 -16 116 18
rect 82 -84 116 -54
rect 82 -88 116 -84
rect 82 -152 116 -126
rect 82 -160 116 -152
rect 82 -220 116 -198
rect 82 -232 116 -220
rect 82 -288 116 -270
rect 82 -304 116 -288
rect 82 -356 116 -342
rect 82 -376 116 -356
rect 82 -424 116 -414
rect 82 -448 116 -424
rect 82 -492 116 -486
rect 82 -520 116 -492
rect 82 -560 116 -558
rect 82 -592 116 -560
rect 180 562 214 594
rect 180 560 214 562
rect 180 494 214 522
rect 180 488 214 494
rect 180 426 214 450
rect 180 416 214 426
rect 180 358 214 378
rect 180 344 214 358
rect 180 290 214 306
rect 180 272 214 290
rect 180 222 214 234
rect 180 200 214 222
rect 180 154 214 162
rect 180 128 214 154
rect 180 86 214 90
rect 180 56 214 86
rect 180 -16 214 18
rect 180 -84 214 -54
rect 180 -88 214 -84
rect 180 -152 214 -126
rect 180 -160 214 -152
rect 180 -220 214 -198
rect 180 -232 214 -220
rect 180 -288 214 -270
rect 180 -304 214 -288
rect 180 -356 214 -342
rect 180 -376 214 -356
rect 180 -424 214 -414
rect 180 -448 214 -424
rect 180 -492 214 -486
rect 180 -520 214 -492
rect 180 -560 214 -558
rect 180 -592 214 -560
rect 278 562 312 594
rect 278 560 312 562
rect 278 494 312 522
rect 278 488 312 494
rect 278 426 312 450
rect 278 416 312 426
rect 278 358 312 378
rect 278 344 312 358
rect 278 290 312 306
rect 278 272 312 290
rect 278 222 312 234
rect 278 200 312 222
rect 278 154 312 162
rect 278 128 312 154
rect 278 86 312 90
rect 278 56 312 86
rect 278 -16 312 18
rect 278 -84 312 -54
rect 278 -88 312 -84
rect 278 -152 312 -126
rect 278 -160 312 -152
rect 278 -220 312 -198
rect 278 -232 312 -220
rect 278 -288 312 -270
rect 278 -304 312 -288
rect 278 -356 312 -342
rect 278 -376 312 -356
rect 278 -424 312 -414
rect 278 -448 312 -424
rect 278 -492 312 -486
rect 278 -520 312 -492
rect 278 -560 312 -558
rect 278 -592 312 -560
rect 376 562 410 594
rect 376 560 410 562
rect 376 494 410 522
rect 376 488 410 494
rect 376 426 410 450
rect 376 416 410 426
rect 376 358 410 378
rect 376 344 410 358
rect 376 290 410 306
rect 376 272 410 290
rect 376 222 410 234
rect 376 200 410 222
rect 376 154 410 162
rect 376 128 410 154
rect 376 86 410 90
rect 376 56 410 86
rect 376 -16 410 18
rect 376 -84 410 -54
rect 376 -88 410 -84
rect 376 -152 410 -126
rect 376 -160 410 -152
rect 376 -220 410 -198
rect 376 -232 410 -220
rect 376 -288 410 -270
rect 376 -304 410 -288
rect 376 -356 410 -342
rect 376 -376 410 -356
rect 376 -424 410 -414
rect 376 -448 410 -424
rect 376 -492 410 -486
rect 376 -520 410 -492
rect 376 -560 410 -558
rect 376 -592 410 -560
rect 474 562 508 594
rect 474 560 508 562
rect 474 494 508 522
rect 474 488 508 494
rect 474 426 508 450
rect 474 416 508 426
rect 474 358 508 378
rect 474 344 508 358
rect 474 290 508 306
rect 474 272 508 290
rect 474 222 508 234
rect 474 200 508 222
rect 474 154 508 162
rect 474 128 508 154
rect 474 86 508 90
rect 474 56 508 86
rect 474 -16 508 18
rect 474 -84 508 -54
rect 474 -88 508 -84
rect 474 -152 508 -126
rect 474 -160 508 -152
rect 474 -220 508 -198
rect 474 -232 508 -220
rect 474 -288 508 -270
rect 474 -304 508 -288
rect 474 -356 508 -342
rect 474 -376 508 -356
rect 474 -424 508 -414
rect 474 -448 508 -424
rect 474 -492 508 -486
rect 474 -520 508 -492
rect 474 -560 508 -558
rect 474 -592 508 -560
rect 572 562 606 594
rect 572 560 606 562
rect 572 494 606 522
rect 572 488 606 494
rect 572 426 606 450
rect 572 416 606 426
rect 572 358 606 378
rect 572 344 606 358
rect 572 290 606 306
rect 572 272 606 290
rect 572 222 606 234
rect 572 200 606 222
rect 572 154 606 162
rect 572 128 606 154
rect 572 86 606 90
rect 572 56 606 86
rect 572 -16 606 18
rect 572 -84 606 -54
rect 572 -88 606 -84
rect 572 -152 606 -126
rect 572 -160 606 -152
rect 572 -220 606 -198
rect 572 -232 606 -220
rect 572 -288 606 -270
rect 572 -304 606 -288
rect 572 -356 606 -342
rect 572 -376 606 -356
rect 572 -424 606 -414
rect 572 -448 606 -424
rect 572 -492 606 -486
rect 572 -520 606 -492
rect 572 -560 606 -558
rect 572 -592 606 -560
rect 670 562 704 594
rect 670 560 704 562
rect 670 494 704 522
rect 670 488 704 494
rect 670 426 704 450
rect 670 416 704 426
rect 670 358 704 378
rect 670 344 704 358
rect 670 290 704 306
rect 670 272 704 290
rect 670 222 704 234
rect 670 200 704 222
rect 670 154 704 162
rect 670 128 704 154
rect 670 86 704 90
rect 670 56 704 86
rect 670 -16 704 18
rect 670 -84 704 -54
rect 670 -88 704 -84
rect 670 -152 704 -126
rect 670 -160 704 -152
rect 670 -220 704 -198
rect 670 -232 704 -220
rect 670 -288 704 -270
rect 670 -304 704 -288
rect 670 -356 704 -342
rect 670 -376 704 -356
rect 670 -424 704 -414
rect 670 -448 704 -424
rect 670 -492 704 -486
rect 670 -520 704 -492
rect 670 -560 704 -558
rect 670 -592 704 -560
rect 768 562 802 594
rect 768 560 802 562
rect 768 494 802 522
rect 768 488 802 494
rect 768 426 802 450
rect 768 416 802 426
rect 768 358 802 378
rect 768 344 802 358
rect 768 290 802 306
rect 768 272 802 290
rect 768 222 802 234
rect 768 200 802 222
rect 768 154 802 162
rect 768 128 802 154
rect 768 86 802 90
rect 768 56 802 86
rect 768 -16 802 18
rect 768 -84 802 -54
rect 768 -88 802 -84
rect 768 -152 802 -126
rect 768 -160 802 -152
rect 768 -220 802 -198
rect 768 -232 802 -220
rect 768 -288 802 -270
rect 768 -304 802 -288
rect 768 -356 802 -342
rect 768 -376 802 -356
rect 768 -424 802 -414
rect 768 -448 802 -424
rect 768 -492 802 -486
rect 768 -520 802 -492
rect 768 -560 802 -558
rect 768 -592 802 -560
<< metal1 >>
rect -702 744 704 778
rect -1088 697 -910 732
rect -1088 591 -1051 697
rect -945 591 -910 697
rect -702 626 -668 744
rect -506 626 -472 744
rect -310 626 -276 744
rect -114 626 -80 744
rect 82 626 116 744
rect 278 626 312 744
rect 474 626 508 744
rect 670 626 704 744
rect -1088 556 -910 591
rect -806 594 -760 626
rect -806 560 -800 594
rect -766 560 -760 594
rect -806 522 -760 560
rect -806 488 -800 522
rect -766 488 -760 522
rect -806 450 -760 488
rect -806 416 -800 450
rect -766 416 -760 450
rect -806 378 -760 416
rect -806 344 -800 378
rect -766 344 -760 378
rect -806 306 -760 344
rect -806 272 -800 306
rect -766 272 -760 306
rect -806 234 -760 272
rect -806 200 -800 234
rect -766 200 -760 234
rect -806 162 -760 200
rect -806 128 -800 162
rect -766 128 -760 162
rect -806 90 -760 128
rect -806 56 -800 90
rect -766 56 -760 90
rect -806 18 -760 56
rect -806 -16 -800 18
rect -766 -16 -760 18
rect -806 -54 -760 -16
rect -806 -88 -800 -54
rect -766 -88 -760 -54
rect -806 -126 -760 -88
rect -806 -160 -800 -126
rect -766 -160 -760 -126
rect -806 -198 -760 -160
rect -806 -232 -800 -198
rect -766 -232 -760 -198
rect -806 -270 -760 -232
rect -806 -304 -800 -270
rect -766 -304 -760 -270
rect -806 -342 -760 -304
rect -806 -376 -800 -342
rect -766 -376 -760 -342
rect -806 -414 -760 -376
rect -806 -448 -800 -414
rect -766 -448 -760 -414
rect -806 -486 -760 -448
rect -806 -520 -800 -486
rect -766 -520 -760 -486
rect -1088 -589 -910 -554
rect -1088 -695 -1051 -589
rect -945 -695 -910 -589
rect -806 -558 -760 -520
rect -806 -592 -800 -558
rect -766 -592 -760 -558
rect -806 -624 -760 -592
rect -708 594 -662 626
rect -708 560 -702 594
rect -668 560 -662 594
rect -708 522 -662 560
rect -708 488 -702 522
rect -668 488 -662 522
rect -708 450 -662 488
rect -708 416 -702 450
rect -668 416 -662 450
rect -708 378 -662 416
rect -708 344 -702 378
rect -668 344 -662 378
rect -708 306 -662 344
rect -708 272 -702 306
rect -668 272 -662 306
rect -708 234 -662 272
rect -708 200 -702 234
rect -668 200 -662 234
rect -708 162 -662 200
rect -708 128 -702 162
rect -668 128 -662 162
rect -708 90 -662 128
rect -708 56 -702 90
rect -668 56 -662 90
rect -708 18 -662 56
rect -708 -16 -702 18
rect -668 -16 -662 18
rect -708 -54 -662 -16
rect -708 -88 -702 -54
rect -668 -88 -662 -54
rect -708 -126 -662 -88
rect -708 -160 -702 -126
rect -668 -160 -662 -126
rect -708 -198 -662 -160
rect -708 -232 -702 -198
rect -668 -232 -662 -198
rect -708 -270 -662 -232
rect -708 -304 -702 -270
rect -668 -304 -662 -270
rect -708 -342 -662 -304
rect -708 -376 -702 -342
rect -668 -376 -662 -342
rect -708 -414 -662 -376
rect -708 -448 -702 -414
rect -668 -448 -662 -414
rect -708 -486 -662 -448
rect -708 -520 -702 -486
rect -668 -520 -662 -486
rect -708 -558 -662 -520
rect -708 -592 -702 -558
rect -668 -592 -662 -558
rect -708 -624 -662 -592
rect -610 594 -564 626
rect -610 560 -604 594
rect -570 560 -564 594
rect -610 522 -564 560
rect -610 488 -604 522
rect -570 488 -564 522
rect -610 450 -564 488
rect -610 416 -604 450
rect -570 416 -564 450
rect -610 378 -564 416
rect -610 344 -604 378
rect -570 344 -564 378
rect -610 306 -564 344
rect -610 272 -604 306
rect -570 272 -564 306
rect -610 234 -564 272
rect -610 200 -604 234
rect -570 200 -564 234
rect -610 162 -564 200
rect -610 128 -604 162
rect -570 128 -564 162
rect -610 90 -564 128
rect -610 56 -604 90
rect -570 56 -564 90
rect -610 18 -564 56
rect -610 -16 -604 18
rect -570 -16 -564 18
rect -610 -54 -564 -16
rect -610 -88 -604 -54
rect -570 -88 -564 -54
rect -610 -126 -564 -88
rect -610 -160 -604 -126
rect -570 -160 -564 -126
rect -610 -198 -564 -160
rect -610 -232 -604 -198
rect -570 -232 -564 -198
rect -610 -270 -564 -232
rect -610 -304 -604 -270
rect -570 -304 -564 -270
rect -610 -342 -564 -304
rect -610 -376 -604 -342
rect -570 -376 -564 -342
rect -610 -414 -564 -376
rect -610 -448 -604 -414
rect -570 -448 -564 -414
rect -610 -486 -564 -448
rect -610 -520 -604 -486
rect -570 -520 -564 -486
rect -610 -558 -564 -520
rect -610 -592 -604 -558
rect -570 -592 -564 -558
rect -1088 -730 -910 -695
rect -800 -838 -766 -624
rect -610 -742 -564 -592
rect -512 594 -466 626
rect -512 560 -506 594
rect -472 560 -466 594
rect -512 522 -466 560
rect -512 488 -506 522
rect -472 488 -466 522
rect -512 450 -466 488
rect -512 416 -506 450
rect -472 416 -466 450
rect -512 378 -466 416
rect -512 344 -506 378
rect -472 344 -466 378
rect -512 306 -466 344
rect -512 272 -506 306
rect -472 272 -466 306
rect -512 234 -466 272
rect -512 200 -506 234
rect -472 200 -466 234
rect -512 162 -466 200
rect -512 128 -506 162
rect -472 128 -466 162
rect -512 90 -466 128
rect -512 56 -506 90
rect -472 56 -466 90
rect -512 18 -466 56
rect -512 -16 -506 18
rect -472 -16 -466 18
rect -512 -54 -466 -16
rect -512 -88 -506 -54
rect -472 -88 -466 -54
rect -512 -126 -466 -88
rect -512 -160 -506 -126
rect -472 -160 -466 -126
rect -512 -198 -466 -160
rect -512 -232 -506 -198
rect -472 -232 -466 -198
rect -512 -270 -466 -232
rect -512 -304 -506 -270
rect -472 -304 -466 -270
rect -512 -342 -466 -304
rect -512 -376 -506 -342
rect -472 -376 -466 -342
rect -512 -414 -466 -376
rect -512 -448 -506 -414
rect -472 -448 -466 -414
rect -512 -486 -466 -448
rect -512 -520 -506 -486
rect -472 -520 -466 -486
rect -512 -558 -466 -520
rect -512 -592 -506 -558
rect -472 -592 -466 -558
rect -512 -624 -466 -592
rect -414 594 -368 626
rect -414 560 -408 594
rect -374 560 -368 594
rect -414 522 -368 560
rect -414 488 -408 522
rect -374 488 -368 522
rect -414 450 -368 488
rect -414 416 -408 450
rect -374 416 -368 450
rect -414 378 -368 416
rect -414 344 -408 378
rect -374 344 -368 378
rect -414 306 -368 344
rect -414 272 -408 306
rect -374 272 -368 306
rect -414 234 -368 272
rect -414 200 -408 234
rect -374 200 -368 234
rect -414 162 -368 200
rect -414 128 -408 162
rect -374 128 -368 162
rect -414 90 -368 128
rect -414 56 -408 90
rect -374 56 -368 90
rect -414 18 -368 56
rect -414 -16 -408 18
rect -374 -16 -368 18
rect -414 -54 -368 -16
rect -414 -88 -408 -54
rect -374 -88 -368 -54
rect -414 -126 -368 -88
rect -414 -160 -408 -126
rect -374 -160 -368 -126
rect -414 -198 -368 -160
rect -414 -232 -408 -198
rect -374 -232 -368 -198
rect -414 -270 -368 -232
rect -414 -304 -408 -270
rect -374 -304 -368 -270
rect -414 -342 -368 -304
rect -414 -376 -408 -342
rect -374 -376 -368 -342
rect -414 -414 -368 -376
rect -414 -448 -408 -414
rect -374 -448 -368 -414
rect -414 -486 -368 -448
rect -414 -520 -408 -486
rect -374 -520 -368 -486
rect -414 -558 -368 -520
rect -414 -592 -408 -558
rect -374 -592 -368 -558
rect -414 -624 -368 -592
rect -316 594 -270 626
rect -316 560 -310 594
rect -276 560 -270 594
rect -316 522 -270 560
rect -316 488 -310 522
rect -276 488 -270 522
rect -316 450 -270 488
rect -316 416 -310 450
rect -276 416 -270 450
rect -316 378 -270 416
rect -316 344 -310 378
rect -276 344 -270 378
rect -316 306 -270 344
rect -316 272 -310 306
rect -276 272 -270 306
rect -316 234 -270 272
rect -316 200 -310 234
rect -276 200 -270 234
rect -316 162 -270 200
rect -316 128 -310 162
rect -276 128 -270 162
rect -316 90 -270 128
rect -316 56 -310 90
rect -276 56 -270 90
rect -316 18 -270 56
rect -316 -16 -310 18
rect -276 -16 -270 18
rect -316 -54 -270 -16
rect -316 -88 -310 -54
rect -276 -88 -270 -54
rect -316 -126 -270 -88
rect -316 -160 -310 -126
rect -276 -160 -270 -126
rect -316 -198 -270 -160
rect -316 -232 -310 -198
rect -276 -232 -270 -198
rect -316 -270 -270 -232
rect -316 -304 -310 -270
rect -276 -304 -270 -270
rect -316 -342 -270 -304
rect -316 -376 -310 -342
rect -276 -376 -270 -342
rect -316 -414 -270 -376
rect -316 -448 -310 -414
rect -276 -448 -270 -414
rect -316 -486 -270 -448
rect -316 -520 -310 -486
rect -276 -520 -270 -486
rect -316 -558 -270 -520
rect -316 -592 -310 -558
rect -276 -592 -270 -558
rect -316 -624 -270 -592
rect -218 594 -172 626
rect -218 560 -212 594
rect -178 560 -172 594
rect -218 522 -172 560
rect -218 488 -212 522
rect -178 488 -172 522
rect -218 450 -172 488
rect -218 416 -212 450
rect -178 416 -172 450
rect -218 378 -172 416
rect -218 344 -212 378
rect -178 344 -172 378
rect -218 306 -172 344
rect -218 272 -212 306
rect -178 272 -172 306
rect -218 234 -172 272
rect -218 200 -212 234
rect -178 200 -172 234
rect -218 162 -172 200
rect -218 128 -212 162
rect -178 128 -172 162
rect -218 90 -172 128
rect -218 56 -212 90
rect -178 56 -172 90
rect -218 18 -172 56
rect -218 -16 -212 18
rect -178 -16 -172 18
rect -218 -54 -172 -16
rect -218 -88 -212 -54
rect -178 -88 -172 -54
rect -218 -126 -172 -88
rect -218 -160 -212 -126
rect -178 -160 -172 -126
rect -218 -198 -172 -160
rect -218 -232 -212 -198
rect -178 -232 -172 -198
rect -218 -270 -172 -232
rect -218 -304 -212 -270
rect -178 -304 -172 -270
rect -218 -342 -172 -304
rect -218 -376 -212 -342
rect -178 -376 -172 -342
rect -218 -414 -172 -376
rect -218 -448 -212 -414
rect -178 -448 -172 -414
rect -218 -486 -172 -448
rect -218 -520 -212 -486
rect -178 -520 -172 -486
rect -218 -558 -172 -520
rect -218 -592 -212 -558
rect -178 -592 -172 -558
rect -636 -748 -536 -742
rect -636 -800 -612 -748
rect -560 -800 -536 -748
rect -636 -806 -536 -800
rect -408 -838 -374 -624
rect -218 -742 -172 -592
rect -120 594 -74 626
rect -120 560 -114 594
rect -80 560 -74 594
rect -120 522 -74 560
rect -120 488 -114 522
rect -80 488 -74 522
rect -120 450 -74 488
rect -120 416 -114 450
rect -80 416 -74 450
rect -120 378 -74 416
rect -120 344 -114 378
rect -80 344 -74 378
rect -120 306 -74 344
rect -120 272 -114 306
rect -80 272 -74 306
rect -120 234 -74 272
rect -120 200 -114 234
rect -80 200 -74 234
rect -120 162 -74 200
rect -120 128 -114 162
rect -80 128 -74 162
rect -120 90 -74 128
rect -120 56 -114 90
rect -80 56 -74 90
rect -120 18 -74 56
rect -120 -16 -114 18
rect -80 -16 -74 18
rect -120 -54 -74 -16
rect -120 -88 -114 -54
rect -80 -88 -74 -54
rect -120 -126 -74 -88
rect -120 -160 -114 -126
rect -80 -160 -74 -126
rect -120 -198 -74 -160
rect -120 -232 -114 -198
rect -80 -232 -74 -198
rect -120 -270 -74 -232
rect -120 -304 -114 -270
rect -80 -304 -74 -270
rect -120 -342 -74 -304
rect -120 -376 -114 -342
rect -80 -376 -74 -342
rect -120 -414 -74 -376
rect -120 -448 -114 -414
rect -80 -448 -74 -414
rect -120 -486 -74 -448
rect -120 -520 -114 -486
rect -80 -520 -74 -486
rect -120 -558 -74 -520
rect -120 -592 -114 -558
rect -80 -592 -74 -558
rect -120 -624 -74 -592
rect -22 594 24 626
rect -22 560 -16 594
rect 18 560 24 594
rect -22 522 24 560
rect -22 488 -16 522
rect 18 488 24 522
rect -22 450 24 488
rect -22 416 -16 450
rect 18 416 24 450
rect -22 378 24 416
rect -22 344 -16 378
rect 18 344 24 378
rect -22 306 24 344
rect -22 272 -16 306
rect 18 272 24 306
rect -22 234 24 272
rect -22 200 -16 234
rect 18 200 24 234
rect -22 162 24 200
rect -22 128 -16 162
rect 18 128 24 162
rect -22 90 24 128
rect -22 56 -16 90
rect 18 56 24 90
rect -22 18 24 56
rect -22 -16 -16 18
rect 18 -16 24 18
rect -22 -54 24 -16
rect -22 -88 -16 -54
rect 18 -88 24 -54
rect -22 -126 24 -88
rect -22 -160 -16 -126
rect 18 -160 24 -126
rect -22 -198 24 -160
rect -22 -232 -16 -198
rect 18 -232 24 -198
rect -22 -270 24 -232
rect -22 -304 -16 -270
rect 18 -304 24 -270
rect -22 -342 24 -304
rect -22 -376 -16 -342
rect 18 -376 24 -342
rect -22 -414 24 -376
rect -22 -448 -16 -414
rect 18 -448 24 -414
rect -22 -486 24 -448
rect -22 -520 -16 -486
rect 18 -520 24 -486
rect -22 -558 24 -520
rect -22 -592 -16 -558
rect 18 -592 24 -558
rect -22 -624 24 -592
rect 76 594 122 626
rect 76 560 82 594
rect 116 560 122 594
rect 76 522 122 560
rect 76 488 82 522
rect 116 488 122 522
rect 76 450 122 488
rect 76 416 82 450
rect 116 416 122 450
rect 76 378 122 416
rect 76 344 82 378
rect 116 344 122 378
rect 76 306 122 344
rect 76 272 82 306
rect 116 272 122 306
rect 76 234 122 272
rect 76 200 82 234
rect 116 200 122 234
rect 76 162 122 200
rect 76 128 82 162
rect 116 128 122 162
rect 76 90 122 128
rect 76 56 82 90
rect 116 56 122 90
rect 76 18 122 56
rect 76 -16 82 18
rect 116 -16 122 18
rect 76 -54 122 -16
rect 76 -88 82 -54
rect 116 -88 122 -54
rect 76 -126 122 -88
rect 76 -160 82 -126
rect 116 -160 122 -126
rect 76 -198 122 -160
rect 76 -232 82 -198
rect 116 -232 122 -198
rect 76 -270 122 -232
rect 76 -304 82 -270
rect 116 -304 122 -270
rect 76 -342 122 -304
rect 76 -376 82 -342
rect 116 -376 122 -342
rect 76 -414 122 -376
rect 76 -448 82 -414
rect 116 -448 122 -414
rect 76 -486 122 -448
rect 76 -520 82 -486
rect 116 -520 122 -486
rect 76 -558 122 -520
rect 76 -592 82 -558
rect 116 -592 122 -558
rect 76 -624 122 -592
rect 174 594 220 626
rect 174 560 180 594
rect 214 560 220 594
rect 174 522 220 560
rect 174 488 180 522
rect 214 488 220 522
rect 174 450 220 488
rect 174 416 180 450
rect 214 416 220 450
rect 174 378 220 416
rect 174 344 180 378
rect 214 344 220 378
rect 174 306 220 344
rect 174 272 180 306
rect 214 272 220 306
rect 174 234 220 272
rect 174 200 180 234
rect 214 200 220 234
rect 174 162 220 200
rect 174 128 180 162
rect 214 128 220 162
rect 174 90 220 128
rect 174 56 180 90
rect 214 56 220 90
rect 174 18 220 56
rect 174 -16 180 18
rect 214 -16 220 18
rect 174 -54 220 -16
rect 174 -88 180 -54
rect 214 -88 220 -54
rect 174 -126 220 -88
rect 174 -160 180 -126
rect 214 -160 220 -126
rect 174 -198 220 -160
rect 174 -232 180 -198
rect 214 -232 220 -198
rect 174 -270 220 -232
rect 174 -304 180 -270
rect 214 -304 220 -270
rect 174 -342 220 -304
rect 174 -376 180 -342
rect 214 -376 220 -342
rect 174 -414 220 -376
rect 174 -448 180 -414
rect 214 -448 220 -414
rect 174 -486 220 -448
rect 174 -520 180 -486
rect 214 -520 220 -486
rect 174 -558 220 -520
rect 174 -592 180 -558
rect 214 -592 220 -558
rect -244 -748 -144 -742
rect -244 -800 -220 -748
rect -168 -800 -144 -748
rect -244 -806 -144 -800
rect -16 -838 18 -624
rect 174 -742 220 -592
rect 272 594 318 626
rect 272 560 278 594
rect 312 560 318 594
rect 272 522 318 560
rect 272 488 278 522
rect 312 488 318 522
rect 272 450 318 488
rect 272 416 278 450
rect 312 416 318 450
rect 272 378 318 416
rect 272 344 278 378
rect 312 344 318 378
rect 272 306 318 344
rect 272 272 278 306
rect 312 272 318 306
rect 272 234 318 272
rect 272 200 278 234
rect 312 200 318 234
rect 272 162 318 200
rect 272 128 278 162
rect 312 128 318 162
rect 272 90 318 128
rect 272 56 278 90
rect 312 56 318 90
rect 272 18 318 56
rect 272 -16 278 18
rect 312 -16 318 18
rect 272 -54 318 -16
rect 272 -88 278 -54
rect 312 -88 318 -54
rect 272 -126 318 -88
rect 272 -160 278 -126
rect 312 -160 318 -126
rect 272 -198 318 -160
rect 272 -232 278 -198
rect 312 -232 318 -198
rect 272 -270 318 -232
rect 272 -304 278 -270
rect 312 -304 318 -270
rect 272 -342 318 -304
rect 272 -376 278 -342
rect 312 -376 318 -342
rect 272 -414 318 -376
rect 272 -448 278 -414
rect 312 -448 318 -414
rect 272 -486 318 -448
rect 272 -520 278 -486
rect 312 -520 318 -486
rect 272 -558 318 -520
rect 272 -592 278 -558
rect 312 -592 318 -558
rect 272 -624 318 -592
rect 370 594 416 626
rect 370 560 376 594
rect 410 560 416 594
rect 370 522 416 560
rect 370 488 376 522
rect 410 488 416 522
rect 370 450 416 488
rect 370 416 376 450
rect 410 416 416 450
rect 370 378 416 416
rect 370 344 376 378
rect 410 344 416 378
rect 370 306 416 344
rect 370 272 376 306
rect 410 272 416 306
rect 370 234 416 272
rect 370 200 376 234
rect 410 200 416 234
rect 370 162 416 200
rect 370 128 376 162
rect 410 128 416 162
rect 370 90 416 128
rect 370 56 376 90
rect 410 56 416 90
rect 370 18 416 56
rect 370 -16 376 18
rect 410 -16 416 18
rect 370 -54 416 -16
rect 370 -88 376 -54
rect 410 -88 416 -54
rect 370 -126 416 -88
rect 370 -160 376 -126
rect 410 -160 416 -126
rect 370 -198 416 -160
rect 370 -232 376 -198
rect 410 -232 416 -198
rect 370 -270 416 -232
rect 370 -304 376 -270
rect 410 -304 416 -270
rect 370 -342 416 -304
rect 370 -376 376 -342
rect 410 -376 416 -342
rect 370 -414 416 -376
rect 370 -448 376 -414
rect 410 -448 416 -414
rect 370 -486 416 -448
rect 370 -520 376 -486
rect 410 -520 416 -486
rect 370 -558 416 -520
rect 370 -592 376 -558
rect 410 -592 416 -558
rect 370 -624 416 -592
rect 468 594 514 626
rect 468 560 474 594
rect 508 560 514 594
rect 468 522 514 560
rect 468 488 474 522
rect 508 488 514 522
rect 468 450 514 488
rect 468 416 474 450
rect 508 416 514 450
rect 468 378 514 416
rect 468 344 474 378
rect 508 344 514 378
rect 468 306 514 344
rect 468 272 474 306
rect 508 272 514 306
rect 468 234 514 272
rect 468 200 474 234
rect 508 200 514 234
rect 468 162 514 200
rect 468 128 474 162
rect 508 128 514 162
rect 468 90 514 128
rect 468 56 474 90
rect 508 56 514 90
rect 468 18 514 56
rect 468 -16 474 18
rect 508 -16 514 18
rect 468 -54 514 -16
rect 468 -88 474 -54
rect 508 -88 514 -54
rect 468 -126 514 -88
rect 468 -160 474 -126
rect 508 -160 514 -126
rect 468 -198 514 -160
rect 468 -232 474 -198
rect 508 -232 514 -198
rect 468 -270 514 -232
rect 468 -304 474 -270
rect 508 -304 514 -270
rect 468 -342 514 -304
rect 468 -376 474 -342
rect 508 -376 514 -342
rect 468 -414 514 -376
rect 468 -448 474 -414
rect 508 -448 514 -414
rect 468 -486 514 -448
rect 468 -520 474 -486
rect 508 -520 514 -486
rect 468 -558 514 -520
rect 468 -592 474 -558
rect 508 -592 514 -558
rect 468 -624 514 -592
rect 566 594 612 626
rect 566 560 572 594
rect 606 560 612 594
rect 566 522 612 560
rect 566 488 572 522
rect 606 488 612 522
rect 566 450 612 488
rect 566 416 572 450
rect 606 416 612 450
rect 566 378 612 416
rect 566 344 572 378
rect 606 344 612 378
rect 566 306 612 344
rect 566 272 572 306
rect 606 272 612 306
rect 566 234 612 272
rect 566 200 572 234
rect 606 200 612 234
rect 566 162 612 200
rect 566 128 572 162
rect 606 128 612 162
rect 566 90 612 128
rect 566 56 572 90
rect 606 56 612 90
rect 566 18 612 56
rect 566 -16 572 18
rect 606 -16 612 18
rect 566 -54 612 -16
rect 566 -88 572 -54
rect 606 -88 612 -54
rect 566 -126 612 -88
rect 566 -160 572 -126
rect 606 -160 612 -126
rect 566 -198 612 -160
rect 566 -232 572 -198
rect 606 -232 612 -198
rect 566 -270 612 -232
rect 566 -304 572 -270
rect 606 -304 612 -270
rect 566 -342 612 -304
rect 566 -376 572 -342
rect 606 -376 612 -342
rect 566 -414 612 -376
rect 566 -448 572 -414
rect 606 -448 612 -414
rect 566 -486 612 -448
rect 566 -520 572 -486
rect 606 -520 612 -486
rect 566 -558 612 -520
rect 566 -592 572 -558
rect 606 -592 612 -558
rect 148 -748 248 -742
rect 148 -800 172 -748
rect 224 -800 248 -748
rect 148 -806 248 -800
rect 376 -838 410 -624
rect 566 -742 612 -592
rect 664 594 710 626
rect 664 560 670 594
rect 704 560 710 594
rect 664 522 710 560
rect 664 488 670 522
rect 704 488 710 522
rect 664 450 710 488
rect 664 416 670 450
rect 704 416 710 450
rect 664 378 710 416
rect 664 344 670 378
rect 704 344 710 378
rect 664 306 710 344
rect 664 272 670 306
rect 704 272 710 306
rect 664 234 710 272
rect 664 200 670 234
rect 704 200 710 234
rect 664 162 710 200
rect 664 128 670 162
rect 704 128 710 162
rect 664 90 710 128
rect 664 56 670 90
rect 704 56 710 90
rect 664 18 710 56
rect 664 -16 670 18
rect 704 -16 710 18
rect 664 -54 710 -16
rect 664 -88 670 -54
rect 704 -88 710 -54
rect 664 -126 710 -88
rect 664 -160 670 -126
rect 704 -160 710 -126
rect 664 -198 710 -160
rect 664 -232 670 -198
rect 704 -232 710 -198
rect 664 -270 710 -232
rect 664 -304 670 -270
rect 704 -304 710 -270
rect 664 -342 710 -304
rect 664 -376 670 -342
rect 704 -376 710 -342
rect 664 -414 710 -376
rect 664 -448 670 -414
rect 704 -448 710 -414
rect 664 -486 710 -448
rect 664 -520 670 -486
rect 704 -520 710 -486
rect 664 -558 710 -520
rect 664 -592 670 -558
rect 704 -592 710 -558
rect 664 -624 710 -592
rect 762 594 808 626
rect 762 560 768 594
rect 802 560 808 594
rect 762 522 808 560
rect 762 488 768 522
rect 802 488 808 522
rect 762 450 808 488
rect 762 416 768 450
rect 802 416 808 450
rect 762 378 808 416
rect 762 344 768 378
rect 802 344 808 378
rect 762 306 808 344
rect 762 272 768 306
rect 802 272 808 306
rect 762 234 808 272
rect 762 200 768 234
rect 802 200 808 234
rect 762 162 808 200
rect 762 128 768 162
rect 802 128 808 162
rect 762 90 808 128
rect 762 56 768 90
rect 802 56 808 90
rect 762 18 808 56
rect 762 -16 768 18
rect 802 -16 808 18
rect 762 -54 808 -16
rect 762 -88 768 -54
rect 802 -88 808 -54
rect 762 -126 808 -88
rect 762 -160 768 -126
rect 802 -160 808 -126
rect 762 -198 808 -160
rect 762 -232 768 -198
rect 802 -232 808 -198
rect 762 -270 808 -232
rect 762 -304 768 -270
rect 802 -304 808 -270
rect 762 -342 808 -304
rect 762 -376 768 -342
rect 802 -376 808 -342
rect 762 -414 808 -376
rect 762 -448 768 -414
rect 802 -448 808 -414
rect 762 -486 808 -448
rect 762 -520 768 -486
rect 802 -520 808 -486
rect 762 -558 808 -520
rect 762 -592 768 -558
rect 802 -592 808 -558
rect 762 -624 808 -592
rect 540 -748 640 -742
rect 540 -800 564 -748
rect 616 -800 640 -748
rect 540 -806 640 -800
rect 768 -838 802 -624
rect -800 -872 802 -838
<< via1 >>
rect -612 -800 -560 -748
rect -220 -800 -168 -748
rect 172 -800 224 -748
rect 564 -800 616 -748
<< metal2 >>
rect -636 -748 640 -742
rect -636 -800 -612 -748
rect -560 -800 -220 -748
rect -168 -800 172 -748
rect 224 -800 564 -748
rect 616 -800 640 -748
rect -636 -806 640 -800
<< end >>
