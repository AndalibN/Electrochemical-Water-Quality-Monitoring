magic
tech sky130A
magscale 1 2
timestamp 1668031433
<< checkpaint >>
rect 426 22098 3020 24148
rect -306 22060 3020 22098
rect -1868 828 3020 22060
rect 4934 3024 7528 26344
rect -1868 -1222 2288 828
rect -1868 -1260 1932 -1222
rect -1418 -1748 1908 -1260
rect -1126 -2274 1908 -1748
rect -1126 -5026 1644 -2274
rect -950 -5582 1644 -5026
<< psubdiff >>
rect -608 3856 -248 3958
rect -608 2854 -522 3856
rect -338 2854 -248 3856
rect -608 2734 -248 2854
<< psubdiffcont >>
rect -522 2854 -338 3856
<< locali >>
rect 284 10046 414 10072
rect 284 9078 312 10046
rect 382 9078 414 10046
rect 284 9052 414 9078
rect -564 3856 -290 3914
rect -564 2854 -522 3856
rect -338 2854 -290 3856
rect -564 2794 -290 2854
rect 264 3080 430 3108
rect 264 2112 308 3080
rect 382 2112 430 3080
rect 264 2084 430 2112
<< viali >>
rect 312 9078 382 10046
rect 308 2112 382 3080
<< metal1 >>
rect 284 10046 414 10072
rect 284 9078 312 10046
rect 382 9078 414 10046
rect 284 9052 414 9078
rect 264 3080 430 3108
rect 264 2112 308 3080
rect 382 2112 430 3080
rect 264 2084 430 2112
use sky130_fd_pr__res_xhigh_po_0p35_RGUCK9  sky130_fd_pr__res_xhigh_po_0p35_RGUCK9_0
timestamp 1668029120
transform 1 0 347 0 1 6078
box -37 -10400 37 10400
<< labels >>
rlabel space 672 6692 672 6692 5 top
rlabel space 30 88 30 88 1 bot
rlabel psubdiffcont -430 3360 -430 3360 7 gnd
<< end >>
