magic
tech sky130A
magscale 1 2
timestamp 1667321908
<< error_p >>
rect -31 6655 31 6661
rect -31 6621 -19 6655
rect -31 6615 31 6621
rect -31 3417 31 3423
rect -31 3383 -19 3417
rect -31 3377 31 3383
rect -31 3309 31 3315
rect -31 3275 -19 3309
rect -31 3269 31 3275
rect -31 71 31 77
rect -31 37 -19 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect -31 -77 31 -71
rect -31 -3275 31 -3269
rect -31 -3309 -19 -3275
rect -31 -3315 31 -3309
rect -31 -3383 31 -3377
rect -31 -3417 -19 -3383
rect -31 -3423 31 -3417
rect -31 -6621 31 -6615
rect -31 -6655 -19 -6621
rect -31 -6661 31 -6655
<< nwell >>
rect -231 -6793 231 6793
<< pmoslvt >>
rect -35 3464 35 6574
rect -35 118 35 3228
rect -35 -3228 35 -118
rect -35 -6574 35 -3464
<< pdiff >>
rect -93 6562 -35 6574
rect -93 3476 -81 6562
rect -47 3476 -35 6562
rect -93 3464 -35 3476
rect 35 6562 93 6574
rect 35 3476 47 6562
rect 81 3476 93 6562
rect 35 3464 93 3476
rect -93 3216 -35 3228
rect -93 130 -81 3216
rect -47 130 -35 3216
rect -93 118 -35 130
rect 35 3216 93 3228
rect 35 130 47 3216
rect 81 130 93 3216
rect 35 118 93 130
rect -93 -130 -35 -118
rect -93 -3216 -81 -130
rect -47 -3216 -35 -130
rect -93 -3228 -35 -3216
rect 35 -130 93 -118
rect 35 -3216 47 -130
rect 81 -3216 93 -130
rect 35 -3228 93 -3216
rect -93 -3476 -35 -3464
rect -93 -6562 -81 -3476
rect -47 -6562 -35 -3476
rect -93 -6574 -35 -6562
rect 35 -3476 93 -3464
rect 35 -6562 47 -3476
rect 81 -6562 93 -3476
rect 35 -6574 93 -6562
<< pdiffc >>
rect -81 3476 -47 6562
rect 47 3476 81 6562
rect -81 130 -47 3216
rect 47 130 81 3216
rect -81 -3216 -47 -130
rect 47 -3216 81 -130
rect -81 -6562 -47 -3476
rect 47 -6562 81 -3476
<< nsubdiff >>
rect -195 6723 -99 6757
rect 99 6723 195 6757
rect -195 6661 -161 6723
rect 161 6661 195 6723
rect -195 -6723 -161 -6661
rect 161 -6723 195 -6661
rect -195 -6757 -99 -6723
rect 99 -6757 195 -6723
<< nsubdiffcont >>
rect -99 6723 99 6757
rect -195 -6661 -161 6661
rect 161 -6661 195 6661
rect -99 -6757 99 -6723
<< poly >>
rect -35 6655 35 6671
rect -35 6621 -19 6655
rect 19 6621 35 6655
rect -35 6574 35 6621
rect -35 3417 35 3464
rect -35 3383 -19 3417
rect 19 3383 35 3417
rect -35 3367 35 3383
rect -35 3309 35 3325
rect -35 3275 -19 3309
rect 19 3275 35 3309
rect -35 3228 35 3275
rect -35 71 35 118
rect -35 37 -19 71
rect 19 37 35 71
rect -35 21 35 37
rect -35 -37 35 -21
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -35 -118 35 -71
rect -35 -3275 35 -3228
rect -35 -3309 -19 -3275
rect 19 -3309 35 -3275
rect -35 -3325 35 -3309
rect -35 -3383 35 -3367
rect -35 -3417 -19 -3383
rect 19 -3417 35 -3383
rect -35 -3464 35 -3417
rect -35 -6621 35 -6574
rect -35 -6655 -19 -6621
rect 19 -6655 35 -6621
rect -35 -6671 35 -6655
<< polycont >>
rect -19 6621 19 6655
rect -19 3383 19 3417
rect -19 3275 19 3309
rect -19 37 19 71
rect -19 -71 19 -37
rect -19 -3309 19 -3275
rect -19 -3417 19 -3383
rect -19 -6655 19 -6621
<< locali >>
rect -195 6723 -99 6757
rect 99 6723 195 6757
rect -195 6661 -161 6723
rect 161 6661 195 6723
rect -35 6621 -19 6655
rect 19 6621 35 6655
rect -81 6562 -47 6578
rect -81 3460 -47 3476
rect 47 6562 81 6578
rect 47 3460 81 3476
rect -35 3383 -19 3417
rect 19 3383 35 3417
rect -35 3275 -19 3309
rect 19 3275 35 3309
rect -81 3216 -47 3232
rect -81 114 -47 130
rect 47 3216 81 3232
rect 47 114 81 130
rect -35 37 -19 71
rect 19 37 35 71
rect -35 -71 -19 -37
rect 19 -71 35 -37
rect -81 -130 -47 -114
rect -81 -3232 -47 -3216
rect 47 -130 81 -114
rect 47 -3232 81 -3216
rect -35 -3309 -19 -3275
rect 19 -3309 35 -3275
rect -35 -3417 -19 -3383
rect 19 -3417 35 -3383
rect -81 -3476 -47 -3460
rect -81 -6578 -47 -6562
rect 47 -3476 81 -3460
rect 47 -6578 81 -6562
rect -35 -6655 -19 -6621
rect 19 -6655 35 -6621
rect -195 -6723 -161 -6661
rect 161 -6723 195 -6661
rect -195 -6757 -99 -6723
rect 99 -6757 195 -6723
<< viali >>
rect -19 6621 19 6655
rect -81 3476 -47 6562
rect 47 3476 81 6562
rect -19 3383 19 3417
rect -19 3275 19 3309
rect -81 130 -47 3216
rect 47 130 81 3216
rect -19 37 19 71
rect -19 -71 19 -37
rect -81 -3216 -47 -130
rect 47 -3216 81 -130
rect -19 -3309 19 -3275
rect -19 -3417 19 -3383
rect -81 -6562 -47 -3476
rect 47 -6562 81 -3476
rect -19 -6655 19 -6621
<< metal1 >>
rect -31 6655 31 6661
rect -31 6621 -19 6655
rect 19 6621 31 6655
rect -31 6615 31 6621
rect -87 6562 -41 6574
rect -87 3476 -81 6562
rect -47 3476 -41 6562
rect -87 3464 -41 3476
rect 41 6562 87 6574
rect 41 3476 47 6562
rect 81 3476 87 6562
rect 41 3464 87 3476
rect -31 3417 31 3423
rect -31 3383 -19 3417
rect 19 3383 31 3417
rect -31 3377 31 3383
rect -31 3309 31 3315
rect -31 3275 -19 3309
rect 19 3275 31 3309
rect -31 3269 31 3275
rect -87 3216 -41 3228
rect -87 130 -81 3216
rect -47 130 -41 3216
rect -87 118 -41 130
rect 41 3216 87 3228
rect 41 130 47 3216
rect 81 130 87 3216
rect 41 118 87 130
rect -31 71 31 77
rect -31 37 -19 71
rect 19 37 31 71
rect -31 31 31 37
rect -31 -37 31 -31
rect -31 -71 -19 -37
rect 19 -71 31 -37
rect -31 -77 31 -71
rect -87 -130 -41 -118
rect -87 -3216 -81 -130
rect -47 -3216 -41 -130
rect -87 -3228 -41 -3216
rect 41 -130 87 -118
rect 41 -3216 47 -130
rect 81 -3216 87 -130
rect 41 -3228 87 -3216
rect -31 -3275 31 -3269
rect -31 -3309 -19 -3275
rect 19 -3309 31 -3275
rect -31 -3315 31 -3309
rect -31 -3383 31 -3377
rect -31 -3417 -19 -3383
rect 19 -3417 31 -3383
rect -31 -3423 31 -3417
rect -87 -3476 -41 -3464
rect -87 -6562 -81 -3476
rect -47 -6562 -41 -3476
rect -87 -6574 -41 -6562
rect 41 -3476 87 -3464
rect 41 -6562 47 -3476
rect 81 -6562 87 -3476
rect 41 -6574 87 -6562
rect -31 -6621 31 -6615
rect -31 -6655 -19 -6621
rect 19 -6655 31 -6621
rect -31 -6661 31 -6655
<< properties >>
string FIXED_BBOX -178 -6740 178 6740
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 15.55 l 0.35 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
