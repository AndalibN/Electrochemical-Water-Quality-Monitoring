magic
tech sky130A
magscale 1 2
timestamp 1668369844
<< error_p >>
rect -1445 9672 -1387 9678
rect -1327 9672 -1269 9678
rect -1209 9672 -1151 9678
rect -1091 9672 -1033 9678
rect -973 9672 -915 9678
rect -855 9672 -797 9678
rect -737 9672 -679 9678
rect -619 9672 -561 9678
rect -501 9672 -443 9678
rect -383 9672 -325 9678
rect -265 9672 -207 9678
rect -147 9672 -89 9678
rect -29 9672 29 9678
rect 89 9672 147 9678
rect 207 9672 265 9678
rect 325 9672 383 9678
rect 443 9672 501 9678
rect 561 9672 619 9678
rect 679 9672 737 9678
rect 797 9672 855 9678
rect 915 9672 973 9678
rect 1033 9672 1091 9678
rect 1151 9672 1209 9678
rect 1269 9672 1327 9678
rect 1387 9672 1445 9678
rect -1445 9638 -1433 9672
rect -1327 9638 -1315 9672
rect -1209 9638 -1197 9672
rect -1091 9638 -1079 9672
rect -973 9638 -961 9672
rect -855 9638 -843 9672
rect -737 9638 -725 9672
rect -619 9638 -607 9672
rect -501 9638 -489 9672
rect -383 9638 -371 9672
rect -265 9638 -253 9672
rect -147 9638 -135 9672
rect -29 9638 -17 9672
rect 89 9638 101 9672
rect 207 9638 219 9672
rect 325 9638 337 9672
rect 443 9638 455 9672
rect 561 9638 573 9672
rect 679 9638 691 9672
rect 797 9638 809 9672
rect 915 9638 927 9672
rect 1033 9638 1045 9672
rect 1151 9638 1163 9672
rect 1269 9638 1281 9672
rect 1387 9638 1399 9672
rect -1445 9632 -1387 9638
rect -1327 9632 -1269 9638
rect -1209 9632 -1151 9638
rect -1091 9632 -1033 9638
rect -973 9632 -915 9638
rect -855 9632 -797 9638
rect -737 9632 -679 9638
rect -619 9632 -561 9638
rect -501 9632 -443 9638
rect -383 9632 -325 9638
rect -265 9632 -207 9638
rect -147 9632 -89 9638
rect -29 9632 29 9638
rect 89 9632 147 9638
rect 207 9632 265 9638
rect 325 9632 383 9638
rect 443 9632 501 9638
rect 561 9632 619 9638
rect 679 9632 737 9638
rect 797 9632 855 9638
rect 915 9632 973 9638
rect 1033 9632 1091 9638
rect 1151 9632 1209 9638
rect 1269 9632 1327 9638
rect 1387 9632 1445 9638
rect -1445 -9638 -1387 -9632
rect -1327 -9638 -1269 -9632
rect -1209 -9638 -1151 -9632
rect -1091 -9638 -1033 -9632
rect -973 -9638 -915 -9632
rect -855 -9638 -797 -9632
rect -737 -9638 -679 -9632
rect -619 -9638 -561 -9632
rect -501 -9638 -443 -9632
rect -383 -9638 -325 -9632
rect -265 -9638 -207 -9632
rect -147 -9638 -89 -9632
rect -29 -9638 29 -9632
rect 89 -9638 147 -9632
rect 207 -9638 265 -9632
rect 325 -9638 383 -9632
rect 443 -9638 501 -9632
rect 561 -9638 619 -9632
rect 679 -9638 737 -9632
rect 797 -9638 855 -9632
rect 915 -9638 973 -9632
rect 1033 -9638 1091 -9632
rect 1151 -9638 1209 -9632
rect 1269 -9638 1327 -9632
rect 1387 -9638 1445 -9632
rect -1445 -9672 -1433 -9638
rect -1327 -9672 -1315 -9638
rect -1209 -9672 -1197 -9638
rect -1091 -9672 -1079 -9638
rect -973 -9672 -961 -9638
rect -855 -9672 -843 -9638
rect -737 -9672 -725 -9638
rect -619 -9672 -607 -9638
rect -501 -9672 -489 -9638
rect -383 -9672 -371 -9638
rect -265 -9672 -253 -9638
rect -147 -9672 -135 -9638
rect -29 -9672 -17 -9638
rect 89 -9672 101 -9638
rect 207 -9672 219 -9638
rect 325 -9672 337 -9638
rect 443 -9672 455 -9638
rect 561 -9672 573 -9638
rect 679 -9672 691 -9638
rect 797 -9672 809 -9638
rect 915 -9672 927 -9638
rect 1033 -9672 1045 -9638
rect 1151 -9672 1163 -9638
rect 1269 -9672 1281 -9638
rect 1387 -9672 1399 -9638
rect -1445 -9678 -1387 -9672
rect -1327 -9678 -1269 -9672
rect -1209 -9678 -1151 -9672
rect -1091 -9678 -1033 -9672
rect -973 -9678 -915 -9672
rect -855 -9678 -797 -9672
rect -737 -9678 -679 -9672
rect -619 -9678 -561 -9672
rect -501 -9678 -443 -9672
rect -383 -9678 -325 -9672
rect -265 -9678 -207 -9672
rect -147 -9678 -89 -9672
rect -29 -9678 29 -9672
rect 89 -9678 147 -9672
rect 207 -9678 265 -9672
rect 325 -9678 383 -9672
rect 443 -9678 501 -9672
rect 561 -9678 619 -9672
rect 679 -9678 737 -9672
rect 797 -9678 855 -9672
rect 915 -9678 973 -9672
rect 1033 -9678 1091 -9672
rect 1151 -9678 1209 -9672
rect 1269 -9678 1327 -9672
rect 1387 -9678 1445 -9672
<< nmos >>
rect -1446 -9600 -1386 9600
rect -1328 -9600 -1268 9600
rect -1210 -9600 -1150 9600
rect -1092 -9600 -1032 9600
rect -974 -9600 -914 9600
rect -856 -9600 -796 9600
rect -738 -9600 -678 9600
rect -620 -9600 -560 9600
rect -502 -9600 -442 9600
rect -384 -9600 -324 9600
rect -266 -9600 -206 9600
rect -148 -9600 -88 9600
rect -30 -9600 30 9600
rect 88 -9600 148 9600
rect 206 -9600 266 9600
rect 324 -9600 384 9600
rect 442 -9600 502 9600
rect 560 -9600 620 9600
rect 678 -9600 738 9600
rect 796 -9600 856 9600
rect 914 -9600 974 9600
rect 1032 -9600 1092 9600
rect 1150 -9600 1210 9600
rect 1268 -9600 1328 9600
rect 1386 -9600 1446 9600
<< ndiff >>
rect -1504 9588 -1446 9600
rect -1504 -9588 -1492 9588
rect -1458 -9588 -1446 9588
rect -1504 -9600 -1446 -9588
rect -1386 9588 -1328 9600
rect -1386 -9588 -1374 9588
rect -1340 -9588 -1328 9588
rect -1386 -9600 -1328 -9588
rect -1268 9588 -1210 9600
rect -1268 -9588 -1256 9588
rect -1222 -9588 -1210 9588
rect -1268 -9600 -1210 -9588
rect -1150 9588 -1092 9600
rect -1150 -9588 -1138 9588
rect -1104 -9588 -1092 9588
rect -1150 -9600 -1092 -9588
rect -1032 9588 -974 9600
rect -1032 -9588 -1020 9588
rect -986 -9588 -974 9588
rect -1032 -9600 -974 -9588
rect -914 9588 -856 9600
rect -914 -9588 -902 9588
rect -868 -9588 -856 9588
rect -914 -9600 -856 -9588
rect -796 9588 -738 9600
rect -796 -9588 -784 9588
rect -750 -9588 -738 9588
rect -796 -9600 -738 -9588
rect -678 9588 -620 9600
rect -678 -9588 -666 9588
rect -632 -9588 -620 9588
rect -678 -9600 -620 -9588
rect -560 9588 -502 9600
rect -560 -9588 -548 9588
rect -514 -9588 -502 9588
rect -560 -9600 -502 -9588
rect -442 9588 -384 9600
rect -442 -9588 -430 9588
rect -396 -9588 -384 9588
rect -442 -9600 -384 -9588
rect -324 9588 -266 9600
rect -324 -9588 -312 9588
rect -278 -9588 -266 9588
rect -324 -9600 -266 -9588
rect -206 9588 -148 9600
rect -206 -9588 -194 9588
rect -160 -9588 -148 9588
rect -206 -9600 -148 -9588
rect -88 9588 -30 9600
rect -88 -9588 -76 9588
rect -42 -9588 -30 9588
rect -88 -9600 -30 -9588
rect 30 9588 88 9600
rect 30 -9588 42 9588
rect 76 -9588 88 9588
rect 30 -9600 88 -9588
rect 148 9588 206 9600
rect 148 -9588 160 9588
rect 194 -9588 206 9588
rect 148 -9600 206 -9588
rect 266 9588 324 9600
rect 266 -9588 278 9588
rect 312 -9588 324 9588
rect 266 -9600 324 -9588
rect 384 9588 442 9600
rect 384 -9588 396 9588
rect 430 -9588 442 9588
rect 384 -9600 442 -9588
rect 502 9588 560 9600
rect 502 -9588 514 9588
rect 548 -9588 560 9588
rect 502 -9600 560 -9588
rect 620 9588 678 9600
rect 620 -9588 632 9588
rect 666 -9588 678 9588
rect 620 -9600 678 -9588
rect 738 9588 796 9600
rect 738 -9588 750 9588
rect 784 -9588 796 9588
rect 738 -9600 796 -9588
rect 856 9588 914 9600
rect 856 -9588 868 9588
rect 902 -9588 914 9588
rect 856 -9600 914 -9588
rect 974 9588 1032 9600
rect 974 -9588 986 9588
rect 1020 -9588 1032 9588
rect 974 -9600 1032 -9588
rect 1092 9588 1150 9600
rect 1092 -9588 1104 9588
rect 1138 -9588 1150 9588
rect 1092 -9600 1150 -9588
rect 1210 9588 1268 9600
rect 1210 -9588 1222 9588
rect 1256 -9588 1268 9588
rect 1210 -9600 1268 -9588
rect 1328 9588 1386 9600
rect 1328 -9588 1340 9588
rect 1374 -9588 1386 9588
rect 1328 -9600 1386 -9588
rect 1446 9588 1504 9600
rect 1446 -9588 1458 9588
rect 1492 -9588 1504 9588
rect 1446 -9600 1504 -9588
<< ndiffc >>
rect -1492 -9588 -1458 9588
rect -1374 -9588 -1340 9588
rect -1256 -9588 -1222 9588
rect -1138 -9588 -1104 9588
rect -1020 -9588 -986 9588
rect -902 -9588 -868 9588
rect -784 -9588 -750 9588
rect -666 -9588 -632 9588
rect -548 -9588 -514 9588
rect -430 -9588 -396 9588
rect -312 -9588 -278 9588
rect -194 -9588 -160 9588
rect -76 -9588 -42 9588
rect 42 -9588 76 9588
rect 160 -9588 194 9588
rect 278 -9588 312 9588
rect 396 -9588 430 9588
rect 514 -9588 548 9588
rect 632 -9588 666 9588
rect 750 -9588 784 9588
rect 868 -9588 902 9588
rect 986 -9588 1020 9588
rect 1104 -9588 1138 9588
rect 1222 -9588 1256 9588
rect 1340 -9588 1374 9588
rect 1458 -9588 1492 9588
<< poly >>
rect -1449 9672 -1383 9688
rect -1449 9638 -1433 9672
rect -1399 9638 -1383 9672
rect -1449 9622 -1383 9638
rect -1331 9672 -1265 9688
rect -1331 9638 -1315 9672
rect -1281 9638 -1265 9672
rect -1331 9622 -1265 9638
rect -1213 9672 -1147 9688
rect -1213 9638 -1197 9672
rect -1163 9638 -1147 9672
rect -1213 9622 -1147 9638
rect -1095 9672 -1029 9688
rect -1095 9638 -1079 9672
rect -1045 9638 -1029 9672
rect -1095 9622 -1029 9638
rect -977 9672 -911 9688
rect -977 9638 -961 9672
rect -927 9638 -911 9672
rect -977 9622 -911 9638
rect -859 9672 -793 9688
rect -859 9638 -843 9672
rect -809 9638 -793 9672
rect -859 9622 -793 9638
rect -741 9672 -675 9688
rect -741 9638 -725 9672
rect -691 9638 -675 9672
rect -741 9622 -675 9638
rect -623 9672 -557 9688
rect -623 9638 -607 9672
rect -573 9638 -557 9672
rect -623 9622 -557 9638
rect -505 9672 -439 9688
rect -505 9638 -489 9672
rect -455 9638 -439 9672
rect -505 9622 -439 9638
rect -387 9672 -321 9688
rect -387 9638 -371 9672
rect -337 9638 -321 9672
rect -387 9622 -321 9638
rect -269 9672 -203 9688
rect -269 9638 -253 9672
rect -219 9638 -203 9672
rect -269 9622 -203 9638
rect -151 9672 -85 9688
rect -151 9638 -135 9672
rect -101 9638 -85 9672
rect -151 9622 -85 9638
rect -33 9672 33 9688
rect -33 9638 -17 9672
rect 17 9638 33 9672
rect -33 9622 33 9638
rect 85 9672 151 9688
rect 85 9638 101 9672
rect 135 9638 151 9672
rect 85 9622 151 9638
rect 203 9672 269 9688
rect 203 9638 219 9672
rect 253 9638 269 9672
rect 203 9622 269 9638
rect 321 9672 387 9688
rect 321 9638 337 9672
rect 371 9638 387 9672
rect 321 9622 387 9638
rect 439 9672 505 9688
rect 439 9638 455 9672
rect 489 9638 505 9672
rect 439 9622 505 9638
rect 557 9672 623 9688
rect 557 9638 573 9672
rect 607 9638 623 9672
rect 557 9622 623 9638
rect 675 9672 741 9688
rect 675 9638 691 9672
rect 725 9638 741 9672
rect 675 9622 741 9638
rect 793 9672 859 9688
rect 793 9638 809 9672
rect 843 9638 859 9672
rect 793 9622 859 9638
rect 911 9672 977 9688
rect 911 9638 927 9672
rect 961 9638 977 9672
rect 911 9622 977 9638
rect 1029 9672 1095 9688
rect 1029 9638 1045 9672
rect 1079 9638 1095 9672
rect 1029 9622 1095 9638
rect 1147 9672 1213 9688
rect 1147 9638 1163 9672
rect 1197 9638 1213 9672
rect 1147 9622 1213 9638
rect 1265 9672 1331 9688
rect 1265 9638 1281 9672
rect 1315 9638 1331 9672
rect 1265 9622 1331 9638
rect 1383 9672 1449 9688
rect 1383 9638 1399 9672
rect 1433 9638 1449 9672
rect 1383 9622 1449 9638
rect -1446 9600 -1386 9622
rect -1328 9600 -1268 9622
rect -1210 9600 -1150 9622
rect -1092 9600 -1032 9622
rect -974 9600 -914 9622
rect -856 9600 -796 9622
rect -738 9600 -678 9622
rect -620 9600 -560 9622
rect -502 9600 -442 9622
rect -384 9600 -324 9622
rect -266 9600 -206 9622
rect -148 9600 -88 9622
rect -30 9600 30 9622
rect 88 9600 148 9622
rect 206 9600 266 9622
rect 324 9600 384 9622
rect 442 9600 502 9622
rect 560 9600 620 9622
rect 678 9600 738 9622
rect 796 9600 856 9622
rect 914 9600 974 9622
rect 1032 9600 1092 9622
rect 1150 9600 1210 9622
rect 1268 9600 1328 9622
rect 1386 9600 1446 9622
rect -1446 -9622 -1386 -9600
rect -1328 -9622 -1268 -9600
rect -1210 -9622 -1150 -9600
rect -1092 -9622 -1032 -9600
rect -974 -9622 -914 -9600
rect -856 -9622 -796 -9600
rect -738 -9622 -678 -9600
rect -620 -9622 -560 -9600
rect -502 -9622 -442 -9600
rect -384 -9622 -324 -9600
rect -266 -9622 -206 -9600
rect -148 -9622 -88 -9600
rect -30 -9622 30 -9600
rect 88 -9622 148 -9600
rect 206 -9622 266 -9600
rect 324 -9622 384 -9600
rect 442 -9622 502 -9600
rect 560 -9622 620 -9600
rect 678 -9622 738 -9600
rect 796 -9622 856 -9600
rect 914 -9622 974 -9600
rect 1032 -9622 1092 -9600
rect 1150 -9622 1210 -9600
rect 1268 -9622 1328 -9600
rect 1386 -9622 1446 -9600
rect -1449 -9638 -1383 -9622
rect -1449 -9672 -1433 -9638
rect -1399 -9672 -1383 -9638
rect -1449 -9688 -1383 -9672
rect -1331 -9638 -1265 -9622
rect -1331 -9672 -1315 -9638
rect -1281 -9672 -1265 -9638
rect -1331 -9688 -1265 -9672
rect -1213 -9638 -1147 -9622
rect -1213 -9672 -1197 -9638
rect -1163 -9672 -1147 -9638
rect -1213 -9688 -1147 -9672
rect -1095 -9638 -1029 -9622
rect -1095 -9672 -1079 -9638
rect -1045 -9672 -1029 -9638
rect -1095 -9688 -1029 -9672
rect -977 -9638 -911 -9622
rect -977 -9672 -961 -9638
rect -927 -9672 -911 -9638
rect -977 -9688 -911 -9672
rect -859 -9638 -793 -9622
rect -859 -9672 -843 -9638
rect -809 -9672 -793 -9638
rect -859 -9688 -793 -9672
rect -741 -9638 -675 -9622
rect -741 -9672 -725 -9638
rect -691 -9672 -675 -9638
rect -741 -9688 -675 -9672
rect -623 -9638 -557 -9622
rect -623 -9672 -607 -9638
rect -573 -9672 -557 -9638
rect -623 -9688 -557 -9672
rect -505 -9638 -439 -9622
rect -505 -9672 -489 -9638
rect -455 -9672 -439 -9638
rect -505 -9688 -439 -9672
rect -387 -9638 -321 -9622
rect -387 -9672 -371 -9638
rect -337 -9672 -321 -9638
rect -387 -9688 -321 -9672
rect -269 -9638 -203 -9622
rect -269 -9672 -253 -9638
rect -219 -9672 -203 -9638
rect -269 -9688 -203 -9672
rect -151 -9638 -85 -9622
rect -151 -9672 -135 -9638
rect -101 -9672 -85 -9638
rect -151 -9688 -85 -9672
rect -33 -9638 33 -9622
rect -33 -9672 -17 -9638
rect 17 -9672 33 -9638
rect -33 -9688 33 -9672
rect 85 -9638 151 -9622
rect 85 -9672 101 -9638
rect 135 -9672 151 -9638
rect 85 -9688 151 -9672
rect 203 -9638 269 -9622
rect 203 -9672 219 -9638
rect 253 -9672 269 -9638
rect 203 -9688 269 -9672
rect 321 -9638 387 -9622
rect 321 -9672 337 -9638
rect 371 -9672 387 -9638
rect 321 -9688 387 -9672
rect 439 -9638 505 -9622
rect 439 -9672 455 -9638
rect 489 -9672 505 -9638
rect 439 -9688 505 -9672
rect 557 -9638 623 -9622
rect 557 -9672 573 -9638
rect 607 -9672 623 -9638
rect 557 -9688 623 -9672
rect 675 -9638 741 -9622
rect 675 -9672 691 -9638
rect 725 -9672 741 -9638
rect 675 -9688 741 -9672
rect 793 -9638 859 -9622
rect 793 -9672 809 -9638
rect 843 -9672 859 -9638
rect 793 -9688 859 -9672
rect 911 -9638 977 -9622
rect 911 -9672 927 -9638
rect 961 -9672 977 -9638
rect 911 -9688 977 -9672
rect 1029 -9638 1095 -9622
rect 1029 -9672 1045 -9638
rect 1079 -9672 1095 -9638
rect 1029 -9688 1095 -9672
rect 1147 -9638 1213 -9622
rect 1147 -9672 1163 -9638
rect 1197 -9672 1213 -9638
rect 1147 -9688 1213 -9672
rect 1265 -9638 1331 -9622
rect 1265 -9672 1281 -9638
rect 1315 -9672 1331 -9638
rect 1265 -9688 1331 -9672
rect 1383 -9638 1449 -9622
rect 1383 -9672 1399 -9638
rect 1433 -9672 1449 -9638
rect 1383 -9688 1449 -9672
<< polycont >>
rect -1433 9638 -1399 9672
rect -1315 9638 -1281 9672
rect -1197 9638 -1163 9672
rect -1079 9638 -1045 9672
rect -961 9638 -927 9672
rect -843 9638 -809 9672
rect -725 9638 -691 9672
rect -607 9638 -573 9672
rect -489 9638 -455 9672
rect -371 9638 -337 9672
rect -253 9638 -219 9672
rect -135 9638 -101 9672
rect -17 9638 17 9672
rect 101 9638 135 9672
rect 219 9638 253 9672
rect 337 9638 371 9672
rect 455 9638 489 9672
rect 573 9638 607 9672
rect 691 9638 725 9672
rect 809 9638 843 9672
rect 927 9638 961 9672
rect 1045 9638 1079 9672
rect 1163 9638 1197 9672
rect 1281 9638 1315 9672
rect 1399 9638 1433 9672
rect -1433 -9672 -1399 -9638
rect -1315 -9672 -1281 -9638
rect -1197 -9672 -1163 -9638
rect -1079 -9672 -1045 -9638
rect -961 -9672 -927 -9638
rect -843 -9672 -809 -9638
rect -725 -9672 -691 -9638
rect -607 -9672 -573 -9638
rect -489 -9672 -455 -9638
rect -371 -9672 -337 -9638
rect -253 -9672 -219 -9638
rect -135 -9672 -101 -9638
rect -17 -9672 17 -9638
rect 101 -9672 135 -9638
rect 219 -9672 253 -9638
rect 337 -9672 371 -9638
rect 455 -9672 489 -9638
rect 573 -9672 607 -9638
rect 691 -9672 725 -9638
rect 809 -9672 843 -9638
rect 927 -9672 961 -9638
rect 1045 -9672 1079 -9638
rect 1163 -9672 1197 -9638
rect 1281 -9672 1315 -9638
rect 1399 -9672 1433 -9638
<< locali >>
rect -1449 9638 -1433 9672
rect -1399 9638 -1383 9672
rect -1331 9638 -1315 9672
rect -1281 9638 -1265 9672
rect -1213 9638 -1197 9672
rect -1163 9638 -1147 9672
rect -1095 9638 -1079 9672
rect -1045 9638 -1029 9672
rect -977 9638 -961 9672
rect -927 9638 -911 9672
rect -859 9638 -843 9672
rect -809 9638 -793 9672
rect -741 9638 -725 9672
rect -691 9638 -675 9672
rect -623 9638 -607 9672
rect -573 9638 -557 9672
rect -505 9638 -489 9672
rect -455 9638 -439 9672
rect -387 9638 -371 9672
rect -337 9638 -321 9672
rect -269 9638 -253 9672
rect -219 9638 -203 9672
rect -151 9638 -135 9672
rect -101 9638 -85 9672
rect -33 9638 -17 9672
rect 17 9638 33 9672
rect 85 9638 101 9672
rect 135 9638 151 9672
rect 203 9638 219 9672
rect 253 9638 269 9672
rect 321 9638 337 9672
rect 371 9638 387 9672
rect 439 9638 455 9672
rect 489 9638 505 9672
rect 557 9638 573 9672
rect 607 9638 623 9672
rect 675 9638 691 9672
rect 725 9638 741 9672
rect 793 9638 809 9672
rect 843 9638 859 9672
rect 911 9638 927 9672
rect 961 9638 977 9672
rect 1029 9638 1045 9672
rect 1079 9638 1095 9672
rect 1147 9638 1163 9672
rect 1197 9638 1213 9672
rect 1265 9638 1281 9672
rect 1315 9638 1331 9672
rect 1383 9638 1399 9672
rect 1433 9638 1449 9672
rect -1492 9588 -1458 9604
rect -1492 -9604 -1458 -9588
rect -1374 9588 -1340 9604
rect -1374 -9604 -1340 -9588
rect -1256 9588 -1222 9604
rect -1256 -9604 -1222 -9588
rect -1138 9588 -1104 9604
rect -1138 -9604 -1104 -9588
rect -1020 9588 -986 9604
rect -1020 -9604 -986 -9588
rect -902 9588 -868 9604
rect -902 -9604 -868 -9588
rect -784 9588 -750 9604
rect -784 -9604 -750 -9588
rect -666 9588 -632 9604
rect -666 -9604 -632 -9588
rect -548 9588 -514 9604
rect -548 -9604 -514 -9588
rect -430 9588 -396 9604
rect -430 -9604 -396 -9588
rect -312 9588 -278 9604
rect -312 -9604 -278 -9588
rect -194 9588 -160 9604
rect -194 -9604 -160 -9588
rect -76 9588 -42 9604
rect -76 -9604 -42 -9588
rect 42 9588 76 9604
rect 42 -9604 76 -9588
rect 160 9588 194 9604
rect 160 -9604 194 -9588
rect 278 9588 312 9604
rect 278 -9604 312 -9588
rect 396 9588 430 9604
rect 396 -9604 430 -9588
rect 514 9588 548 9604
rect 514 -9604 548 -9588
rect 632 9588 666 9604
rect 632 -9604 666 -9588
rect 750 9588 784 9604
rect 750 -9604 784 -9588
rect 868 9588 902 9604
rect 868 -9604 902 -9588
rect 986 9588 1020 9604
rect 986 -9604 1020 -9588
rect 1104 9588 1138 9604
rect 1104 -9604 1138 -9588
rect 1222 9588 1256 9604
rect 1222 -9604 1256 -9588
rect 1340 9588 1374 9604
rect 1340 -9604 1374 -9588
rect 1458 9588 1492 9604
rect 1458 -9604 1492 -9588
rect -1449 -9672 -1433 -9638
rect -1399 -9672 -1383 -9638
rect -1331 -9672 -1315 -9638
rect -1281 -9672 -1265 -9638
rect -1213 -9672 -1197 -9638
rect -1163 -9672 -1147 -9638
rect -1095 -9672 -1079 -9638
rect -1045 -9672 -1029 -9638
rect -977 -9672 -961 -9638
rect -927 -9672 -911 -9638
rect -859 -9672 -843 -9638
rect -809 -9672 -793 -9638
rect -741 -9672 -725 -9638
rect -691 -9672 -675 -9638
rect -623 -9672 -607 -9638
rect -573 -9672 -557 -9638
rect -505 -9672 -489 -9638
rect -455 -9672 -439 -9638
rect -387 -9672 -371 -9638
rect -337 -9672 -321 -9638
rect -269 -9672 -253 -9638
rect -219 -9672 -203 -9638
rect -151 -9672 -135 -9638
rect -101 -9672 -85 -9638
rect -33 -9672 -17 -9638
rect 17 -9672 33 -9638
rect 85 -9672 101 -9638
rect 135 -9672 151 -9638
rect 203 -9672 219 -9638
rect 253 -9672 269 -9638
rect 321 -9672 337 -9638
rect 371 -9672 387 -9638
rect 439 -9672 455 -9638
rect 489 -9672 505 -9638
rect 557 -9672 573 -9638
rect 607 -9672 623 -9638
rect 675 -9672 691 -9638
rect 725 -9672 741 -9638
rect 793 -9672 809 -9638
rect 843 -9672 859 -9638
rect 911 -9672 927 -9638
rect 961 -9672 977 -9638
rect 1029 -9672 1045 -9638
rect 1079 -9672 1095 -9638
rect 1147 -9672 1163 -9638
rect 1197 -9672 1213 -9638
rect 1265 -9672 1281 -9638
rect 1315 -9672 1331 -9638
rect 1383 -9672 1399 -9638
rect 1433 -9672 1449 -9638
<< viali >>
rect -1433 9638 -1399 9672
rect -1315 9638 -1281 9672
rect -1197 9638 -1163 9672
rect -1079 9638 -1045 9672
rect -961 9638 -927 9672
rect -843 9638 -809 9672
rect -725 9638 -691 9672
rect -607 9638 -573 9672
rect -489 9638 -455 9672
rect -371 9638 -337 9672
rect -253 9638 -219 9672
rect -135 9638 -101 9672
rect -17 9638 17 9672
rect 101 9638 135 9672
rect 219 9638 253 9672
rect 337 9638 371 9672
rect 455 9638 489 9672
rect 573 9638 607 9672
rect 691 9638 725 9672
rect 809 9638 843 9672
rect 927 9638 961 9672
rect 1045 9638 1079 9672
rect 1163 9638 1197 9672
rect 1281 9638 1315 9672
rect 1399 9638 1433 9672
rect -1492 -9588 -1458 9588
rect -1374 -9588 -1340 9588
rect -1256 -9588 -1222 9588
rect -1138 -9588 -1104 9588
rect -1020 -9588 -986 9588
rect -902 -9588 -868 9588
rect -784 -9588 -750 9588
rect -666 -9588 -632 9588
rect -548 -9588 -514 9588
rect -430 -9588 -396 9588
rect -312 -9588 -278 9588
rect -194 -9588 -160 9588
rect -76 -9588 -42 9588
rect 42 -9588 76 9588
rect 160 -9588 194 9588
rect 278 -9588 312 9588
rect 396 -9588 430 9588
rect 514 -9588 548 9588
rect 632 -9588 666 9588
rect 750 -9588 784 9588
rect 868 -9588 902 9588
rect 986 -9588 1020 9588
rect 1104 -9588 1138 9588
rect 1222 -9588 1256 9588
rect 1340 -9588 1374 9588
rect 1458 -9588 1492 9588
rect -1433 -9672 -1399 -9638
rect -1315 -9672 -1281 -9638
rect -1197 -9672 -1163 -9638
rect -1079 -9672 -1045 -9638
rect -961 -9672 -927 -9638
rect -843 -9672 -809 -9638
rect -725 -9672 -691 -9638
rect -607 -9672 -573 -9638
rect -489 -9672 -455 -9638
rect -371 -9672 -337 -9638
rect -253 -9672 -219 -9638
rect -135 -9672 -101 -9638
rect -17 -9672 17 -9638
rect 101 -9672 135 -9638
rect 219 -9672 253 -9638
rect 337 -9672 371 -9638
rect 455 -9672 489 -9638
rect 573 -9672 607 -9638
rect 691 -9672 725 -9638
rect 809 -9672 843 -9638
rect 927 -9672 961 -9638
rect 1045 -9672 1079 -9638
rect 1163 -9672 1197 -9638
rect 1281 -9672 1315 -9638
rect 1399 -9672 1433 -9638
<< metal1 >>
rect -1445 9672 -1387 9678
rect -1445 9638 -1433 9672
rect -1399 9638 -1387 9672
rect -1445 9632 -1387 9638
rect -1327 9672 -1269 9678
rect -1327 9638 -1315 9672
rect -1281 9638 -1269 9672
rect -1327 9632 -1269 9638
rect -1209 9672 -1151 9678
rect -1209 9638 -1197 9672
rect -1163 9638 -1151 9672
rect -1209 9632 -1151 9638
rect -1091 9672 -1033 9678
rect -1091 9638 -1079 9672
rect -1045 9638 -1033 9672
rect -1091 9632 -1033 9638
rect -973 9672 -915 9678
rect -973 9638 -961 9672
rect -927 9638 -915 9672
rect -973 9632 -915 9638
rect -855 9672 -797 9678
rect -855 9638 -843 9672
rect -809 9638 -797 9672
rect -855 9632 -797 9638
rect -737 9672 -679 9678
rect -737 9638 -725 9672
rect -691 9638 -679 9672
rect -737 9632 -679 9638
rect -619 9672 -561 9678
rect -619 9638 -607 9672
rect -573 9638 -561 9672
rect -619 9632 -561 9638
rect -501 9672 -443 9678
rect -501 9638 -489 9672
rect -455 9638 -443 9672
rect -501 9632 -443 9638
rect -383 9672 -325 9678
rect -383 9638 -371 9672
rect -337 9638 -325 9672
rect -383 9632 -325 9638
rect -265 9672 -207 9678
rect -265 9638 -253 9672
rect -219 9638 -207 9672
rect -265 9632 -207 9638
rect -147 9672 -89 9678
rect -147 9638 -135 9672
rect -101 9638 -89 9672
rect -147 9632 -89 9638
rect -29 9672 29 9678
rect -29 9638 -17 9672
rect 17 9638 29 9672
rect -29 9632 29 9638
rect 89 9672 147 9678
rect 89 9638 101 9672
rect 135 9638 147 9672
rect 89 9632 147 9638
rect 207 9672 265 9678
rect 207 9638 219 9672
rect 253 9638 265 9672
rect 207 9632 265 9638
rect 325 9672 383 9678
rect 325 9638 337 9672
rect 371 9638 383 9672
rect 325 9632 383 9638
rect 443 9672 501 9678
rect 443 9638 455 9672
rect 489 9638 501 9672
rect 443 9632 501 9638
rect 561 9672 619 9678
rect 561 9638 573 9672
rect 607 9638 619 9672
rect 561 9632 619 9638
rect 679 9672 737 9678
rect 679 9638 691 9672
rect 725 9638 737 9672
rect 679 9632 737 9638
rect 797 9672 855 9678
rect 797 9638 809 9672
rect 843 9638 855 9672
rect 797 9632 855 9638
rect 915 9672 973 9678
rect 915 9638 927 9672
rect 961 9638 973 9672
rect 915 9632 973 9638
rect 1033 9672 1091 9678
rect 1033 9638 1045 9672
rect 1079 9638 1091 9672
rect 1033 9632 1091 9638
rect 1151 9672 1209 9678
rect 1151 9638 1163 9672
rect 1197 9638 1209 9672
rect 1151 9632 1209 9638
rect 1269 9672 1327 9678
rect 1269 9638 1281 9672
rect 1315 9638 1327 9672
rect 1269 9632 1327 9638
rect 1387 9672 1445 9678
rect 1387 9638 1399 9672
rect 1433 9638 1445 9672
rect 1387 9632 1445 9638
rect -1498 9588 -1452 9600
rect -1498 -9588 -1492 9588
rect -1458 -9588 -1452 9588
rect -1498 -9600 -1452 -9588
rect -1380 9588 -1334 9600
rect -1380 -9588 -1374 9588
rect -1340 -9588 -1334 9588
rect -1380 -9600 -1334 -9588
rect -1262 9588 -1216 9600
rect -1262 -9588 -1256 9588
rect -1222 -9588 -1216 9588
rect -1262 -9600 -1216 -9588
rect -1144 9588 -1098 9600
rect -1144 -9588 -1138 9588
rect -1104 -9588 -1098 9588
rect -1144 -9600 -1098 -9588
rect -1026 9588 -980 9600
rect -1026 -9588 -1020 9588
rect -986 -9588 -980 9588
rect -1026 -9600 -980 -9588
rect -908 9588 -862 9600
rect -908 -9588 -902 9588
rect -868 -9588 -862 9588
rect -908 -9600 -862 -9588
rect -790 9588 -744 9600
rect -790 -9588 -784 9588
rect -750 -9588 -744 9588
rect -790 -9600 -744 -9588
rect -672 9588 -626 9600
rect -672 -9588 -666 9588
rect -632 -9588 -626 9588
rect -672 -9600 -626 -9588
rect -554 9588 -508 9600
rect -554 -9588 -548 9588
rect -514 -9588 -508 9588
rect -554 -9600 -508 -9588
rect -436 9588 -390 9600
rect -436 -9588 -430 9588
rect -396 -9588 -390 9588
rect -436 -9600 -390 -9588
rect -318 9588 -272 9600
rect -318 -9588 -312 9588
rect -278 -9588 -272 9588
rect -318 -9600 -272 -9588
rect -200 9588 -154 9600
rect -200 -9588 -194 9588
rect -160 -9588 -154 9588
rect -200 -9600 -154 -9588
rect -82 9588 -36 9600
rect -82 -9588 -76 9588
rect -42 -9588 -36 9588
rect -82 -9600 -36 -9588
rect 36 9588 82 9600
rect 36 -9588 42 9588
rect 76 -9588 82 9588
rect 36 -9600 82 -9588
rect 154 9588 200 9600
rect 154 -9588 160 9588
rect 194 -9588 200 9588
rect 154 -9600 200 -9588
rect 272 9588 318 9600
rect 272 -9588 278 9588
rect 312 -9588 318 9588
rect 272 -9600 318 -9588
rect 390 9588 436 9600
rect 390 -9588 396 9588
rect 430 -9588 436 9588
rect 390 -9600 436 -9588
rect 508 9588 554 9600
rect 508 -9588 514 9588
rect 548 -9588 554 9588
rect 508 -9600 554 -9588
rect 626 9588 672 9600
rect 626 -9588 632 9588
rect 666 -9588 672 9588
rect 626 -9600 672 -9588
rect 744 9588 790 9600
rect 744 -9588 750 9588
rect 784 -9588 790 9588
rect 744 -9600 790 -9588
rect 862 9588 908 9600
rect 862 -9588 868 9588
rect 902 -9588 908 9588
rect 862 -9600 908 -9588
rect 980 9588 1026 9600
rect 980 -9588 986 9588
rect 1020 -9588 1026 9588
rect 980 -9600 1026 -9588
rect 1098 9588 1144 9600
rect 1098 -9588 1104 9588
rect 1138 -9588 1144 9588
rect 1098 -9600 1144 -9588
rect 1216 9588 1262 9600
rect 1216 -9588 1222 9588
rect 1256 -9588 1262 9588
rect 1216 -9600 1262 -9588
rect 1334 9588 1380 9600
rect 1334 -9588 1340 9588
rect 1374 -9588 1380 9588
rect 1334 -9600 1380 -9588
rect 1452 9588 1498 9600
rect 1452 -9588 1458 9588
rect 1492 -9588 1498 9588
rect 1452 -9600 1498 -9588
rect -1445 -9638 -1387 -9632
rect -1445 -9672 -1433 -9638
rect -1399 -9672 -1387 -9638
rect -1445 -9678 -1387 -9672
rect -1327 -9638 -1269 -9632
rect -1327 -9672 -1315 -9638
rect -1281 -9672 -1269 -9638
rect -1327 -9678 -1269 -9672
rect -1209 -9638 -1151 -9632
rect -1209 -9672 -1197 -9638
rect -1163 -9672 -1151 -9638
rect -1209 -9678 -1151 -9672
rect -1091 -9638 -1033 -9632
rect -1091 -9672 -1079 -9638
rect -1045 -9672 -1033 -9638
rect -1091 -9678 -1033 -9672
rect -973 -9638 -915 -9632
rect -973 -9672 -961 -9638
rect -927 -9672 -915 -9638
rect -973 -9678 -915 -9672
rect -855 -9638 -797 -9632
rect -855 -9672 -843 -9638
rect -809 -9672 -797 -9638
rect -855 -9678 -797 -9672
rect -737 -9638 -679 -9632
rect -737 -9672 -725 -9638
rect -691 -9672 -679 -9638
rect -737 -9678 -679 -9672
rect -619 -9638 -561 -9632
rect -619 -9672 -607 -9638
rect -573 -9672 -561 -9638
rect -619 -9678 -561 -9672
rect -501 -9638 -443 -9632
rect -501 -9672 -489 -9638
rect -455 -9672 -443 -9638
rect -501 -9678 -443 -9672
rect -383 -9638 -325 -9632
rect -383 -9672 -371 -9638
rect -337 -9672 -325 -9638
rect -383 -9678 -325 -9672
rect -265 -9638 -207 -9632
rect -265 -9672 -253 -9638
rect -219 -9672 -207 -9638
rect -265 -9678 -207 -9672
rect -147 -9638 -89 -9632
rect -147 -9672 -135 -9638
rect -101 -9672 -89 -9638
rect -147 -9678 -89 -9672
rect -29 -9638 29 -9632
rect -29 -9672 -17 -9638
rect 17 -9672 29 -9638
rect -29 -9678 29 -9672
rect 89 -9638 147 -9632
rect 89 -9672 101 -9638
rect 135 -9672 147 -9638
rect 89 -9678 147 -9672
rect 207 -9638 265 -9632
rect 207 -9672 219 -9638
rect 253 -9672 265 -9638
rect 207 -9678 265 -9672
rect 325 -9638 383 -9632
rect 325 -9672 337 -9638
rect 371 -9672 383 -9638
rect 325 -9678 383 -9672
rect 443 -9638 501 -9632
rect 443 -9672 455 -9638
rect 489 -9672 501 -9638
rect 443 -9678 501 -9672
rect 561 -9638 619 -9632
rect 561 -9672 573 -9638
rect 607 -9672 619 -9638
rect 561 -9678 619 -9672
rect 679 -9638 737 -9632
rect 679 -9672 691 -9638
rect 725 -9672 737 -9638
rect 679 -9678 737 -9672
rect 797 -9638 855 -9632
rect 797 -9672 809 -9638
rect 843 -9672 855 -9638
rect 797 -9678 855 -9672
rect 915 -9638 973 -9632
rect 915 -9672 927 -9638
rect 961 -9672 973 -9638
rect 915 -9678 973 -9672
rect 1033 -9638 1091 -9632
rect 1033 -9672 1045 -9638
rect 1079 -9672 1091 -9638
rect 1033 -9678 1091 -9672
rect 1151 -9638 1209 -9632
rect 1151 -9672 1163 -9638
rect 1197 -9672 1209 -9638
rect 1151 -9678 1209 -9672
rect 1269 -9638 1327 -9632
rect 1269 -9672 1281 -9638
rect 1315 -9672 1327 -9638
rect 1269 -9678 1327 -9672
rect 1387 -9638 1445 -9632
rect 1387 -9672 1399 -9638
rect 1433 -9672 1445 -9638
rect 1387 -9678 1445 -9672
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 96 l 0.3 m 1 nf 25 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
