magic
tech sky130A
magscale 1 2
timestamp 1667831724
<< error_p >>
rect -527 1018 -463 1024
rect -527 984 -515 1018
rect -527 978 -463 984
<< nmos >>
rect -531 -903 -459 903
rect -361 -903 -289 903
rect -231 -903 -159 903
rect -101 -903 -29 903
rect 29 -903 101 903
rect 159 -903 231 903
rect 289 -903 361 903
rect 419 -903 491 903
<< ndiff >>
rect -589 891 -531 903
rect -589 -891 -577 891
rect -543 -891 -531 891
rect -589 -903 -531 -891
rect -459 891 -361 903
rect -459 -891 -445 891
rect -373 -891 -361 891
rect -459 -903 -361 -891
rect -289 891 -231 903
rect -289 -891 -277 891
rect -243 -891 -231 891
rect -289 -903 -231 -891
rect -159 891 -101 903
rect -159 -891 -147 891
rect -113 -891 -101 891
rect -159 -903 -101 -891
rect -29 891 29 903
rect -29 -891 -17 891
rect 17 -891 29 891
rect -29 -903 29 -891
rect 101 891 159 903
rect 101 -891 113 891
rect 147 -891 159 891
rect 101 -903 159 -891
rect 231 891 289 903
rect 231 -891 243 891
rect 277 -891 289 891
rect 231 -903 289 -891
rect 361 891 419 903
rect 361 -891 373 891
rect 407 -891 419 891
rect 361 -903 419 -891
rect 491 891 549 903
rect 491 -891 503 891
rect 537 -891 549 891
rect 491 -903 549 -891
<< ndiffc >>
rect -577 -891 -543 891
rect -445 -891 -373 891
rect -277 -891 -243 891
rect -147 -891 -113 891
rect -17 -891 17 891
rect 113 -891 147 891
rect 243 -891 277 891
rect 373 -891 407 891
rect 503 -891 537 891
<< poly >>
rect -531 1018 -459 1034
rect -531 984 -515 1018
rect -475 984 -459 1018
rect -531 903 -459 984
rect -361 927 -159 979
rect -361 903 -289 927
rect -231 903 -159 927
rect -101 927 101 979
rect -101 903 -29 927
rect 29 903 101 927
rect 159 927 361 979
rect 159 903 231 927
rect 289 903 361 927
rect 419 903 491 930
rect -531 -931 -459 -903
rect -361 -931 -289 -903
rect -531 -983 -289 -931
rect -231 -931 -159 -903
rect -101 -931 -29 -903
rect -231 -983 -29 -931
rect 29 -931 101 -903
rect 159 -931 231 -903
rect 29 -983 231 -931
rect 289 -931 361 -903
rect 419 -931 491 -903
rect 289 -983 491 -931
<< polycont >>
rect -515 984 -475 1018
<< locali >>
rect -531 984 -515 1018
rect -475 984 -459 1018
rect -577 891 -543 907
rect -577 -907 -543 -891
rect -445 891 -373 907
rect -445 -907 -373 -891
rect -277 891 -243 907
rect -277 -907 -243 -891
rect -147 891 -113 907
rect -147 -907 -113 -891
rect -17 891 17 907
rect -17 -907 17 -891
rect 113 891 147 907
rect 113 -907 147 -891
rect 243 891 277 907
rect 243 -907 277 -891
rect 373 891 407 907
rect 373 -907 407 -891
rect 503 891 537 907
rect 503 -907 537 -891
<< viali >>
rect -515 984 -475 1018
rect -577 -891 -543 891
rect -445 -891 -373 891
rect -277 -891 -243 891
rect -147 -891 -113 891
rect -17 -891 17 891
rect 113 -891 147 891
rect 243 -891 277 891
rect 373 -891 407 891
rect 503 -891 537 891
<< metal1 >>
rect -527 1018 -463 1024
rect -527 984 -515 1018
rect -475 984 -463 1018
rect -527 978 -463 984
rect -583 891 -537 903
rect -583 -891 -577 891
rect -543 -891 -537 891
rect -583 -903 -537 -891
rect -453 891 -367 903
rect -453 -891 -445 891
rect -373 -891 -367 891
rect -453 -903 -367 -891
rect -283 891 -237 903
rect -283 -891 -277 891
rect -243 -891 -237 891
rect -283 -903 -237 -891
rect -153 891 -107 903
rect -153 -891 -147 891
rect -113 -891 -107 891
rect -153 -903 -107 -891
rect -23 891 23 903
rect -23 -891 -17 891
rect 17 -891 23 891
rect -23 -903 23 -891
rect 107 891 153 903
rect 107 -891 113 891
rect 147 -891 153 891
rect 107 -903 153 -891
rect 237 891 283 903
rect 237 -891 243 891
rect 277 -891 283 891
rect 237 -903 283 -891
rect 367 891 413 903
rect 367 -891 373 891
rect 407 -891 413 891
rect 367 -903 413 -891
rect 497 891 543 903
rect 497 -891 503 891
rect 537 -891 543 891
rect 497 -903 543 -891
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 9.03 l 0.361 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
