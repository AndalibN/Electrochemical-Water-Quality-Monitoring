magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -323 -1498 323 1464
<< pmos >>
rect -229 -1436 -29 1364
rect 29 -1436 229 1364
<< pdiff >>
rect -287 1341 -229 1364
rect -287 1307 -275 1341
rect -241 1307 -229 1341
rect -287 1273 -229 1307
rect -287 1239 -275 1273
rect -241 1239 -229 1273
rect -287 1205 -229 1239
rect -287 1171 -275 1205
rect -241 1171 -229 1205
rect -287 1137 -229 1171
rect -287 1103 -275 1137
rect -241 1103 -229 1137
rect -287 1069 -229 1103
rect -287 1035 -275 1069
rect -241 1035 -229 1069
rect -287 1001 -229 1035
rect -287 967 -275 1001
rect -241 967 -229 1001
rect -287 933 -229 967
rect -287 899 -275 933
rect -241 899 -229 933
rect -287 865 -229 899
rect -287 831 -275 865
rect -241 831 -229 865
rect -287 797 -229 831
rect -287 763 -275 797
rect -241 763 -229 797
rect -287 729 -229 763
rect -287 695 -275 729
rect -241 695 -229 729
rect -287 661 -229 695
rect -287 627 -275 661
rect -241 627 -229 661
rect -287 593 -229 627
rect -287 559 -275 593
rect -241 559 -229 593
rect -287 525 -229 559
rect -287 491 -275 525
rect -241 491 -229 525
rect -287 457 -229 491
rect -287 423 -275 457
rect -241 423 -229 457
rect -287 389 -229 423
rect -287 355 -275 389
rect -241 355 -229 389
rect -287 321 -229 355
rect -287 287 -275 321
rect -241 287 -229 321
rect -287 253 -229 287
rect -287 219 -275 253
rect -241 219 -229 253
rect -287 185 -229 219
rect -287 151 -275 185
rect -241 151 -229 185
rect -287 117 -229 151
rect -287 83 -275 117
rect -241 83 -229 117
rect -287 49 -229 83
rect -287 15 -275 49
rect -241 15 -229 49
rect -287 -19 -229 15
rect -287 -53 -275 -19
rect -241 -53 -229 -19
rect -287 -87 -229 -53
rect -287 -121 -275 -87
rect -241 -121 -229 -87
rect -287 -155 -229 -121
rect -287 -189 -275 -155
rect -241 -189 -229 -155
rect -287 -223 -229 -189
rect -287 -257 -275 -223
rect -241 -257 -229 -223
rect -287 -291 -229 -257
rect -287 -325 -275 -291
rect -241 -325 -229 -291
rect -287 -359 -229 -325
rect -287 -393 -275 -359
rect -241 -393 -229 -359
rect -287 -427 -229 -393
rect -287 -461 -275 -427
rect -241 -461 -229 -427
rect -287 -495 -229 -461
rect -287 -529 -275 -495
rect -241 -529 -229 -495
rect -287 -563 -229 -529
rect -287 -597 -275 -563
rect -241 -597 -229 -563
rect -287 -631 -229 -597
rect -287 -665 -275 -631
rect -241 -665 -229 -631
rect -287 -699 -229 -665
rect -287 -733 -275 -699
rect -241 -733 -229 -699
rect -287 -767 -229 -733
rect -287 -801 -275 -767
rect -241 -801 -229 -767
rect -287 -835 -229 -801
rect -287 -869 -275 -835
rect -241 -869 -229 -835
rect -287 -903 -229 -869
rect -287 -937 -275 -903
rect -241 -937 -229 -903
rect -287 -971 -229 -937
rect -287 -1005 -275 -971
rect -241 -1005 -229 -971
rect -287 -1039 -229 -1005
rect -287 -1073 -275 -1039
rect -241 -1073 -229 -1039
rect -287 -1107 -229 -1073
rect -287 -1141 -275 -1107
rect -241 -1141 -229 -1107
rect -287 -1175 -229 -1141
rect -287 -1209 -275 -1175
rect -241 -1209 -229 -1175
rect -287 -1243 -229 -1209
rect -287 -1277 -275 -1243
rect -241 -1277 -229 -1243
rect -287 -1311 -229 -1277
rect -287 -1345 -275 -1311
rect -241 -1345 -229 -1311
rect -287 -1379 -229 -1345
rect -287 -1413 -275 -1379
rect -241 -1413 -229 -1379
rect -287 -1436 -229 -1413
rect -29 1341 29 1364
rect -29 1307 -17 1341
rect 17 1307 29 1341
rect -29 1273 29 1307
rect -29 1239 -17 1273
rect 17 1239 29 1273
rect -29 1205 29 1239
rect -29 1171 -17 1205
rect 17 1171 29 1205
rect -29 1137 29 1171
rect -29 1103 -17 1137
rect 17 1103 29 1137
rect -29 1069 29 1103
rect -29 1035 -17 1069
rect 17 1035 29 1069
rect -29 1001 29 1035
rect -29 967 -17 1001
rect 17 967 29 1001
rect -29 933 29 967
rect -29 899 -17 933
rect 17 899 29 933
rect -29 865 29 899
rect -29 831 -17 865
rect 17 831 29 865
rect -29 797 29 831
rect -29 763 -17 797
rect 17 763 29 797
rect -29 729 29 763
rect -29 695 -17 729
rect 17 695 29 729
rect -29 661 29 695
rect -29 627 -17 661
rect 17 627 29 661
rect -29 593 29 627
rect -29 559 -17 593
rect 17 559 29 593
rect -29 525 29 559
rect -29 491 -17 525
rect 17 491 29 525
rect -29 457 29 491
rect -29 423 -17 457
rect 17 423 29 457
rect -29 389 29 423
rect -29 355 -17 389
rect 17 355 29 389
rect -29 321 29 355
rect -29 287 -17 321
rect 17 287 29 321
rect -29 253 29 287
rect -29 219 -17 253
rect 17 219 29 253
rect -29 185 29 219
rect -29 151 -17 185
rect 17 151 29 185
rect -29 117 29 151
rect -29 83 -17 117
rect 17 83 29 117
rect -29 49 29 83
rect -29 15 -17 49
rect 17 15 29 49
rect -29 -19 29 15
rect -29 -53 -17 -19
rect 17 -53 29 -19
rect -29 -87 29 -53
rect -29 -121 -17 -87
rect 17 -121 29 -87
rect -29 -155 29 -121
rect -29 -189 -17 -155
rect 17 -189 29 -155
rect -29 -223 29 -189
rect -29 -257 -17 -223
rect 17 -257 29 -223
rect -29 -291 29 -257
rect -29 -325 -17 -291
rect 17 -325 29 -291
rect -29 -359 29 -325
rect -29 -393 -17 -359
rect 17 -393 29 -359
rect -29 -427 29 -393
rect -29 -461 -17 -427
rect 17 -461 29 -427
rect -29 -495 29 -461
rect -29 -529 -17 -495
rect 17 -529 29 -495
rect -29 -563 29 -529
rect -29 -597 -17 -563
rect 17 -597 29 -563
rect -29 -631 29 -597
rect -29 -665 -17 -631
rect 17 -665 29 -631
rect -29 -699 29 -665
rect -29 -733 -17 -699
rect 17 -733 29 -699
rect -29 -767 29 -733
rect -29 -801 -17 -767
rect 17 -801 29 -767
rect -29 -835 29 -801
rect -29 -869 -17 -835
rect 17 -869 29 -835
rect -29 -903 29 -869
rect -29 -937 -17 -903
rect 17 -937 29 -903
rect -29 -971 29 -937
rect -29 -1005 -17 -971
rect 17 -1005 29 -971
rect -29 -1039 29 -1005
rect -29 -1073 -17 -1039
rect 17 -1073 29 -1039
rect -29 -1107 29 -1073
rect -29 -1141 -17 -1107
rect 17 -1141 29 -1107
rect -29 -1175 29 -1141
rect -29 -1209 -17 -1175
rect 17 -1209 29 -1175
rect -29 -1243 29 -1209
rect -29 -1277 -17 -1243
rect 17 -1277 29 -1243
rect -29 -1311 29 -1277
rect -29 -1345 -17 -1311
rect 17 -1345 29 -1311
rect -29 -1379 29 -1345
rect -29 -1413 -17 -1379
rect 17 -1413 29 -1379
rect -29 -1436 29 -1413
rect 229 1341 287 1364
rect 229 1307 241 1341
rect 275 1307 287 1341
rect 229 1273 287 1307
rect 229 1239 241 1273
rect 275 1239 287 1273
rect 229 1205 287 1239
rect 229 1171 241 1205
rect 275 1171 287 1205
rect 229 1137 287 1171
rect 229 1103 241 1137
rect 275 1103 287 1137
rect 229 1069 287 1103
rect 229 1035 241 1069
rect 275 1035 287 1069
rect 229 1001 287 1035
rect 229 967 241 1001
rect 275 967 287 1001
rect 229 933 287 967
rect 229 899 241 933
rect 275 899 287 933
rect 229 865 287 899
rect 229 831 241 865
rect 275 831 287 865
rect 229 797 287 831
rect 229 763 241 797
rect 275 763 287 797
rect 229 729 287 763
rect 229 695 241 729
rect 275 695 287 729
rect 229 661 287 695
rect 229 627 241 661
rect 275 627 287 661
rect 229 593 287 627
rect 229 559 241 593
rect 275 559 287 593
rect 229 525 287 559
rect 229 491 241 525
rect 275 491 287 525
rect 229 457 287 491
rect 229 423 241 457
rect 275 423 287 457
rect 229 389 287 423
rect 229 355 241 389
rect 275 355 287 389
rect 229 321 287 355
rect 229 287 241 321
rect 275 287 287 321
rect 229 253 287 287
rect 229 219 241 253
rect 275 219 287 253
rect 229 185 287 219
rect 229 151 241 185
rect 275 151 287 185
rect 229 117 287 151
rect 229 83 241 117
rect 275 83 287 117
rect 229 49 287 83
rect 229 15 241 49
rect 275 15 287 49
rect 229 -19 287 15
rect 229 -53 241 -19
rect 275 -53 287 -19
rect 229 -87 287 -53
rect 229 -121 241 -87
rect 275 -121 287 -87
rect 229 -155 287 -121
rect 229 -189 241 -155
rect 275 -189 287 -155
rect 229 -223 287 -189
rect 229 -257 241 -223
rect 275 -257 287 -223
rect 229 -291 287 -257
rect 229 -325 241 -291
rect 275 -325 287 -291
rect 229 -359 287 -325
rect 229 -393 241 -359
rect 275 -393 287 -359
rect 229 -427 287 -393
rect 229 -461 241 -427
rect 275 -461 287 -427
rect 229 -495 287 -461
rect 229 -529 241 -495
rect 275 -529 287 -495
rect 229 -563 287 -529
rect 229 -597 241 -563
rect 275 -597 287 -563
rect 229 -631 287 -597
rect 229 -665 241 -631
rect 275 -665 287 -631
rect 229 -699 287 -665
rect 229 -733 241 -699
rect 275 -733 287 -699
rect 229 -767 287 -733
rect 229 -801 241 -767
rect 275 -801 287 -767
rect 229 -835 287 -801
rect 229 -869 241 -835
rect 275 -869 287 -835
rect 229 -903 287 -869
rect 229 -937 241 -903
rect 275 -937 287 -903
rect 229 -971 287 -937
rect 229 -1005 241 -971
rect 275 -1005 287 -971
rect 229 -1039 287 -1005
rect 229 -1073 241 -1039
rect 275 -1073 287 -1039
rect 229 -1107 287 -1073
rect 229 -1141 241 -1107
rect 275 -1141 287 -1107
rect 229 -1175 287 -1141
rect 229 -1209 241 -1175
rect 275 -1209 287 -1175
rect 229 -1243 287 -1209
rect 229 -1277 241 -1243
rect 275 -1277 287 -1243
rect 229 -1311 287 -1277
rect 229 -1345 241 -1311
rect 275 -1345 287 -1311
rect 229 -1379 287 -1345
rect 229 -1413 241 -1379
rect 275 -1413 287 -1379
rect 229 -1436 287 -1413
<< pdiffc >>
rect -275 1307 -241 1341
rect -275 1239 -241 1273
rect -275 1171 -241 1205
rect -275 1103 -241 1137
rect -275 1035 -241 1069
rect -275 967 -241 1001
rect -275 899 -241 933
rect -275 831 -241 865
rect -275 763 -241 797
rect -275 695 -241 729
rect -275 627 -241 661
rect -275 559 -241 593
rect -275 491 -241 525
rect -275 423 -241 457
rect -275 355 -241 389
rect -275 287 -241 321
rect -275 219 -241 253
rect -275 151 -241 185
rect -275 83 -241 117
rect -275 15 -241 49
rect -275 -53 -241 -19
rect -275 -121 -241 -87
rect -275 -189 -241 -155
rect -275 -257 -241 -223
rect -275 -325 -241 -291
rect -275 -393 -241 -359
rect -275 -461 -241 -427
rect -275 -529 -241 -495
rect -275 -597 -241 -563
rect -275 -665 -241 -631
rect -275 -733 -241 -699
rect -275 -801 -241 -767
rect -275 -869 -241 -835
rect -275 -937 -241 -903
rect -275 -1005 -241 -971
rect -275 -1073 -241 -1039
rect -275 -1141 -241 -1107
rect -275 -1209 -241 -1175
rect -275 -1277 -241 -1243
rect -275 -1345 -241 -1311
rect -275 -1413 -241 -1379
rect -17 1307 17 1341
rect -17 1239 17 1273
rect -17 1171 17 1205
rect -17 1103 17 1137
rect -17 1035 17 1069
rect -17 967 17 1001
rect -17 899 17 933
rect -17 831 17 865
rect -17 763 17 797
rect -17 695 17 729
rect -17 627 17 661
rect -17 559 17 593
rect -17 491 17 525
rect -17 423 17 457
rect -17 355 17 389
rect -17 287 17 321
rect -17 219 17 253
rect -17 151 17 185
rect -17 83 17 117
rect -17 15 17 49
rect -17 -53 17 -19
rect -17 -121 17 -87
rect -17 -189 17 -155
rect -17 -257 17 -223
rect -17 -325 17 -291
rect -17 -393 17 -359
rect -17 -461 17 -427
rect -17 -529 17 -495
rect -17 -597 17 -563
rect -17 -665 17 -631
rect -17 -733 17 -699
rect -17 -801 17 -767
rect -17 -869 17 -835
rect -17 -937 17 -903
rect -17 -1005 17 -971
rect -17 -1073 17 -1039
rect -17 -1141 17 -1107
rect -17 -1209 17 -1175
rect -17 -1277 17 -1243
rect -17 -1345 17 -1311
rect -17 -1413 17 -1379
rect 241 1307 275 1341
rect 241 1239 275 1273
rect 241 1171 275 1205
rect 241 1103 275 1137
rect 241 1035 275 1069
rect 241 967 275 1001
rect 241 899 275 933
rect 241 831 275 865
rect 241 763 275 797
rect 241 695 275 729
rect 241 627 275 661
rect 241 559 275 593
rect 241 491 275 525
rect 241 423 275 457
rect 241 355 275 389
rect 241 287 275 321
rect 241 219 275 253
rect 241 151 275 185
rect 241 83 275 117
rect 241 15 275 49
rect 241 -53 275 -19
rect 241 -121 275 -87
rect 241 -189 275 -155
rect 241 -257 275 -223
rect 241 -325 275 -291
rect 241 -393 275 -359
rect 241 -461 275 -427
rect 241 -529 275 -495
rect 241 -597 275 -563
rect 241 -665 275 -631
rect 241 -733 275 -699
rect 241 -801 275 -767
rect 241 -869 275 -835
rect 241 -937 275 -903
rect 241 -1005 275 -971
rect 241 -1073 275 -1039
rect 241 -1141 275 -1107
rect 241 -1209 275 -1175
rect 241 -1277 275 -1243
rect 241 -1345 275 -1311
rect 241 -1413 275 -1379
<< poly >>
rect -229 1445 -29 1461
rect -229 1411 -180 1445
rect -146 1411 -112 1445
rect -78 1411 -29 1445
rect -229 1364 -29 1411
rect 29 1445 229 1461
rect 29 1411 78 1445
rect 112 1411 146 1445
rect 180 1411 229 1445
rect 29 1364 229 1411
rect -229 -1451 -29 -1436
rect 29 -1451 229 -1436
rect -229 -1495 229 -1451
<< polycont >>
rect -180 1411 -146 1445
rect -112 1411 -78 1445
rect 78 1411 112 1445
rect 146 1411 180 1445
<< locali >>
rect -229 1411 -182 1445
rect -146 1411 -112 1445
rect -76 1411 -29 1445
rect 29 1411 76 1445
rect 112 1411 146 1445
rect 182 1411 229 1445
rect -275 1349 -241 1368
rect -275 1277 -241 1307
rect -275 1205 -241 1239
rect -275 1137 -241 1171
rect -275 1069 -241 1099
rect -275 1001 -241 1027
rect -275 933 -241 955
rect -275 865 -241 883
rect -275 797 -241 811
rect -275 729 -241 739
rect -275 661 -241 667
rect -275 593 -241 595
rect -275 557 -241 559
rect -275 485 -241 491
rect -275 413 -241 423
rect -275 341 -241 355
rect -275 269 -241 287
rect -275 197 -241 219
rect -275 125 -241 151
rect -275 53 -241 83
rect -275 -19 -241 15
rect -275 -87 -241 -53
rect -275 -155 -241 -125
rect -275 -223 -241 -197
rect -275 -291 -241 -269
rect -275 -359 -241 -341
rect -275 -427 -241 -413
rect -275 -495 -241 -485
rect -275 -563 -241 -557
rect -275 -631 -241 -629
rect -275 -667 -241 -665
rect -275 -739 -241 -733
rect -275 -811 -241 -801
rect -275 -883 -241 -869
rect -275 -955 -241 -937
rect -275 -1027 -241 -1005
rect -275 -1099 -241 -1073
rect -275 -1171 -241 -1141
rect -275 -1243 -241 -1209
rect -275 -1311 -241 -1277
rect -275 -1379 -241 -1349
rect -275 -1440 -241 -1421
rect -17 1349 17 1368
rect -17 1277 17 1307
rect -17 1205 17 1239
rect -17 1137 17 1171
rect -17 1069 17 1099
rect -17 1001 17 1027
rect -17 933 17 955
rect -17 865 17 883
rect -17 797 17 811
rect -17 729 17 739
rect -17 661 17 667
rect -17 593 17 595
rect -17 557 17 559
rect -17 485 17 491
rect -17 413 17 423
rect -17 341 17 355
rect -17 269 17 287
rect -17 197 17 219
rect -17 125 17 151
rect -17 53 17 83
rect -17 -19 17 15
rect -17 -87 17 -53
rect -17 -155 17 -125
rect -17 -223 17 -197
rect -17 -291 17 -269
rect -17 -359 17 -341
rect -17 -427 17 -413
rect -17 -495 17 -485
rect -17 -563 17 -557
rect -17 -631 17 -629
rect -17 -667 17 -665
rect -17 -739 17 -733
rect -17 -811 17 -801
rect -17 -883 17 -869
rect -17 -955 17 -937
rect -17 -1027 17 -1005
rect -17 -1099 17 -1073
rect -17 -1171 17 -1141
rect -17 -1243 17 -1209
rect -17 -1311 17 -1277
rect -17 -1379 17 -1349
rect -17 -1440 17 -1421
rect 241 1349 275 1368
rect 241 1277 275 1307
rect 241 1205 275 1239
rect 241 1137 275 1171
rect 241 1069 275 1099
rect 241 1001 275 1027
rect 241 933 275 955
rect 241 865 275 883
rect 241 797 275 811
rect 241 729 275 739
rect 241 661 275 667
rect 241 593 275 595
rect 241 557 275 559
rect 241 485 275 491
rect 241 413 275 423
rect 241 341 275 355
rect 241 269 275 287
rect 241 197 275 219
rect 241 125 275 151
rect 241 53 275 83
rect 241 -19 275 15
rect 241 -87 275 -53
rect 241 -155 275 -125
rect 241 -223 275 -197
rect 241 -291 275 -269
rect 241 -359 275 -341
rect 241 -427 275 -413
rect 241 -495 275 -485
rect 241 -563 275 -557
rect 241 -631 275 -629
rect 241 -667 275 -665
rect 241 -739 275 -733
rect 241 -811 275 -801
rect 241 -883 275 -869
rect 241 -955 275 -937
rect 241 -1027 275 -1005
rect 241 -1099 275 -1073
rect 241 -1171 275 -1141
rect 241 -1243 275 -1209
rect 241 -1311 275 -1277
rect 241 -1379 275 -1349
rect 241 -1440 275 -1421
<< viali >>
rect -182 1411 -180 1445
rect -180 1411 -148 1445
rect -110 1411 -78 1445
rect -78 1411 -76 1445
rect 76 1411 78 1445
rect 78 1411 110 1445
rect 148 1411 180 1445
rect 180 1411 182 1445
rect -275 1341 -241 1349
rect -275 1315 -241 1341
rect -275 1273 -241 1277
rect -275 1243 -241 1273
rect -275 1171 -241 1205
rect -275 1103 -241 1133
rect -275 1099 -241 1103
rect -275 1035 -241 1061
rect -275 1027 -241 1035
rect -275 967 -241 989
rect -275 955 -241 967
rect -275 899 -241 917
rect -275 883 -241 899
rect -275 831 -241 845
rect -275 811 -241 831
rect -275 763 -241 773
rect -275 739 -241 763
rect -275 695 -241 701
rect -275 667 -241 695
rect -275 627 -241 629
rect -275 595 -241 627
rect -275 525 -241 557
rect -275 523 -241 525
rect -275 457 -241 485
rect -275 451 -241 457
rect -275 389 -241 413
rect -275 379 -241 389
rect -275 321 -241 341
rect -275 307 -241 321
rect -275 253 -241 269
rect -275 235 -241 253
rect -275 185 -241 197
rect -275 163 -241 185
rect -275 117 -241 125
rect -275 91 -241 117
rect -275 49 -241 53
rect -275 19 -241 49
rect -275 -53 -241 -19
rect -275 -121 -241 -91
rect -275 -125 -241 -121
rect -275 -189 -241 -163
rect -275 -197 -241 -189
rect -275 -257 -241 -235
rect -275 -269 -241 -257
rect -275 -325 -241 -307
rect -275 -341 -241 -325
rect -275 -393 -241 -379
rect -275 -413 -241 -393
rect -275 -461 -241 -451
rect -275 -485 -241 -461
rect -275 -529 -241 -523
rect -275 -557 -241 -529
rect -275 -597 -241 -595
rect -275 -629 -241 -597
rect -275 -699 -241 -667
rect -275 -701 -241 -699
rect -275 -767 -241 -739
rect -275 -773 -241 -767
rect -275 -835 -241 -811
rect -275 -845 -241 -835
rect -275 -903 -241 -883
rect -275 -917 -241 -903
rect -275 -971 -241 -955
rect -275 -989 -241 -971
rect -275 -1039 -241 -1027
rect -275 -1061 -241 -1039
rect -275 -1107 -241 -1099
rect -275 -1133 -241 -1107
rect -275 -1175 -241 -1171
rect -275 -1205 -241 -1175
rect -275 -1277 -241 -1243
rect -275 -1345 -241 -1315
rect -275 -1349 -241 -1345
rect -275 -1413 -241 -1387
rect -275 -1421 -241 -1413
rect -17 1341 17 1349
rect -17 1315 17 1341
rect -17 1273 17 1277
rect -17 1243 17 1273
rect -17 1171 17 1205
rect -17 1103 17 1133
rect -17 1099 17 1103
rect -17 1035 17 1061
rect -17 1027 17 1035
rect -17 967 17 989
rect -17 955 17 967
rect -17 899 17 917
rect -17 883 17 899
rect -17 831 17 845
rect -17 811 17 831
rect -17 763 17 773
rect -17 739 17 763
rect -17 695 17 701
rect -17 667 17 695
rect -17 627 17 629
rect -17 595 17 627
rect -17 525 17 557
rect -17 523 17 525
rect -17 457 17 485
rect -17 451 17 457
rect -17 389 17 413
rect -17 379 17 389
rect -17 321 17 341
rect -17 307 17 321
rect -17 253 17 269
rect -17 235 17 253
rect -17 185 17 197
rect -17 163 17 185
rect -17 117 17 125
rect -17 91 17 117
rect -17 49 17 53
rect -17 19 17 49
rect -17 -53 17 -19
rect -17 -121 17 -91
rect -17 -125 17 -121
rect -17 -189 17 -163
rect -17 -197 17 -189
rect -17 -257 17 -235
rect -17 -269 17 -257
rect -17 -325 17 -307
rect -17 -341 17 -325
rect -17 -393 17 -379
rect -17 -413 17 -393
rect -17 -461 17 -451
rect -17 -485 17 -461
rect -17 -529 17 -523
rect -17 -557 17 -529
rect -17 -597 17 -595
rect -17 -629 17 -597
rect -17 -699 17 -667
rect -17 -701 17 -699
rect -17 -767 17 -739
rect -17 -773 17 -767
rect -17 -835 17 -811
rect -17 -845 17 -835
rect -17 -903 17 -883
rect -17 -917 17 -903
rect -17 -971 17 -955
rect -17 -989 17 -971
rect -17 -1039 17 -1027
rect -17 -1061 17 -1039
rect -17 -1107 17 -1099
rect -17 -1133 17 -1107
rect -17 -1175 17 -1171
rect -17 -1205 17 -1175
rect -17 -1277 17 -1243
rect -17 -1345 17 -1315
rect -17 -1349 17 -1345
rect -17 -1413 17 -1387
rect -17 -1421 17 -1413
rect 241 1341 275 1349
rect 241 1315 275 1341
rect 241 1273 275 1277
rect 241 1243 275 1273
rect 241 1171 275 1205
rect 241 1103 275 1133
rect 241 1099 275 1103
rect 241 1035 275 1061
rect 241 1027 275 1035
rect 241 967 275 989
rect 241 955 275 967
rect 241 899 275 917
rect 241 883 275 899
rect 241 831 275 845
rect 241 811 275 831
rect 241 763 275 773
rect 241 739 275 763
rect 241 695 275 701
rect 241 667 275 695
rect 241 627 275 629
rect 241 595 275 627
rect 241 525 275 557
rect 241 523 275 525
rect 241 457 275 485
rect 241 451 275 457
rect 241 389 275 413
rect 241 379 275 389
rect 241 321 275 341
rect 241 307 275 321
rect 241 253 275 269
rect 241 235 275 253
rect 241 185 275 197
rect 241 163 275 185
rect 241 117 275 125
rect 241 91 275 117
rect 241 49 275 53
rect 241 19 275 49
rect 241 -53 275 -19
rect 241 -121 275 -91
rect 241 -125 275 -121
rect 241 -189 275 -163
rect 241 -197 275 -189
rect 241 -257 275 -235
rect 241 -269 275 -257
rect 241 -325 275 -307
rect 241 -341 275 -325
rect 241 -393 275 -379
rect 241 -413 275 -393
rect 241 -461 275 -451
rect 241 -485 275 -461
rect 241 -529 275 -523
rect 241 -557 275 -529
rect 241 -597 275 -595
rect 241 -629 275 -597
rect 241 -699 275 -667
rect 241 -701 275 -699
rect 241 -767 275 -739
rect 241 -773 275 -767
rect 241 -835 275 -811
rect 241 -845 275 -835
rect 241 -903 275 -883
rect 241 -917 275 -903
rect 241 -971 275 -955
rect 241 -989 275 -971
rect 241 -1039 275 -1027
rect 241 -1061 275 -1039
rect 241 -1107 275 -1099
rect 241 -1133 275 -1107
rect 241 -1175 275 -1171
rect 241 -1205 275 -1175
rect 241 -1277 275 -1243
rect 241 -1345 275 -1315
rect 241 -1349 275 -1345
rect 241 -1413 275 -1387
rect 241 -1421 275 -1413
<< metal1 >>
rect -225 1445 -33 1451
rect -225 1411 -182 1445
rect -148 1411 -110 1445
rect -76 1411 -33 1445
rect -225 1405 -33 1411
rect 33 1445 225 1451
rect 33 1411 76 1445
rect 110 1411 148 1445
rect 182 1411 225 1445
rect 33 1405 225 1411
rect -281 1349 -235 1364
rect -281 1315 -275 1349
rect -241 1315 -235 1349
rect -281 1277 -235 1315
rect -281 1243 -275 1277
rect -241 1243 -235 1277
rect -281 1205 -235 1243
rect -281 1171 -275 1205
rect -241 1171 -235 1205
rect -281 1133 -235 1171
rect -281 1099 -275 1133
rect -241 1099 -235 1133
rect -281 1061 -235 1099
rect -281 1027 -275 1061
rect -241 1027 -235 1061
rect -281 989 -235 1027
rect -281 955 -275 989
rect -241 955 -235 989
rect -281 917 -235 955
rect -281 883 -275 917
rect -241 883 -235 917
rect -281 845 -235 883
rect -281 811 -275 845
rect -241 811 -235 845
rect -281 773 -235 811
rect -281 739 -275 773
rect -241 739 -235 773
rect -281 701 -235 739
rect -281 667 -275 701
rect -241 667 -235 701
rect -281 629 -235 667
rect -281 595 -275 629
rect -241 595 -235 629
rect -281 557 -235 595
rect -281 523 -275 557
rect -241 523 -235 557
rect -281 485 -235 523
rect -281 451 -275 485
rect -241 451 -235 485
rect -281 413 -235 451
rect -281 379 -275 413
rect -241 379 -235 413
rect -281 341 -235 379
rect -281 307 -275 341
rect -241 307 -235 341
rect -281 269 -235 307
rect -281 235 -275 269
rect -241 235 -235 269
rect -281 197 -235 235
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -163 -235 -125
rect -281 -197 -275 -163
rect -241 -197 -235 -163
rect -281 -235 -235 -197
rect -281 -269 -275 -235
rect -241 -269 -235 -235
rect -281 -307 -235 -269
rect -281 -341 -275 -307
rect -241 -341 -235 -307
rect -281 -379 -235 -341
rect -281 -413 -275 -379
rect -241 -413 -235 -379
rect -281 -451 -235 -413
rect -281 -485 -275 -451
rect -241 -485 -235 -451
rect -281 -523 -235 -485
rect -281 -557 -275 -523
rect -241 -557 -235 -523
rect -281 -595 -235 -557
rect -281 -629 -275 -595
rect -241 -629 -235 -595
rect -281 -667 -235 -629
rect -281 -701 -275 -667
rect -241 -701 -235 -667
rect -281 -739 -235 -701
rect -281 -773 -275 -739
rect -241 -773 -235 -739
rect -281 -811 -235 -773
rect -281 -845 -275 -811
rect -241 -845 -235 -811
rect -281 -883 -235 -845
rect -281 -917 -275 -883
rect -241 -917 -235 -883
rect -281 -955 -235 -917
rect -281 -989 -275 -955
rect -241 -989 -235 -955
rect -281 -1027 -235 -989
rect -281 -1061 -275 -1027
rect -241 -1061 -235 -1027
rect -281 -1099 -235 -1061
rect -281 -1133 -275 -1099
rect -241 -1133 -235 -1099
rect -281 -1171 -235 -1133
rect -281 -1205 -275 -1171
rect -241 -1205 -235 -1171
rect -281 -1243 -235 -1205
rect -281 -1277 -275 -1243
rect -241 -1277 -235 -1243
rect -281 -1315 -235 -1277
rect -281 -1349 -275 -1315
rect -241 -1349 -235 -1315
rect -281 -1387 -235 -1349
rect -281 -1421 -275 -1387
rect -241 -1421 -235 -1387
rect -281 -1436 -235 -1421
rect -23 1349 23 1364
rect -23 1315 -17 1349
rect 17 1315 23 1349
rect -23 1277 23 1315
rect -23 1243 -17 1277
rect 17 1243 23 1277
rect -23 1205 23 1243
rect -23 1171 -17 1205
rect 17 1171 23 1205
rect -23 1133 23 1171
rect -23 1099 -17 1133
rect 17 1099 23 1133
rect -23 1061 23 1099
rect -23 1027 -17 1061
rect 17 1027 23 1061
rect -23 989 23 1027
rect -23 955 -17 989
rect 17 955 23 989
rect -23 917 23 955
rect -23 883 -17 917
rect 17 883 23 917
rect -23 845 23 883
rect -23 811 -17 845
rect 17 811 23 845
rect -23 773 23 811
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -811 23 -773
rect -23 -845 -17 -811
rect 17 -845 23 -811
rect -23 -883 23 -845
rect -23 -917 -17 -883
rect 17 -917 23 -883
rect -23 -955 23 -917
rect -23 -989 -17 -955
rect 17 -989 23 -955
rect -23 -1027 23 -989
rect -23 -1061 -17 -1027
rect 17 -1061 23 -1027
rect -23 -1099 23 -1061
rect -23 -1133 -17 -1099
rect 17 -1133 23 -1099
rect -23 -1171 23 -1133
rect -23 -1205 -17 -1171
rect 17 -1205 23 -1171
rect -23 -1243 23 -1205
rect -23 -1277 -17 -1243
rect 17 -1277 23 -1243
rect -23 -1315 23 -1277
rect -23 -1349 -17 -1315
rect 17 -1349 23 -1315
rect -23 -1387 23 -1349
rect -23 -1421 -17 -1387
rect 17 -1421 23 -1387
rect -23 -1436 23 -1421
rect 235 1349 281 1364
rect 235 1315 241 1349
rect 275 1315 281 1349
rect 235 1277 281 1315
rect 235 1243 241 1277
rect 275 1243 281 1277
rect 235 1205 281 1243
rect 235 1171 241 1205
rect 275 1171 281 1205
rect 235 1133 281 1171
rect 235 1099 241 1133
rect 275 1099 281 1133
rect 235 1061 281 1099
rect 235 1027 241 1061
rect 275 1027 281 1061
rect 235 989 281 1027
rect 235 955 241 989
rect 275 955 281 989
rect 235 917 281 955
rect 235 883 241 917
rect 275 883 281 917
rect 235 845 281 883
rect 235 811 241 845
rect 275 811 281 845
rect 235 773 281 811
rect 235 739 241 773
rect 275 739 281 773
rect 235 701 281 739
rect 235 667 241 701
rect 275 667 281 701
rect 235 629 281 667
rect 235 595 241 629
rect 275 595 281 629
rect 235 557 281 595
rect 235 523 241 557
rect 275 523 281 557
rect 235 485 281 523
rect 235 451 241 485
rect 275 451 281 485
rect 235 413 281 451
rect 235 379 241 413
rect 275 379 281 413
rect 235 341 281 379
rect 235 307 241 341
rect 275 307 281 341
rect 235 269 281 307
rect 235 235 241 269
rect 275 235 281 269
rect 235 197 281 235
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -163 281 -125
rect 235 -197 241 -163
rect 275 -197 281 -163
rect 235 -235 281 -197
rect 235 -269 241 -235
rect 275 -269 281 -235
rect 235 -307 281 -269
rect 235 -341 241 -307
rect 275 -341 281 -307
rect 235 -379 281 -341
rect 235 -413 241 -379
rect 275 -413 281 -379
rect 235 -451 281 -413
rect 235 -485 241 -451
rect 275 -485 281 -451
rect 235 -523 281 -485
rect 235 -557 241 -523
rect 275 -557 281 -523
rect 235 -595 281 -557
rect 235 -629 241 -595
rect 275 -629 281 -595
rect 235 -667 281 -629
rect 235 -701 241 -667
rect 275 -701 281 -667
rect 235 -739 281 -701
rect 235 -773 241 -739
rect 275 -773 281 -739
rect 235 -811 281 -773
rect 235 -845 241 -811
rect 275 -845 281 -811
rect 235 -883 281 -845
rect 235 -917 241 -883
rect 275 -917 281 -883
rect 235 -955 281 -917
rect 235 -989 241 -955
rect 275 -989 281 -955
rect 235 -1027 281 -989
rect 235 -1061 241 -1027
rect 275 -1061 281 -1027
rect 235 -1099 281 -1061
rect 235 -1133 241 -1099
rect 275 -1133 281 -1099
rect 235 -1171 281 -1133
rect 235 -1205 241 -1171
rect 275 -1205 281 -1171
rect 235 -1243 281 -1205
rect 235 -1277 241 -1243
rect 275 -1277 281 -1243
rect 235 -1315 281 -1277
rect 235 -1349 241 -1315
rect 275 -1349 281 -1315
rect 235 -1387 281 -1349
rect 235 -1421 241 -1387
rect 275 -1421 281 -1387
rect 235 -1436 281 -1421
<< end >>
