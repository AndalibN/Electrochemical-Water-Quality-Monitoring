magic
tech sky130A
magscale 1 2
timestamp 1667956596
<< error_p >>
rect -29 321 29 327
rect -29 287 -17 321
rect -29 281 29 287
rect -29 -287 29 -281
rect -29 -321 -17 -287
rect -29 -327 29 -321
<< nwell >>
rect -226 -459 226 459
<< pmos >>
rect -30 -240 30 240
<< pdiff >>
rect -88 228 -30 240
rect -88 -228 -76 228
rect -42 -228 -30 228
rect -88 -240 -30 -228
rect 30 228 88 240
rect 30 -228 42 228
rect 76 -228 88 228
rect 30 -240 88 -228
<< pdiffc >>
rect -76 -228 -42 228
rect 42 -228 76 228
<< nsubdiff >>
rect -190 389 -94 423
rect 94 389 190 423
rect -190 327 -156 389
rect 156 327 190 389
rect -190 -389 -156 -327
rect 156 -389 190 -327
rect -190 -423 -94 -389
rect 94 -423 190 -389
<< nsubdiffcont >>
rect -94 389 94 423
rect -190 -327 -156 327
rect 156 -327 190 327
rect -94 -423 94 -389
<< poly >>
rect -33 321 33 337
rect -33 287 -17 321
rect 17 287 33 321
rect -33 271 33 287
rect -30 240 30 271
rect -30 -271 30 -240
rect -33 -287 33 -271
rect -33 -321 -17 -287
rect 17 -321 33 -287
rect -33 -337 33 -321
<< polycont >>
rect -17 287 17 321
rect -17 -321 17 -287
<< locali >>
rect -190 389 -94 423
rect 94 389 190 423
rect -190 327 -156 389
rect 156 327 190 389
rect -33 287 -17 321
rect 17 287 33 321
rect -76 228 -42 244
rect -76 -244 -42 -228
rect 42 228 76 244
rect 42 -244 76 -228
rect -33 -321 -17 -287
rect 17 -321 33 -287
rect -190 -389 -156 -327
rect 156 -389 190 -327
rect -190 -423 -94 -389
rect 94 -423 190 -389
<< viali >>
rect -17 287 17 321
rect -76 -228 -42 228
rect 42 -228 76 228
rect -17 -321 17 -287
<< metal1 >>
rect -29 321 29 327
rect -29 287 -17 321
rect 17 287 29 321
rect -29 281 29 287
rect -82 228 -36 240
rect -82 -228 -76 228
rect -42 -228 -36 228
rect -82 -240 -36 -228
rect 36 228 82 240
rect 36 -228 42 228
rect 76 -228 82 228
rect 36 -240 82 -228
rect -29 -287 29 -281
rect -29 -321 -17 -287
rect 17 -321 29 -287
rect -29 -327 29 -321
<< properties >>
string FIXED_BBOX -173 -406 173 406
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.4 l 0.30 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
