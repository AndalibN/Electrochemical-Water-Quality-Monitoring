magic
tech sky130A
magscale 1 2
timestamp 1666811438
<< error_p >>
rect -32 3683 32 3689
rect -32 3649 -20 3683
rect -32 3643 32 3649
rect -32 -3649 32 -3643
rect -32 -3683 -20 -3649
rect -32 -3689 32 -3683
<< nmos >>
rect -36 -3611 36 3611
<< ndiff >>
rect -94 3599 -36 3611
rect -94 -3599 -82 3599
rect -48 -3599 -36 3599
rect -94 -3611 -36 -3599
rect 36 3599 94 3611
rect 36 -3599 48 3599
rect 82 -3599 94 3599
rect 36 -3611 94 -3599
<< ndiffc >>
rect -82 -3599 -48 3599
rect 48 -3599 82 3599
<< poly >>
rect -36 3683 36 3699
rect -36 3649 -20 3683
rect 20 3649 36 3683
rect -36 3611 36 3649
rect -36 -3649 36 -3611
rect -36 -3683 -20 -3649
rect 20 -3683 36 -3649
rect -36 -3699 36 -3683
<< polycont >>
rect -20 3649 20 3683
rect -20 -3683 20 -3649
<< locali >>
rect -36 3649 -20 3683
rect 20 3649 36 3683
rect -82 3599 -48 3615
rect -82 -3615 -48 -3599
rect 48 3599 82 3615
rect 48 -3615 82 -3599
rect -36 -3683 -20 -3649
rect 20 -3683 36 -3649
<< viali >>
rect -20 3649 20 3683
rect -82 -3599 -48 3599
rect 48 -3599 82 3599
rect -20 -3683 20 -3649
<< metal1 >>
rect -32 3683 32 3689
rect -32 3649 -20 3683
rect 20 3649 32 3683
rect -32 3643 32 3649
rect -88 3599 -42 3611
rect -88 -3599 -82 3599
rect -48 -3599 -42 3599
rect -88 -3611 -42 -3599
rect 42 3599 88 3611
rect 42 -3599 48 3599
rect 82 -3599 88 3599
rect 42 -3611 88 -3599
rect -32 -3649 32 -3643
rect -32 -3683 -20 -3649
rect 20 -3683 32 -3649
rect -32 -3689 32 -3683
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 36.112 l 0.361 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
