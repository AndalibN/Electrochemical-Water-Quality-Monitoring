magic
tech sky130A
magscale 1 2
timestamp 1669756519
<< psubdiff >>
rect 9902 15418 9942 15442
rect 10240 15414 10284 15438
rect 9902 15328 9916 15352
rect 19254 15310 19278 15352
rect 19404 15248 19428 15352
rect 18998 14654 19024 14678
rect 19422 14594 19446 14654
rect 18998 14556 19020 14580
rect 11140 10144 11228 10168
rect 11626 10162 11702 10186
rect 11670 9954 11702 9978
rect 21276 10012 21342 10036
rect 18988 9606 19020 9630
rect 21312 9870 21342 9894
rect 18988 9494 19066 9518
rect 9862 9382 9886 9442
rect 9948 9382 9972 9408
rect 20918 4398 20942 4586
rect 18972 4254 18996 4398
rect 20918 4250 20942 4254
rect 21318 4250 21342 4586
rect 18998 3936 19002 3960
rect 19248 3936 19256 3960
rect 19248 -402 19320 -378
rect 13716 -488 13790 -464
rect 11496 -884 11548 -860
rect 13692 -1000 13716 -956
rect 13790 -1000 13814 -964
rect 11496 -1024 11598 -1000
rect 19220 -1044 19320 -1020
<< psubdiffcont >>
rect 9902 15386 9942 15418
rect 10240 15386 10284 15414
rect 9902 15352 10284 15386
rect 9916 15310 10284 15352
rect 19278 15310 19404 15352
rect 9916 15248 19404 15310
rect 9916 14902 19354 15248
rect 9916 10070 10246 14902
rect 19024 14654 19354 14902
rect 18998 14594 19422 14654
rect 18998 14580 19376 14594
rect 11140 10070 11228 10144
rect 9916 10068 11228 10070
rect 11626 10068 11702 10162
rect 9916 9978 11702 10068
rect 9916 9442 11670 9978
rect 19020 9940 19376 14580
rect 21276 9940 21342 10012
rect 19020 9894 21342 9940
rect 19020 9606 21312 9894
rect 18988 9552 21312 9606
rect 18988 9518 19066 9552
rect 9886 9408 11670 9442
rect 9886 9382 9948 9408
rect 11548 -674 11670 9408
rect 20994 4586 21312 9552
rect 20942 4398 21318 4586
rect 18996 4254 21318 4398
rect 18998 3960 19256 4254
rect 20942 4250 21318 4254
rect 19002 -402 19248 3960
rect 13716 -532 13790 -488
rect 19002 -532 19320 -402
rect 13716 -674 19320 -532
rect 11548 -884 19320 -674
rect 11496 -956 19320 -884
rect 11496 -1000 11598 -956
rect 13716 -964 19320 -956
rect 13716 -1000 13790 -964
rect 19220 -1020 19320 -964
<< poly >>
rect 19761 4590 20048 4656
rect 20217 4598 20479 4655
rect 20217 4590 20296 4598
rect 20272 4552 20296 4590
rect 20350 4590 20479 4598
rect 20350 4552 20376 4590
rect 20272 4540 20376 4552
rect 16573 423 16693 546
rect 17452 441 17569 579
rect 17006 423 17134 424
rect 17452 423 17469 441
rect 16572 384 17469 423
rect 17555 384 17569 441
rect 16572 354 17569 384
rect 17452 353 17569 354
<< polycont >>
rect 20296 4552 20350 4598
rect 17469 384 17555 441
<< locali >>
rect 9902 15418 9942 15434
rect 10240 15414 10284 15430
rect 9902 15336 9916 15352
rect 19262 15310 19278 15352
rect 19404 15248 19420 15352
rect 18998 14654 19024 14670
rect 14747 14609 16550 14610
rect 14747 14607 16917 14609
rect 14747 14575 18448 14607
rect 10532 14574 18448 14575
rect 10532 14572 16561 14574
rect 16882 14573 18448 14574
rect 10532 14539 14781 14572
rect 10532 11798 10589 14539
rect 14747 14458 14781 14539
rect 15103 14458 15137 14572
rect 15459 14459 15493 14572
rect 15815 14459 15849 14572
rect 16171 14458 16205 14572
rect 16527 14459 16561 14572
rect 16883 14459 16917 14573
rect 17316 14571 18448 14573
rect 19422 14594 19438 14654
rect 17316 14473 17351 14571
rect 17672 14473 17706 14571
rect 18028 14473 18062 14571
rect 18384 14473 18418 14571
rect 18998 14564 19020 14580
rect 10506 11773 10615 11798
rect 10506 11733 10538 11773
rect 10585 11733 10615 11773
rect 10506 11714 10615 11733
rect 11626 10162 11702 10178
rect 11140 10144 11228 10160
rect 11670 9962 11702 9978
rect 21276 10012 21342 10028
rect 18988 9606 19020 9622
rect 21312 9878 21342 9894
rect 18988 9502 19066 9518
rect 9870 9382 9886 9442
rect 9948 9382 9964 9408
rect 7702 5946 8068 5980
rect 7874 5618 7908 5946
rect 8510 5670 11548 5716
rect 7842 5600 7948 5618
rect 7842 5564 7876 5600
rect 7912 5564 7948 5600
rect 7842 5554 7948 5564
rect 19991 9017 20261 9053
rect 19991 8932 20025 9017
rect 19790 8892 20025 8932
rect 19790 7477 19824 8892
rect 19991 8880 20025 8892
rect 20227 8880 20261 9017
rect 19035 7473 19824 7477
rect 18734 7463 19824 7473
rect 18734 7381 18746 7463
rect 18836 7381 19824 7463
rect 18734 7373 19824 7381
rect 18734 7370 19050 7373
rect 19790 5028 19824 7373
rect 20276 4598 20368 4616
rect 20276 4552 20296 4598
rect 20350 4552 20368 4598
rect 20276 4520 20368 4552
rect 20276 4470 20296 4520
rect 20350 4470 20368 4520
rect 20276 4452 20368 4470
rect 20926 4398 20942 4586
rect 18980 4254 18996 4398
rect 20926 4250 20942 4254
rect 21318 4250 21334 4586
rect 18998 3944 19002 3960
rect 11926 516 11960 686
rect 12162 516 12196 686
rect 12398 516 12432 685
rect 12634 516 12668 686
rect 11926 498 12668 516
rect 11925 482 12668 498
rect 13271 501 13305 687
rect 13507 501 13541 686
rect 13743 501 13777 687
rect 11925 348 12016 482
rect 13271 467 13931 501
rect 11917 335 12024 348
rect 11876 333 12024 335
rect 11876 270 11927 333
rect 11989 270 12024 333
rect 11876 258 12024 270
rect 11876 248 12016 258
rect 13876 144 13926 467
rect 17494 463 17528 634
rect 17849 463 17884 634
rect 18206 464 18240 635
rect 18086 463 18240 464
rect 17451 450 18240 463
rect 17451 441 17990 450
rect 17451 384 17469 441
rect 17555 384 17990 441
rect 17451 380 17990 384
rect 18080 380 18240 450
rect 17451 363 18240 380
rect 14233 150 14947 152
rect 13960 144 14947 150
rect 13876 140 14947 144
rect 13876 102 14875 140
rect 13960 77 14875 102
rect 14937 77 14947 140
rect 13960 63 14947 77
rect 13960 26 14051 63
rect 14233 62 14947 63
rect 19248 3944 19256 3960
rect 19248 -402 19320 -386
rect 13716 -488 13790 -472
rect 11496 -884 11548 -868
rect 13700 -1000 13716 -956
rect 13790 -1000 13806 -964
rect 11496 -1016 11598 -1000
rect 19220 -1036 19320 -1020
<< viali >>
rect 10538 11733 10585 11773
rect 7876 5564 7912 5600
rect 18746 7381 18836 7463
rect 20296 4470 20350 4520
rect 11927 270 11989 333
rect 17990 380 18080 450
rect 14875 77 14937 140
<< metal1 >>
rect 13861 14642 16935 14675
rect 10506 11773 10615 11783
rect 10506 11733 10538 11773
rect 10585 11733 10615 11773
rect 10506 11688 10615 11733
rect 10511 11448 10611 11688
rect 10511 11395 10524 11448
rect 10601 11395 10611 11448
rect 11850 11432 13598 11504
rect 10511 11378 10611 11395
rect 11851 11096 11917 11432
rect 12398 11254 13262 11295
rect 1954 6156 2204 6258
rect 1940 6134 2916 6156
rect 1940 6064 7502 6134
rect 8256 6112 11008 6120
rect 8256 6102 11440 6112
rect 8256 6078 11442 6102
rect 1940 6040 7512 6064
rect 1940 5918 2916 6040
rect 1954 4270 2204 5918
rect 7442 5854 7512 6040
rect 8258 5852 8328 6078
rect 10936 6070 11442 6078
rect 4632 4994 5236 5418
rect 7342 4994 7376 5794
rect 7866 5600 7922 5612
rect 7866 5564 7876 5600
rect 7912 5564 7922 5600
rect 7866 5190 7922 5564
rect 7866 5188 7936 5190
rect 7866 5184 7872 5188
rect 7858 5134 7872 5184
rect 7924 5134 7936 5188
rect 7858 5122 7936 5134
rect 8158 4994 8192 5793
rect 4632 4928 8192 4994
rect 4632 4918 7388 4928
rect 8158 4920 8192 4928
rect 4632 4728 5236 4918
rect 1952 -1272 2204 4270
rect 3651 2325 3751 2342
rect 3651 2272 3661 2325
rect 3738 2272 3751 2325
rect 3651 2072 3751 2272
rect 3653 -234 3750 2072
rect 11322 1060 11442 6070
rect 11332 520 11428 1060
rect 11808 571 11842 11052
rect 11926 700 11960 11052
rect 12044 571 12078 11052
rect 12162 700 12196 11052
rect 12280 571 12314 11052
rect 12398 700 12432 11254
rect 13196 11097 13262 11254
rect 12516 571 12550 11052
rect 12634 700 12668 11052
rect 12752 571 12786 11052
rect 11808 570 12786 571
rect 13153 573 13187 11053
rect 13271 701 13305 11053
rect 13389 573 13423 11053
rect 13507 701 13541 11432
rect 13625 573 13659 11053
rect 13743 701 13777 11212
rect 13861 573 13895 14642
rect 13979 1305 14013 11053
rect 13979 701 14013 1020
rect 14097 573 14131 11053
rect 14747 634 14781 14444
rect 14925 634 14959 14642
rect 15103 634 15137 14444
rect 15281 634 15315 14642
rect 15459 634 15493 14444
rect 15637 634 15671 14642
rect 15815 634 15849 14444
rect 15993 634 16027 14642
rect 16171 634 16205 14444
rect 16349 634 16383 14642
rect 16527 634 16561 14444
rect 16705 634 16739 14642
rect 16883 634 16917 14444
rect 20480 10991 21484 11045
rect 20480 10904 21490 10991
rect 20483 9309 20571 10904
rect 21390 10842 21490 10904
rect 21390 10789 21403 10842
rect 21480 10789 21490 10842
rect 21390 10772 21490 10789
rect 20483 9306 20588 9309
rect 19670 9207 20588 9306
rect 19672 9123 19707 9207
rect 18717 7463 18855 7514
rect 18717 7381 18746 7463
rect 18836 7381 18855 7463
rect 18717 4143 18855 7381
rect 19672 4703 19706 9123
rect 20109 9092 20470 9160
rect 20109 4690 20143 9092
rect 20436 5604 20470 9092
rect 20375 5558 20526 5604
rect 20375 5474 20397 5558
rect 20498 5474 20526 5558
rect 20375 5425 20526 5474
rect 20436 4717 20470 5425
rect 20554 4717 20588 9207
rect 20284 4520 20364 4532
rect 20284 4470 20296 4520
rect 20350 4472 20364 4520
rect 27316 4472 27826 4764
rect 20350 4470 27826 4472
rect 20284 4424 27826 4470
rect 13153 570 14131 573
rect 11808 545 14131 570
rect 11808 543 13180 545
rect 12774 542 13180 543
rect 11190 518 11458 520
rect 10964 516 11458 518
rect 10962 460 11458 516
rect 10962 458 11232 460
rect 10962 360 10992 458
rect 17980 450 18086 464
rect 17980 380 17990 450
rect 18080 380 18086 450
rect 10962 342 11020 360
rect 11896 342 12005 346
rect 10962 334 12005 342
rect 10832 333 12005 334
rect 10832 320 11927 333
rect 10832 260 10839 320
rect 10899 270 11927 320
rect 11989 270 12005 333
rect 10899 260 12005 270
rect 17980 324 18086 380
rect 17980 262 17994 324
rect 18076 262 18086 324
rect 10832 248 11994 260
rect 10994 246 11994 248
rect 17980 234 18086 262
rect 14859 140 15144 150
rect 14859 77 14875 140
rect 14937 138 15144 140
rect 14937 78 15077 138
rect 15137 78 15144 138
rect 14937 77 15144 78
rect 14859 64 15144 77
rect 18717 -234 18876 4143
rect 27316 4138 27826 4424
rect 3653 -357 18876 -234
rect 3653 -364 12265 -357
rect 18717 -364 18876 -357
rect 3653 -841 3750 -364
rect 1952 -2274 2202 -1272
rect 1952 -2310 15146 -2274
rect 1952 -2506 14876 -2310
rect 2892 -2518 14876 -2506
rect 15098 -2518 15146 -2310
rect 2892 -2540 15146 -2518
<< via1 >>
rect 10524 11395 10601 11448
rect 7872 5134 7924 5188
rect 3661 2272 3738 2325
rect 21403 10789 21480 10842
rect 20397 5474 20498 5558
rect 10839 260 10899 320
rect 17994 262 18076 324
rect 15077 78 15137 138
rect 14876 -2518 15098 -2310
<< metal2 >>
rect 10513 11448 10609 11460
rect 10513 11395 10524 11448
rect 10601 11395 10609 11448
rect 10513 11274 10609 11395
rect 10513 11217 10527 11274
rect 10596 11217 10609 11274
rect 10513 11200 10609 11217
rect 21392 10842 21488 10854
rect 21392 10789 21403 10842
rect 21480 10789 21488 10842
rect 21392 10668 21488 10789
rect 21392 10611 21406 10668
rect 21475 10611 21488 10668
rect 21392 10594 21488 10611
rect 27871 8749 27955 8760
rect 27871 8689 27884 8749
rect 27943 8689 27955 8749
rect 27871 8650 27955 8689
rect 27871 8630 27958 8650
rect 27872 8386 27958 8630
rect 27878 8224 27950 8386
rect 31084 8224 31830 8638
rect 27770 7934 31830 8224
rect 24949 5607 25222 5669
rect 20389 5559 20534 5566
rect 22097 5560 23603 5564
rect 24949 5560 25004 5607
rect 22097 5559 25004 5560
rect 20389 5558 25004 5559
rect 20389 5474 20397 5558
rect 20498 5485 25004 5558
rect 20498 5480 22163 5485
rect 23566 5481 25004 5485
rect 20498 5479 20690 5480
rect 20498 5474 20534 5479
rect 20389 5467 20534 5474
rect 24949 5459 25004 5481
rect 25165 5459 25222 5607
rect 24949 5402 25222 5459
rect 8656 5212 8754 5252
rect 8656 5196 8670 5212
rect 8478 5194 8670 5196
rect 7866 5188 8670 5194
rect 7866 5134 7872 5188
rect 7924 5134 8670 5188
rect 7866 5130 8670 5134
rect 7866 5128 8492 5130
rect 8656 5124 8670 5130
rect 8744 5124 8754 5212
rect 8656 5094 8754 5124
rect 3653 2503 3749 2520
rect 3653 2446 3666 2503
rect 3735 2446 3749 2503
rect 3653 2325 3749 2446
rect 3653 2272 3661 2325
rect 3738 2272 3749 2325
rect 3653 2260 3749 2272
rect 10672 321 10915 333
rect 10672 262 10683 321
rect 10743 320 10915 321
rect 10743 262 10839 320
rect 10672 260 10839 262
rect 10899 260 10915 320
rect 10672 249 10915 260
rect 17982 324 18086 340
rect 17982 262 17994 324
rect 18076 262 18086 324
rect 15061 138 15304 149
rect 15061 78 15077 138
rect 15137 136 15304 138
rect 15137 78 15233 136
rect 15061 77 15233 78
rect 15293 77 15304 136
rect 15061 65 15304 77
rect 14916 -36 15088 -30
rect 15166 -36 15198 65
rect 17982 38 18086 262
rect 17982 -4 18090 38
rect 14904 -90 15212 -36
rect 14916 -1572 15088 -90
rect 17998 -1132 18090 -4
rect 14858 -1858 15138 -1572
rect 14858 -1938 15140 -1858
rect 14860 -2310 15140 -1938
rect 14860 -2518 14876 -2310
rect 15098 -2518 15140 -2310
rect 14860 -2538 15140 -2518
rect 17984 -2280 18090 -1132
rect 27884 -1968 29388 -1328
rect 31084 -1968 31830 7934
rect 27884 -2280 32036 -1968
rect 17984 -2714 32036 -2280
rect 17984 -2716 29388 -2714
rect 17984 -2812 18090 -2716
rect 27884 -2766 29388 -2716
<< via2 >>
rect 10527 11217 10596 11274
rect 21406 10611 21475 10668
rect 27884 8689 27943 8749
rect 25004 5459 25165 5607
rect 8670 5124 8744 5212
rect 3666 2446 3735 2503
rect 10683 262 10743 321
rect 15233 77 15293 136
<< metal3 >>
rect 10511 11274 10609 11282
rect 10511 11217 10527 11274
rect 10596 11217 10609 11274
rect 10511 11145 10609 11217
rect 10510 11127 10609 11145
rect 10510 11070 10608 11127
rect 10510 11004 10524 11070
rect 10595 11004 10608 11070
rect 10510 10990 10608 11004
rect 21390 10668 21488 10676
rect 21390 10611 21406 10668
rect 21475 10611 21488 10668
rect 21390 10539 21488 10611
rect 21389 10521 21488 10539
rect 21389 10464 21487 10521
rect 21389 10398 21403 10464
rect 21474 10398 21487 10464
rect 21389 10384 21487 10398
rect 27872 9007 27954 9014
rect 27872 8941 27880 9007
rect 27946 8941 27954 9007
rect 27872 8749 27954 8941
rect 27872 8689 27884 8749
rect 27943 8689 27954 8749
rect 27872 8675 27954 8689
rect 24976 5607 25186 5626
rect 24976 5459 25004 5607
rect 25165 5459 25186 5607
rect 24976 5396 25186 5459
rect 24975 5377 25186 5396
rect 24975 5251 25185 5377
rect 8920 5220 9504 5222
rect 8662 5212 9504 5220
rect 8662 5124 8670 5212
rect 8744 5202 9504 5212
rect 8744 5132 9426 5202
rect 9492 5132 9504 5202
rect 8744 5124 9504 5132
rect 8662 5112 9504 5124
rect 8662 5110 9050 5112
rect 24975 5108 25014 5251
rect 25147 5108 25185 5251
rect 24975 5054 25185 5108
rect 3654 2716 3752 2730
rect 3654 2650 3667 2716
rect 3738 2650 3752 2716
rect 3654 2593 3752 2650
rect 3653 2575 3752 2593
rect 3653 2503 3751 2575
rect 3653 2446 3666 2503
rect 3735 2446 3751 2503
rect 3653 2438 3751 2446
rect 10418 324 10757 332
rect 10418 258 10425 324
rect 10491 321 10757 324
rect 10491 262 10683 321
rect 10743 262 10757 321
rect 10491 258 10757 262
rect 10418 250 10757 258
rect 15219 140 15558 148
rect 15219 136 15485 140
rect 15219 77 15233 136
rect 15293 77 15485 136
rect 15219 74 15485 77
rect 15551 74 15558 140
rect 15219 66 15558 74
<< via3 >>
rect 10524 11004 10595 11070
rect 21403 10398 21474 10464
rect 27880 8941 27946 9007
rect 9426 5132 9492 5202
rect 25014 5108 25147 5251
rect 3667 2650 3738 2716
rect 10425 258 10491 324
rect 15485 74 15551 140
<< metal4 >>
rect 6868 26648 7320 27642
rect 6838 26618 26490 26648
rect 6838 26316 27998 26618
rect 6868 25324 7320 26316
rect 25190 26286 27998 26316
rect 27818 26194 27998 26286
rect 6718 25232 7496 25324
rect 6694 25144 9300 25232
rect 6694 24354 8120 25144
rect 9164 24354 9300 25144
rect 6694 24220 9300 24354
rect 6718 16028 7496 24220
rect 9286 17408 9938 17502
rect 9286 16636 9336 17408
rect 9844 16636 9938 17408
rect 9286 16504 9938 16636
rect 9606 15054 9814 16504
rect 11484 15800 11784 18366
rect 11480 15568 11816 15800
rect 26520 15570 26700 15598
rect 23712 15568 26730 15570
rect 11480 15474 26730 15568
rect 11504 15456 26730 15474
rect 11578 15448 26730 15456
rect 11578 15440 11746 15448
rect 23712 15418 26730 15448
rect 312 6846 804 7080
rect 9608 6846 9774 15054
rect 19296 14878 22118 14880
rect 10102 14806 22118 14878
rect 10102 14804 20162 14806
rect 10102 11550 10164 14804
rect 10102 11452 10168 11550
rect 10106 10400 10168 11452
rect 10514 11070 10605 11084
rect 10514 11004 10524 11070
rect 10595 11004 10605 11070
rect 10514 10927 10605 11004
rect 10509 10400 10605 10927
rect 10106 10300 10605 10400
rect 21393 10464 21484 10478
rect 21393 10398 21403 10464
rect 21474 10398 21484 10464
rect 21393 10321 21484 10398
rect 10132 10288 10605 10300
rect 312 6732 9774 6846
rect 312 6468 804 6732
rect 9608 6658 9774 6732
rect 3100 6446 10092 6658
rect 3130 -1290 3222 6446
rect 10509 5214 10605 10288
rect 9560 5208 10605 5214
rect 9416 5202 10605 5208
rect 9416 5132 9426 5202
rect 9492 5132 10605 5202
rect 9416 5124 10605 5132
rect 9560 5118 10605 5124
rect 3670 4042 5265 4050
rect 10509 4045 10605 5118
rect 21388 9504 21484 10321
rect 22028 9504 22118 14806
rect 24486 9504 25170 10282
rect 21388 9430 25170 9504
rect 21388 4131 21484 9430
rect 24486 9102 25170 9430
rect 24992 5251 25171 5264
rect 24992 5108 25014 5251
rect 25147 5108 25171 5251
rect 24992 4964 25171 5108
rect 21387 4089 21484 4131
rect 3670 4041 6842 4042
rect 3670 4027 7469 4041
rect 3657 3979 7469 4027
rect 9237 3980 11061 4045
rect 3657 3977 6842 3979
rect 3657 3974 5265 3977
rect 3657 3530 3752 3974
rect 5745 3595 5849 3977
rect 7363 3591 7467 3979
rect 9238 3783 9342 3980
rect 10957 3785 11061 3980
rect 20838 3990 22663 4089
rect 25035 4041 25128 4964
rect 20838 3730 20942 3990
rect 22558 3734 22662 3990
rect 24384 3942 26209 4041
rect 22558 3728 22684 3734
rect 22660 3668 22684 3728
rect 24466 3558 24569 3942
rect 26085 3556 26188 3942
rect 3657 2793 3753 3530
rect 3657 2716 3748 2793
rect 3657 2650 3667 2716
rect 3738 2650 3748 2716
rect 3657 2636 3748 2650
rect 5023 348 5127 604
rect 6642 348 6746 619
rect 8468 354 8572 595
rect 6904 348 8572 354
rect 4999 337 8572 348
rect 10187 348 10291 595
rect 10187 337 10507 348
rect 4999 324 10507 337
rect 4999 258 10425 324
rect 10491 258 10507 324
rect 20067 283 20172 550
rect 20537 283 20783 360
rect 21787 283 21892 553
rect 20067 281 21895 283
rect 23746 281 23850 569
rect 25365 281 25469 571
rect 20067 267 25469 281
rect 4999 241 10507 258
rect 6904 239 10507 241
rect 8467 230 10507 239
rect 9369 -596 9615 230
rect 10290 229 10507 230
rect 20071 201 25469 267
rect 20071 186 25466 201
rect 15566 176 25466 186
rect 15566 169 20783 176
rect 21663 173 25466 176
rect 15469 140 20783 169
rect 15469 74 15485 140
rect 15551 74 20783 140
rect 15469 50 20783 74
rect 15566 48 20783 50
rect 20537 -130 20783 48
rect 26520 -130 26700 15418
rect 27818 9230 28030 26194
rect 27834 9022 27972 9230
rect 27851 9007 27970 9022
rect 27851 8941 27880 9007
rect 27946 8941 27970 9007
rect 27851 8925 27970 8941
rect 30080 -130 30702 186
rect 20537 -208 30702 -130
rect 20632 -250 30702 -208
rect 9410 -1290 9592 -596
rect 30080 -630 30702 -250
rect 2964 -1472 9592 -1290
rect 9440 -1714 9592 -1472
<< via4 >>
rect 8120 24354 9164 25144
rect 9336 16636 9844 17408
<< metal5 >>
rect 9936 25220 10452 25262
rect 8074 25144 10452 25220
rect 8074 24354 8120 25144
rect 9164 24354 10452 25144
rect 8074 24276 10452 24354
rect 8074 24268 10402 24276
rect 9940 24246 10402 24268
use sky130_fd_pr__cap_var_lvt_HDS5MT  XC1
timestamp 1668702877
transform 1 0 7477 0 1 5717
box -293 -301 293 301
use sky130_fd_pr__cap_mim_m3_1_UTEGVV  XC4
timestamp 1668708426
transform 1 0 9379 0 1 2187
box -1609 -1600 1709 1600
use sky130_fd_pr__cap_mim_m3_1_R9ELCP  XC5
timestamp 1668714113
transform 1 0 5886 0 1 2097
box -1509 -1500 1609 1500
use sky130_fd_pr__cap_var_lvt_HDS5MT  XC6
timestamp 1668702877
transform 1 0 8293 0 1 5715
box -293 -301 293 301
use sky130_fd_pr__nfet_01v8_4E7PL2  XM2
timestamp 1668722322
transform 1 0 19748 0 1 4858
box -88 -255 88 255
use sky130_fd_pr__nfet_01v8_ALQQLP  XM3
timestamp 1668722322
transform 1 0 20126 0 1 6778
box -147 -2188 147 2188
use sky130_fd_pr__nfet_01v8_54NRFS  XM5
timestamp 1668714756
transform 1 0 15832 0 1 7539
box -1097 -7005 1097 7005
use sky130_fd_pr__nfet_01v8_QT5LHM  XM6
timestamp 1668718364
transform 1 0 17867 0 1 7553
box -563 -7005 563 7005
use sky130_fd_pr__nfet_01v8_YNDJ8L  XM8
timestamp 1669755697
transform 1 0 12297 0 1 5876
box -501 -5276 501 5276
use ind_PA  ind_PA_0
timestamp 1669522153
transform 0 -1 8096 1 0 14272
box 1200 -12000 11600 -2200
use ind_PA  ind_PA_1
timestamp 1669522153
transform -1 0 11140 0 1 19702
box 1200 -12000 11600 -2200
use sky130_fd_pr__cap_mim_m3_1_R9ELCP  sky130_fd_pr__cap_mim_m3_1_R9ELCP_0
timestamp 1668714113
transform 1 0 24607 0 1 2067
box -1509 -1500 1609 1500
use sky130_fd_pr__cap_mim_m3_1_UTEGVV  sky130_fd_pr__cap_mim_m3_1_UTEGVV_0
timestamp 1668708426
transform 1 0 20979 0 1 2137
box -1609 -1600 1709 1600
use sky130_fd_pr__nfet_01v8_4E7PL2  sky130_fd_pr__nfet_01v8_4E7PL2_0
timestamp 1668722322
transform 1 0 20512 0 1 4872
box -88 -255 88 255
use sky130_fd_pr__nfet_01v8_YNDJ8L  sky130_fd_pr__nfet_01v8_YNDJ8L_0
timestamp 1669755697
transform 1 0 13642 0 1 5877
box -501 -5276 501 5276
<< labels >>
rlabel metal4 312 6468 804 7080 1 Vy
port 1 n
rlabel metal4 30080 -630 30702 186 1 Vx
port 2 n
rlabel metal1 4632 4728 5236 5418 1 Vctr
port 4 n
rlabel metal4 24486 9102 25170 10282 1 GND
port 6 n
rlabel metal2 27884 -2766 29388 -1328 1 VDD
port 5 n
rlabel metal1 27316 4138 27826 4764 1 Vband
port 3 n
<< end >>
