magic
tech sky130A
magscale 1 2
timestamp 1666402782
<< metal3 >>
rect -1150 772 1149 800
rect -1150 -772 1065 772
rect 1129 -772 1149 772
rect -1150 -800 1149 -772
<< via3 >>
rect 1065 -772 1129 772
<< mimcap >>
rect -1050 660 950 700
rect -1050 -660 -1010 660
rect 910 -660 950 660
rect -1050 -700 950 -660
<< mimcapcontact >>
rect -1010 -660 910 660
<< metal4 >>
rect 1049 772 1145 788
rect -1011 660 911 661
rect -1011 -660 -1010 660
rect 910 -660 911 660
rect -1011 -661 911 -660
rect 1049 -772 1065 772
rect 1129 -772 1145 772
rect 1049 -788 1145 -772
<< properties >>
string FIXED_BBOX -1150 -800 1050 800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 7.0 val 146.46 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
