magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -228 1130 -92 1502
<< psubdiff >>
rect -202 1435 -118 1476
rect -202 1401 -176 1435
rect -142 1401 -118 1435
rect -202 1367 -118 1401
rect -202 1333 -176 1367
rect -142 1333 -118 1367
rect -202 1299 -118 1333
rect -202 1265 -176 1299
rect -142 1265 -118 1299
rect -202 1231 -118 1265
rect -202 1197 -176 1231
rect -142 1197 -118 1231
rect -202 1156 -118 1197
<< psubdiffcont >>
rect -176 1401 -142 1435
rect -176 1333 -142 1367
rect -176 1265 -142 1299
rect -176 1197 -142 1231
<< locali >>
rect -188 1435 -132 1460
rect -188 1401 -176 1435
rect -142 1401 -132 1435
rect -188 1367 -132 1401
rect -188 1333 -176 1367
rect -142 1333 -132 1367
rect -188 1299 -132 1333
rect -188 1265 -176 1299
rect -142 1265 -132 1299
rect -188 1231 -132 1265
rect -188 1197 -176 1231
rect -142 1197 -132 1231
rect -188 1174 -132 1197
use sky130_fd_pr__res_xhigh_po_0p35_YXA95U  sky130_fd_pr__res_xhigh_po_0p35_YXA95U_0
timestamp 1669522153
transform 1 0 15 0 1 1394
box -35 -732 35 732
<< labels >>
rlabel locali s -163 1248 -163 1248 4 gnd
port 1 nsew
<< end >>
