magic
tech sky130A
magscale 1 2
timestamp 1667020045
<< xpolycontact >>
rect -512 2100 -442 2532
rect -512 -2532 -442 -2100
rect -194 2100 -124 2532
rect -194 -2532 -124 -2100
rect 124 2100 194 2532
rect 124 -2532 194 -2100
rect 442 2100 512 2532
rect 442 -2532 512 -2100
<< xpolyres >>
rect -512 -2100 -442 2100
rect -194 -2100 -124 2100
rect 124 -2100 194 2100
rect 442 -2100 512 2100
<< locali >>
rect -124 2106 124 2526
rect -442 -2524 -194 -2104
rect 194 -2526 442 -2106
<< viali >>
rect -496 2117 -458 2514
rect -178 2117 -140 2514
rect 140 2117 178 2514
rect 458 2117 496 2514
rect -496 -2514 -458 -2117
rect -178 -2514 -140 -2117
rect 140 -2514 178 -2117
rect 458 -2514 496 -2117
<< metal1 >>
rect -502 2514 -452 2526
rect -502 2117 -496 2514
rect -458 2117 -452 2514
rect -502 2105 -452 2117
rect -184 2514 -134 2526
rect -184 2117 -178 2514
rect -140 2117 -134 2514
rect -184 2105 -134 2117
rect 134 2514 184 2526
rect 134 2117 140 2514
rect 178 2117 184 2514
rect 134 2105 184 2117
rect 452 2514 502 2526
rect 452 2117 458 2514
rect 496 2117 502 2514
rect 452 2105 502 2117
rect -502 -2117 -452 -2105
rect -502 -2514 -496 -2117
rect -458 -2514 -452 -2117
rect -502 -2526 -452 -2514
rect -184 -2117 -134 -2105
rect -184 -2514 -178 -2117
rect -140 -2514 -134 -2117
rect -184 -2526 -134 -2514
rect 134 -2117 184 -2105
rect 134 -2514 140 -2117
rect 178 -2514 184 -2117
rect 134 -2526 184 -2514
rect 452 -2117 502 -2105
rect 452 -2514 458 -2117
rect 496 -2514 502 -2117
rect 452 -2526 502 -2514
<< res0p35 >>
rect -514 -2102 -440 2102
rect -196 -2102 -122 2102
rect 122 -2102 196 2102
rect 440 -2102 514 2102
<< labels >>
rlabel viali -482 2316 -482 2316 1 top
rlabel viali 474 2258 474 2258 1 bot
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 21 m 1 nx 4 wmin 0.350 lmin 0.50 rho 2000 val 121.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
