magic
tech sky130A
magscale 1 2
timestamp 1666910672
<< nwell >>
rect -144 18 144 1218
rect 406 12 694 1212
<< pmos >>
rect -50 118 50 1118
rect 500 112 600 1112
<< pdiff >>
rect -108 1106 -50 1118
rect -108 130 -96 1106
rect -62 130 -50 1106
rect -108 118 -50 130
rect 50 1106 108 1118
rect 50 130 62 1106
rect 96 130 108 1106
rect 50 118 108 130
rect 442 1100 500 1112
rect 442 124 454 1100
rect 488 124 500 1100
rect 442 112 500 124
rect 600 1100 658 1112
rect 600 124 612 1100
rect 646 124 658 1100
rect 600 112 658 124
<< pdiffc >>
rect -96 130 -62 1106
rect 62 130 96 1106
rect 454 124 488 1100
rect 612 124 646 1100
<< poly >>
rect -50 1199 50 1215
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -50 1118 50 1165
rect 500 1193 600 1209
rect 500 1159 516 1193
rect 584 1159 600 1193
rect 500 1112 600 1159
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect 500 65 600 112
rect 500 31 516 65
rect 584 31 600 65
rect 500 15 600 31
<< polycont >>
rect -34 1165 34 1199
rect 516 1159 584 1193
rect -34 37 34 71
rect 516 31 584 65
<< locali >>
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect 500 1159 516 1193
rect 584 1159 600 1193
rect -96 1106 -62 1122
rect -96 114 -62 130
rect 62 1106 96 1122
rect 62 114 96 130
rect 454 1100 488 1116
rect 454 108 488 124
rect 612 1100 646 1116
rect 612 108 646 124
rect -50 37 -34 71
rect 34 37 50 71
rect 500 31 516 65
rect 584 31 600 65
<< viali >>
rect -34 1165 34 1199
rect 516 1159 584 1193
rect -96 130 -62 1106
rect 62 130 96 1106
rect 454 124 488 1100
rect 612 124 646 1100
rect -34 37 34 71
rect 516 31 584 65
<< metal1 >>
rect -46 1199 46 1205
rect -46 1165 -34 1199
rect 34 1165 46 1199
rect -46 1159 46 1165
rect 504 1193 596 1199
rect 504 1159 516 1193
rect 584 1159 596 1193
rect 504 1153 596 1159
rect -102 1106 -56 1118
rect -102 130 -96 1106
rect -62 130 -56 1106
rect -102 118 -56 130
rect 56 1106 102 1118
rect 56 130 62 1106
rect 96 130 102 1106
rect 56 118 102 130
rect 448 1100 494 1112
rect 448 124 454 1100
rect 488 124 494 1100
rect 448 112 494 124
rect 606 1100 652 1112
rect 606 124 612 1100
rect 646 124 652 1100
rect 606 112 652 124
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect 504 65 596 71
rect 504 31 516 65
rect 584 31 596 65
rect 504 25 596 31
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
