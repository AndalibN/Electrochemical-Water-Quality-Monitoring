magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 195 35 627
rect -35 -627 35 -195
<< ppolyres >>
rect -35 -195 35 195
<< viali >>
rect -17 573 17 607
rect -17 501 17 535
rect -17 429 17 463
rect -17 357 17 391
rect -17 285 17 319
rect -17 213 17 247
rect -17 -248 17 -214
rect -17 -320 17 -286
rect -17 -392 17 -358
rect -17 -464 17 -430
rect -17 -536 17 -502
rect -17 -608 17 -574
<< metal1 >>
rect -25 607 25 621
rect -25 573 -17 607
rect 17 573 25 607
rect -25 535 25 573
rect -25 501 -17 535
rect 17 501 25 535
rect -25 463 25 501
rect -25 429 -17 463
rect 17 429 25 463
rect -25 391 25 429
rect -25 357 -17 391
rect 17 357 25 391
rect -25 319 25 357
rect -25 285 -17 319
rect 17 285 25 319
rect -25 247 25 285
rect -25 213 -17 247
rect 17 213 25 247
rect -25 200 25 213
rect -25 -214 25 -200
rect -25 -248 -17 -214
rect 17 -248 25 -214
rect -25 -286 25 -248
rect -25 -320 -17 -286
rect 17 -320 25 -286
rect -25 -358 25 -320
rect -25 -392 -17 -358
rect 17 -392 25 -358
rect -25 -430 25 -392
rect -25 -464 -17 -430
rect 17 -464 25 -430
rect -25 -502 25 -464
rect -25 -536 -17 -502
rect 17 -536 25 -502
rect -25 -574 25 -536
rect -25 -608 -17 -574
rect 17 -608 25 -574
rect -25 -621 25 -608
<< end >>
