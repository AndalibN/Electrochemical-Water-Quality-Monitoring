magic
tech sky130A
timestamp 1664679546
<< nmos >>
rect -15 -21 15 21
<< ndiff >>
rect -44 15 -15 21
rect -44 -15 -38 15
rect -21 -15 -15 15
rect -44 -21 -15 -15
rect 15 15 44 21
rect 15 -15 21 15
rect 38 -15 44 15
rect 15 -21 44 -15
<< ndiffc >>
rect -38 -15 -21 15
rect 21 -15 38 15
<< poly >>
rect -15 21 15 34
rect -15 -34 15 -21
<< locali >>
rect -38 15 -21 23
rect -38 -23 -21 -15
rect 21 15 38 23
rect 21 -23 38 -15
<< viali >>
rect -38 -15 -21 15
rect 21 -15 38 15
<< metal1 >>
rect -41 15 -18 21
rect -41 -15 -38 15
rect -21 -15 -18 15
rect -41 -21 -18 -15
rect 18 15 41 21
rect 18 -15 21 15
rect 38 -15 41 15
rect 18 -21 41 -15
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
