magic
tech sky130A
magscale 1 2
timestamp 1667590273
<< xpolycontact >>
rect -35 4545 35 4977
rect -35 -4977 35 -4545
<< xpolyres >>
rect -35 -4545 35 4545
<< viali >>
rect -19 4562 19 4959
rect -19 -4959 19 -4562
<< metal1 >>
rect -25 4959 25 4971
rect -25 4562 -19 4959
rect 19 4562 25 4959
rect -25 4550 25 4562
rect -25 -4562 25 -4550
rect -25 -4959 -19 -4562
rect 19 -4959 25 -4562
rect -25 -4971 25 -4959
<< res0p35 >>
rect -37 -4547 37 4547
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 45.45 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 260.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
