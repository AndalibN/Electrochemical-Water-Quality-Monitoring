magic
tech sky130A
magscale 1 2
timestamp 1666829797
<< nmos >>
rect -1274 55 -1174 1055
rect -1002 55 -902 1055
rect -730 55 -630 1055
rect -458 55 -358 1055
rect -186 55 -86 1055
rect 86 55 186 1055
rect 358 55 458 1055
rect 630 55 730 1055
rect 902 55 1002 1055
rect 1174 55 1274 1055
rect -1274 -1055 -1174 -55
rect -1002 -1055 -902 -55
rect -730 -1055 -630 -55
rect -458 -1055 -358 -55
rect -186 -1055 -86 -55
rect 86 -1055 186 -55
rect 358 -1055 458 -55
rect 630 -1055 730 -55
rect 902 -1055 1002 -55
rect 1174 -1055 1274 -55
<< ndiff >>
rect -1332 1043 -1274 1055
rect -1332 67 -1320 1043
rect -1286 67 -1274 1043
rect -1332 55 -1274 67
rect -1174 1043 -1116 1055
rect -1174 67 -1162 1043
rect -1128 67 -1116 1043
rect -1174 55 -1116 67
rect -1060 1043 -1002 1055
rect -1060 67 -1048 1043
rect -1014 67 -1002 1043
rect -1060 55 -1002 67
rect -902 1043 -844 1055
rect -902 67 -890 1043
rect -856 67 -844 1043
rect -902 55 -844 67
rect -788 1043 -730 1055
rect -788 67 -776 1043
rect -742 67 -730 1043
rect -788 55 -730 67
rect -630 1043 -572 1055
rect -630 67 -618 1043
rect -584 67 -572 1043
rect -630 55 -572 67
rect -516 1043 -458 1055
rect -516 67 -504 1043
rect -470 67 -458 1043
rect -516 55 -458 67
rect -358 1043 -300 1055
rect -358 67 -346 1043
rect -312 67 -300 1043
rect -358 55 -300 67
rect -244 1043 -186 1055
rect -244 67 -232 1043
rect -198 67 -186 1043
rect -244 55 -186 67
rect -86 1043 -28 1055
rect -86 67 -74 1043
rect -40 67 -28 1043
rect -86 55 -28 67
rect 28 1043 86 1055
rect 28 67 40 1043
rect 74 67 86 1043
rect 28 55 86 67
rect 186 1043 244 1055
rect 186 67 198 1043
rect 232 67 244 1043
rect 186 55 244 67
rect 300 1043 358 1055
rect 300 67 312 1043
rect 346 67 358 1043
rect 300 55 358 67
rect 458 1043 516 1055
rect 458 67 470 1043
rect 504 67 516 1043
rect 458 55 516 67
rect 572 1043 630 1055
rect 572 67 584 1043
rect 618 67 630 1043
rect 572 55 630 67
rect 730 1043 788 1055
rect 730 67 742 1043
rect 776 67 788 1043
rect 730 55 788 67
rect 844 1043 902 1055
rect 844 67 856 1043
rect 890 67 902 1043
rect 844 55 902 67
rect 1002 1043 1060 1055
rect 1002 67 1014 1043
rect 1048 67 1060 1043
rect 1002 55 1060 67
rect 1116 1043 1174 1055
rect 1116 67 1128 1043
rect 1162 67 1174 1043
rect 1116 55 1174 67
rect 1274 1043 1332 1055
rect 1274 67 1286 1043
rect 1320 67 1332 1043
rect 1274 55 1332 67
rect -1332 -67 -1274 -55
rect -1332 -1043 -1320 -67
rect -1286 -1043 -1274 -67
rect -1332 -1055 -1274 -1043
rect -1174 -67 -1116 -55
rect -1174 -1043 -1162 -67
rect -1128 -1043 -1116 -67
rect -1174 -1055 -1116 -1043
rect -1060 -67 -1002 -55
rect -1060 -1043 -1048 -67
rect -1014 -1043 -1002 -67
rect -1060 -1055 -1002 -1043
rect -902 -67 -844 -55
rect -902 -1043 -890 -67
rect -856 -1043 -844 -67
rect -902 -1055 -844 -1043
rect -788 -67 -730 -55
rect -788 -1043 -776 -67
rect -742 -1043 -730 -67
rect -788 -1055 -730 -1043
rect -630 -67 -572 -55
rect -630 -1043 -618 -67
rect -584 -1043 -572 -67
rect -630 -1055 -572 -1043
rect -516 -67 -458 -55
rect -516 -1043 -504 -67
rect -470 -1043 -458 -67
rect -516 -1055 -458 -1043
rect -358 -67 -300 -55
rect -358 -1043 -346 -67
rect -312 -1043 -300 -67
rect -358 -1055 -300 -1043
rect -244 -67 -186 -55
rect -244 -1043 -232 -67
rect -198 -1043 -186 -67
rect -244 -1055 -186 -1043
rect -86 -67 -28 -55
rect -86 -1043 -74 -67
rect -40 -1043 -28 -67
rect -86 -1055 -28 -1043
rect 28 -67 86 -55
rect 28 -1043 40 -67
rect 74 -1043 86 -67
rect 28 -1055 86 -1043
rect 186 -67 244 -55
rect 186 -1043 198 -67
rect 232 -1043 244 -67
rect 186 -1055 244 -1043
rect 300 -67 358 -55
rect 300 -1043 312 -67
rect 346 -1043 358 -67
rect 300 -1055 358 -1043
rect 458 -67 516 -55
rect 458 -1043 470 -67
rect 504 -1043 516 -67
rect 458 -1055 516 -1043
rect 572 -67 630 -55
rect 572 -1043 584 -67
rect 618 -1043 630 -67
rect 572 -1055 630 -1043
rect 730 -67 788 -55
rect 730 -1043 742 -67
rect 776 -1043 788 -67
rect 730 -1055 788 -1043
rect 844 -67 902 -55
rect 844 -1043 856 -67
rect 890 -1043 902 -67
rect 844 -1055 902 -1043
rect 1002 -67 1060 -55
rect 1002 -1043 1014 -67
rect 1048 -1043 1060 -67
rect 1002 -1055 1060 -1043
rect 1116 -67 1174 -55
rect 1116 -1043 1128 -67
rect 1162 -1043 1174 -67
rect 1116 -1055 1174 -1043
rect 1274 -67 1332 -55
rect 1274 -1043 1286 -67
rect 1320 -1043 1332 -67
rect 1274 -1055 1332 -1043
<< ndiffc >>
rect -1320 67 -1286 1043
rect -1162 67 -1128 1043
rect -1048 67 -1014 1043
rect -890 67 -856 1043
rect -776 67 -742 1043
rect -618 67 -584 1043
rect -504 67 -470 1043
rect -346 67 -312 1043
rect -232 67 -198 1043
rect -74 67 -40 1043
rect 40 67 74 1043
rect 198 67 232 1043
rect 312 67 346 1043
rect 470 67 504 1043
rect 584 67 618 1043
rect 742 67 776 1043
rect 856 67 890 1043
rect 1014 67 1048 1043
rect 1128 67 1162 1043
rect 1286 67 1320 1043
rect -1320 -1043 -1286 -67
rect -1162 -1043 -1128 -67
rect -1048 -1043 -1014 -67
rect -890 -1043 -856 -67
rect -776 -1043 -742 -67
rect -618 -1043 -584 -67
rect -504 -1043 -470 -67
rect -346 -1043 -312 -67
rect -232 -1043 -198 -67
rect -74 -1043 -40 -67
rect 40 -1043 74 -67
rect 198 -1043 232 -67
rect 312 -1043 346 -67
rect 470 -1043 504 -67
rect 584 -1043 618 -67
rect 742 -1043 776 -67
rect 856 -1043 890 -67
rect 1014 -1043 1048 -67
rect 1128 -1043 1162 -67
rect 1286 -1043 1320 -67
<< poly >>
rect -1274 1127 -1174 1143
rect -1274 1093 -1258 1127
rect -1190 1093 -1174 1127
rect -1274 1055 -1174 1093
rect -1002 1127 -902 1143
rect -1002 1093 -986 1127
rect -918 1093 -902 1127
rect -1002 1055 -902 1093
rect -730 1127 -630 1143
rect -730 1093 -714 1127
rect -646 1093 -630 1127
rect -730 1055 -630 1093
rect -458 1127 -358 1143
rect -458 1093 -442 1127
rect -374 1093 -358 1127
rect -458 1055 -358 1093
rect -186 1127 -86 1143
rect -186 1093 -170 1127
rect -102 1093 -86 1127
rect -186 1055 -86 1093
rect 86 1127 186 1143
rect 86 1093 102 1127
rect 170 1093 186 1127
rect 86 1055 186 1093
rect 358 1127 458 1143
rect 358 1093 374 1127
rect 442 1093 458 1127
rect 358 1055 458 1093
rect 630 1127 730 1143
rect 630 1093 646 1127
rect 714 1093 730 1127
rect 630 1055 730 1093
rect 902 1127 1002 1143
rect 902 1093 918 1127
rect 986 1093 1002 1127
rect 902 1055 1002 1093
rect 1174 1127 1274 1143
rect 1174 1093 1190 1127
rect 1258 1093 1274 1127
rect 1174 1055 1274 1093
rect -1274 17 -1174 55
rect -1274 -17 -1258 17
rect -1190 -17 -1174 17
rect -1274 -55 -1174 -17
rect -1002 17 -902 55
rect -1002 -17 -986 17
rect -918 -17 -902 17
rect -1002 -55 -902 -17
rect -730 17 -630 55
rect -730 -17 -714 17
rect -646 -17 -630 17
rect -730 -55 -630 -17
rect -458 17 -358 55
rect -458 -17 -442 17
rect -374 -17 -358 17
rect -458 -55 -358 -17
rect -186 17 -86 55
rect -186 -17 -170 17
rect -102 -17 -86 17
rect -186 -55 -86 -17
rect 86 17 186 55
rect 86 -17 102 17
rect 170 -17 186 17
rect 86 -55 186 -17
rect 358 17 458 55
rect 358 -17 374 17
rect 442 -17 458 17
rect 358 -55 458 -17
rect 630 17 730 55
rect 630 -17 646 17
rect 714 -17 730 17
rect 630 -55 730 -17
rect 902 17 1002 55
rect 902 -17 918 17
rect 986 -17 1002 17
rect 902 -55 1002 -17
rect 1174 17 1274 55
rect 1174 -17 1190 17
rect 1258 -17 1274 17
rect 1174 -55 1274 -17
rect -1274 -1093 -1174 -1055
rect -1274 -1127 -1258 -1093
rect -1190 -1127 -1174 -1093
rect -1274 -1143 -1174 -1127
rect -1002 -1093 -902 -1055
rect -1002 -1127 -986 -1093
rect -918 -1127 -902 -1093
rect -1002 -1143 -902 -1127
rect -730 -1093 -630 -1055
rect -730 -1127 -714 -1093
rect -646 -1127 -630 -1093
rect -730 -1143 -630 -1127
rect -458 -1093 -358 -1055
rect -458 -1127 -442 -1093
rect -374 -1127 -358 -1093
rect -458 -1143 -358 -1127
rect -186 -1093 -86 -1055
rect -186 -1127 -170 -1093
rect -102 -1127 -86 -1093
rect -186 -1143 -86 -1127
rect 86 -1093 186 -1055
rect 86 -1127 102 -1093
rect 170 -1127 186 -1093
rect 86 -1143 186 -1127
rect 358 -1093 458 -1055
rect 358 -1127 374 -1093
rect 442 -1127 458 -1093
rect 358 -1143 458 -1127
rect 630 -1093 730 -1055
rect 630 -1127 646 -1093
rect 714 -1127 730 -1093
rect 630 -1143 730 -1127
rect 902 -1093 1002 -1055
rect 902 -1127 918 -1093
rect 986 -1127 1002 -1093
rect 902 -1143 1002 -1127
rect 1174 -1093 1274 -1055
rect 1174 -1127 1190 -1093
rect 1258 -1127 1274 -1093
rect 1174 -1143 1274 -1127
<< polycont >>
rect -1258 1093 -1190 1127
rect -986 1093 -918 1127
rect -714 1093 -646 1127
rect -442 1093 -374 1127
rect -170 1093 -102 1127
rect 102 1093 170 1127
rect 374 1093 442 1127
rect 646 1093 714 1127
rect 918 1093 986 1127
rect 1190 1093 1258 1127
rect -1258 -17 -1190 17
rect -986 -17 -918 17
rect -714 -17 -646 17
rect -442 -17 -374 17
rect -170 -17 -102 17
rect 102 -17 170 17
rect 374 -17 442 17
rect 646 -17 714 17
rect 918 -17 986 17
rect 1190 -17 1258 17
rect -1258 -1127 -1190 -1093
rect -986 -1127 -918 -1093
rect -714 -1127 -646 -1093
rect -442 -1127 -374 -1093
rect -170 -1127 -102 -1093
rect 102 -1127 170 -1093
rect 374 -1127 442 -1093
rect 646 -1127 714 -1093
rect 918 -1127 986 -1093
rect 1190 -1127 1258 -1093
<< locali >>
rect -1274 1093 -1258 1127
rect -1190 1093 -1174 1127
rect -1002 1093 -986 1127
rect -918 1093 -902 1127
rect -730 1093 -714 1127
rect -646 1093 -630 1127
rect -458 1093 -442 1127
rect -374 1093 -358 1127
rect -186 1093 -170 1127
rect -102 1093 -86 1127
rect 86 1093 102 1127
rect 170 1093 186 1127
rect 358 1093 374 1127
rect 442 1093 458 1127
rect 630 1093 646 1127
rect 714 1093 730 1127
rect 902 1093 918 1127
rect 986 1093 1002 1127
rect 1174 1093 1190 1127
rect 1258 1093 1274 1127
rect -1320 1043 -1286 1059
rect -1320 51 -1286 67
rect -1162 1043 -1128 1059
rect -1162 51 -1128 67
rect -1048 1043 -1014 1059
rect -1048 51 -1014 67
rect -890 1043 -856 1059
rect -890 51 -856 67
rect -776 1043 -742 1059
rect -776 51 -742 67
rect -618 1043 -584 1059
rect -618 51 -584 67
rect -504 1043 -470 1059
rect -504 51 -470 67
rect -346 1043 -312 1059
rect -346 51 -312 67
rect -232 1043 -198 1059
rect -232 51 -198 67
rect -74 1043 -40 1059
rect -74 51 -40 67
rect 40 1043 74 1059
rect 40 51 74 67
rect 198 1043 232 1059
rect 198 51 232 67
rect 312 1043 346 1059
rect 312 51 346 67
rect 470 1043 504 1059
rect 470 51 504 67
rect 584 1043 618 1059
rect 584 51 618 67
rect 742 1043 776 1059
rect 742 51 776 67
rect 856 1043 890 1059
rect 856 51 890 67
rect 1014 1043 1048 1059
rect 1014 51 1048 67
rect 1128 1043 1162 1059
rect 1128 51 1162 67
rect 1286 1043 1320 1059
rect 1286 51 1320 67
rect -1274 -17 -1258 17
rect -1190 -17 -1174 17
rect -1002 -17 -986 17
rect -918 -17 -902 17
rect -730 -17 -714 17
rect -646 -17 -630 17
rect -458 -17 -442 17
rect -374 -17 -358 17
rect -186 -17 -170 17
rect -102 -17 -86 17
rect 86 -17 102 17
rect 170 -17 186 17
rect 358 -17 374 17
rect 442 -17 458 17
rect 630 -17 646 17
rect 714 -17 730 17
rect 902 -17 918 17
rect 986 -17 1002 17
rect 1174 -17 1190 17
rect 1258 -17 1274 17
rect -1320 -67 -1286 -51
rect -1320 -1059 -1286 -1043
rect -1162 -67 -1128 -51
rect -1162 -1059 -1128 -1043
rect -1048 -67 -1014 -51
rect -1048 -1059 -1014 -1043
rect -890 -67 -856 -51
rect -890 -1059 -856 -1043
rect -776 -67 -742 -51
rect -776 -1059 -742 -1043
rect -618 -67 -584 -51
rect -618 -1059 -584 -1043
rect -504 -67 -470 -51
rect -504 -1059 -470 -1043
rect -346 -67 -312 -51
rect -346 -1059 -312 -1043
rect -232 -67 -198 -51
rect -232 -1059 -198 -1043
rect -74 -67 -40 -51
rect -74 -1059 -40 -1043
rect 40 -67 74 -51
rect 40 -1059 74 -1043
rect 198 -67 232 -51
rect 198 -1059 232 -1043
rect 312 -67 346 -51
rect 312 -1059 346 -1043
rect 470 -67 504 -51
rect 470 -1059 504 -1043
rect 584 -67 618 -51
rect 584 -1059 618 -1043
rect 742 -67 776 -51
rect 742 -1059 776 -1043
rect 856 -67 890 -51
rect 856 -1059 890 -1043
rect 1014 -67 1048 -51
rect 1014 -1059 1048 -1043
rect 1128 -67 1162 -51
rect 1128 -1059 1162 -1043
rect 1286 -67 1320 -51
rect 1286 -1059 1320 -1043
rect -1274 -1127 -1258 -1093
rect -1190 -1127 -1174 -1093
rect -1002 -1127 -986 -1093
rect -918 -1127 -902 -1093
rect -730 -1127 -714 -1093
rect -646 -1127 -630 -1093
rect -458 -1127 -442 -1093
rect -374 -1127 -358 -1093
rect -186 -1127 -170 -1093
rect -102 -1127 -86 -1093
rect 86 -1127 102 -1093
rect 170 -1127 186 -1093
rect 358 -1127 374 -1093
rect 442 -1127 458 -1093
rect 630 -1127 646 -1093
rect 714 -1127 730 -1093
rect 902 -1127 918 -1093
rect 986 -1127 1002 -1093
rect 1174 -1127 1190 -1093
rect 1258 -1127 1274 -1093
<< viali >>
rect -1258 1093 -1190 1127
rect -986 1093 -918 1127
rect -714 1093 -646 1127
rect -442 1093 -374 1127
rect -170 1093 -102 1127
rect 102 1093 170 1127
rect 374 1093 442 1127
rect 646 1093 714 1127
rect 918 1093 986 1127
rect 1190 1093 1258 1127
rect -1320 67 -1286 1043
rect -1162 67 -1128 1043
rect -1048 67 -1014 1043
rect -890 67 -856 1043
rect -776 67 -742 1043
rect -618 67 -584 1043
rect -504 67 -470 1043
rect -346 67 -312 1043
rect -232 67 -198 1043
rect -74 67 -40 1043
rect 40 67 74 1043
rect 198 67 232 1043
rect 312 67 346 1043
rect 470 67 504 1043
rect 584 67 618 1043
rect 742 67 776 1043
rect 856 67 890 1043
rect 1014 67 1048 1043
rect 1128 67 1162 1043
rect 1286 67 1320 1043
rect -1258 -17 -1190 17
rect -986 -17 -918 17
rect -714 -17 -646 17
rect -442 -17 -374 17
rect -170 -17 -102 17
rect 102 -17 170 17
rect 374 -17 442 17
rect 646 -17 714 17
rect 918 -17 986 17
rect 1190 -17 1258 17
rect -1320 -1043 -1286 -67
rect -1162 -1043 -1128 -67
rect -1048 -1043 -1014 -67
rect -890 -1043 -856 -67
rect -776 -1043 -742 -67
rect -618 -1043 -584 -67
rect -504 -1043 -470 -67
rect -346 -1043 -312 -67
rect -232 -1043 -198 -67
rect -74 -1043 -40 -67
rect 40 -1043 74 -67
rect 198 -1043 232 -67
rect 312 -1043 346 -67
rect 470 -1043 504 -67
rect 584 -1043 618 -67
rect 742 -1043 776 -67
rect 856 -1043 890 -67
rect 1014 -1043 1048 -67
rect 1128 -1043 1162 -67
rect 1286 -1043 1320 -67
rect -1258 -1127 -1190 -1093
rect -986 -1127 -918 -1093
rect -714 -1127 -646 -1093
rect -442 -1127 -374 -1093
rect -170 -1127 -102 -1093
rect 102 -1127 170 -1093
rect 374 -1127 442 -1093
rect 646 -1127 714 -1093
rect 918 -1127 986 -1093
rect 1190 -1127 1258 -1093
<< metal1 >>
rect -1270 1127 -1178 1133
rect -1270 1093 -1258 1127
rect -1190 1093 -1178 1127
rect -1270 1087 -1178 1093
rect -998 1127 -906 1133
rect -998 1093 -986 1127
rect -918 1093 -906 1127
rect -998 1087 -906 1093
rect -726 1127 -634 1133
rect -726 1093 -714 1127
rect -646 1093 -634 1127
rect -726 1087 -634 1093
rect -454 1127 -362 1133
rect -454 1093 -442 1127
rect -374 1093 -362 1127
rect -454 1087 -362 1093
rect -182 1127 -90 1133
rect -182 1093 -170 1127
rect -102 1093 -90 1127
rect -182 1087 -90 1093
rect 90 1127 182 1133
rect 90 1093 102 1127
rect 170 1093 182 1127
rect 90 1087 182 1093
rect 362 1127 454 1133
rect 362 1093 374 1127
rect 442 1093 454 1127
rect 362 1087 454 1093
rect 634 1127 726 1133
rect 634 1093 646 1127
rect 714 1093 726 1127
rect 634 1087 726 1093
rect 906 1127 998 1133
rect 906 1093 918 1127
rect 986 1093 998 1127
rect 906 1087 998 1093
rect 1178 1127 1270 1133
rect 1178 1093 1190 1127
rect 1258 1093 1270 1127
rect 1178 1087 1270 1093
rect -1326 1043 -1280 1055
rect -1326 67 -1320 1043
rect -1286 67 -1280 1043
rect -1326 55 -1280 67
rect -1168 1043 -1122 1055
rect -1168 67 -1162 1043
rect -1128 67 -1122 1043
rect -1168 55 -1122 67
rect -1054 1043 -1008 1055
rect -1054 67 -1048 1043
rect -1014 67 -1008 1043
rect -1054 55 -1008 67
rect -896 1043 -850 1055
rect -896 67 -890 1043
rect -856 67 -850 1043
rect -896 55 -850 67
rect -782 1043 -736 1055
rect -782 67 -776 1043
rect -742 67 -736 1043
rect -782 55 -736 67
rect -624 1043 -578 1055
rect -624 67 -618 1043
rect -584 67 -578 1043
rect -624 55 -578 67
rect -510 1043 -464 1055
rect -510 67 -504 1043
rect -470 67 -464 1043
rect -510 55 -464 67
rect -352 1043 -306 1055
rect -352 67 -346 1043
rect -312 67 -306 1043
rect -352 55 -306 67
rect -238 1043 -192 1055
rect -238 67 -232 1043
rect -198 67 -192 1043
rect -238 55 -192 67
rect -80 1043 -34 1055
rect -80 67 -74 1043
rect -40 67 -34 1043
rect -80 55 -34 67
rect 34 1043 80 1055
rect 34 67 40 1043
rect 74 67 80 1043
rect 34 55 80 67
rect 192 1043 238 1055
rect 192 67 198 1043
rect 232 67 238 1043
rect 192 55 238 67
rect 306 1043 352 1055
rect 306 67 312 1043
rect 346 67 352 1043
rect 306 55 352 67
rect 464 1043 510 1055
rect 464 67 470 1043
rect 504 67 510 1043
rect 464 55 510 67
rect 578 1043 624 1055
rect 578 67 584 1043
rect 618 67 624 1043
rect 578 55 624 67
rect 736 1043 782 1055
rect 736 67 742 1043
rect 776 67 782 1043
rect 736 55 782 67
rect 850 1043 896 1055
rect 850 67 856 1043
rect 890 67 896 1043
rect 850 55 896 67
rect 1008 1043 1054 1055
rect 1008 67 1014 1043
rect 1048 67 1054 1043
rect 1008 55 1054 67
rect 1122 1043 1168 1055
rect 1122 67 1128 1043
rect 1162 67 1168 1043
rect 1122 55 1168 67
rect 1280 1043 1326 1055
rect 1280 67 1286 1043
rect 1320 67 1326 1043
rect 1280 55 1326 67
rect -1270 17 -1178 23
rect -1270 -17 -1258 17
rect -1190 -17 -1178 17
rect -1270 -23 -1178 -17
rect -998 17 -906 23
rect -998 -17 -986 17
rect -918 -17 -906 17
rect -998 -23 -906 -17
rect -726 17 -634 23
rect -726 -17 -714 17
rect -646 -17 -634 17
rect -726 -23 -634 -17
rect -454 17 -362 23
rect -454 -17 -442 17
rect -374 -17 -362 17
rect -454 -23 -362 -17
rect -182 17 -90 23
rect -182 -17 -170 17
rect -102 -17 -90 17
rect -182 -23 -90 -17
rect 90 17 182 23
rect 90 -17 102 17
rect 170 -17 182 17
rect 90 -23 182 -17
rect 362 17 454 23
rect 362 -17 374 17
rect 442 -17 454 17
rect 362 -23 454 -17
rect 634 17 726 23
rect 634 -17 646 17
rect 714 -17 726 17
rect 634 -23 726 -17
rect 906 17 998 23
rect 906 -17 918 17
rect 986 -17 998 17
rect 906 -23 998 -17
rect 1178 17 1270 23
rect 1178 -17 1190 17
rect 1258 -17 1270 17
rect 1178 -23 1270 -17
rect -1326 -67 -1280 -55
rect -1326 -1043 -1320 -67
rect -1286 -1043 -1280 -67
rect -1326 -1055 -1280 -1043
rect -1168 -67 -1122 -55
rect -1168 -1043 -1162 -67
rect -1128 -1043 -1122 -67
rect -1168 -1055 -1122 -1043
rect -1054 -67 -1008 -55
rect -1054 -1043 -1048 -67
rect -1014 -1043 -1008 -67
rect -1054 -1055 -1008 -1043
rect -896 -67 -850 -55
rect -896 -1043 -890 -67
rect -856 -1043 -850 -67
rect -896 -1055 -850 -1043
rect -782 -67 -736 -55
rect -782 -1043 -776 -67
rect -742 -1043 -736 -67
rect -782 -1055 -736 -1043
rect -624 -67 -578 -55
rect -624 -1043 -618 -67
rect -584 -1043 -578 -67
rect -624 -1055 -578 -1043
rect -510 -67 -464 -55
rect -510 -1043 -504 -67
rect -470 -1043 -464 -67
rect -510 -1055 -464 -1043
rect -352 -67 -306 -55
rect -352 -1043 -346 -67
rect -312 -1043 -306 -67
rect -352 -1055 -306 -1043
rect -238 -67 -192 -55
rect -238 -1043 -232 -67
rect -198 -1043 -192 -67
rect -238 -1055 -192 -1043
rect -80 -67 -34 -55
rect -80 -1043 -74 -67
rect -40 -1043 -34 -67
rect -80 -1055 -34 -1043
rect 34 -67 80 -55
rect 34 -1043 40 -67
rect 74 -1043 80 -67
rect 34 -1055 80 -1043
rect 192 -67 238 -55
rect 192 -1043 198 -67
rect 232 -1043 238 -67
rect 192 -1055 238 -1043
rect 306 -67 352 -55
rect 306 -1043 312 -67
rect 346 -1043 352 -67
rect 306 -1055 352 -1043
rect 464 -67 510 -55
rect 464 -1043 470 -67
rect 504 -1043 510 -67
rect 464 -1055 510 -1043
rect 578 -67 624 -55
rect 578 -1043 584 -67
rect 618 -1043 624 -67
rect 578 -1055 624 -1043
rect 736 -67 782 -55
rect 736 -1043 742 -67
rect 776 -1043 782 -67
rect 736 -1055 782 -1043
rect 850 -67 896 -55
rect 850 -1043 856 -67
rect 890 -1043 896 -67
rect 850 -1055 896 -1043
rect 1008 -67 1054 -55
rect 1008 -1043 1014 -67
rect 1048 -1043 1054 -67
rect 1008 -1055 1054 -1043
rect 1122 -67 1168 -55
rect 1122 -1043 1128 -67
rect 1162 -1043 1168 -67
rect 1122 -1055 1168 -1043
rect 1280 -67 1326 -55
rect 1280 -1043 1286 -67
rect 1320 -1043 1326 -67
rect 1280 -1055 1326 -1043
rect -1270 -1093 -1178 -1087
rect -1270 -1127 -1258 -1093
rect -1190 -1127 -1178 -1093
rect -1270 -1133 -1178 -1127
rect -998 -1093 -906 -1087
rect -998 -1127 -986 -1093
rect -918 -1127 -906 -1093
rect -998 -1133 -906 -1127
rect -726 -1093 -634 -1087
rect -726 -1127 -714 -1093
rect -646 -1127 -634 -1093
rect -726 -1133 -634 -1127
rect -454 -1093 -362 -1087
rect -454 -1127 -442 -1093
rect -374 -1127 -362 -1093
rect -454 -1133 -362 -1127
rect -182 -1093 -90 -1087
rect -182 -1127 -170 -1093
rect -102 -1127 -90 -1093
rect -182 -1133 -90 -1127
rect 90 -1093 182 -1087
rect 90 -1127 102 -1093
rect 170 -1127 182 -1093
rect 90 -1133 182 -1127
rect 362 -1093 454 -1087
rect 362 -1127 374 -1093
rect 442 -1127 454 -1093
rect 362 -1133 454 -1127
rect 634 -1093 726 -1087
rect 634 -1127 646 -1093
rect 714 -1127 726 -1093
rect 634 -1133 726 -1127
rect 906 -1093 998 -1087
rect 906 -1127 918 -1093
rect 986 -1127 998 -1093
rect 906 -1133 998 -1127
rect 1178 -1093 1270 -1087
rect 1178 -1127 1190 -1093
rect 1258 -1127 1270 -1093
rect 1178 -1133 1270 -1127
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
