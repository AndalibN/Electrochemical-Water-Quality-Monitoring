magic
tech sky130B
timestamp 1658694498
<< metal4 >>
rect 2700 -3550 3200 700
rect 2700 -3700 2750 -3550
rect 2900 -3700 2950 -3550
rect 3100 -3700 3200 -3550
rect 2700 -3750 3200 -3700
rect 2700 -3900 2800 -3750
rect 2950 -3900 3000 -3750
rect 3150 -3900 3200 -3750
rect 2700 -4000 3200 -3900
<< via4 >>
rect 2750 -3700 2900 -3550
rect 2950 -3700 3100 -3550
rect 2800 -3900 2950 -3750
rect 3000 -3900 3150 -3750
<< metal5 >>
rect -500 0 11500 500
rect -500 -800 10700 -300
rect -500 -11000 0 -800
rect 300 -1600 9900 -1100
rect 300 -10200 800 -1600
rect 1100 -2400 9100 -1900
rect 1100 -9400 1600 -2400
rect 1900 -3200 8300 -2700
rect 1900 -8600 2400 -3200
rect 2700 -3550 3200 -3500
rect 2700 -3700 2750 -3550
rect 2900 -3700 2950 -3550
rect 3100 -3700 3200 -3550
rect 2700 -3750 3200 -3700
rect 2700 -3900 2800 -3750
rect 2950 -3900 3000 -3750
rect 3150 -3900 3200 -3750
rect 2700 -7800 3200 -3900
rect 7800 -7800 8300 -3200
rect 2700 -8300 8300 -7800
rect 8600 -8600 9100 -2400
rect 1900 -9100 9100 -8600
rect 9400 -9400 9900 -1600
rect 1100 -9900 9900 -9400
rect 10200 -10200 10700 -800
rect 300 -10700 10700 -10200
rect 11000 -11000 11500 0
rect -500 -11500 11500 -11000
<< end >>
