magic
tech sky130A
magscale 1 2
timestamp 1668708426
<< metal3 >>
rect -1609 1522 -10 1550
rect -1609 78 -94 1522
rect -30 78 -10 1522
rect -1609 50 -10 78
rect 110 1522 1709 1550
rect 110 78 1625 1522
rect 1689 78 1709 1522
rect 110 50 1709 78
rect -1609 -78 -10 -50
rect -1609 -1522 -94 -78
rect -30 -1522 -10 -78
rect -1609 -1550 -10 -1522
rect 110 -78 1709 -50
rect 110 -1522 1625 -78
rect 1689 -1522 1709 -78
rect 110 -1550 1709 -1522
<< via3 >>
rect -94 78 -30 1522
rect 1625 78 1689 1522
rect -94 -1522 -30 -78
rect 1625 -1522 1689 -78
<< mimcap >>
rect -1509 1410 -209 1450
rect -1509 190 -1469 1410
rect -249 190 -209 1410
rect -1509 150 -209 190
rect 210 1410 1510 1450
rect 210 190 250 1410
rect 1470 190 1510 1410
rect 210 150 1510 190
rect -1509 -190 -209 -150
rect -1509 -1410 -1469 -190
rect -249 -1410 -209 -190
rect -1509 -1450 -209 -1410
rect 210 -190 1510 -150
rect 210 -1410 250 -190
rect 1470 -1410 1510 -190
rect 210 -1450 1510 -1410
<< mimcapcontact >>
rect -1469 190 -249 1410
rect 250 190 1470 1410
rect -1469 -1410 -249 -190
rect 250 -1410 1470 -190
<< metal4 >>
rect -911 1411 -807 1600
rect -141 1538 -37 1600
rect -141 1522 -14 1538
rect -1470 1410 -248 1411
rect -1470 190 -1469 1410
rect -249 190 -248 1410
rect -1470 189 -248 190
rect -911 -189 -807 189
rect -141 78 -94 1522
rect -30 78 -14 1522
rect 808 1411 912 1600
rect 1578 1538 1682 1600
rect 1578 1522 1705 1538
rect 249 1410 1471 1411
rect 249 190 250 1410
rect 1470 190 1471 1410
rect 249 189 1471 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -1470 -190 -248 -189
rect -1470 -1410 -1469 -190
rect -249 -1410 -248 -190
rect -1470 -1411 -248 -1410
rect -911 -1600 -807 -1411
rect -141 -1522 -94 -78
rect -30 -1522 -14 -78
rect 808 -189 912 189
rect 1578 78 1625 1522
rect 1689 78 1705 1522
rect 1578 62 1705 78
rect 1578 -62 1682 62
rect 1578 -78 1705 -62
rect 249 -190 1471 -189
rect 249 -1410 250 -190
rect 1470 -1410 1471 -190
rect 249 -1411 1471 -1410
rect -141 -1538 -14 -1522
rect -141 -1600 -37 -1538
rect 808 -1600 912 -1411
rect 1578 -1522 1625 -78
rect 1689 -1522 1705 -78
rect 1578 -1538 1705 -1522
rect 1578 -1600 1682 -1538
<< properties >>
string FIXED_BBOX 10 50 1510 1550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6.5 l 6.5 val 89.44 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
