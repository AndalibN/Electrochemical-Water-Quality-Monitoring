magic
tech sky130A
magscale 1 2
timestamp 1668226266
<< error_p >>
rect -35 693 35 837
rect -35 -589 35 -445
<< xpolycontact >>
rect -35 1439 35 1871
rect -35 693 35 1125
rect -35 157 35 589
rect -35 -589 35 -157
rect -35 -1125 35 -693
rect -35 -1871 35 -1439
<< xpolyres >>
rect -35 1125 35 1439
rect -35 -157 35 157
rect -35 -1439 35 -1125
<< viali >>
rect -19 1456 19 1853
rect -19 711 19 1108
rect -19 174 19 571
rect -19 -571 19 -174
rect -19 -1108 19 -711
rect -19 -1853 19 -1456
<< metal1 >>
rect -25 1853 25 1865
rect -25 1456 -19 1853
rect 19 1456 25 1853
rect -25 1444 25 1456
rect -25 1108 25 1120
rect -25 711 -19 1108
rect 19 711 25 1108
rect -25 699 25 711
rect -25 571 25 583
rect -25 174 -19 571
rect 19 174 25 571
rect -25 162 25 174
rect -25 -174 25 -162
rect -25 -571 -19 -174
rect 19 -571 25 -174
rect -25 -583 25 -571
rect -25 -711 25 -699
rect -25 -1108 -19 -711
rect 19 -1108 25 -711
rect -25 -1120 25 -1108
rect -25 -1456 25 -1444
rect -25 -1853 -19 -1456
rect 19 -1853 25 -1456
rect -25 -1865 25 -1853
<< res0p35 >>
rect -37 1123 37 1441
rect -37 -159 37 159
rect -37 -1441 37 -1123
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 1.57 m 3 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 10.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
