magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -2890 2792 2889 2840
rect -2890 2728 2805 2792
rect 2869 2728 2889 2792
rect -2890 2712 2889 2728
rect -2890 2648 2805 2712
rect 2869 2648 2889 2712
rect -2890 2632 2889 2648
rect -2890 2568 2805 2632
rect 2869 2568 2889 2632
rect -2890 2552 2889 2568
rect -2890 2488 2805 2552
rect 2869 2488 2889 2552
rect -2890 2472 2889 2488
rect -2890 2408 2805 2472
rect 2869 2408 2889 2472
rect -2890 2392 2889 2408
rect -2890 2328 2805 2392
rect 2869 2328 2889 2392
rect -2890 2312 2889 2328
rect -2890 2248 2805 2312
rect 2869 2248 2889 2312
rect -2890 2232 2889 2248
rect -2890 2168 2805 2232
rect 2869 2168 2889 2232
rect -2890 2152 2889 2168
rect -2890 2088 2805 2152
rect 2869 2088 2889 2152
rect -2890 2072 2889 2088
rect -2890 2008 2805 2072
rect 2869 2008 2889 2072
rect -2890 1992 2889 2008
rect -2890 1928 2805 1992
rect 2869 1928 2889 1992
rect -2890 1912 2889 1928
rect -2890 1848 2805 1912
rect 2869 1848 2889 1912
rect -2890 1832 2889 1848
rect -2890 1768 2805 1832
rect 2869 1768 2889 1832
rect -2890 1752 2889 1768
rect -2890 1688 2805 1752
rect 2869 1688 2889 1752
rect -2890 1672 2889 1688
rect -2890 1608 2805 1672
rect 2869 1608 2889 1672
rect -2890 1592 2889 1608
rect -2890 1528 2805 1592
rect 2869 1528 2889 1592
rect -2890 1512 2889 1528
rect -2890 1448 2805 1512
rect 2869 1448 2889 1512
rect -2890 1432 2889 1448
rect -2890 1368 2805 1432
rect 2869 1368 2889 1432
rect -2890 1352 2889 1368
rect -2890 1288 2805 1352
rect 2869 1288 2889 1352
rect -2890 1272 2889 1288
rect -2890 1208 2805 1272
rect 2869 1208 2889 1272
rect -2890 1192 2889 1208
rect -2890 1128 2805 1192
rect 2869 1128 2889 1192
rect -2890 1112 2889 1128
rect -2890 1048 2805 1112
rect 2869 1048 2889 1112
rect -2890 1032 2889 1048
rect -2890 968 2805 1032
rect 2869 968 2889 1032
rect -2890 952 2889 968
rect -2890 888 2805 952
rect 2869 888 2889 952
rect -2890 872 2889 888
rect -2890 808 2805 872
rect 2869 808 2889 872
rect -2890 792 2889 808
rect -2890 728 2805 792
rect 2869 728 2889 792
rect -2890 712 2889 728
rect -2890 648 2805 712
rect 2869 648 2889 712
rect -2890 632 2889 648
rect -2890 568 2805 632
rect 2869 568 2889 632
rect -2890 552 2889 568
rect -2890 488 2805 552
rect 2869 488 2889 552
rect -2890 472 2889 488
rect -2890 408 2805 472
rect 2869 408 2889 472
rect -2890 392 2889 408
rect -2890 328 2805 392
rect 2869 328 2889 392
rect -2890 312 2889 328
rect -2890 248 2805 312
rect 2869 248 2889 312
rect -2890 232 2889 248
rect -2890 168 2805 232
rect 2869 168 2889 232
rect -2890 152 2889 168
rect -2890 88 2805 152
rect 2869 88 2889 152
rect -2890 72 2889 88
rect -2890 8 2805 72
rect 2869 8 2889 72
rect -2890 -8 2889 8
rect -2890 -72 2805 -8
rect 2869 -72 2889 -8
rect -2890 -88 2889 -72
rect -2890 -152 2805 -88
rect 2869 -152 2889 -88
rect -2890 -168 2889 -152
rect -2890 -232 2805 -168
rect 2869 -232 2889 -168
rect -2890 -248 2889 -232
rect -2890 -312 2805 -248
rect 2869 -312 2889 -248
rect -2890 -328 2889 -312
rect -2890 -392 2805 -328
rect 2869 -392 2889 -328
rect -2890 -408 2889 -392
rect -2890 -472 2805 -408
rect 2869 -472 2889 -408
rect -2890 -488 2889 -472
rect -2890 -552 2805 -488
rect 2869 -552 2889 -488
rect -2890 -568 2889 -552
rect -2890 -632 2805 -568
rect 2869 -632 2889 -568
rect -2890 -648 2889 -632
rect -2890 -712 2805 -648
rect 2869 -712 2889 -648
rect -2890 -728 2889 -712
rect -2890 -792 2805 -728
rect 2869 -792 2889 -728
rect -2890 -808 2889 -792
rect -2890 -872 2805 -808
rect 2869 -872 2889 -808
rect -2890 -888 2889 -872
rect -2890 -952 2805 -888
rect 2869 -952 2889 -888
rect -2890 -968 2889 -952
rect -2890 -1032 2805 -968
rect 2869 -1032 2889 -968
rect -2890 -1048 2889 -1032
rect -2890 -1112 2805 -1048
rect 2869 -1112 2889 -1048
rect -2890 -1128 2889 -1112
rect -2890 -1192 2805 -1128
rect 2869 -1192 2889 -1128
rect -2890 -1208 2889 -1192
rect -2890 -1272 2805 -1208
rect 2869 -1272 2889 -1208
rect -2890 -1288 2889 -1272
rect -2890 -1352 2805 -1288
rect 2869 -1352 2889 -1288
rect -2890 -1368 2889 -1352
rect -2890 -1432 2805 -1368
rect 2869 -1432 2889 -1368
rect -2890 -1448 2889 -1432
rect -2890 -1512 2805 -1448
rect 2869 -1512 2889 -1448
rect -2890 -1528 2889 -1512
rect -2890 -1592 2805 -1528
rect 2869 -1592 2889 -1528
rect -2890 -1608 2889 -1592
rect -2890 -1672 2805 -1608
rect 2869 -1672 2889 -1608
rect -2890 -1688 2889 -1672
rect -2890 -1752 2805 -1688
rect 2869 -1752 2889 -1688
rect -2890 -1768 2889 -1752
rect -2890 -1832 2805 -1768
rect 2869 -1832 2889 -1768
rect -2890 -1848 2889 -1832
rect -2890 -1912 2805 -1848
rect 2869 -1912 2889 -1848
rect -2890 -1928 2889 -1912
rect -2890 -1992 2805 -1928
rect 2869 -1992 2889 -1928
rect -2890 -2008 2889 -1992
rect -2890 -2072 2805 -2008
rect 2869 -2072 2889 -2008
rect -2890 -2088 2889 -2072
rect -2890 -2152 2805 -2088
rect 2869 -2152 2889 -2088
rect -2890 -2168 2889 -2152
rect -2890 -2232 2805 -2168
rect 2869 -2232 2889 -2168
rect -2890 -2248 2889 -2232
rect -2890 -2312 2805 -2248
rect 2869 -2312 2889 -2248
rect -2890 -2328 2889 -2312
rect -2890 -2392 2805 -2328
rect 2869 -2392 2889 -2328
rect -2890 -2408 2889 -2392
rect -2890 -2472 2805 -2408
rect 2869 -2472 2889 -2408
rect -2890 -2488 2889 -2472
rect -2890 -2552 2805 -2488
rect 2869 -2552 2889 -2488
rect -2890 -2568 2889 -2552
rect -2890 -2632 2805 -2568
rect 2869 -2632 2889 -2568
rect -2890 -2648 2889 -2632
rect -2890 -2712 2805 -2648
rect 2869 -2712 2889 -2648
rect -2890 -2728 2889 -2712
rect -2890 -2792 2805 -2728
rect 2869 -2792 2889 -2728
rect -2890 -2840 2889 -2792
<< via3 >>
rect 2805 2728 2869 2792
rect 2805 2648 2869 2712
rect 2805 2568 2869 2632
rect 2805 2488 2869 2552
rect 2805 2408 2869 2472
rect 2805 2328 2869 2392
rect 2805 2248 2869 2312
rect 2805 2168 2869 2232
rect 2805 2088 2869 2152
rect 2805 2008 2869 2072
rect 2805 1928 2869 1992
rect 2805 1848 2869 1912
rect 2805 1768 2869 1832
rect 2805 1688 2869 1752
rect 2805 1608 2869 1672
rect 2805 1528 2869 1592
rect 2805 1448 2869 1512
rect 2805 1368 2869 1432
rect 2805 1288 2869 1352
rect 2805 1208 2869 1272
rect 2805 1128 2869 1192
rect 2805 1048 2869 1112
rect 2805 968 2869 1032
rect 2805 888 2869 952
rect 2805 808 2869 872
rect 2805 728 2869 792
rect 2805 648 2869 712
rect 2805 568 2869 632
rect 2805 488 2869 552
rect 2805 408 2869 472
rect 2805 328 2869 392
rect 2805 248 2869 312
rect 2805 168 2869 232
rect 2805 88 2869 152
rect 2805 8 2869 72
rect 2805 -72 2869 -8
rect 2805 -152 2869 -88
rect 2805 -232 2869 -168
rect 2805 -312 2869 -248
rect 2805 -392 2869 -328
rect 2805 -472 2869 -408
rect 2805 -552 2869 -488
rect 2805 -632 2869 -568
rect 2805 -712 2869 -648
rect 2805 -792 2869 -728
rect 2805 -872 2869 -808
rect 2805 -952 2869 -888
rect 2805 -1032 2869 -968
rect 2805 -1112 2869 -1048
rect 2805 -1192 2869 -1128
rect 2805 -1272 2869 -1208
rect 2805 -1352 2869 -1288
rect 2805 -1432 2869 -1368
rect 2805 -1512 2869 -1448
rect 2805 -1592 2869 -1528
rect 2805 -1672 2869 -1608
rect 2805 -1752 2869 -1688
rect 2805 -1832 2869 -1768
rect 2805 -1912 2869 -1848
rect 2805 -1992 2869 -1928
rect 2805 -2072 2869 -2008
rect 2805 -2152 2869 -2088
rect 2805 -2232 2869 -2168
rect 2805 -2312 2869 -2248
rect 2805 -2392 2869 -2328
rect 2805 -2472 2869 -2408
rect 2805 -2552 2869 -2488
rect 2805 -2632 2869 -2568
rect 2805 -2712 2869 -2648
rect 2805 -2792 2869 -2728
<< mimcap >>
rect -2790 2672 2690 2740
rect -2790 -2672 -2722 2672
rect 2622 -2672 2690 2672
rect -2790 -2740 2690 -2672
<< mimcapcontact >>
rect -2722 -2672 2622 2672
<< metal4 >>
rect 2789 2792 2885 2828
rect 2789 2728 2805 2792
rect 2869 2728 2885 2792
rect 2789 2712 2885 2728
rect -2751 2672 2651 2701
rect -2751 -2672 -2722 2672
rect 2622 -2672 2651 2672
rect -2751 -2701 2651 -2672
rect 2789 2648 2805 2712
rect 2869 2648 2885 2712
rect 2789 2632 2885 2648
rect 2789 2568 2805 2632
rect 2869 2568 2885 2632
rect 2789 2552 2885 2568
rect 2789 2488 2805 2552
rect 2869 2488 2885 2552
rect 2789 2472 2885 2488
rect 2789 2408 2805 2472
rect 2869 2408 2885 2472
rect 2789 2392 2885 2408
rect 2789 2328 2805 2392
rect 2869 2328 2885 2392
rect 2789 2312 2885 2328
rect 2789 2248 2805 2312
rect 2869 2248 2885 2312
rect 2789 2232 2885 2248
rect 2789 2168 2805 2232
rect 2869 2168 2885 2232
rect 2789 2152 2885 2168
rect 2789 2088 2805 2152
rect 2869 2088 2885 2152
rect 2789 2072 2885 2088
rect 2789 2008 2805 2072
rect 2869 2008 2885 2072
rect 2789 1992 2885 2008
rect 2789 1928 2805 1992
rect 2869 1928 2885 1992
rect 2789 1912 2885 1928
rect 2789 1848 2805 1912
rect 2869 1848 2885 1912
rect 2789 1832 2885 1848
rect 2789 1768 2805 1832
rect 2869 1768 2885 1832
rect 2789 1752 2885 1768
rect 2789 1688 2805 1752
rect 2869 1688 2885 1752
rect 2789 1672 2885 1688
rect 2789 1608 2805 1672
rect 2869 1608 2885 1672
rect 2789 1592 2885 1608
rect 2789 1528 2805 1592
rect 2869 1528 2885 1592
rect 2789 1512 2885 1528
rect 2789 1448 2805 1512
rect 2869 1448 2885 1512
rect 2789 1432 2885 1448
rect 2789 1368 2805 1432
rect 2869 1368 2885 1432
rect 2789 1352 2885 1368
rect 2789 1288 2805 1352
rect 2869 1288 2885 1352
rect 2789 1272 2885 1288
rect 2789 1208 2805 1272
rect 2869 1208 2885 1272
rect 2789 1192 2885 1208
rect 2789 1128 2805 1192
rect 2869 1128 2885 1192
rect 2789 1112 2885 1128
rect 2789 1048 2805 1112
rect 2869 1048 2885 1112
rect 2789 1032 2885 1048
rect 2789 968 2805 1032
rect 2869 968 2885 1032
rect 2789 952 2885 968
rect 2789 888 2805 952
rect 2869 888 2885 952
rect 2789 872 2885 888
rect 2789 808 2805 872
rect 2869 808 2885 872
rect 2789 792 2885 808
rect 2789 728 2805 792
rect 2869 728 2885 792
rect 2789 712 2885 728
rect 2789 648 2805 712
rect 2869 648 2885 712
rect 2789 632 2885 648
rect 2789 568 2805 632
rect 2869 568 2885 632
rect 2789 552 2885 568
rect 2789 488 2805 552
rect 2869 488 2885 552
rect 2789 472 2885 488
rect 2789 408 2805 472
rect 2869 408 2885 472
rect 2789 392 2885 408
rect 2789 328 2805 392
rect 2869 328 2885 392
rect 2789 312 2885 328
rect 2789 248 2805 312
rect 2869 248 2885 312
rect 2789 232 2885 248
rect 2789 168 2805 232
rect 2869 168 2885 232
rect 2789 152 2885 168
rect 2789 88 2805 152
rect 2869 88 2885 152
rect 2789 72 2885 88
rect 2789 8 2805 72
rect 2869 8 2885 72
rect 2789 -8 2885 8
rect 2789 -72 2805 -8
rect 2869 -72 2885 -8
rect 2789 -88 2885 -72
rect 2789 -152 2805 -88
rect 2869 -152 2885 -88
rect 2789 -168 2885 -152
rect 2789 -232 2805 -168
rect 2869 -232 2885 -168
rect 2789 -248 2885 -232
rect 2789 -312 2805 -248
rect 2869 -312 2885 -248
rect 2789 -328 2885 -312
rect 2789 -392 2805 -328
rect 2869 -392 2885 -328
rect 2789 -408 2885 -392
rect 2789 -472 2805 -408
rect 2869 -472 2885 -408
rect 2789 -488 2885 -472
rect 2789 -552 2805 -488
rect 2869 -552 2885 -488
rect 2789 -568 2885 -552
rect 2789 -632 2805 -568
rect 2869 -632 2885 -568
rect 2789 -648 2885 -632
rect 2789 -712 2805 -648
rect 2869 -712 2885 -648
rect 2789 -728 2885 -712
rect 2789 -792 2805 -728
rect 2869 -792 2885 -728
rect 2789 -808 2885 -792
rect 2789 -872 2805 -808
rect 2869 -872 2885 -808
rect 2789 -888 2885 -872
rect 2789 -952 2805 -888
rect 2869 -952 2885 -888
rect 2789 -968 2885 -952
rect 2789 -1032 2805 -968
rect 2869 -1032 2885 -968
rect 2789 -1048 2885 -1032
rect 2789 -1112 2805 -1048
rect 2869 -1112 2885 -1048
rect 2789 -1128 2885 -1112
rect 2789 -1192 2805 -1128
rect 2869 -1192 2885 -1128
rect 2789 -1208 2885 -1192
rect 2789 -1272 2805 -1208
rect 2869 -1272 2885 -1208
rect 2789 -1288 2885 -1272
rect 2789 -1352 2805 -1288
rect 2869 -1352 2885 -1288
rect 2789 -1368 2885 -1352
rect 2789 -1432 2805 -1368
rect 2869 -1432 2885 -1368
rect 2789 -1448 2885 -1432
rect 2789 -1512 2805 -1448
rect 2869 -1512 2885 -1448
rect 2789 -1528 2885 -1512
rect 2789 -1592 2805 -1528
rect 2869 -1592 2885 -1528
rect 2789 -1608 2885 -1592
rect 2789 -1672 2805 -1608
rect 2869 -1672 2885 -1608
rect 2789 -1688 2885 -1672
rect 2789 -1752 2805 -1688
rect 2869 -1752 2885 -1688
rect 2789 -1768 2885 -1752
rect 2789 -1832 2805 -1768
rect 2869 -1832 2885 -1768
rect 2789 -1848 2885 -1832
rect 2789 -1912 2805 -1848
rect 2869 -1912 2885 -1848
rect 2789 -1928 2885 -1912
rect 2789 -1992 2805 -1928
rect 2869 -1992 2885 -1928
rect 2789 -2008 2885 -1992
rect 2789 -2072 2805 -2008
rect 2869 -2072 2885 -2008
rect 2789 -2088 2885 -2072
rect 2789 -2152 2805 -2088
rect 2869 -2152 2885 -2088
rect 2789 -2168 2885 -2152
rect 2789 -2232 2805 -2168
rect 2869 -2232 2885 -2168
rect 2789 -2248 2885 -2232
rect 2789 -2312 2805 -2248
rect 2869 -2312 2885 -2248
rect 2789 -2328 2885 -2312
rect 2789 -2392 2805 -2328
rect 2869 -2392 2885 -2328
rect 2789 -2408 2885 -2392
rect 2789 -2472 2805 -2408
rect 2869 -2472 2885 -2408
rect 2789 -2488 2885 -2472
rect 2789 -2552 2805 -2488
rect 2869 -2552 2885 -2488
rect 2789 -2568 2885 -2552
rect 2789 -2632 2805 -2568
rect 2869 -2632 2885 -2568
rect 2789 -2648 2885 -2632
rect 2789 -2712 2805 -2648
rect 2869 -2712 2885 -2648
rect 2789 -2728 2885 -2712
rect 2789 -2792 2805 -2728
rect 2869 -2792 2885 -2728
rect 2789 -2828 2885 -2792
<< properties >>
string FIXED_BBOX -2890 -2840 2790 2840
<< end >>
