magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -844 -994 846 1058
<< nmos >>
rect -760 -968 -660 1032
rect -602 -968 -502 1032
rect -444 -968 -344 1032
rect -286 -968 -186 1032
rect -128 -968 -28 1032
rect 30 -968 130 1032
rect 188 -968 288 1032
rect 346 -968 446 1032
rect 504 -968 604 1032
rect 662 -968 762 1032
<< ndiff >>
rect -818 1001 -760 1032
rect -818 967 -806 1001
rect -772 967 -760 1001
rect -818 933 -760 967
rect -818 899 -806 933
rect -772 899 -760 933
rect -818 865 -760 899
rect -818 831 -806 865
rect -772 831 -760 865
rect -818 797 -760 831
rect -818 763 -806 797
rect -772 763 -760 797
rect -818 729 -760 763
rect -818 695 -806 729
rect -772 695 -760 729
rect -818 661 -760 695
rect -818 627 -806 661
rect -772 627 -760 661
rect -818 593 -760 627
rect -818 559 -806 593
rect -772 559 -760 593
rect -818 525 -760 559
rect -818 491 -806 525
rect -772 491 -760 525
rect -818 457 -760 491
rect -818 423 -806 457
rect -772 423 -760 457
rect -818 389 -760 423
rect -818 355 -806 389
rect -772 355 -760 389
rect -818 321 -760 355
rect -818 287 -806 321
rect -772 287 -760 321
rect -818 253 -760 287
rect -818 219 -806 253
rect -772 219 -760 253
rect -818 185 -760 219
rect -818 151 -806 185
rect -772 151 -760 185
rect -818 117 -760 151
rect -818 83 -806 117
rect -772 83 -760 117
rect -818 49 -760 83
rect -818 15 -806 49
rect -772 15 -760 49
rect -818 -19 -760 15
rect -818 -53 -806 -19
rect -772 -53 -760 -19
rect -818 -87 -760 -53
rect -818 -121 -806 -87
rect -772 -121 -760 -87
rect -818 -155 -760 -121
rect -818 -189 -806 -155
rect -772 -189 -760 -155
rect -818 -223 -760 -189
rect -818 -257 -806 -223
rect -772 -257 -760 -223
rect -818 -291 -760 -257
rect -818 -325 -806 -291
rect -772 -325 -760 -291
rect -818 -359 -760 -325
rect -818 -393 -806 -359
rect -772 -393 -760 -359
rect -818 -427 -760 -393
rect -818 -461 -806 -427
rect -772 -461 -760 -427
rect -818 -495 -760 -461
rect -818 -529 -806 -495
rect -772 -529 -760 -495
rect -818 -563 -760 -529
rect -818 -597 -806 -563
rect -772 -597 -760 -563
rect -818 -631 -760 -597
rect -818 -665 -806 -631
rect -772 -665 -760 -631
rect -818 -699 -760 -665
rect -818 -733 -806 -699
rect -772 -733 -760 -699
rect -818 -767 -760 -733
rect -818 -801 -806 -767
rect -772 -801 -760 -767
rect -818 -835 -760 -801
rect -818 -869 -806 -835
rect -772 -869 -760 -835
rect -818 -903 -760 -869
rect -818 -937 -806 -903
rect -772 -937 -760 -903
rect -818 -968 -760 -937
rect -660 1001 -602 1032
rect -660 967 -648 1001
rect -614 967 -602 1001
rect -660 933 -602 967
rect -660 899 -648 933
rect -614 899 -602 933
rect -660 865 -602 899
rect -660 831 -648 865
rect -614 831 -602 865
rect -660 797 -602 831
rect -660 763 -648 797
rect -614 763 -602 797
rect -660 729 -602 763
rect -660 695 -648 729
rect -614 695 -602 729
rect -660 661 -602 695
rect -660 627 -648 661
rect -614 627 -602 661
rect -660 593 -602 627
rect -660 559 -648 593
rect -614 559 -602 593
rect -660 525 -602 559
rect -660 491 -648 525
rect -614 491 -602 525
rect -660 457 -602 491
rect -660 423 -648 457
rect -614 423 -602 457
rect -660 389 -602 423
rect -660 355 -648 389
rect -614 355 -602 389
rect -660 321 -602 355
rect -660 287 -648 321
rect -614 287 -602 321
rect -660 253 -602 287
rect -660 219 -648 253
rect -614 219 -602 253
rect -660 185 -602 219
rect -660 151 -648 185
rect -614 151 -602 185
rect -660 117 -602 151
rect -660 83 -648 117
rect -614 83 -602 117
rect -660 49 -602 83
rect -660 15 -648 49
rect -614 15 -602 49
rect -660 -19 -602 15
rect -660 -53 -648 -19
rect -614 -53 -602 -19
rect -660 -87 -602 -53
rect -660 -121 -648 -87
rect -614 -121 -602 -87
rect -660 -155 -602 -121
rect -660 -189 -648 -155
rect -614 -189 -602 -155
rect -660 -223 -602 -189
rect -660 -257 -648 -223
rect -614 -257 -602 -223
rect -660 -291 -602 -257
rect -660 -325 -648 -291
rect -614 -325 -602 -291
rect -660 -359 -602 -325
rect -660 -393 -648 -359
rect -614 -393 -602 -359
rect -660 -427 -602 -393
rect -660 -461 -648 -427
rect -614 -461 -602 -427
rect -660 -495 -602 -461
rect -660 -529 -648 -495
rect -614 -529 -602 -495
rect -660 -563 -602 -529
rect -660 -597 -648 -563
rect -614 -597 -602 -563
rect -660 -631 -602 -597
rect -660 -665 -648 -631
rect -614 -665 -602 -631
rect -660 -699 -602 -665
rect -660 -733 -648 -699
rect -614 -733 -602 -699
rect -660 -767 -602 -733
rect -660 -801 -648 -767
rect -614 -801 -602 -767
rect -660 -835 -602 -801
rect -660 -869 -648 -835
rect -614 -869 -602 -835
rect -660 -903 -602 -869
rect -660 -937 -648 -903
rect -614 -937 -602 -903
rect -660 -968 -602 -937
rect -502 1001 -444 1032
rect -502 967 -490 1001
rect -456 967 -444 1001
rect -502 933 -444 967
rect -502 899 -490 933
rect -456 899 -444 933
rect -502 865 -444 899
rect -502 831 -490 865
rect -456 831 -444 865
rect -502 797 -444 831
rect -502 763 -490 797
rect -456 763 -444 797
rect -502 729 -444 763
rect -502 695 -490 729
rect -456 695 -444 729
rect -502 661 -444 695
rect -502 627 -490 661
rect -456 627 -444 661
rect -502 593 -444 627
rect -502 559 -490 593
rect -456 559 -444 593
rect -502 525 -444 559
rect -502 491 -490 525
rect -456 491 -444 525
rect -502 457 -444 491
rect -502 423 -490 457
rect -456 423 -444 457
rect -502 389 -444 423
rect -502 355 -490 389
rect -456 355 -444 389
rect -502 321 -444 355
rect -502 287 -490 321
rect -456 287 -444 321
rect -502 253 -444 287
rect -502 219 -490 253
rect -456 219 -444 253
rect -502 185 -444 219
rect -502 151 -490 185
rect -456 151 -444 185
rect -502 117 -444 151
rect -502 83 -490 117
rect -456 83 -444 117
rect -502 49 -444 83
rect -502 15 -490 49
rect -456 15 -444 49
rect -502 -19 -444 15
rect -502 -53 -490 -19
rect -456 -53 -444 -19
rect -502 -87 -444 -53
rect -502 -121 -490 -87
rect -456 -121 -444 -87
rect -502 -155 -444 -121
rect -502 -189 -490 -155
rect -456 -189 -444 -155
rect -502 -223 -444 -189
rect -502 -257 -490 -223
rect -456 -257 -444 -223
rect -502 -291 -444 -257
rect -502 -325 -490 -291
rect -456 -325 -444 -291
rect -502 -359 -444 -325
rect -502 -393 -490 -359
rect -456 -393 -444 -359
rect -502 -427 -444 -393
rect -502 -461 -490 -427
rect -456 -461 -444 -427
rect -502 -495 -444 -461
rect -502 -529 -490 -495
rect -456 -529 -444 -495
rect -502 -563 -444 -529
rect -502 -597 -490 -563
rect -456 -597 -444 -563
rect -502 -631 -444 -597
rect -502 -665 -490 -631
rect -456 -665 -444 -631
rect -502 -699 -444 -665
rect -502 -733 -490 -699
rect -456 -733 -444 -699
rect -502 -767 -444 -733
rect -502 -801 -490 -767
rect -456 -801 -444 -767
rect -502 -835 -444 -801
rect -502 -869 -490 -835
rect -456 -869 -444 -835
rect -502 -903 -444 -869
rect -502 -937 -490 -903
rect -456 -937 -444 -903
rect -502 -968 -444 -937
rect -344 1001 -286 1032
rect -344 967 -332 1001
rect -298 967 -286 1001
rect -344 933 -286 967
rect -344 899 -332 933
rect -298 899 -286 933
rect -344 865 -286 899
rect -344 831 -332 865
rect -298 831 -286 865
rect -344 797 -286 831
rect -344 763 -332 797
rect -298 763 -286 797
rect -344 729 -286 763
rect -344 695 -332 729
rect -298 695 -286 729
rect -344 661 -286 695
rect -344 627 -332 661
rect -298 627 -286 661
rect -344 593 -286 627
rect -344 559 -332 593
rect -298 559 -286 593
rect -344 525 -286 559
rect -344 491 -332 525
rect -298 491 -286 525
rect -344 457 -286 491
rect -344 423 -332 457
rect -298 423 -286 457
rect -344 389 -286 423
rect -344 355 -332 389
rect -298 355 -286 389
rect -344 321 -286 355
rect -344 287 -332 321
rect -298 287 -286 321
rect -344 253 -286 287
rect -344 219 -332 253
rect -298 219 -286 253
rect -344 185 -286 219
rect -344 151 -332 185
rect -298 151 -286 185
rect -344 117 -286 151
rect -344 83 -332 117
rect -298 83 -286 117
rect -344 49 -286 83
rect -344 15 -332 49
rect -298 15 -286 49
rect -344 -19 -286 15
rect -344 -53 -332 -19
rect -298 -53 -286 -19
rect -344 -87 -286 -53
rect -344 -121 -332 -87
rect -298 -121 -286 -87
rect -344 -155 -286 -121
rect -344 -189 -332 -155
rect -298 -189 -286 -155
rect -344 -223 -286 -189
rect -344 -257 -332 -223
rect -298 -257 -286 -223
rect -344 -291 -286 -257
rect -344 -325 -332 -291
rect -298 -325 -286 -291
rect -344 -359 -286 -325
rect -344 -393 -332 -359
rect -298 -393 -286 -359
rect -344 -427 -286 -393
rect -344 -461 -332 -427
rect -298 -461 -286 -427
rect -344 -495 -286 -461
rect -344 -529 -332 -495
rect -298 -529 -286 -495
rect -344 -563 -286 -529
rect -344 -597 -332 -563
rect -298 -597 -286 -563
rect -344 -631 -286 -597
rect -344 -665 -332 -631
rect -298 -665 -286 -631
rect -344 -699 -286 -665
rect -344 -733 -332 -699
rect -298 -733 -286 -699
rect -344 -767 -286 -733
rect -344 -801 -332 -767
rect -298 -801 -286 -767
rect -344 -835 -286 -801
rect -344 -869 -332 -835
rect -298 -869 -286 -835
rect -344 -903 -286 -869
rect -344 -937 -332 -903
rect -298 -937 -286 -903
rect -344 -968 -286 -937
rect -186 1001 -128 1032
rect -186 967 -174 1001
rect -140 967 -128 1001
rect -186 933 -128 967
rect -186 899 -174 933
rect -140 899 -128 933
rect -186 865 -128 899
rect -186 831 -174 865
rect -140 831 -128 865
rect -186 797 -128 831
rect -186 763 -174 797
rect -140 763 -128 797
rect -186 729 -128 763
rect -186 695 -174 729
rect -140 695 -128 729
rect -186 661 -128 695
rect -186 627 -174 661
rect -140 627 -128 661
rect -186 593 -128 627
rect -186 559 -174 593
rect -140 559 -128 593
rect -186 525 -128 559
rect -186 491 -174 525
rect -140 491 -128 525
rect -186 457 -128 491
rect -186 423 -174 457
rect -140 423 -128 457
rect -186 389 -128 423
rect -186 355 -174 389
rect -140 355 -128 389
rect -186 321 -128 355
rect -186 287 -174 321
rect -140 287 -128 321
rect -186 253 -128 287
rect -186 219 -174 253
rect -140 219 -128 253
rect -186 185 -128 219
rect -186 151 -174 185
rect -140 151 -128 185
rect -186 117 -128 151
rect -186 83 -174 117
rect -140 83 -128 117
rect -186 49 -128 83
rect -186 15 -174 49
rect -140 15 -128 49
rect -186 -19 -128 15
rect -186 -53 -174 -19
rect -140 -53 -128 -19
rect -186 -87 -128 -53
rect -186 -121 -174 -87
rect -140 -121 -128 -87
rect -186 -155 -128 -121
rect -186 -189 -174 -155
rect -140 -189 -128 -155
rect -186 -223 -128 -189
rect -186 -257 -174 -223
rect -140 -257 -128 -223
rect -186 -291 -128 -257
rect -186 -325 -174 -291
rect -140 -325 -128 -291
rect -186 -359 -128 -325
rect -186 -393 -174 -359
rect -140 -393 -128 -359
rect -186 -427 -128 -393
rect -186 -461 -174 -427
rect -140 -461 -128 -427
rect -186 -495 -128 -461
rect -186 -529 -174 -495
rect -140 -529 -128 -495
rect -186 -563 -128 -529
rect -186 -597 -174 -563
rect -140 -597 -128 -563
rect -186 -631 -128 -597
rect -186 -665 -174 -631
rect -140 -665 -128 -631
rect -186 -699 -128 -665
rect -186 -733 -174 -699
rect -140 -733 -128 -699
rect -186 -767 -128 -733
rect -186 -801 -174 -767
rect -140 -801 -128 -767
rect -186 -835 -128 -801
rect -186 -869 -174 -835
rect -140 -869 -128 -835
rect -186 -903 -128 -869
rect -186 -937 -174 -903
rect -140 -937 -128 -903
rect -186 -968 -128 -937
rect -28 1001 30 1032
rect -28 967 -16 1001
rect 18 967 30 1001
rect -28 933 30 967
rect -28 899 -16 933
rect 18 899 30 933
rect -28 865 30 899
rect -28 831 -16 865
rect 18 831 30 865
rect -28 797 30 831
rect -28 763 -16 797
rect 18 763 30 797
rect -28 729 30 763
rect -28 695 -16 729
rect 18 695 30 729
rect -28 661 30 695
rect -28 627 -16 661
rect 18 627 30 661
rect -28 593 30 627
rect -28 559 -16 593
rect 18 559 30 593
rect -28 525 30 559
rect -28 491 -16 525
rect 18 491 30 525
rect -28 457 30 491
rect -28 423 -16 457
rect 18 423 30 457
rect -28 389 30 423
rect -28 355 -16 389
rect 18 355 30 389
rect -28 321 30 355
rect -28 287 -16 321
rect 18 287 30 321
rect -28 253 30 287
rect -28 219 -16 253
rect 18 219 30 253
rect -28 185 30 219
rect -28 151 -16 185
rect 18 151 30 185
rect -28 117 30 151
rect -28 83 -16 117
rect 18 83 30 117
rect -28 49 30 83
rect -28 15 -16 49
rect 18 15 30 49
rect -28 -19 30 15
rect -28 -53 -16 -19
rect 18 -53 30 -19
rect -28 -87 30 -53
rect -28 -121 -16 -87
rect 18 -121 30 -87
rect -28 -155 30 -121
rect -28 -189 -16 -155
rect 18 -189 30 -155
rect -28 -223 30 -189
rect -28 -257 -16 -223
rect 18 -257 30 -223
rect -28 -291 30 -257
rect -28 -325 -16 -291
rect 18 -325 30 -291
rect -28 -359 30 -325
rect -28 -393 -16 -359
rect 18 -393 30 -359
rect -28 -427 30 -393
rect -28 -461 -16 -427
rect 18 -461 30 -427
rect -28 -495 30 -461
rect -28 -529 -16 -495
rect 18 -529 30 -495
rect -28 -563 30 -529
rect -28 -597 -16 -563
rect 18 -597 30 -563
rect -28 -631 30 -597
rect -28 -665 -16 -631
rect 18 -665 30 -631
rect -28 -699 30 -665
rect -28 -733 -16 -699
rect 18 -733 30 -699
rect -28 -767 30 -733
rect -28 -801 -16 -767
rect 18 -801 30 -767
rect -28 -835 30 -801
rect -28 -869 -16 -835
rect 18 -869 30 -835
rect -28 -903 30 -869
rect -28 -937 -16 -903
rect 18 -937 30 -903
rect -28 -968 30 -937
rect 130 1001 188 1032
rect 130 967 142 1001
rect 176 967 188 1001
rect 130 933 188 967
rect 130 899 142 933
rect 176 899 188 933
rect 130 865 188 899
rect 130 831 142 865
rect 176 831 188 865
rect 130 797 188 831
rect 130 763 142 797
rect 176 763 188 797
rect 130 729 188 763
rect 130 695 142 729
rect 176 695 188 729
rect 130 661 188 695
rect 130 627 142 661
rect 176 627 188 661
rect 130 593 188 627
rect 130 559 142 593
rect 176 559 188 593
rect 130 525 188 559
rect 130 491 142 525
rect 176 491 188 525
rect 130 457 188 491
rect 130 423 142 457
rect 176 423 188 457
rect 130 389 188 423
rect 130 355 142 389
rect 176 355 188 389
rect 130 321 188 355
rect 130 287 142 321
rect 176 287 188 321
rect 130 253 188 287
rect 130 219 142 253
rect 176 219 188 253
rect 130 185 188 219
rect 130 151 142 185
rect 176 151 188 185
rect 130 117 188 151
rect 130 83 142 117
rect 176 83 188 117
rect 130 49 188 83
rect 130 15 142 49
rect 176 15 188 49
rect 130 -19 188 15
rect 130 -53 142 -19
rect 176 -53 188 -19
rect 130 -87 188 -53
rect 130 -121 142 -87
rect 176 -121 188 -87
rect 130 -155 188 -121
rect 130 -189 142 -155
rect 176 -189 188 -155
rect 130 -223 188 -189
rect 130 -257 142 -223
rect 176 -257 188 -223
rect 130 -291 188 -257
rect 130 -325 142 -291
rect 176 -325 188 -291
rect 130 -359 188 -325
rect 130 -393 142 -359
rect 176 -393 188 -359
rect 130 -427 188 -393
rect 130 -461 142 -427
rect 176 -461 188 -427
rect 130 -495 188 -461
rect 130 -529 142 -495
rect 176 -529 188 -495
rect 130 -563 188 -529
rect 130 -597 142 -563
rect 176 -597 188 -563
rect 130 -631 188 -597
rect 130 -665 142 -631
rect 176 -665 188 -631
rect 130 -699 188 -665
rect 130 -733 142 -699
rect 176 -733 188 -699
rect 130 -767 188 -733
rect 130 -801 142 -767
rect 176 -801 188 -767
rect 130 -835 188 -801
rect 130 -869 142 -835
rect 176 -869 188 -835
rect 130 -903 188 -869
rect 130 -937 142 -903
rect 176 -937 188 -903
rect 130 -968 188 -937
rect 288 1001 346 1032
rect 288 967 300 1001
rect 334 967 346 1001
rect 288 933 346 967
rect 288 899 300 933
rect 334 899 346 933
rect 288 865 346 899
rect 288 831 300 865
rect 334 831 346 865
rect 288 797 346 831
rect 288 763 300 797
rect 334 763 346 797
rect 288 729 346 763
rect 288 695 300 729
rect 334 695 346 729
rect 288 661 346 695
rect 288 627 300 661
rect 334 627 346 661
rect 288 593 346 627
rect 288 559 300 593
rect 334 559 346 593
rect 288 525 346 559
rect 288 491 300 525
rect 334 491 346 525
rect 288 457 346 491
rect 288 423 300 457
rect 334 423 346 457
rect 288 389 346 423
rect 288 355 300 389
rect 334 355 346 389
rect 288 321 346 355
rect 288 287 300 321
rect 334 287 346 321
rect 288 253 346 287
rect 288 219 300 253
rect 334 219 346 253
rect 288 185 346 219
rect 288 151 300 185
rect 334 151 346 185
rect 288 117 346 151
rect 288 83 300 117
rect 334 83 346 117
rect 288 49 346 83
rect 288 15 300 49
rect 334 15 346 49
rect 288 -19 346 15
rect 288 -53 300 -19
rect 334 -53 346 -19
rect 288 -87 346 -53
rect 288 -121 300 -87
rect 334 -121 346 -87
rect 288 -155 346 -121
rect 288 -189 300 -155
rect 334 -189 346 -155
rect 288 -223 346 -189
rect 288 -257 300 -223
rect 334 -257 346 -223
rect 288 -291 346 -257
rect 288 -325 300 -291
rect 334 -325 346 -291
rect 288 -359 346 -325
rect 288 -393 300 -359
rect 334 -393 346 -359
rect 288 -427 346 -393
rect 288 -461 300 -427
rect 334 -461 346 -427
rect 288 -495 346 -461
rect 288 -529 300 -495
rect 334 -529 346 -495
rect 288 -563 346 -529
rect 288 -597 300 -563
rect 334 -597 346 -563
rect 288 -631 346 -597
rect 288 -665 300 -631
rect 334 -665 346 -631
rect 288 -699 346 -665
rect 288 -733 300 -699
rect 334 -733 346 -699
rect 288 -767 346 -733
rect 288 -801 300 -767
rect 334 -801 346 -767
rect 288 -835 346 -801
rect 288 -869 300 -835
rect 334 -869 346 -835
rect 288 -903 346 -869
rect 288 -937 300 -903
rect 334 -937 346 -903
rect 288 -968 346 -937
rect 446 1001 504 1032
rect 446 967 458 1001
rect 492 967 504 1001
rect 446 933 504 967
rect 446 899 458 933
rect 492 899 504 933
rect 446 865 504 899
rect 446 831 458 865
rect 492 831 504 865
rect 446 797 504 831
rect 446 763 458 797
rect 492 763 504 797
rect 446 729 504 763
rect 446 695 458 729
rect 492 695 504 729
rect 446 661 504 695
rect 446 627 458 661
rect 492 627 504 661
rect 446 593 504 627
rect 446 559 458 593
rect 492 559 504 593
rect 446 525 504 559
rect 446 491 458 525
rect 492 491 504 525
rect 446 457 504 491
rect 446 423 458 457
rect 492 423 504 457
rect 446 389 504 423
rect 446 355 458 389
rect 492 355 504 389
rect 446 321 504 355
rect 446 287 458 321
rect 492 287 504 321
rect 446 253 504 287
rect 446 219 458 253
rect 492 219 504 253
rect 446 185 504 219
rect 446 151 458 185
rect 492 151 504 185
rect 446 117 504 151
rect 446 83 458 117
rect 492 83 504 117
rect 446 49 504 83
rect 446 15 458 49
rect 492 15 504 49
rect 446 -19 504 15
rect 446 -53 458 -19
rect 492 -53 504 -19
rect 446 -87 504 -53
rect 446 -121 458 -87
rect 492 -121 504 -87
rect 446 -155 504 -121
rect 446 -189 458 -155
rect 492 -189 504 -155
rect 446 -223 504 -189
rect 446 -257 458 -223
rect 492 -257 504 -223
rect 446 -291 504 -257
rect 446 -325 458 -291
rect 492 -325 504 -291
rect 446 -359 504 -325
rect 446 -393 458 -359
rect 492 -393 504 -359
rect 446 -427 504 -393
rect 446 -461 458 -427
rect 492 -461 504 -427
rect 446 -495 504 -461
rect 446 -529 458 -495
rect 492 -529 504 -495
rect 446 -563 504 -529
rect 446 -597 458 -563
rect 492 -597 504 -563
rect 446 -631 504 -597
rect 446 -665 458 -631
rect 492 -665 504 -631
rect 446 -699 504 -665
rect 446 -733 458 -699
rect 492 -733 504 -699
rect 446 -767 504 -733
rect 446 -801 458 -767
rect 492 -801 504 -767
rect 446 -835 504 -801
rect 446 -869 458 -835
rect 492 -869 504 -835
rect 446 -903 504 -869
rect 446 -937 458 -903
rect 492 -937 504 -903
rect 446 -968 504 -937
rect 604 1001 662 1032
rect 604 967 616 1001
rect 650 967 662 1001
rect 604 933 662 967
rect 604 899 616 933
rect 650 899 662 933
rect 604 865 662 899
rect 604 831 616 865
rect 650 831 662 865
rect 604 797 662 831
rect 604 763 616 797
rect 650 763 662 797
rect 604 729 662 763
rect 604 695 616 729
rect 650 695 662 729
rect 604 661 662 695
rect 604 627 616 661
rect 650 627 662 661
rect 604 593 662 627
rect 604 559 616 593
rect 650 559 662 593
rect 604 525 662 559
rect 604 491 616 525
rect 650 491 662 525
rect 604 457 662 491
rect 604 423 616 457
rect 650 423 662 457
rect 604 389 662 423
rect 604 355 616 389
rect 650 355 662 389
rect 604 321 662 355
rect 604 287 616 321
rect 650 287 662 321
rect 604 253 662 287
rect 604 219 616 253
rect 650 219 662 253
rect 604 185 662 219
rect 604 151 616 185
rect 650 151 662 185
rect 604 117 662 151
rect 604 83 616 117
rect 650 83 662 117
rect 604 49 662 83
rect 604 15 616 49
rect 650 15 662 49
rect 604 -19 662 15
rect 604 -53 616 -19
rect 650 -53 662 -19
rect 604 -87 662 -53
rect 604 -121 616 -87
rect 650 -121 662 -87
rect 604 -155 662 -121
rect 604 -189 616 -155
rect 650 -189 662 -155
rect 604 -223 662 -189
rect 604 -257 616 -223
rect 650 -257 662 -223
rect 604 -291 662 -257
rect 604 -325 616 -291
rect 650 -325 662 -291
rect 604 -359 662 -325
rect 604 -393 616 -359
rect 650 -393 662 -359
rect 604 -427 662 -393
rect 604 -461 616 -427
rect 650 -461 662 -427
rect 604 -495 662 -461
rect 604 -529 616 -495
rect 650 -529 662 -495
rect 604 -563 662 -529
rect 604 -597 616 -563
rect 650 -597 662 -563
rect 604 -631 662 -597
rect 604 -665 616 -631
rect 650 -665 662 -631
rect 604 -699 662 -665
rect 604 -733 616 -699
rect 650 -733 662 -699
rect 604 -767 662 -733
rect 604 -801 616 -767
rect 650 -801 662 -767
rect 604 -835 662 -801
rect 604 -869 616 -835
rect 650 -869 662 -835
rect 604 -903 662 -869
rect 604 -937 616 -903
rect 650 -937 662 -903
rect 604 -968 662 -937
rect 762 1001 820 1032
rect 762 967 774 1001
rect 808 967 820 1001
rect 762 933 820 967
rect 762 899 774 933
rect 808 899 820 933
rect 762 865 820 899
rect 762 831 774 865
rect 808 831 820 865
rect 762 797 820 831
rect 762 763 774 797
rect 808 763 820 797
rect 762 729 820 763
rect 762 695 774 729
rect 808 695 820 729
rect 762 661 820 695
rect 762 627 774 661
rect 808 627 820 661
rect 762 593 820 627
rect 762 559 774 593
rect 808 559 820 593
rect 762 525 820 559
rect 762 491 774 525
rect 808 491 820 525
rect 762 457 820 491
rect 762 423 774 457
rect 808 423 820 457
rect 762 389 820 423
rect 762 355 774 389
rect 808 355 820 389
rect 762 321 820 355
rect 762 287 774 321
rect 808 287 820 321
rect 762 253 820 287
rect 762 219 774 253
rect 808 219 820 253
rect 762 185 820 219
rect 762 151 774 185
rect 808 151 820 185
rect 762 117 820 151
rect 762 83 774 117
rect 808 83 820 117
rect 762 49 820 83
rect 762 15 774 49
rect 808 15 820 49
rect 762 -19 820 15
rect 762 -53 774 -19
rect 808 -53 820 -19
rect 762 -87 820 -53
rect 762 -121 774 -87
rect 808 -121 820 -87
rect 762 -155 820 -121
rect 762 -189 774 -155
rect 808 -189 820 -155
rect 762 -223 820 -189
rect 762 -257 774 -223
rect 808 -257 820 -223
rect 762 -291 820 -257
rect 762 -325 774 -291
rect 808 -325 820 -291
rect 762 -359 820 -325
rect 762 -393 774 -359
rect 808 -393 820 -359
rect 762 -427 820 -393
rect 762 -461 774 -427
rect 808 -461 820 -427
rect 762 -495 820 -461
rect 762 -529 774 -495
rect 808 -529 820 -495
rect 762 -563 820 -529
rect 762 -597 774 -563
rect 808 -597 820 -563
rect 762 -631 820 -597
rect 762 -665 774 -631
rect 808 -665 820 -631
rect 762 -699 820 -665
rect 762 -733 774 -699
rect 808 -733 820 -699
rect 762 -767 820 -733
rect 762 -801 774 -767
rect 808 -801 820 -767
rect 762 -835 820 -801
rect 762 -869 774 -835
rect 808 -869 820 -835
rect 762 -903 820 -869
rect 762 -937 774 -903
rect 808 -937 820 -903
rect 762 -968 820 -937
<< ndiffc >>
rect -806 967 -772 1001
rect -806 899 -772 933
rect -806 831 -772 865
rect -806 763 -772 797
rect -806 695 -772 729
rect -806 627 -772 661
rect -806 559 -772 593
rect -806 491 -772 525
rect -806 423 -772 457
rect -806 355 -772 389
rect -806 287 -772 321
rect -806 219 -772 253
rect -806 151 -772 185
rect -806 83 -772 117
rect -806 15 -772 49
rect -806 -53 -772 -19
rect -806 -121 -772 -87
rect -806 -189 -772 -155
rect -806 -257 -772 -223
rect -806 -325 -772 -291
rect -806 -393 -772 -359
rect -806 -461 -772 -427
rect -806 -529 -772 -495
rect -806 -597 -772 -563
rect -806 -665 -772 -631
rect -806 -733 -772 -699
rect -806 -801 -772 -767
rect -806 -869 -772 -835
rect -806 -937 -772 -903
rect -648 967 -614 1001
rect -648 899 -614 933
rect -648 831 -614 865
rect -648 763 -614 797
rect -648 695 -614 729
rect -648 627 -614 661
rect -648 559 -614 593
rect -648 491 -614 525
rect -648 423 -614 457
rect -648 355 -614 389
rect -648 287 -614 321
rect -648 219 -614 253
rect -648 151 -614 185
rect -648 83 -614 117
rect -648 15 -614 49
rect -648 -53 -614 -19
rect -648 -121 -614 -87
rect -648 -189 -614 -155
rect -648 -257 -614 -223
rect -648 -325 -614 -291
rect -648 -393 -614 -359
rect -648 -461 -614 -427
rect -648 -529 -614 -495
rect -648 -597 -614 -563
rect -648 -665 -614 -631
rect -648 -733 -614 -699
rect -648 -801 -614 -767
rect -648 -869 -614 -835
rect -648 -937 -614 -903
rect -490 967 -456 1001
rect -490 899 -456 933
rect -490 831 -456 865
rect -490 763 -456 797
rect -490 695 -456 729
rect -490 627 -456 661
rect -490 559 -456 593
rect -490 491 -456 525
rect -490 423 -456 457
rect -490 355 -456 389
rect -490 287 -456 321
rect -490 219 -456 253
rect -490 151 -456 185
rect -490 83 -456 117
rect -490 15 -456 49
rect -490 -53 -456 -19
rect -490 -121 -456 -87
rect -490 -189 -456 -155
rect -490 -257 -456 -223
rect -490 -325 -456 -291
rect -490 -393 -456 -359
rect -490 -461 -456 -427
rect -490 -529 -456 -495
rect -490 -597 -456 -563
rect -490 -665 -456 -631
rect -490 -733 -456 -699
rect -490 -801 -456 -767
rect -490 -869 -456 -835
rect -490 -937 -456 -903
rect -332 967 -298 1001
rect -332 899 -298 933
rect -332 831 -298 865
rect -332 763 -298 797
rect -332 695 -298 729
rect -332 627 -298 661
rect -332 559 -298 593
rect -332 491 -298 525
rect -332 423 -298 457
rect -332 355 -298 389
rect -332 287 -298 321
rect -332 219 -298 253
rect -332 151 -298 185
rect -332 83 -298 117
rect -332 15 -298 49
rect -332 -53 -298 -19
rect -332 -121 -298 -87
rect -332 -189 -298 -155
rect -332 -257 -298 -223
rect -332 -325 -298 -291
rect -332 -393 -298 -359
rect -332 -461 -298 -427
rect -332 -529 -298 -495
rect -332 -597 -298 -563
rect -332 -665 -298 -631
rect -332 -733 -298 -699
rect -332 -801 -298 -767
rect -332 -869 -298 -835
rect -332 -937 -298 -903
rect -174 967 -140 1001
rect -174 899 -140 933
rect -174 831 -140 865
rect -174 763 -140 797
rect -174 695 -140 729
rect -174 627 -140 661
rect -174 559 -140 593
rect -174 491 -140 525
rect -174 423 -140 457
rect -174 355 -140 389
rect -174 287 -140 321
rect -174 219 -140 253
rect -174 151 -140 185
rect -174 83 -140 117
rect -174 15 -140 49
rect -174 -53 -140 -19
rect -174 -121 -140 -87
rect -174 -189 -140 -155
rect -174 -257 -140 -223
rect -174 -325 -140 -291
rect -174 -393 -140 -359
rect -174 -461 -140 -427
rect -174 -529 -140 -495
rect -174 -597 -140 -563
rect -174 -665 -140 -631
rect -174 -733 -140 -699
rect -174 -801 -140 -767
rect -174 -869 -140 -835
rect -174 -937 -140 -903
rect -16 967 18 1001
rect -16 899 18 933
rect -16 831 18 865
rect -16 763 18 797
rect -16 695 18 729
rect -16 627 18 661
rect -16 559 18 593
rect -16 491 18 525
rect -16 423 18 457
rect -16 355 18 389
rect -16 287 18 321
rect -16 219 18 253
rect -16 151 18 185
rect -16 83 18 117
rect -16 15 18 49
rect -16 -53 18 -19
rect -16 -121 18 -87
rect -16 -189 18 -155
rect -16 -257 18 -223
rect -16 -325 18 -291
rect -16 -393 18 -359
rect -16 -461 18 -427
rect -16 -529 18 -495
rect -16 -597 18 -563
rect -16 -665 18 -631
rect -16 -733 18 -699
rect -16 -801 18 -767
rect -16 -869 18 -835
rect -16 -937 18 -903
rect 142 967 176 1001
rect 142 899 176 933
rect 142 831 176 865
rect 142 763 176 797
rect 142 695 176 729
rect 142 627 176 661
rect 142 559 176 593
rect 142 491 176 525
rect 142 423 176 457
rect 142 355 176 389
rect 142 287 176 321
rect 142 219 176 253
rect 142 151 176 185
rect 142 83 176 117
rect 142 15 176 49
rect 142 -53 176 -19
rect 142 -121 176 -87
rect 142 -189 176 -155
rect 142 -257 176 -223
rect 142 -325 176 -291
rect 142 -393 176 -359
rect 142 -461 176 -427
rect 142 -529 176 -495
rect 142 -597 176 -563
rect 142 -665 176 -631
rect 142 -733 176 -699
rect 142 -801 176 -767
rect 142 -869 176 -835
rect 142 -937 176 -903
rect 300 967 334 1001
rect 300 899 334 933
rect 300 831 334 865
rect 300 763 334 797
rect 300 695 334 729
rect 300 627 334 661
rect 300 559 334 593
rect 300 491 334 525
rect 300 423 334 457
rect 300 355 334 389
rect 300 287 334 321
rect 300 219 334 253
rect 300 151 334 185
rect 300 83 334 117
rect 300 15 334 49
rect 300 -53 334 -19
rect 300 -121 334 -87
rect 300 -189 334 -155
rect 300 -257 334 -223
rect 300 -325 334 -291
rect 300 -393 334 -359
rect 300 -461 334 -427
rect 300 -529 334 -495
rect 300 -597 334 -563
rect 300 -665 334 -631
rect 300 -733 334 -699
rect 300 -801 334 -767
rect 300 -869 334 -835
rect 300 -937 334 -903
rect 458 967 492 1001
rect 458 899 492 933
rect 458 831 492 865
rect 458 763 492 797
rect 458 695 492 729
rect 458 627 492 661
rect 458 559 492 593
rect 458 491 492 525
rect 458 423 492 457
rect 458 355 492 389
rect 458 287 492 321
rect 458 219 492 253
rect 458 151 492 185
rect 458 83 492 117
rect 458 15 492 49
rect 458 -53 492 -19
rect 458 -121 492 -87
rect 458 -189 492 -155
rect 458 -257 492 -223
rect 458 -325 492 -291
rect 458 -393 492 -359
rect 458 -461 492 -427
rect 458 -529 492 -495
rect 458 -597 492 -563
rect 458 -665 492 -631
rect 458 -733 492 -699
rect 458 -801 492 -767
rect 458 -869 492 -835
rect 458 -937 492 -903
rect 616 967 650 1001
rect 616 899 650 933
rect 616 831 650 865
rect 616 763 650 797
rect 616 695 650 729
rect 616 627 650 661
rect 616 559 650 593
rect 616 491 650 525
rect 616 423 650 457
rect 616 355 650 389
rect 616 287 650 321
rect 616 219 650 253
rect 616 151 650 185
rect 616 83 650 117
rect 616 15 650 49
rect 616 -53 650 -19
rect 616 -121 650 -87
rect 616 -189 650 -155
rect 616 -257 650 -223
rect 616 -325 650 -291
rect 616 -393 650 -359
rect 616 -461 650 -427
rect 616 -529 650 -495
rect 616 -597 650 -563
rect 616 -665 650 -631
rect 616 -733 650 -699
rect 616 -801 650 -767
rect 616 -869 650 -835
rect 616 -937 650 -903
rect 774 967 808 1001
rect 774 899 808 933
rect 774 831 808 865
rect 774 763 808 797
rect 774 695 808 729
rect 774 627 808 661
rect 774 559 808 593
rect 774 491 808 525
rect 774 423 808 457
rect 774 355 808 389
rect 774 287 808 321
rect 774 219 808 253
rect 774 151 808 185
rect 774 83 808 117
rect 774 15 808 49
rect 774 -53 808 -19
rect 774 -121 808 -87
rect 774 -189 808 -155
rect 774 -257 808 -223
rect 774 -325 808 -291
rect 774 -393 808 -359
rect 774 -461 808 -427
rect 774 -529 808 -495
rect 774 -597 808 -563
rect 774 -665 808 -631
rect 774 -733 808 -699
rect 774 -801 808 -767
rect 774 -869 808 -835
rect 774 -937 808 -903
<< poly >>
rect -760 1058 762 1108
rect -760 1032 -660 1058
rect -602 1032 -502 1058
rect -444 1032 -344 1058
rect -286 1032 -186 1058
rect -128 1032 -28 1058
rect 30 1032 130 1058
rect 188 1032 288 1058
rect 346 1032 446 1058
rect 504 1032 604 1058
rect 662 1032 762 1058
rect -760 -1006 -660 -968
rect -602 -1006 -502 -968
rect -444 -1006 -344 -968
rect -286 -1006 -186 -968
rect -128 -1006 -28 -968
rect 30 -1006 130 -968
rect 188 -1006 288 -968
rect 346 -1006 446 -968
rect 504 -1006 604 -968
rect 662 -1006 762 -968
rect -760 -1040 -736 -1006
rect -702 -1040 762 -1006
rect -760 -1056 762 -1040
<< polycont >>
rect -736 -1040 -702 -1006
<< locali >>
rect -806 1001 -772 1036
rect -806 933 -772 951
rect -806 865 -772 879
rect -806 797 -772 807
rect -806 729 -772 735
rect -806 661 -772 663
rect -806 625 -772 627
rect -806 553 -772 559
rect -806 481 -772 491
rect -806 409 -772 423
rect -806 337 -772 355
rect -806 265 -772 287
rect -806 193 -772 219
rect -806 121 -772 151
rect -806 49 -772 83
rect -806 -19 -772 15
rect -806 -87 -772 -57
rect -806 -155 -772 -129
rect -806 -223 -772 -201
rect -806 -291 -772 -273
rect -806 -359 -772 -345
rect -806 -427 -772 -417
rect -806 -495 -772 -489
rect -806 -563 -772 -561
rect -806 -599 -772 -597
rect -806 -671 -772 -665
rect -806 -743 -772 -733
rect -806 -815 -772 -801
rect -806 -887 -772 -869
rect -806 -972 -772 -937
rect -648 1001 -614 1036
rect -648 933 -614 951
rect -648 865 -614 879
rect -648 797 -614 807
rect -648 729 -614 735
rect -648 661 -614 663
rect -648 625 -614 627
rect -648 553 -614 559
rect -648 481 -614 491
rect -648 409 -614 423
rect -648 337 -614 355
rect -648 265 -614 287
rect -648 193 -614 219
rect -648 121 -614 151
rect -648 49 -614 83
rect -648 -19 -614 15
rect -648 -87 -614 -57
rect -648 -155 -614 -129
rect -648 -223 -614 -201
rect -648 -291 -614 -273
rect -648 -359 -614 -345
rect -648 -427 -614 -417
rect -648 -495 -614 -489
rect -648 -563 -614 -561
rect -648 -599 -614 -597
rect -648 -671 -614 -665
rect -648 -743 -614 -733
rect -648 -815 -614 -801
rect -648 -887 -614 -869
rect -648 -972 -614 -937
rect -490 1001 -456 1036
rect -490 933 -456 951
rect -490 865 -456 879
rect -490 797 -456 807
rect -490 729 -456 735
rect -490 661 -456 663
rect -490 625 -456 627
rect -490 553 -456 559
rect -490 481 -456 491
rect -490 409 -456 423
rect -490 337 -456 355
rect -490 265 -456 287
rect -490 193 -456 219
rect -490 121 -456 151
rect -490 49 -456 83
rect -490 -19 -456 15
rect -490 -87 -456 -57
rect -490 -155 -456 -129
rect -490 -223 -456 -201
rect -490 -291 -456 -273
rect -490 -359 -456 -345
rect -490 -427 -456 -417
rect -490 -495 -456 -489
rect -490 -563 -456 -561
rect -490 -599 -456 -597
rect -490 -671 -456 -665
rect -490 -743 -456 -733
rect -490 -815 -456 -801
rect -490 -887 -456 -869
rect -490 -972 -456 -937
rect -332 1001 -298 1036
rect -332 933 -298 951
rect -332 865 -298 879
rect -332 797 -298 807
rect -332 729 -298 735
rect -332 661 -298 663
rect -332 625 -298 627
rect -332 553 -298 559
rect -332 481 -298 491
rect -332 409 -298 423
rect -332 337 -298 355
rect -332 265 -298 287
rect -332 193 -298 219
rect -332 121 -298 151
rect -332 49 -298 83
rect -332 -19 -298 15
rect -332 -87 -298 -57
rect -332 -155 -298 -129
rect -332 -223 -298 -201
rect -332 -291 -298 -273
rect -332 -359 -298 -345
rect -332 -427 -298 -417
rect -332 -495 -298 -489
rect -332 -563 -298 -561
rect -332 -599 -298 -597
rect -332 -671 -298 -665
rect -332 -743 -298 -733
rect -332 -815 -298 -801
rect -332 -887 -298 -869
rect -332 -972 -298 -937
rect -174 1001 -140 1036
rect -174 933 -140 951
rect -174 865 -140 879
rect -174 797 -140 807
rect -174 729 -140 735
rect -174 661 -140 663
rect -174 625 -140 627
rect -174 553 -140 559
rect -174 481 -140 491
rect -174 409 -140 423
rect -174 337 -140 355
rect -174 265 -140 287
rect -174 193 -140 219
rect -174 121 -140 151
rect -174 49 -140 83
rect -174 -19 -140 15
rect -174 -87 -140 -57
rect -174 -155 -140 -129
rect -174 -223 -140 -201
rect -174 -291 -140 -273
rect -174 -359 -140 -345
rect -174 -427 -140 -417
rect -174 -495 -140 -489
rect -174 -563 -140 -561
rect -174 -599 -140 -597
rect -174 -671 -140 -665
rect -174 -743 -140 -733
rect -174 -815 -140 -801
rect -174 -887 -140 -869
rect -174 -972 -140 -937
rect -16 1001 18 1036
rect -16 933 18 951
rect -16 865 18 879
rect -16 797 18 807
rect -16 729 18 735
rect -16 661 18 663
rect -16 625 18 627
rect -16 553 18 559
rect -16 481 18 491
rect -16 409 18 423
rect -16 337 18 355
rect -16 265 18 287
rect -16 193 18 219
rect -16 121 18 151
rect -16 49 18 83
rect -16 -19 18 15
rect -16 -87 18 -57
rect -16 -155 18 -129
rect -16 -223 18 -201
rect -16 -291 18 -273
rect -16 -359 18 -345
rect -16 -427 18 -417
rect -16 -495 18 -489
rect -16 -563 18 -561
rect -16 -599 18 -597
rect -16 -671 18 -665
rect -16 -743 18 -733
rect -16 -815 18 -801
rect -16 -887 18 -869
rect -16 -972 18 -937
rect 142 1001 176 1036
rect 142 933 176 951
rect 142 865 176 879
rect 142 797 176 807
rect 142 729 176 735
rect 142 661 176 663
rect 142 625 176 627
rect 142 553 176 559
rect 142 481 176 491
rect 142 409 176 423
rect 142 337 176 355
rect 142 265 176 287
rect 142 193 176 219
rect 142 121 176 151
rect 142 49 176 83
rect 142 -19 176 15
rect 142 -87 176 -57
rect 142 -155 176 -129
rect 142 -223 176 -201
rect 142 -291 176 -273
rect 142 -359 176 -345
rect 142 -427 176 -417
rect 142 -495 176 -489
rect 142 -563 176 -561
rect 142 -599 176 -597
rect 142 -671 176 -665
rect 142 -743 176 -733
rect 142 -815 176 -801
rect 142 -887 176 -869
rect 142 -972 176 -937
rect 300 1001 334 1036
rect 300 933 334 951
rect 300 865 334 879
rect 300 797 334 807
rect 300 729 334 735
rect 300 661 334 663
rect 300 625 334 627
rect 300 553 334 559
rect 300 481 334 491
rect 300 409 334 423
rect 300 337 334 355
rect 300 265 334 287
rect 300 193 334 219
rect 300 121 334 151
rect 300 49 334 83
rect 300 -19 334 15
rect 300 -87 334 -57
rect 300 -155 334 -129
rect 300 -223 334 -201
rect 300 -291 334 -273
rect 300 -359 334 -345
rect 300 -427 334 -417
rect 300 -495 334 -489
rect 300 -563 334 -561
rect 300 -599 334 -597
rect 300 -671 334 -665
rect 300 -743 334 -733
rect 300 -815 334 -801
rect 300 -887 334 -869
rect 300 -972 334 -937
rect 458 1001 492 1036
rect 458 933 492 951
rect 458 865 492 879
rect 458 797 492 807
rect 458 729 492 735
rect 458 661 492 663
rect 458 625 492 627
rect 458 553 492 559
rect 458 481 492 491
rect 458 409 492 423
rect 458 337 492 355
rect 458 265 492 287
rect 458 193 492 219
rect 458 121 492 151
rect 458 49 492 83
rect 458 -19 492 15
rect 458 -87 492 -57
rect 458 -155 492 -129
rect 458 -223 492 -201
rect 458 -291 492 -273
rect 458 -359 492 -345
rect 458 -427 492 -417
rect 458 -495 492 -489
rect 458 -563 492 -561
rect 458 -599 492 -597
rect 458 -671 492 -665
rect 458 -743 492 -733
rect 458 -815 492 -801
rect 458 -887 492 -869
rect 458 -972 492 -937
rect 616 1001 650 1036
rect 616 933 650 951
rect 616 865 650 879
rect 616 797 650 807
rect 616 729 650 735
rect 616 661 650 663
rect 616 625 650 627
rect 616 553 650 559
rect 616 481 650 491
rect 616 409 650 423
rect 616 337 650 355
rect 616 265 650 287
rect 616 193 650 219
rect 616 121 650 151
rect 616 49 650 83
rect 616 -19 650 15
rect 616 -87 650 -57
rect 616 -155 650 -129
rect 616 -223 650 -201
rect 616 -291 650 -273
rect 616 -359 650 -345
rect 616 -427 650 -417
rect 616 -495 650 -489
rect 616 -563 650 -561
rect 616 -599 650 -597
rect 616 -671 650 -665
rect 616 -743 650 -733
rect 616 -815 650 -801
rect 616 -887 650 -869
rect 616 -972 650 -937
rect 774 1001 808 1036
rect 774 933 808 951
rect 774 865 808 879
rect 774 797 808 807
rect 774 729 808 735
rect 774 661 808 663
rect 774 625 808 627
rect 774 553 808 559
rect 774 481 808 491
rect 774 409 808 423
rect 774 337 808 355
rect 774 265 808 287
rect 774 193 808 219
rect 774 121 808 151
rect 774 49 808 83
rect 774 -19 808 15
rect 774 -87 808 -57
rect 774 -155 808 -129
rect 774 -223 808 -201
rect 774 -291 808 -273
rect 774 -359 808 -345
rect 774 -427 808 -417
rect 774 -495 808 -489
rect 774 -563 808 -561
rect 774 -599 808 -597
rect 774 -671 808 -665
rect 774 -743 808 -733
rect 774 -815 808 -801
rect 774 -887 808 -869
rect 774 -972 808 -937
rect -760 -1040 -736 -1006
rect -702 -1040 -678 -1006
<< viali >>
rect -806 967 -772 985
rect -806 951 -772 967
rect -806 899 -772 913
rect -806 879 -772 899
rect -806 831 -772 841
rect -806 807 -772 831
rect -806 763 -772 769
rect -806 735 -772 763
rect -806 695 -772 697
rect -806 663 -772 695
rect -806 593 -772 625
rect -806 591 -772 593
rect -806 525 -772 553
rect -806 519 -772 525
rect -806 457 -772 481
rect -806 447 -772 457
rect -806 389 -772 409
rect -806 375 -772 389
rect -806 321 -772 337
rect -806 303 -772 321
rect -806 253 -772 265
rect -806 231 -772 253
rect -806 185 -772 193
rect -806 159 -772 185
rect -806 117 -772 121
rect -806 87 -772 117
rect -806 15 -772 49
rect -806 -53 -772 -23
rect -806 -57 -772 -53
rect -806 -121 -772 -95
rect -806 -129 -772 -121
rect -806 -189 -772 -167
rect -806 -201 -772 -189
rect -806 -257 -772 -239
rect -806 -273 -772 -257
rect -806 -325 -772 -311
rect -806 -345 -772 -325
rect -806 -393 -772 -383
rect -806 -417 -772 -393
rect -806 -461 -772 -455
rect -806 -489 -772 -461
rect -806 -529 -772 -527
rect -806 -561 -772 -529
rect -806 -631 -772 -599
rect -806 -633 -772 -631
rect -806 -699 -772 -671
rect -806 -705 -772 -699
rect -806 -767 -772 -743
rect -806 -777 -772 -767
rect -806 -835 -772 -815
rect -806 -849 -772 -835
rect -806 -903 -772 -887
rect -806 -921 -772 -903
rect -648 967 -614 985
rect -648 951 -614 967
rect -648 899 -614 913
rect -648 879 -614 899
rect -648 831 -614 841
rect -648 807 -614 831
rect -648 763 -614 769
rect -648 735 -614 763
rect -648 695 -614 697
rect -648 663 -614 695
rect -648 593 -614 625
rect -648 591 -614 593
rect -648 525 -614 553
rect -648 519 -614 525
rect -648 457 -614 481
rect -648 447 -614 457
rect -648 389 -614 409
rect -648 375 -614 389
rect -648 321 -614 337
rect -648 303 -614 321
rect -648 253 -614 265
rect -648 231 -614 253
rect -648 185 -614 193
rect -648 159 -614 185
rect -648 117 -614 121
rect -648 87 -614 117
rect -648 15 -614 49
rect -648 -53 -614 -23
rect -648 -57 -614 -53
rect -648 -121 -614 -95
rect -648 -129 -614 -121
rect -648 -189 -614 -167
rect -648 -201 -614 -189
rect -648 -257 -614 -239
rect -648 -273 -614 -257
rect -648 -325 -614 -311
rect -648 -345 -614 -325
rect -648 -393 -614 -383
rect -648 -417 -614 -393
rect -648 -461 -614 -455
rect -648 -489 -614 -461
rect -648 -529 -614 -527
rect -648 -561 -614 -529
rect -648 -631 -614 -599
rect -648 -633 -614 -631
rect -648 -699 -614 -671
rect -648 -705 -614 -699
rect -648 -767 -614 -743
rect -648 -777 -614 -767
rect -648 -835 -614 -815
rect -648 -849 -614 -835
rect -648 -903 -614 -887
rect -648 -921 -614 -903
rect -490 967 -456 985
rect -490 951 -456 967
rect -490 899 -456 913
rect -490 879 -456 899
rect -490 831 -456 841
rect -490 807 -456 831
rect -490 763 -456 769
rect -490 735 -456 763
rect -490 695 -456 697
rect -490 663 -456 695
rect -490 593 -456 625
rect -490 591 -456 593
rect -490 525 -456 553
rect -490 519 -456 525
rect -490 457 -456 481
rect -490 447 -456 457
rect -490 389 -456 409
rect -490 375 -456 389
rect -490 321 -456 337
rect -490 303 -456 321
rect -490 253 -456 265
rect -490 231 -456 253
rect -490 185 -456 193
rect -490 159 -456 185
rect -490 117 -456 121
rect -490 87 -456 117
rect -490 15 -456 49
rect -490 -53 -456 -23
rect -490 -57 -456 -53
rect -490 -121 -456 -95
rect -490 -129 -456 -121
rect -490 -189 -456 -167
rect -490 -201 -456 -189
rect -490 -257 -456 -239
rect -490 -273 -456 -257
rect -490 -325 -456 -311
rect -490 -345 -456 -325
rect -490 -393 -456 -383
rect -490 -417 -456 -393
rect -490 -461 -456 -455
rect -490 -489 -456 -461
rect -490 -529 -456 -527
rect -490 -561 -456 -529
rect -490 -631 -456 -599
rect -490 -633 -456 -631
rect -490 -699 -456 -671
rect -490 -705 -456 -699
rect -490 -767 -456 -743
rect -490 -777 -456 -767
rect -490 -835 -456 -815
rect -490 -849 -456 -835
rect -490 -903 -456 -887
rect -490 -921 -456 -903
rect -332 967 -298 985
rect -332 951 -298 967
rect -332 899 -298 913
rect -332 879 -298 899
rect -332 831 -298 841
rect -332 807 -298 831
rect -332 763 -298 769
rect -332 735 -298 763
rect -332 695 -298 697
rect -332 663 -298 695
rect -332 593 -298 625
rect -332 591 -298 593
rect -332 525 -298 553
rect -332 519 -298 525
rect -332 457 -298 481
rect -332 447 -298 457
rect -332 389 -298 409
rect -332 375 -298 389
rect -332 321 -298 337
rect -332 303 -298 321
rect -332 253 -298 265
rect -332 231 -298 253
rect -332 185 -298 193
rect -332 159 -298 185
rect -332 117 -298 121
rect -332 87 -298 117
rect -332 15 -298 49
rect -332 -53 -298 -23
rect -332 -57 -298 -53
rect -332 -121 -298 -95
rect -332 -129 -298 -121
rect -332 -189 -298 -167
rect -332 -201 -298 -189
rect -332 -257 -298 -239
rect -332 -273 -298 -257
rect -332 -325 -298 -311
rect -332 -345 -298 -325
rect -332 -393 -298 -383
rect -332 -417 -298 -393
rect -332 -461 -298 -455
rect -332 -489 -298 -461
rect -332 -529 -298 -527
rect -332 -561 -298 -529
rect -332 -631 -298 -599
rect -332 -633 -298 -631
rect -332 -699 -298 -671
rect -332 -705 -298 -699
rect -332 -767 -298 -743
rect -332 -777 -298 -767
rect -332 -835 -298 -815
rect -332 -849 -298 -835
rect -332 -903 -298 -887
rect -332 -921 -298 -903
rect -174 967 -140 985
rect -174 951 -140 967
rect -174 899 -140 913
rect -174 879 -140 899
rect -174 831 -140 841
rect -174 807 -140 831
rect -174 763 -140 769
rect -174 735 -140 763
rect -174 695 -140 697
rect -174 663 -140 695
rect -174 593 -140 625
rect -174 591 -140 593
rect -174 525 -140 553
rect -174 519 -140 525
rect -174 457 -140 481
rect -174 447 -140 457
rect -174 389 -140 409
rect -174 375 -140 389
rect -174 321 -140 337
rect -174 303 -140 321
rect -174 253 -140 265
rect -174 231 -140 253
rect -174 185 -140 193
rect -174 159 -140 185
rect -174 117 -140 121
rect -174 87 -140 117
rect -174 15 -140 49
rect -174 -53 -140 -23
rect -174 -57 -140 -53
rect -174 -121 -140 -95
rect -174 -129 -140 -121
rect -174 -189 -140 -167
rect -174 -201 -140 -189
rect -174 -257 -140 -239
rect -174 -273 -140 -257
rect -174 -325 -140 -311
rect -174 -345 -140 -325
rect -174 -393 -140 -383
rect -174 -417 -140 -393
rect -174 -461 -140 -455
rect -174 -489 -140 -461
rect -174 -529 -140 -527
rect -174 -561 -140 -529
rect -174 -631 -140 -599
rect -174 -633 -140 -631
rect -174 -699 -140 -671
rect -174 -705 -140 -699
rect -174 -767 -140 -743
rect -174 -777 -140 -767
rect -174 -835 -140 -815
rect -174 -849 -140 -835
rect -174 -903 -140 -887
rect -174 -921 -140 -903
rect -16 967 18 985
rect -16 951 18 967
rect -16 899 18 913
rect -16 879 18 899
rect -16 831 18 841
rect -16 807 18 831
rect -16 763 18 769
rect -16 735 18 763
rect -16 695 18 697
rect -16 663 18 695
rect -16 593 18 625
rect -16 591 18 593
rect -16 525 18 553
rect -16 519 18 525
rect -16 457 18 481
rect -16 447 18 457
rect -16 389 18 409
rect -16 375 18 389
rect -16 321 18 337
rect -16 303 18 321
rect -16 253 18 265
rect -16 231 18 253
rect -16 185 18 193
rect -16 159 18 185
rect -16 117 18 121
rect -16 87 18 117
rect -16 15 18 49
rect -16 -53 18 -23
rect -16 -57 18 -53
rect -16 -121 18 -95
rect -16 -129 18 -121
rect -16 -189 18 -167
rect -16 -201 18 -189
rect -16 -257 18 -239
rect -16 -273 18 -257
rect -16 -325 18 -311
rect -16 -345 18 -325
rect -16 -393 18 -383
rect -16 -417 18 -393
rect -16 -461 18 -455
rect -16 -489 18 -461
rect -16 -529 18 -527
rect -16 -561 18 -529
rect -16 -631 18 -599
rect -16 -633 18 -631
rect -16 -699 18 -671
rect -16 -705 18 -699
rect -16 -767 18 -743
rect -16 -777 18 -767
rect -16 -835 18 -815
rect -16 -849 18 -835
rect -16 -903 18 -887
rect -16 -921 18 -903
rect 142 967 176 985
rect 142 951 176 967
rect 142 899 176 913
rect 142 879 176 899
rect 142 831 176 841
rect 142 807 176 831
rect 142 763 176 769
rect 142 735 176 763
rect 142 695 176 697
rect 142 663 176 695
rect 142 593 176 625
rect 142 591 176 593
rect 142 525 176 553
rect 142 519 176 525
rect 142 457 176 481
rect 142 447 176 457
rect 142 389 176 409
rect 142 375 176 389
rect 142 321 176 337
rect 142 303 176 321
rect 142 253 176 265
rect 142 231 176 253
rect 142 185 176 193
rect 142 159 176 185
rect 142 117 176 121
rect 142 87 176 117
rect 142 15 176 49
rect 142 -53 176 -23
rect 142 -57 176 -53
rect 142 -121 176 -95
rect 142 -129 176 -121
rect 142 -189 176 -167
rect 142 -201 176 -189
rect 142 -257 176 -239
rect 142 -273 176 -257
rect 142 -325 176 -311
rect 142 -345 176 -325
rect 142 -393 176 -383
rect 142 -417 176 -393
rect 142 -461 176 -455
rect 142 -489 176 -461
rect 142 -529 176 -527
rect 142 -561 176 -529
rect 142 -631 176 -599
rect 142 -633 176 -631
rect 142 -699 176 -671
rect 142 -705 176 -699
rect 142 -767 176 -743
rect 142 -777 176 -767
rect 142 -835 176 -815
rect 142 -849 176 -835
rect 142 -903 176 -887
rect 142 -921 176 -903
rect 300 967 334 985
rect 300 951 334 967
rect 300 899 334 913
rect 300 879 334 899
rect 300 831 334 841
rect 300 807 334 831
rect 300 763 334 769
rect 300 735 334 763
rect 300 695 334 697
rect 300 663 334 695
rect 300 593 334 625
rect 300 591 334 593
rect 300 525 334 553
rect 300 519 334 525
rect 300 457 334 481
rect 300 447 334 457
rect 300 389 334 409
rect 300 375 334 389
rect 300 321 334 337
rect 300 303 334 321
rect 300 253 334 265
rect 300 231 334 253
rect 300 185 334 193
rect 300 159 334 185
rect 300 117 334 121
rect 300 87 334 117
rect 300 15 334 49
rect 300 -53 334 -23
rect 300 -57 334 -53
rect 300 -121 334 -95
rect 300 -129 334 -121
rect 300 -189 334 -167
rect 300 -201 334 -189
rect 300 -257 334 -239
rect 300 -273 334 -257
rect 300 -325 334 -311
rect 300 -345 334 -325
rect 300 -393 334 -383
rect 300 -417 334 -393
rect 300 -461 334 -455
rect 300 -489 334 -461
rect 300 -529 334 -527
rect 300 -561 334 -529
rect 300 -631 334 -599
rect 300 -633 334 -631
rect 300 -699 334 -671
rect 300 -705 334 -699
rect 300 -767 334 -743
rect 300 -777 334 -767
rect 300 -835 334 -815
rect 300 -849 334 -835
rect 300 -903 334 -887
rect 300 -921 334 -903
rect 458 967 492 985
rect 458 951 492 967
rect 458 899 492 913
rect 458 879 492 899
rect 458 831 492 841
rect 458 807 492 831
rect 458 763 492 769
rect 458 735 492 763
rect 458 695 492 697
rect 458 663 492 695
rect 458 593 492 625
rect 458 591 492 593
rect 458 525 492 553
rect 458 519 492 525
rect 458 457 492 481
rect 458 447 492 457
rect 458 389 492 409
rect 458 375 492 389
rect 458 321 492 337
rect 458 303 492 321
rect 458 253 492 265
rect 458 231 492 253
rect 458 185 492 193
rect 458 159 492 185
rect 458 117 492 121
rect 458 87 492 117
rect 458 15 492 49
rect 458 -53 492 -23
rect 458 -57 492 -53
rect 458 -121 492 -95
rect 458 -129 492 -121
rect 458 -189 492 -167
rect 458 -201 492 -189
rect 458 -257 492 -239
rect 458 -273 492 -257
rect 458 -325 492 -311
rect 458 -345 492 -325
rect 458 -393 492 -383
rect 458 -417 492 -393
rect 458 -461 492 -455
rect 458 -489 492 -461
rect 458 -529 492 -527
rect 458 -561 492 -529
rect 458 -631 492 -599
rect 458 -633 492 -631
rect 458 -699 492 -671
rect 458 -705 492 -699
rect 458 -767 492 -743
rect 458 -777 492 -767
rect 458 -835 492 -815
rect 458 -849 492 -835
rect 458 -903 492 -887
rect 458 -921 492 -903
rect 616 967 650 985
rect 616 951 650 967
rect 616 899 650 913
rect 616 879 650 899
rect 616 831 650 841
rect 616 807 650 831
rect 616 763 650 769
rect 616 735 650 763
rect 616 695 650 697
rect 616 663 650 695
rect 616 593 650 625
rect 616 591 650 593
rect 616 525 650 553
rect 616 519 650 525
rect 616 457 650 481
rect 616 447 650 457
rect 616 389 650 409
rect 616 375 650 389
rect 616 321 650 337
rect 616 303 650 321
rect 616 253 650 265
rect 616 231 650 253
rect 616 185 650 193
rect 616 159 650 185
rect 616 117 650 121
rect 616 87 650 117
rect 616 15 650 49
rect 616 -53 650 -23
rect 616 -57 650 -53
rect 616 -121 650 -95
rect 616 -129 650 -121
rect 616 -189 650 -167
rect 616 -201 650 -189
rect 616 -257 650 -239
rect 616 -273 650 -257
rect 616 -325 650 -311
rect 616 -345 650 -325
rect 616 -393 650 -383
rect 616 -417 650 -393
rect 616 -461 650 -455
rect 616 -489 650 -461
rect 616 -529 650 -527
rect 616 -561 650 -529
rect 616 -631 650 -599
rect 616 -633 650 -631
rect 616 -699 650 -671
rect 616 -705 650 -699
rect 616 -767 650 -743
rect 616 -777 650 -767
rect 616 -835 650 -815
rect 616 -849 650 -835
rect 616 -903 650 -887
rect 616 -921 650 -903
rect 774 967 808 985
rect 774 951 808 967
rect 774 899 808 913
rect 774 879 808 899
rect 774 831 808 841
rect 774 807 808 831
rect 774 763 808 769
rect 774 735 808 763
rect 774 695 808 697
rect 774 663 808 695
rect 774 593 808 625
rect 774 591 808 593
rect 774 525 808 553
rect 774 519 808 525
rect 774 457 808 481
rect 774 447 808 457
rect 774 389 808 409
rect 774 375 808 389
rect 774 321 808 337
rect 774 303 808 321
rect 774 253 808 265
rect 774 231 808 253
rect 774 185 808 193
rect 774 159 808 185
rect 774 117 808 121
rect 774 87 808 117
rect 774 15 808 49
rect 774 -53 808 -23
rect 774 -57 808 -53
rect 774 -121 808 -95
rect 774 -129 808 -121
rect 774 -189 808 -167
rect 774 -201 808 -189
rect 774 -257 808 -239
rect 774 -273 808 -257
rect 774 -325 808 -311
rect 774 -345 808 -325
rect 774 -393 808 -383
rect 774 -417 808 -393
rect 774 -461 808 -455
rect 774 -489 808 -461
rect 774 -529 808 -527
rect 774 -561 808 -529
rect 774 -631 808 -599
rect 774 -633 808 -631
rect 774 -699 808 -671
rect 774 -705 808 -699
rect 774 -767 808 -743
rect 774 -777 808 -767
rect 774 -835 808 -815
rect 774 -849 808 -835
rect 774 -903 808 -887
rect 774 -921 808 -903
rect -736 -1040 -702 -1006
<< metal1 >>
rect -22 1160 24 1186
rect -812 1114 814 1160
rect -812 985 -766 1114
rect -812 951 -806 985
rect -772 951 -766 985
rect -812 913 -766 951
rect -812 879 -806 913
rect -772 879 -766 913
rect -812 841 -766 879
rect -812 807 -806 841
rect -772 807 -766 841
rect -812 769 -766 807
rect -812 735 -806 769
rect -772 735 -766 769
rect -812 697 -766 735
rect -812 663 -806 697
rect -772 663 -766 697
rect -812 625 -766 663
rect -812 591 -806 625
rect -772 591 -766 625
rect -812 553 -766 591
rect -812 519 -806 553
rect -772 519 -766 553
rect -812 481 -766 519
rect -812 447 -806 481
rect -772 447 -766 481
rect -812 409 -766 447
rect -812 375 -806 409
rect -772 375 -766 409
rect -812 337 -766 375
rect -812 303 -806 337
rect -772 303 -766 337
rect -812 265 -766 303
rect -812 231 -806 265
rect -772 231 -766 265
rect -812 193 -766 231
rect -812 159 -806 193
rect -772 159 -766 193
rect -812 121 -766 159
rect -812 87 -806 121
rect -772 87 -766 121
rect -812 49 -766 87
rect -812 15 -806 49
rect -772 15 -766 49
rect -812 -23 -766 15
rect -812 -57 -806 -23
rect -772 -57 -766 -23
rect -812 -95 -766 -57
rect -812 -129 -806 -95
rect -772 -129 -766 -95
rect -812 -167 -766 -129
rect -812 -201 -806 -167
rect -772 -201 -766 -167
rect -812 -239 -766 -201
rect -812 -273 -806 -239
rect -772 -273 -766 -239
rect -812 -311 -766 -273
rect -812 -345 -806 -311
rect -772 -345 -766 -311
rect -812 -383 -766 -345
rect -812 -417 -806 -383
rect -772 -417 -766 -383
rect -812 -455 -766 -417
rect -812 -489 -806 -455
rect -772 -489 -766 -455
rect -812 -527 -766 -489
rect -812 -561 -806 -527
rect -772 -561 -766 -527
rect -812 -599 -766 -561
rect -812 -633 -806 -599
rect -772 -633 -766 -599
rect -812 -671 -766 -633
rect -812 -705 -806 -671
rect -772 -705 -766 -671
rect -812 -743 -766 -705
rect -812 -777 -806 -743
rect -772 -777 -766 -743
rect -812 -815 -766 -777
rect -812 -849 -806 -815
rect -772 -849 -766 -815
rect -812 -887 -766 -849
rect -812 -921 -806 -887
rect -772 -921 -766 -887
rect -812 -968 -766 -921
rect -654 985 -608 1032
rect -654 951 -648 985
rect -614 951 -608 985
rect -654 913 -608 951
rect -654 879 -648 913
rect -614 879 -608 913
rect -654 841 -608 879
rect -654 807 -648 841
rect -614 807 -608 841
rect -654 769 -608 807
rect -654 735 -648 769
rect -614 735 -608 769
rect -654 697 -608 735
rect -654 663 -648 697
rect -614 663 -608 697
rect -654 625 -608 663
rect -654 591 -648 625
rect -614 591 -608 625
rect -654 553 -608 591
rect -654 519 -648 553
rect -614 519 -608 553
rect -654 481 -608 519
rect -654 447 -648 481
rect -614 447 -608 481
rect -654 409 -608 447
rect -654 375 -648 409
rect -614 375 -608 409
rect -654 337 -608 375
rect -654 303 -648 337
rect -614 303 -608 337
rect -654 265 -608 303
rect -654 231 -648 265
rect -614 231 -608 265
rect -654 193 -608 231
rect -654 159 -648 193
rect -614 159 -608 193
rect -654 121 -608 159
rect -654 87 -648 121
rect -614 87 -608 121
rect -654 49 -608 87
rect -654 15 -648 49
rect -614 15 -608 49
rect -654 -23 -608 15
rect -654 -57 -648 -23
rect -614 -57 -608 -23
rect -654 -95 -608 -57
rect -654 -129 -648 -95
rect -614 -129 -608 -95
rect -654 -167 -608 -129
rect -654 -201 -648 -167
rect -614 -201 -608 -167
rect -654 -239 -608 -201
rect -654 -273 -648 -239
rect -614 -273 -608 -239
rect -654 -311 -608 -273
rect -654 -345 -648 -311
rect -614 -345 -608 -311
rect -654 -383 -608 -345
rect -654 -417 -648 -383
rect -614 -417 -608 -383
rect -654 -455 -608 -417
rect -654 -489 -648 -455
rect -614 -489 -608 -455
rect -654 -527 -608 -489
rect -654 -561 -648 -527
rect -614 -561 -608 -527
rect -654 -599 -608 -561
rect -654 -633 -648 -599
rect -614 -633 -608 -599
rect -654 -671 -608 -633
rect -654 -705 -648 -671
rect -614 -705 -608 -671
rect -654 -743 -608 -705
rect -654 -777 -648 -743
rect -614 -777 -608 -743
rect -654 -815 -608 -777
rect -654 -849 -648 -815
rect -614 -849 -608 -815
rect -654 -887 -608 -849
rect -654 -921 -648 -887
rect -614 -921 -608 -887
rect -756 -1006 -682 -1000
rect -756 -1040 -736 -1006
rect -702 -1040 -682 -1006
rect -756 -1046 -682 -1040
rect -654 -1062 -608 -921
rect -496 985 -450 1114
rect -496 951 -490 985
rect -456 951 -450 985
rect -496 913 -450 951
rect -496 879 -490 913
rect -456 879 -450 913
rect -496 841 -450 879
rect -496 807 -490 841
rect -456 807 -450 841
rect -496 769 -450 807
rect -496 735 -490 769
rect -456 735 -450 769
rect -496 697 -450 735
rect -496 663 -490 697
rect -456 663 -450 697
rect -496 625 -450 663
rect -496 591 -490 625
rect -456 591 -450 625
rect -496 553 -450 591
rect -496 519 -490 553
rect -456 519 -450 553
rect -496 481 -450 519
rect -496 447 -490 481
rect -456 447 -450 481
rect -496 409 -450 447
rect -496 375 -490 409
rect -456 375 -450 409
rect -496 337 -450 375
rect -496 303 -490 337
rect -456 303 -450 337
rect -496 265 -450 303
rect -496 231 -490 265
rect -456 231 -450 265
rect -496 193 -450 231
rect -496 159 -490 193
rect -456 159 -450 193
rect -496 121 -450 159
rect -496 87 -490 121
rect -456 87 -450 121
rect -496 49 -450 87
rect -496 15 -490 49
rect -456 15 -450 49
rect -496 -23 -450 15
rect -496 -57 -490 -23
rect -456 -57 -450 -23
rect -496 -95 -450 -57
rect -496 -129 -490 -95
rect -456 -129 -450 -95
rect -496 -167 -450 -129
rect -496 -201 -490 -167
rect -456 -201 -450 -167
rect -496 -239 -450 -201
rect -496 -273 -490 -239
rect -456 -273 -450 -239
rect -496 -311 -450 -273
rect -496 -345 -490 -311
rect -456 -345 -450 -311
rect -496 -383 -450 -345
rect -496 -417 -490 -383
rect -456 -417 -450 -383
rect -496 -455 -450 -417
rect -496 -489 -490 -455
rect -456 -489 -450 -455
rect -496 -527 -450 -489
rect -496 -561 -490 -527
rect -456 -561 -450 -527
rect -496 -599 -450 -561
rect -496 -633 -490 -599
rect -456 -633 -450 -599
rect -496 -671 -450 -633
rect -496 -705 -490 -671
rect -456 -705 -450 -671
rect -496 -743 -450 -705
rect -496 -777 -490 -743
rect -456 -777 -450 -743
rect -496 -815 -450 -777
rect -496 -849 -490 -815
rect -456 -849 -450 -815
rect -496 -887 -450 -849
rect -496 -921 -490 -887
rect -456 -921 -450 -887
rect -496 -968 -450 -921
rect -338 985 -292 1032
rect -338 951 -332 985
rect -298 951 -292 985
rect -338 913 -292 951
rect -338 879 -332 913
rect -298 879 -292 913
rect -338 841 -292 879
rect -338 807 -332 841
rect -298 807 -292 841
rect -338 769 -292 807
rect -338 735 -332 769
rect -298 735 -292 769
rect -338 697 -292 735
rect -338 663 -332 697
rect -298 663 -292 697
rect -338 625 -292 663
rect -338 591 -332 625
rect -298 591 -292 625
rect -338 553 -292 591
rect -338 519 -332 553
rect -298 519 -292 553
rect -338 481 -292 519
rect -338 447 -332 481
rect -298 447 -292 481
rect -338 409 -292 447
rect -338 375 -332 409
rect -298 375 -292 409
rect -338 337 -292 375
rect -338 303 -332 337
rect -298 303 -292 337
rect -338 265 -292 303
rect -338 231 -332 265
rect -298 231 -292 265
rect -338 193 -292 231
rect -338 159 -332 193
rect -298 159 -292 193
rect -338 121 -292 159
rect -338 87 -332 121
rect -298 87 -292 121
rect -338 49 -292 87
rect -338 15 -332 49
rect -298 15 -292 49
rect -338 -23 -292 15
rect -338 -57 -332 -23
rect -298 -57 -292 -23
rect -338 -95 -292 -57
rect -338 -129 -332 -95
rect -298 -129 -292 -95
rect -338 -167 -292 -129
rect -338 -201 -332 -167
rect -298 -201 -292 -167
rect -338 -239 -292 -201
rect -338 -273 -332 -239
rect -298 -273 -292 -239
rect -338 -311 -292 -273
rect -338 -345 -332 -311
rect -298 -345 -292 -311
rect -338 -383 -292 -345
rect -338 -417 -332 -383
rect -298 -417 -292 -383
rect -338 -455 -292 -417
rect -338 -489 -332 -455
rect -298 -489 -292 -455
rect -338 -527 -292 -489
rect -338 -561 -332 -527
rect -298 -561 -292 -527
rect -338 -599 -292 -561
rect -338 -633 -332 -599
rect -298 -633 -292 -599
rect -338 -671 -292 -633
rect -338 -705 -332 -671
rect -298 -705 -292 -671
rect -338 -743 -292 -705
rect -338 -777 -332 -743
rect -298 -777 -292 -743
rect -338 -815 -292 -777
rect -338 -849 -332 -815
rect -298 -849 -292 -815
rect -338 -887 -292 -849
rect -338 -921 -332 -887
rect -298 -921 -292 -887
rect -338 -1062 -292 -921
rect -180 985 -134 1114
rect -180 951 -174 985
rect -140 951 -134 985
rect -180 913 -134 951
rect -180 879 -174 913
rect -140 879 -134 913
rect -180 841 -134 879
rect -180 807 -174 841
rect -140 807 -134 841
rect -180 769 -134 807
rect -180 735 -174 769
rect -140 735 -134 769
rect -180 697 -134 735
rect -180 663 -174 697
rect -140 663 -134 697
rect -180 625 -134 663
rect -180 591 -174 625
rect -140 591 -134 625
rect -180 553 -134 591
rect -180 519 -174 553
rect -140 519 -134 553
rect -180 481 -134 519
rect -180 447 -174 481
rect -140 447 -134 481
rect -180 409 -134 447
rect -180 375 -174 409
rect -140 375 -134 409
rect -180 337 -134 375
rect -180 303 -174 337
rect -140 303 -134 337
rect -180 265 -134 303
rect -180 231 -174 265
rect -140 231 -134 265
rect -180 193 -134 231
rect -180 159 -174 193
rect -140 159 -134 193
rect -180 121 -134 159
rect -180 87 -174 121
rect -140 87 -134 121
rect -180 49 -134 87
rect -180 15 -174 49
rect -140 15 -134 49
rect -180 -23 -134 15
rect -180 -57 -174 -23
rect -140 -57 -134 -23
rect -180 -95 -134 -57
rect -180 -129 -174 -95
rect -140 -129 -134 -95
rect -180 -167 -134 -129
rect -180 -201 -174 -167
rect -140 -201 -134 -167
rect -180 -239 -134 -201
rect -180 -273 -174 -239
rect -140 -273 -134 -239
rect -180 -311 -134 -273
rect -180 -345 -174 -311
rect -140 -345 -134 -311
rect -180 -383 -134 -345
rect -180 -417 -174 -383
rect -140 -417 -134 -383
rect -180 -455 -134 -417
rect -180 -489 -174 -455
rect -140 -489 -134 -455
rect -180 -527 -134 -489
rect -180 -561 -174 -527
rect -140 -561 -134 -527
rect -180 -599 -134 -561
rect -180 -633 -174 -599
rect -140 -633 -134 -599
rect -180 -671 -134 -633
rect -180 -705 -174 -671
rect -140 -705 -134 -671
rect -180 -743 -134 -705
rect -180 -777 -174 -743
rect -140 -777 -134 -743
rect -180 -815 -134 -777
rect -180 -849 -174 -815
rect -140 -849 -134 -815
rect -180 -887 -134 -849
rect -180 -921 -174 -887
rect -140 -921 -134 -887
rect -180 -968 -134 -921
rect -22 985 24 1032
rect -22 951 -16 985
rect 18 951 24 985
rect -22 913 24 951
rect -22 879 -16 913
rect 18 879 24 913
rect -22 841 24 879
rect -22 807 -16 841
rect 18 807 24 841
rect -22 769 24 807
rect -22 735 -16 769
rect 18 735 24 769
rect -22 697 24 735
rect -22 663 -16 697
rect 18 663 24 697
rect -22 625 24 663
rect -22 591 -16 625
rect 18 591 24 625
rect -22 553 24 591
rect -22 519 -16 553
rect 18 519 24 553
rect -22 481 24 519
rect -22 447 -16 481
rect 18 447 24 481
rect -22 409 24 447
rect -22 375 -16 409
rect 18 375 24 409
rect -22 337 24 375
rect -22 303 -16 337
rect 18 303 24 337
rect -22 265 24 303
rect -22 231 -16 265
rect 18 231 24 265
rect -22 193 24 231
rect -22 159 -16 193
rect 18 159 24 193
rect -22 121 24 159
rect -22 87 -16 121
rect 18 87 24 121
rect -22 49 24 87
rect -22 15 -16 49
rect 18 15 24 49
rect -22 -23 24 15
rect -22 -57 -16 -23
rect 18 -57 24 -23
rect -22 -95 24 -57
rect -22 -129 -16 -95
rect 18 -129 24 -95
rect -22 -167 24 -129
rect -22 -201 -16 -167
rect 18 -201 24 -167
rect -22 -239 24 -201
rect -22 -273 -16 -239
rect 18 -273 24 -239
rect -22 -311 24 -273
rect -22 -345 -16 -311
rect 18 -345 24 -311
rect -22 -383 24 -345
rect -22 -417 -16 -383
rect 18 -417 24 -383
rect -22 -455 24 -417
rect -22 -489 -16 -455
rect 18 -489 24 -455
rect -22 -527 24 -489
rect -22 -561 -16 -527
rect 18 -561 24 -527
rect -22 -599 24 -561
rect -22 -633 -16 -599
rect 18 -633 24 -599
rect -22 -671 24 -633
rect -22 -705 -16 -671
rect 18 -705 24 -671
rect -22 -743 24 -705
rect -22 -777 -16 -743
rect 18 -777 24 -743
rect -22 -815 24 -777
rect -22 -849 -16 -815
rect 18 -849 24 -815
rect -22 -887 24 -849
rect -22 -921 -16 -887
rect 18 -921 24 -887
rect -22 -1062 24 -921
rect 136 985 182 1114
rect 136 951 142 985
rect 176 951 182 985
rect 136 913 182 951
rect 136 879 142 913
rect 176 879 182 913
rect 136 841 182 879
rect 136 807 142 841
rect 176 807 182 841
rect 136 769 182 807
rect 136 735 142 769
rect 176 735 182 769
rect 136 697 182 735
rect 136 663 142 697
rect 176 663 182 697
rect 136 625 182 663
rect 136 591 142 625
rect 176 591 182 625
rect 136 553 182 591
rect 136 519 142 553
rect 176 519 182 553
rect 136 481 182 519
rect 136 447 142 481
rect 176 447 182 481
rect 136 409 182 447
rect 136 375 142 409
rect 176 375 182 409
rect 136 337 182 375
rect 136 303 142 337
rect 176 303 182 337
rect 136 265 182 303
rect 136 231 142 265
rect 176 231 182 265
rect 136 193 182 231
rect 136 159 142 193
rect 176 159 182 193
rect 136 121 182 159
rect 136 87 142 121
rect 176 87 182 121
rect 136 49 182 87
rect 136 15 142 49
rect 176 15 182 49
rect 136 -23 182 15
rect 136 -57 142 -23
rect 176 -57 182 -23
rect 136 -95 182 -57
rect 136 -129 142 -95
rect 176 -129 182 -95
rect 136 -167 182 -129
rect 136 -201 142 -167
rect 176 -201 182 -167
rect 136 -239 182 -201
rect 136 -273 142 -239
rect 176 -273 182 -239
rect 136 -311 182 -273
rect 136 -345 142 -311
rect 176 -345 182 -311
rect 136 -383 182 -345
rect 136 -417 142 -383
rect 176 -417 182 -383
rect 136 -455 182 -417
rect 136 -489 142 -455
rect 176 -489 182 -455
rect 136 -527 182 -489
rect 136 -561 142 -527
rect 176 -561 182 -527
rect 136 -599 182 -561
rect 136 -633 142 -599
rect 176 -633 182 -599
rect 136 -671 182 -633
rect 136 -705 142 -671
rect 176 -705 182 -671
rect 136 -743 182 -705
rect 136 -777 142 -743
rect 176 -777 182 -743
rect 136 -815 182 -777
rect 136 -849 142 -815
rect 176 -849 182 -815
rect 136 -887 182 -849
rect 136 -921 142 -887
rect 176 -921 182 -887
rect 136 -968 182 -921
rect 294 985 340 1032
rect 294 951 300 985
rect 334 951 340 985
rect 294 913 340 951
rect 294 879 300 913
rect 334 879 340 913
rect 294 841 340 879
rect 294 807 300 841
rect 334 807 340 841
rect 294 769 340 807
rect 294 735 300 769
rect 334 735 340 769
rect 294 697 340 735
rect 294 663 300 697
rect 334 663 340 697
rect 294 625 340 663
rect 294 591 300 625
rect 334 591 340 625
rect 294 553 340 591
rect 294 519 300 553
rect 334 519 340 553
rect 294 481 340 519
rect 294 447 300 481
rect 334 447 340 481
rect 294 409 340 447
rect 294 375 300 409
rect 334 375 340 409
rect 294 337 340 375
rect 294 303 300 337
rect 334 303 340 337
rect 294 265 340 303
rect 294 231 300 265
rect 334 231 340 265
rect 294 193 340 231
rect 294 159 300 193
rect 334 159 340 193
rect 294 121 340 159
rect 294 87 300 121
rect 334 87 340 121
rect 294 49 340 87
rect 294 15 300 49
rect 334 15 340 49
rect 294 -23 340 15
rect 294 -57 300 -23
rect 334 -57 340 -23
rect 294 -95 340 -57
rect 294 -129 300 -95
rect 334 -129 340 -95
rect 294 -167 340 -129
rect 294 -201 300 -167
rect 334 -201 340 -167
rect 294 -239 340 -201
rect 294 -273 300 -239
rect 334 -273 340 -239
rect 294 -311 340 -273
rect 294 -345 300 -311
rect 334 -345 340 -311
rect 294 -383 340 -345
rect 294 -417 300 -383
rect 334 -417 340 -383
rect 294 -455 340 -417
rect 294 -489 300 -455
rect 334 -489 340 -455
rect 294 -527 340 -489
rect 294 -561 300 -527
rect 334 -561 340 -527
rect 294 -599 340 -561
rect 294 -633 300 -599
rect 334 -633 340 -599
rect 294 -671 340 -633
rect 294 -705 300 -671
rect 334 -705 340 -671
rect 294 -743 340 -705
rect 294 -777 300 -743
rect 334 -777 340 -743
rect 294 -815 340 -777
rect 294 -849 300 -815
rect 334 -849 340 -815
rect 294 -887 340 -849
rect 294 -921 300 -887
rect 334 -921 340 -887
rect 294 -1062 340 -921
rect 452 985 498 1114
rect 452 951 458 985
rect 492 951 498 985
rect 452 913 498 951
rect 452 879 458 913
rect 492 879 498 913
rect 452 841 498 879
rect 452 807 458 841
rect 492 807 498 841
rect 452 769 498 807
rect 452 735 458 769
rect 492 735 498 769
rect 452 697 498 735
rect 452 663 458 697
rect 492 663 498 697
rect 452 625 498 663
rect 452 591 458 625
rect 492 591 498 625
rect 452 553 498 591
rect 452 519 458 553
rect 492 519 498 553
rect 452 481 498 519
rect 452 447 458 481
rect 492 447 498 481
rect 452 409 498 447
rect 452 375 458 409
rect 492 375 498 409
rect 452 337 498 375
rect 452 303 458 337
rect 492 303 498 337
rect 452 265 498 303
rect 452 231 458 265
rect 492 231 498 265
rect 452 193 498 231
rect 452 159 458 193
rect 492 159 498 193
rect 452 121 498 159
rect 452 87 458 121
rect 492 87 498 121
rect 452 49 498 87
rect 452 15 458 49
rect 492 15 498 49
rect 452 -23 498 15
rect 452 -57 458 -23
rect 492 -57 498 -23
rect 452 -95 498 -57
rect 452 -129 458 -95
rect 492 -129 498 -95
rect 452 -167 498 -129
rect 452 -201 458 -167
rect 492 -201 498 -167
rect 452 -239 498 -201
rect 452 -273 458 -239
rect 492 -273 498 -239
rect 452 -311 498 -273
rect 452 -345 458 -311
rect 492 -345 498 -311
rect 452 -383 498 -345
rect 452 -417 458 -383
rect 492 -417 498 -383
rect 452 -455 498 -417
rect 452 -489 458 -455
rect 492 -489 498 -455
rect 452 -527 498 -489
rect 452 -561 458 -527
rect 492 -561 498 -527
rect 452 -599 498 -561
rect 452 -633 458 -599
rect 492 -633 498 -599
rect 452 -671 498 -633
rect 452 -705 458 -671
rect 492 -705 498 -671
rect 452 -743 498 -705
rect 452 -777 458 -743
rect 492 -777 498 -743
rect 452 -815 498 -777
rect 452 -849 458 -815
rect 492 -849 498 -815
rect 452 -887 498 -849
rect 452 -921 458 -887
rect 492 -921 498 -887
rect 452 -968 498 -921
rect 610 985 656 1032
rect 610 951 616 985
rect 650 951 656 985
rect 610 913 656 951
rect 610 879 616 913
rect 650 879 656 913
rect 610 841 656 879
rect 610 807 616 841
rect 650 807 656 841
rect 610 769 656 807
rect 610 735 616 769
rect 650 735 656 769
rect 610 697 656 735
rect 610 663 616 697
rect 650 663 656 697
rect 610 625 656 663
rect 610 591 616 625
rect 650 591 656 625
rect 610 553 656 591
rect 610 519 616 553
rect 650 519 656 553
rect 610 481 656 519
rect 610 447 616 481
rect 650 447 656 481
rect 610 409 656 447
rect 610 375 616 409
rect 650 375 656 409
rect 610 337 656 375
rect 610 303 616 337
rect 650 303 656 337
rect 610 265 656 303
rect 610 231 616 265
rect 650 231 656 265
rect 610 193 656 231
rect 610 159 616 193
rect 650 159 656 193
rect 610 121 656 159
rect 610 87 616 121
rect 650 87 656 121
rect 610 49 656 87
rect 610 15 616 49
rect 650 15 656 49
rect 610 -23 656 15
rect 610 -57 616 -23
rect 650 -57 656 -23
rect 610 -95 656 -57
rect 610 -129 616 -95
rect 650 -129 656 -95
rect 610 -167 656 -129
rect 610 -201 616 -167
rect 650 -201 656 -167
rect 610 -239 656 -201
rect 610 -273 616 -239
rect 650 -273 656 -239
rect 610 -311 656 -273
rect 610 -345 616 -311
rect 650 -345 656 -311
rect 610 -383 656 -345
rect 610 -417 616 -383
rect 650 -417 656 -383
rect 610 -455 656 -417
rect 610 -489 616 -455
rect 650 -489 656 -455
rect 610 -527 656 -489
rect 610 -561 616 -527
rect 650 -561 656 -527
rect 610 -599 656 -561
rect 610 -633 616 -599
rect 650 -633 656 -599
rect 610 -671 656 -633
rect 610 -705 616 -671
rect 650 -705 656 -671
rect 610 -743 656 -705
rect 610 -777 616 -743
rect 650 -777 656 -743
rect 610 -815 656 -777
rect 610 -849 616 -815
rect 650 -849 656 -815
rect 610 -887 656 -849
rect 610 -921 616 -887
rect 650 -921 656 -887
rect 610 -1062 656 -921
rect 768 985 814 1114
rect 768 951 774 985
rect 808 951 814 985
rect 768 913 814 951
rect 768 879 774 913
rect 808 879 814 913
rect 768 841 814 879
rect 768 807 774 841
rect 808 807 814 841
rect 768 769 814 807
rect 768 735 774 769
rect 808 735 814 769
rect 768 697 814 735
rect 768 663 774 697
rect 808 663 814 697
rect 768 625 814 663
rect 768 591 774 625
rect 808 591 814 625
rect 768 553 814 591
rect 768 519 774 553
rect 808 519 814 553
rect 768 481 814 519
rect 768 447 774 481
rect 808 447 814 481
rect 768 409 814 447
rect 768 375 774 409
rect 808 375 814 409
rect 768 337 814 375
rect 768 303 774 337
rect 808 303 814 337
rect 768 265 814 303
rect 768 231 774 265
rect 808 231 814 265
rect 768 193 814 231
rect 768 159 774 193
rect 808 159 814 193
rect 768 121 814 159
rect 768 87 774 121
rect 808 87 814 121
rect 768 49 814 87
rect 768 15 774 49
rect 808 15 814 49
rect 768 -23 814 15
rect 768 -57 774 -23
rect 808 -57 814 -23
rect 768 -95 814 -57
rect 768 -129 774 -95
rect 808 -129 814 -95
rect 768 -167 814 -129
rect 768 -201 774 -167
rect 808 -201 814 -167
rect 768 -239 814 -201
rect 768 -273 774 -239
rect 808 -273 814 -239
rect 768 -311 814 -273
rect 768 -345 774 -311
rect 808 -345 814 -311
rect 768 -383 814 -345
rect 768 -417 774 -383
rect 808 -417 814 -383
rect 768 -455 814 -417
rect 768 -489 774 -455
rect 808 -489 814 -455
rect 768 -527 814 -489
rect 768 -561 774 -527
rect 808 -561 814 -527
rect 768 -599 814 -561
rect 768 -633 774 -599
rect 808 -633 814 -599
rect 768 -671 814 -633
rect 768 -705 774 -671
rect 808 -705 814 -671
rect 768 -743 814 -705
rect 768 -777 774 -743
rect 808 -777 814 -743
rect 768 -815 814 -777
rect 768 -849 774 -815
rect 808 -849 814 -815
rect 768 -887 814 -849
rect 768 -921 774 -887
rect 808 -921 814 -887
rect 768 -968 814 -921
rect -654 -1108 656 -1062
rect -22 -1136 24 -1108
<< end >>
