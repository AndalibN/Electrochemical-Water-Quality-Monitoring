magic
tech sky130A
magscale 1 2
timestamp 1666625676
<< xpolycontact >>
rect -7826 85 -7756 517
rect -7826 -517 -7756 -85
rect -7508 85 -7438 517
rect -7508 -517 -7438 -85
rect -7190 85 -7120 517
rect -7190 -517 -7120 -85
rect -6872 85 -6802 517
rect -6872 -517 -6802 -85
rect -6554 85 -6484 517
rect -6554 -517 -6484 -85
rect -6236 85 -6166 517
rect -6236 -517 -6166 -85
rect -5918 85 -5848 517
rect -5918 -517 -5848 -85
rect -5600 85 -5530 517
rect -5600 -517 -5530 -85
rect -5282 85 -5212 517
rect -5282 -517 -5212 -85
rect -4964 85 -4894 517
rect -4964 -517 -4894 -85
rect -4646 85 -4576 517
rect -4646 -517 -4576 -85
rect -4328 85 -4258 517
rect -4328 -517 -4258 -85
rect -4010 85 -3940 517
rect -4010 -517 -3940 -85
rect -3692 85 -3622 517
rect -3692 -517 -3622 -85
rect -3374 85 -3304 517
rect -3374 -517 -3304 -85
rect -3056 85 -2986 517
rect -3056 -517 -2986 -85
rect -2738 85 -2668 517
rect -2738 -517 -2668 -85
rect -2420 85 -2350 517
rect -2420 -517 -2350 -85
rect -2102 85 -2032 517
rect -2102 -517 -2032 -85
rect -1784 85 -1714 517
rect -1784 -517 -1714 -85
rect -1466 85 -1396 517
rect -1466 -517 -1396 -85
rect -1148 85 -1078 517
rect -1148 -517 -1078 -85
rect -830 85 -760 517
rect -830 -517 -760 -85
rect -512 85 -442 517
rect -512 -517 -442 -85
rect -194 85 -124 517
rect -194 -517 -124 -85
rect 124 85 194 517
rect 124 -517 194 -85
rect 442 85 512 517
rect 442 -517 512 -85
rect 760 85 830 517
rect 760 -517 830 -85
rect 1078 85 1148 517
rect 1078 -517 1148 -85
rect 1396 85 1466 517
rect 1396 -517 1466 -85
rect 1714 85 1784 517
rect 1714 -517 1784 -85
rect 2032 85 2102 517
rect 2032 -517 2102 -85
rect 2350 85 2420 517
rect 2350 -517 2420 -85
rect 2668 85 2738 517
rect 2668 -517 2738 -85
rect 2986 85 3056 517
rect 2986 -517 3056 -85
rect 3304 85 3374 517
rect 3304 -517 3374 -85
rect 3622 85 3692 517
rect 3622 -517 3692 -85
rect 3940 85 4010 517
rect 3940 -517 4010 -85
rect 4258 85 4328 517
rect 4258 -517 4328 -85
rect 4576 85 4646 517
rect 4576 -517 4646 -85
rect 4894 85 4964 517
rect 4894 -517 4964 -85
rect 5212 85 5282 517
rect 5212 -517 5282 -85
rect 5530 85 5600 517
rect 5530 -517 5600 -85
rect 5848 85 5918 517
rect 5848 -517 5918 -85
rect 6166 85 6236 517
rect 6166 -517 6236 -85
rect 6484 85 6554 517
rect 6484 -517 6554 -85
rect 6802 85 6872 517
rect 6802 -517 6872 -85
rect 7120 85 7190 517
rect 7120 -517 7190 -85
rect 7438 85 7508 517
rect 7438 -517 7508 -85
rect 7756 85 7826 517
rect 7756 -517 7826 -85
<< xpolyres >>
rect -7826 -85 -7756 85
rect -7508 -85 -7438 85
rect -7190 -85 -7120 85
rect -6872 -85 -6802 85
rect -6554 -85 -6484 85
rect -6236 -85 -6166 85
rect -5918 -85 -5848 85
rect -5600 -85 -5530 85
rect -5282 -85 -5212 85
rect -4964 -85 -4894 85
rect -4646 -85 -4576 85
rect -4328 -85 -4258 85
rect -4010 -85 -3940 85
rect -3692 -85 -3622 85
rect -3374 -85 -3304 85
rect -3056 -85 -2986 85
rect -2738 -85 -2668 85
rect -2420 -85 -2350 85
rect -2102 -85 -2032 85
rect -1784 -85 -1714 85
rect -1466 -85 -1396 85
rect -1148 -85 -1078 85
rect -830 -85 -760 85
rect -512 -85 -442 85
rect -194 -85 -124 85
rect 124 -85 194 85
rect 442 -85 512 85
rect 760 -85 830 85
rect 1078 -85 1148 85
rect 1396 -85 1466 85
rect 1714 -85 1784 85
rect 2032 -85 2102 85
rect 2350 -85 2420 85
rect 2668 -85 2738 85
rect 2986 -85 3056 85
rect 3304 -85 3374 85
rect 3622 -85 3692 85
rect 3940 -85 4010 85
rect 4258 -85 4328 85
rect 4576 -85 4646 85
rect 4894 -85 4964 85
rect 5212 -85 5282 85
rect 5530 -85 5600 85
rect 5848 -85 5918 85
rect 6166 -85 6236 85
rect 6484 -85 6554 85
rect 6802 -85 6872 85
rect 7120 -85 7190 85
rect 7438 -85 7508 85
rect 7756 -85 7826 85
<< viali >>
rect -7810 102 -7772 499
rect -7492 102 -7454 499
rect -7174 102 -7136 499
rect -6856 102 -6818 499
rect -6538 102 -6500 499
rect -6220 102 -6182 499
rect -5902 102 -5864 499
rect -5584 102 -5546 499
rect -5266 102 -5228 499
rect -4948 102 -4910 499
rect -4630 102 -4592 499
rect -4312 102 -4274 499
rect -3994 102 -3956 499
rect -3676 102 -3638 499
rect -3358 102 -3320 499
rect -3040 102 -3002 499
rect -2722 102 -2684 499
rect -2404 102 -2366 499
rect -2086 102 -2048 499
rect -1768 102 -1730 499
rect -1450 102 -1412 499
rect -1132 102 -1094 499
rect -814 102 -776 499
rect -496 102 -458 499
rect -178 102 -140 499
rect 140 102 178 499
rect 458 102 496 499
rect 776 102 814 499
rect 1094 102 1132 499
rect 1412 102 1450 499
rect 1730 102 1768 499
rect 2048 102 2086 499
rect 2366 102 2404 499
rect 2684 102 2722 499
rect 3002 102 3040 499
rect 3320 102 3358 499
rect 3638 102 3676 499
rect 3956 102 3994 499
rect 4274 102 4312 499
rect 4592 102 4630 499
rect 4910 102 4948 499
rect 5228 102 5266 499
rect 5546 102 5584 499
rect 5864 102 5902 499
rect 6182 102 6220 499
rect 6500 102 6538 499
rect 6818 102 6856 499
rect 7136 102 7174 499
rect 7454 102 7492 499
rect 7772 102 7810 499
rect -7810 -499 -7772 -102
rect -7492 -499 -7454 -102
rect -7174 -499 -7136 -102
rect -6856 -499 -6818 -102
rect -6538 -499 -6500 -102
rect -6220 -499 -6182 -102
rect -5902 -499 -5864 -102
rect -5584 -499 -5546 -102
rect -5266 -499 -5228 -102
rect -4948 -499 -4910 -102
rect -4630 -499 -4592 -102
rect -4312 -499 -4274 -102
rect -3994 -499 -3956 -102
rect -3676 -499 -3638 -102
rect -3358 -499 -3320 -102
rect -3040 -499 -3002 -102
rect -2722 -499 -2684 -102
rect -2404 -499 -2366 -102
rect -2086 -499 -2048 -102
rect -1768 -499 -1730 -102
rect -1450 -499 -1412 -102
rect -1132 -499 -1094 -102
rect -814 -499 -776 -102
rect -496 -499 -458 -102
rect -178 -499 -140 -102
rect 140 -499 178 -102
rect 458 -499 496 -102
rect 776 -499 814 -102
rect 1094 -499 1132 -102
rect 1412 -499 1450 -102
rect 1730 -499 1768 -102
rect 2048 -499 2086 -102
rect 2366 -499 2404 -102
rect 2684 -499 2722 -102
rect 3002 -499 3040 -102
rect 3320 -499 3358 -102
rect 3638 -499 3676 -102
rect 3956 -499 3994 -102
rect 4274 -499 4312 -102
rect 4592 -499 4630 -102
rect 4910 -499 4948 -102
rect 5228 -499 5266 -102
rect 5546 -499 5584 -102
rect 5864 -499 5902 -102
rect 6182 -499 6220 -102
rect 6500 -499 6538 -102
rect 6818 -499 6856 -102
rect 7136 -499 7174 -102
rect 7454 -499 7492 -102
rect 7772 -499 7810 -102
<< metal1 >>
rect -7816 499 -7766 511
rect -7816 102 -7810 499
rect -7772 102 -7766 499
rect -7816 90 -7766 102
rect -7498 499 -7448 511
rect -7498 102 -7492 499
rect -7454 102 -7448 499
rect -7498 90 -7448 102
rect -7180 499 -7130 511
rect -7180 102 -7174 499
rect -7136 102 -7130 499
rect -7180 90 -7130 102
rect -6862 499 -6812 511
rect -6862 102 -6856 499
rect -6818 102 -6812 499
rect -6862 90 -6812 102
rect -6544 499 -6494 511
rect -6544 102 -6538 499
rect -6500 102 -6494 499
rect -6544 90 -6494 102
rect -6226 499 -6176 511
rect -6226 102 -6220 499
rect -6182 102 -6176 499
rect -6226 90 -6176 102
rect -5908 499 -5858 511
rect -5908 102 -5902 499
rect -5864 102 -5858 499
rect -5908 90 -5858 102
rect -5590 499 -5540 511
rect -5590 102 -5584 499
rect -5546 102 -5540 499
rect -5590 90 -5540 102
rect -5272 499 -5222 511
rect -5272 102 -5266 499
rect -5228 102 -5222 499
rect -5272 90 -5222 102
rect -4954 499 -4904 511
rect -4954 102 -4948 499
rect -4910 102 -4904 499
rect -4954 90 -4904 102
rect -4636 499 -4586 511
rect -4636 102 -4630 499
rect -4592 102 -4586 499
rect -4636 90 -4586 102
rect -4318 499 -4268 511
rect -4318 102 -4312 499
rect -4274 102 -4268 499
rect -4318 90 -4268 102
rect -4000 499 -3950 511
rect -4000 102 -3994 499
rect -3956 102 -3950 499
rect -4000 90 -3950 102
rect -3682 499 -3632 511
rect -3682 102 -3676 499
rect -3638 102 -3632 499
rect -3682 90 -3632 102
rect -3364 499 -3314 511
rect -3364 102 -3358 499
rect -3320 102 -3314 499
rect -3364 90 -3314 102
rect -3046 499 -2996 511
rect -3046 102 -3040 499
rect -3002 102 -2996 499
rect -3046 90 -2996 102
rect -2728 499 -2678 511
rect -2728 102 -2722 499
rect -2684 102 -2678 499
rect -2728 90 -2678 102
rect -2410 499 -2360 511
rect -2410 102 -2404 499
rect -2366 102 -2360 499
rect -2410 90 -2360 102
rect -2092 499 -2042 511
rect -2092 102 -2086 499
rect -2048 102 -2042 499
rect -2092 90 -2042 102
rect -1774 499 -1724 511
rect -1774 102 -1768 499
rect -1730 102 -1724 499
rect -1774 90 -1724 102
rect -1456 499 -1406 511
rect -1456 102 -1450 499
rect -1412 102 -1406 499
rect -1456 90 -1406 102
rect -1138 499 -1088 511
rect -1138 102 -1132 499
rect -1094 102 -1088 499
rect -1138 90 -1088 102
rect -820 499 -770 511
rect -820 102 -814 499
rect -776 102 -770 499
rect -820 90 -770 102
rect -502 499 -452 511
rect -502 102 -496 499
rect -458 102 -452 499
rect -502 90 -452 102
rect -184 499 -134 511
rect -184 102 -178 499
rect -140 102 -134 499
rect -184 90 -134 102
rect 134 499 184 511
rect 134 102 140 499
rect 178 102 184 499
rect 134 90 184 102
rect 452 499 502 511
rect 452 102 458 499
rect 496 102 502 499
rect 452 90 502 102
rect 770 499 820 511
rect 770 102 776 499
rect 814 102 820 499
rect 770 90 820 102
rect 1088 499 1138 511
rect 1088 102 1094 499
rect 1132 102 1138 499
rect 1088 90 1138 102
rect 1406 499 1456 511
rect 1406 102 1412 499
rect 1450 102 1456 499
rect 1406 90 1456 102
rect 1724 499 1774 511
rect 1724 102 1730 499
rect 1768 102 1774 499
rect 1724 90 1774 102
rect 2042 499 2092 511
rect 2042 102 2048 499
rect 2086 102 2092 499
rect 2042 90 2092 102
rect 2360 499 2410 511
rect 2360 102 2366 499
rect 2404 102 2410 499
rect 2360 90 2410 102
rect 2678 499 2728 511
rect 2678 102 2684 499
rect 2722 102 2728 499
rect 2678 90 2728 102
rect 2996 499 3046 511
rect 2996 102 3002 499
rect 3040 102 3046 499
rect 2996 90 3046 102
rect 3314 499 3364 511
rect 3314 102 3320 499
rect 3358 102 3364 499
rect 3314 90 3364 102
rect 3632 499 3682 511
rect 3632 102 3638 499
rect 3676 102 3682 499
rect 3632 90 3682 102
rect 3950 499 4000 511
rect 3950 102 3956 499
rect 3994 102 4000 499
rect 3950 90 4000 102
rect 4268 499 4318 511
rect 4268 102 4274 499
rect 4312 102 4318 499
rect 4268 90 4318 102
rect 4586 499 4636 511
rect 4586 102 4592 499
rect 4630 102 4636 499
rect 4586 90 4636 102
rect 4904 499 4954 511
rect 4904 102 4910 499
rect 4948 102 4954 499
rect 4904 90 4954 102
rect 5222 499 5272 511
rect 5222 102 5228 499
rect 5266 102 5272 499
rect 5222 90 5272 102
rect 5540 499 5590 511
rect 5540 102 5546 499
rect 5584 102 5590 499
rect 5540 90 5590 102
rect 5858 499 5908 511
rect 5858 102 5864 499
rect 5902 102 5908 499
rect 5858 90 5908 102
rect 6176 499 6226 511
rect 6176 102 6182 499
rect 6220 102 6226 499
rect 6176 90 6226 102
rect 6494 499 6544 511
rect 6494 102 6500 499
rect 6538 102 6544 499
rect 6494 90 6544 102
rect 6812 499 6862 511
rect 6812 102 6818 499
rect 6856 102 6862 499
rect 6812 90 6862 102
rect 7130 499 7180 511
rect 7130 102 7136 499
rect 7174 102 7180 499
rect 7130 90 7180 102
rect 7448 499 7498 511
rect 7448 102 7454 499
rect 7492 102 7498 499
rect 7448 90 7498 102
rect 7766 499 7816 511
rect 7766 102 7772 499
rect 7810 102 7816 499
rect 7766 90 7816 102
rect -7816 -102 -7766 -90
rect -7816 -499 -7810 -102
rect -7772 -499 -7766 -102
rect -7816 -511 -7766 -499
rect -7498 -102 -7448 -90
rect -7498 -499 -7492 -102
rect -7454 -499 -7448 -102
rect -7498 -511 -7448 -499
rect -7180 -102 -7130 -90
rect -7180 -499 -7174 -102
rect -7136 -499 -7130 -102
rect -7180 -511 -7130 -499
rect -6862 -102 -6812 -90
rect -6862 -499 -6856 -102
rect -6818 -499 -6812 -102
rect -6862 -511 -6812 -499
rect -6544 -102 -6494 -90
rect -6544 -499 -6538 -102
rect -6500 -499 -6494 -102
rect -6544 -511 -6494 -499
rect -6226 -102 -6176 -90
rect -6226 -499 -6220 -102
rect -6182 -499 -6176 -102
rect -6226 -511 -6176 -499
rect -5908 -102 -5858 -90
rect -5908 -499 -5902 -102
rect -5864 -499 -5858 -102
rect -5908 -511 -5858 -499
rect -5590 -102 -5540 -90
rect -5590 -499 -5584 -102
rect -5546 -499 -5540 -102
rect -5590 -511 -5540 -499
rect -5272 -102 -5222 -90
rect -5272 -499 -5266 -102
rect -5228 -499 -5222 -102
rect -5272 -511 -5222 -499
rect -4954 -102 -4904 -90
rect -4954 -499 -4948 -102
rect -4910 -499 -4904 -102
rect -4954 -511 -4904 -499
rect -4636 -102 -4586 -90
rect -4636 -499 -4630 -102
rect -4592 -499 -4586 -102
rect -4636 -511 -4586 -499
rect -4318 -102 -4268 -90
rect -4318 -499 -4312 -102
rect -4274 -499 -4268 -102
rect -4318 -511 -4268 -499
rect -4000 -102 -3950 -90
rect -4000 -499 -3994 -102
rect -3956 -499 -3950 -102
rect -4000 -511 -3950 -499
rect -3682 -102 -3632 -90
rect -3682 -499 -3676 -102
rect -3638 -499 -3632 -102
rect -3682 -511 -3632 -499
rect -3364 -102 -3314 -90
rect -3364 -499 -3358 -102
rect -3320 -499 -3314 -102
rect -3364 -511 -3314 -499
rect -3046 -102 -2996 -90
rect -3046 -499 -3040 -102
rect -3002 -499 -2996 -102
rect -3046 -511 -2996 -499
rect -2728 -102 -2678 -90
rect -2728 -499 -2722 -102
rect -2684 -499 -2678 -102
rect -2728 -511 -2678 -499
rect -2410 -102 -2360 -90
rect -2410 -499 -2404 -102
rect -2366 -499 -2360 -102
rect -2410 -511 -2360 -499
rect -2092 -102 -2042 -90
rect -2092 -499 -2086 -102
rect -2048 -499 -2042 -102
rect -2092 -511 -2042 -499
rect -1774 -102 -1724 -90
rect -1774 -499 -1768 -102
rect -1730 -499 -1724 -102
rect -1774 -511 -1724 -499
rect -1456 -102 -1406 -90
rect -1456 -499 -1450 -102
rect -1412 -499 -1406 -102
rect -1456 -511 -1406 -499
rect -1138 -102 -1088 -90
rect -1138 -499 -1132 -102
rect -1094 -499 -1088 -102
rect -1138 -511 -1088 -499
rect -820 -102 -770 -90
rect -820 -499 -814 -102
rect -776 -499 -770 -102
rect -820 -511 -770 -499
rect -502 -102 -452 -90
rect -502 -499 -496 -102
rect -458 -499 -452 -102
rect -502 -511 -452 -499
rect -184 -102 -134 -90
rect -184 -499 -178 -102
rect -140 -499 -134 -102
rect -184 -511 -134 -499
rect 134 -102 184 -90
rect 134 -499 140 -102
rect 178 -499 184 -102
rect 134 -511 184 -499
rect 452 -102 502 -90
rect 452 -499 458 -102
rect 496 -499 502 -102
rect 452 -511 502 -499
rect 770 -102 820 -90
rect 770 -499 776 -102
rect 814 -499 820 -102
rect 770 -511 820 -499
rect 1088 -102 1138 -90
rect 1088 -499 1094 -102
rect 1132 -499 1138 -102
rect 1088 -511 1138 -499
rect 1406 -102 1456 -90
rect 1406 -499 1412 -102
rect 1450 -499 1456 -102
rect 1406 -511 1456 -499
rect 1724 -102 1774 -90
rect 1724 -499 1730 -102
rect 1768 -499 1774 -102
rect 1724 -511 1774 -499
rect 2042 -102 2092 -90
rect 2042 -499 2048 -102
rect 2086 -499 2092 -102
rect 2042 -511 2092 -499
rect 2360 -102 2410 -90
rect 2360 -499 2366 -102
rect 2404 -499 2410 -102
rect 2360 -511 2410 -499
rect 2678 -102 2728 -90
rect 2678 -499 2684 -102
rect 2722 -499 2728 -102
rect 2678 -511 2728 -499
rect 2996 -102 3046 -90
rect 2996 -499 3002 -102
rect 3040 -499 3046 -102
rect 2996 -511 3046 -499
rect 3314 -102 3364 -90
rect 3314 -499 3320 -102
rect 3358 -499 3364 -102
rect 3314 -511 3364 -499
rect 3632 -102 3682 -90
rect 3632 -499 3638 -102
rect 3676 -499 3682 -102
rect 3632 -511 3682 -499
rect 3950 -102 4000 -90
rect 3950 -499 3956 -102
rect 3994 -499 4000 -102
rect 3950 -511 4000 -499
rect 4268 -102 4318 -90
rect 4268 -499 4274 -102
rect 4312 -499 4318 -102
rect 4268 -511 4318 -499
rect 4586 -102 4636 -90
rect 4586 -499 4592 -102
rect 4630 -499 4636 -102
rect 4586 -511 4636 -499
rect 4904 -102 4954 -90
rect 4904 -499 4910 -102
rect 4948 -499 4954 -102
rect 4904 -511 4954 -499
rect 5222 -102 5272 -90
rect 5222 -499 5228 -102
rect 5266 -499 5272 -102
rect 5222 -511 5272 -499
rect 5540 -102 5590 -90
rect 5540 -499 5546 -102
rect 5584 -499 5590 -102
rect 5540 -511 5590 -499
rect 5858 -102 5908 -90
rect 5858 -499 5864 -102
rect 5902 -499 5908 -102
rect 5858 -511 5908 -499
rect 6176 -102 6226 -90
rect 6176 -499 6182 -102
rect 6220 -499 6226 -102
rect 6176 -511 6226 -499
rect 6494 -102 6544 -90
rect 6494 -499 6500 -102
rect 6538 -499 6544 -102
rect 6494 -511 6544 -499
rect 6812 -102 6862 -90
rect 6812 -499 6818 -102
rect 6856 -499 6862 -102
rect 6812 -511 6862 -499
rect 7130 -102 7180 -90
rect 7130 -499 7136 -102
rect 7174 -499 7180 -102
rect 7130 -511 7180 -499
rect 7448 -102 7498 -90
rect 7448 -499 7454 -102
rect 7492 -499 7498 -102
rect 7448 -511 7498 -499
rect 7766 -102 7816 -90
rect 7766 -499 7772 -102
rect 7810 -499 7816 -102
rect 7766 -511 7816 -499
<< res0p35 >>
rect -7828 -87 -7754 87
rect -7510 -87 -7436 87
rect -7192 -87 -7118 87
rect -6874 -87 -6800 87
rect -6556 -87 -6482 87
rect -6238 -87 -6164 87
rect -5920 -87 -5846 87
rect -5602 -87 -5528 87
rect -5284 -87 -5210 87
rect -4966 -87 -4892 87
rect -4648 -87 -4574 87
rect -4330 -87 -4256 87
rect -4012 -87 -3938 87
rect -3694 -87 -3620 87
rect -3376 -87 -3302 87
rect -3058 -87 -2984 87
rect -2740 -87 -2666 87
rect -2422 -87 -2348 87
rect -2104 -87 -2030 87
rect -1786 -87 -1712 87
rect -1468 -87 -1394 87
rect -1150 -87 -1076 87
rect -832 -87 -758 87
rect -514 -87 -440 87
rect -196 -87 -122 87
rect 122 -87 196 87
rect 440 -87 514 87
rect 758 -87 832 87
rect 1076 -87 1150 87
rect 1394 -87 1468 87
rect 1712 -87 1786 87
rect 2030 -87 2104 87
rect 2348 -87 2422 87
rect 2666 -87 2740 87
rect 2984 -87 3058 87
rect 3302 -87 3376 87
rect 3620 -87 3694 87
rect 3938 -87 4012 87
rect 4256 -87 4330 87
rect 4574 -87 4648 87
rect 4892 -87 4966 87
rect 5210 -87 5284 87
rect 5528 -87 5602 87
rect 5846 -87 5920 87
rect 6164 -87 6238 87
rect 6482 -87 6556 87
rect 6800 -87 6874 87
rect 7118 -87 7192 87
rect 7436 -87 7510 87
rect 7754 -87 7828 87
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.85 m 1 nx 50 wmin 0.350 lmin 0.50 rho 2000 val 5.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
