magic
tech sky130A
magscale 1 2
timestamp 1676693800
<< metal1 >>
rect -5921 738 -5424 790
rect -5921 344 -5870 738
rect -5484 642 -5424 738
rect -5484 508 -4608 642
rect -5484 344 -5424 508
rect -5921 293 -5424 344
<< via1 >>
rect -5870 344 -5484 738
<< metal2 >>
rect -5921 738 -5424 790
rect -5921 344 -5870 738
rect -5484 344 -5424 738
rect -5921 293 -5424 344
<< via2 >>
rect -5870 344 -5484 738
<< metal3 >>
rect -5921 738 -5424 790
rect -5921 344 -5870 738
rect -5484 344 -5424 738
rect -5921 293 -5424 344
<< via3 >>
rect -5870 344 -5484 738
<< metal4 >>
rect -56060 738 -5424 790
rect -56060 344 -5870 738
rect -5484 344 -5424 738
rect -56060 293 -5424 344
use VCO  VCO_0
timestamp 1671232119
transform 1 0 -4102 0 1 806
box -808 -1396 2776 990
use tia  tia_0
timestamp 1670179985
transform 1 0 -73806 0 1 -3591
box -1768 -1627 18245 8897
<< end >>
