magic
tech sky130A
magscale 1 2
timestamp 1668226266
<< xpolycontact >>
rect -353 157 -283 589
rect -353 -589 -283 -157
rect -35 157 35 589
rect -35 -589 35 -157
rect 283 157 353 589
rect 283 -589 353 -157
<< xpolyres >>
rect -353 -157 -283 157
rect -35 -157 35 157
rect 283 -157 353 157
<< viali >>
rect -337 174 -299 571
rect -19 174 19 571
rect 299 174 337 571
rect -337 -571 -299 -174
rect -19 -571 19 -174
rect 299 -571 337 -174
<< metal1 >>
rect -343 571 -293 583
rect -343 174 -337 571
rect -299 174 -293 571
rect -343 162 -293 174
rect -25 571 25 583
rect -25 174 -19 571
rect 19 174 25 571
rect -25 162 25 174
rect 293 571 343 583
rect 293 174 299 571
rect 337 174 343 571
rect 293 162 343 174
rect -343 -174 -293 -162
rect -343 -571 -337 -174
rect -299 -571 -293 -174
rect -343 -583 -293 -571
rect -25 -174 25 -162
rect -25 -571 -19 -174
rect 19 -571 25 -174
rect -25 -583 25 -571
rect 293 -174 343 -162
rect 293 -571 299 -174
rect 337 -571 343 -174
rect 293 -583 343 -571
<< res0p35 >>
rect -355 -159 -281 159
rect -37 -159 37 159
rect 281 -159 355 159
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 1.57 m 1 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 10.046k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
