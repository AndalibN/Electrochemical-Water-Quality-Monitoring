magic
tech sky130A
timestamp 1668374365
<< nmos >>
rect -1407 -4800 -1377 4800
rect -1291 -4800 -1261 4800
rect -1175 -4800 -1145 4800
rect -1059 -4800 -1029 4800
rect -943 -4800 -913 4800
rect -827 -4800 -797 4800
rect -711 -4800 -681 4800
rect -595 -4800 -565 4800
rect -479 -4800 -449 4800
rect -363 -4800 -333 4800
rect -247 -4800 -217 4800
rect -131 -4800 -101 4800
rect -15 -4800 15 4800
rect 101 -4800 131 4800
rect 217 -4800 247 4800
rect 333 -4800 363 4800
rect 449 -4800 479 4800
rect 565 -4800 595 4800
rect 681 -4800 711 4800
rect 797 -4800 827 4800
rect 913 -4800 943 4800
rect 1029 -4800 1059 4800
rect 1145 -4800 1175 4800
rect 1261 -4800 1291 4800
rect 1377 -4800 1407 4800
<< ndiff >>
rect -1436 4794 -1407 4800
rect -1436 -4794 -1430 4794
rect -1413 -4794 -1407 4794
rect -1436 -4800 -1407 -4794
rect -1377 4794 -1348 4800
rect -1377 -4794 -1371 4794
rect -1354 -4794 -1348 4794
rect -1377 -4800 -1348 -4794
rect -1320 4794 -1291 4800
rect -1320 -4794 -1314 4794
rect -1297 -4794 -1291 4794
rect -1320 -4800 -1291 -4794
rect -1261 4794 -1232 4800
rect -1261 -4794 -1255 4794
rect -1238 -4794 -1232 4794
rect -1261 -4800 -1232 -4794
rect -1204 4794 -1175 4800
rect -1204 -4794 -1198 4794
rect -1181 -4794 -1175 4794
rect -1204 -4800 -1175 -4794
rect -1145 4794 -1116 4800
rect -1145 -4794 -1139 4794
rect -1122 -4794 -1116 4794
rect -1145 -4800 -1116 -4794
rect -1088 4794 -1059 4800
rect -1088 -4794 -1082 4794
rect -1065 -4794 -1059 4794
rect -1088 -4800 -1059 -4794
rect -1029 4794 -1000 4800
rect -1029 -4794 -1023 4794
rect -1006 -4794 -1000 4794
rect -1029 -4800 -1000 -4794
rect -972 4794 -943 4800
rect -972 -4794 -966 4794
rect -949 -4794 -943 4794
rect -972 -4800 -943 -4794
rect -913 4794 -884 4800
rect -913 -4794 -907 4794
rect -890 -4794 -884 4794
rect -913 -4800 -884 -4794
rect -856 4794 -827 4800
rect -856 -4794 -850 4794
rect -833 -4794 -827 4794
rect -856 -4800 -827 -4794
rect -797 4794 -768 4800
rect -797 -4794 -791 4794
rect -774 -4794 -768 4794
rect -797 -4800 -768 -4794
rect -740 4794 -711 4800
rect -740 -4794 -734 4794
rect -717 -4794 -711 4794
rect -740 -4800 -711 -4794
rect -681 4794 -652 4800
rect -681 -4794 -675 4794
rect -658 -4794 -652 4794
rect -681 -4800 -652 -4794
rect -624 4794 -595 4800
rect -624 -4794 -618 4794
rect -601 -4794 -595 4794
rect -624 -4800 -595 -4794
rect -565 4794 -536 4800
rect -565 -4794 -559 4794
rect -542 -4794 -536 4794
rect -565 -4800 -536 -4794
rect -508 4794 -479 4800
rect -508 -4794 -502 4794
rect -485 -4794 -479 4794
rect -508 -4800 -479 -4794
rect -449 4794 -420 4800
rect -449 -4794 -443 4794
rect -426 -4794 -420 4794
rect -449 -4800 -420 -4794
rect -392 4794 -363 4800
rect -392 -4794 -386 4794
rect -369 -4794 -363 4794
rect -392 -4800 -363 -4794
rect -333 4794 -304 4800
rect -333 -4794 -327 4794
rect -310 -4794 -304 4794
rect -333 -4800 -304 -4794
rect -276 4794 -247 4800
rect -276 -4794 -270 4794
rect -253 -4794 -247 4794
rect -276 -4800 -247 -4794
rect -217 4794 -188 4800
rect -217 -4794 -211 4794
rect -194 -4794 -188 4794
rect -217 -4800 -188 -4794
rect -160 4794 -131 4800
rect -160 -4794 -154 4794
rect -137 -4794 -131 4794
rect -160 -4800 -131 -4794
rect -101 4794 -72 4800
rect -101 -4794 -95 4794
rect -78 -4794 -72 4794
rect -101 -4800 -72 -4794
rect -44 4794 -15 4800
rect -44 -4794 -38 4794
rect -21 -4794 -15 4794
rect -44 -4800 -15 -4794
rect 15 4794 44 4800
rect 15 -4794 21 4794
rect 38 -4794 44 4794
rect 15 -4800 44 -4794
rect 72 4794 101 4800
rect 72 -4794 78 4794
rect 95 -4794 101 4794
rect 72 -4800 101 -4794
rect 131 4794 160 4800
rect 131 -4794 137 4794
rect 154 -4794 160 4794
rect 131 -4800 160 -4794
rect 188 4794 217 4800
rect 188 -4794 194 4794
rect 211 -4794 217 4794
rect 188 -4800 217 -4794
rect 247 4794 276 4800
rect 247 -4794 253 4794
rect 270 -4794 276 4794
rect 247 -4800 276 -4794
rect 304 4794 333 4800
rect 304 -4794 310 4794
rect 327 -4794 333 4794
rect 304 -4800 333 -4794
rect 363 4794 392 4800
rect 363 -4794 369 4794
rect 386 -4794 392 4794
rect 363 -4800 392 -4794
rect 420 4794 449 4800
rect 420 -4794 426 4794
rect 443 -4794 449 4794
rect 420 -4800 449 -4794
rect 479 4794 508 4800
rect 479 -4794 485 4794
rect 502 -4794 508 4794
rect 479 -4800 508 -4794
rect 536 4794 565 4800
rect 536 -4794 542 4794
rect 559 -4794 565 4794
rect 536 -4800 565 -4794
rect 595 4794 624 4800
rect 595 -4794 601 4794
rect 618 -4794 624 4794
rect 595 -4800 624 -4794
rect 652 4794 681 4800
rect 652 -4794 658 4794
rect 675 -4794 681 4794
rect 652 -4800 681 -4794
rect 711 4794 740 4800
rect 711 -4794 717 4794
rect 734 -4794 740 4794
rect 711 -4800 740 -4794
rect 768 4794 797 4800
rect 768 -4794 774 4794
rect 791 -4794 797 4794
rect 768 -4800 797 -4794
rect 827 4794 856 4800
rect 827 -4794 833 4794
rect 850 -4794 856 4794
rect 827 -4800 856 -4794
rect 884 4794 913 4800
rect 884 -4794 890 4794
rect 907 -4794 913 4794
rect 884 -4800 913 -4794
rect 943 4794 972 4800
rect 943 -4794 949 4794
rect 966 -4794 972 4794
rect 943 -4800 972 -4794
rect 1000 4794 1029 4800
rect 1000 -4794 1006 4794
rect 1023 -4794 1029 4794
rect 1000 -4800 1029 -4794
rect 1059 4794 1088 4800
rect 1059 -4794 1065 4794
rect 1082 -4794 1088 4794
rect 1059 -4800 1088 -4794
rect 1116 4794 1145 4800
rect 1116 -4794 1122 4794
rect 1139 -4794 1145 4794
rect 1116 -4800 1145 -4794
rect 1175 4794 1204 4800
rect 1175 -4794 1181 4794
rect 1198 -4794 1204 4794
rect 1175 -4800 1204 -4794
rect 1232 4794 1261 4800
rect 1232 -4794 1238 4794
rect 1255 -4794 1261 4794
rect 1232 -4800 1261 -4794
rect 1291 4794 1320 4800
rect 1291 -4794 1297 4794
rect 1314 -4794 1320 4794
rect 1291 -4800 1320 -4794
rect 1348 4794 1377 4800
rect 1348 -4794 1354 4794
rect 1371 -4794 1377 4794
rect 1348 -4800 1377 -4794
rect 1407 4794 1436 4800
rect 1407 -4794 1413 4794
rect 1430 -4794 1436 4794
rect 1407 -4800 1436 -4794
<< ndiffc >>
rect -1430 -4794 -1413 4794
rect -1371 -4794 -1354 4794
rect -1314 -4794 -1297 4794
rect -1255 -4794 -1238 4794
rect -1198 -4794 -1181 4794
rect -1139 -4794 -1122 4794
rect -1082 -4794 -1065 4794
rect -1023 -4794 -1006 4794
rect -966 -4794 -949 4794
rect -907 -4794 -890 4794
rect -850 -4794 -833 4794
rect -791 -4794 -774 4794
rect -734 -4794 -717 4794
rect -675 -4794 -658 4794
rect -618 -4794 -601 4794
rect -559 -4794 -542 4794
rect -502 -4794 -485 4794
rect -443 -4794 -426 4794
rect -386 -4794 -369 4794
rect -327 -4794 -310 4794
rect -270 -4794 -253 4794
rect -211 -4794 -194 4794
rect -154 -4794 -137 4794
rect -95 -4794 -78 4794
rect -38 -4794 -21 4794
rect 21 -4794 38 4794
rect 78 -4794 95 4794
rect 137 -4794 154 4794
rect 194 -4794 211 4794
rect 253 -4794 270 4794
rect 310 -4794 327 4794
rect 369 -4794 386 4794
rect 426 -4794 443 4794
rect 485 -4794 502 4794
rect 542 -4794 559 4794
rect 601 -4794 618 4794
rect 658 -4794 675 4794
rect 717 -4794 734 4794
rect 774 -4794 791 4794
rect 833 -4794 850 4794
rect 890 -4794 907 4794
rect 949 -4794 966 4794
rect 1006 -4794 1023 4794
rect 1065 -4794 1082 4794
rect 1122 -4794 1139 4794
rect 1181 -4794 1198 4794
rect 1238 -4794 1255 4794
rect 1297 -4794 1314 4794
rect 1354 -4794 1371 4794
rect 1413 -4794 1430 4794
<< poly >>
rect -1407 4800 -1377 4813
rect -1291 4800 -1261 4813
rect -1175 4800 -1145 4813
rect -1059 4800 -1029 4813
rect -943 4800 -913 4813
rect -827 4800 -797 4813
rect -711 4800 -681 4813
rect -595 4800 -565 4813
rect -479 4800 -449 4813
rect -363 4800 -333 4813
rect -247 4800 -217 4813
rect -131 4800 -101 4813
rect -15 4800 15 4813
rect 101 4800 131 4813
rect 217 4800 247 4813
rect 333 4800 363 4813
rect 449 4800 479 4813
rect 565 4800 595 4813
rect 681 4800 711 4813
rect 797 4800 827 4813
rect 913 4800 943 4813
rect 1029 4800 1059 4813
rect 1145 4800 1175 4813
rect 1261 4800 1291 4813
rect 1377 4800 1407 4813
rect -1407 -4813 -1377 -4800
rect -1291 -4813 -1261 -4800
rect -1175 -4813 -1145 -4800
rect -1059 -4813 -1029 -4800
rect -943 -4813 -913 -4800
rect -827 -4813 -797 -4800
rect -711 -4813 -681 -4800
rect -595 -4813 -565 -4800
rect -479 -4813 -449 -4800
rect -363 -4813 -333 -4800
rect -247 -4813 -217 -4800
rect -131 -4813 -101 -4800
rect -15 -4813 15 -4800
rect 101 -4813 131 -4800
rect 217 -4813 247 -4800
rect 333 -4813 363 -4800
rect 449 -4813 479 -4800
rect 565 -4813 595 -4800
rect 681 -4813 711 -4800
rect 797 -4813 827 -4800
rect 913 -4813 943 -4800
rect 1029 -4813 1059 -4800
rect 1145 -4813 1175 -4800
rect 1261 -4813 1291 -4800
rect 1377 -4813 1407 -4800
<< locali >>
rect -1430 4794 -1413 4802
rect -1430 -4802 -1413 -4794
rect -1371 4794 -1354 4802
rect -1371 -4802 -1354 -4794
rect -1314 4794 -1297 4802
rect -1314 -4802 -1297 -4794
rect -1255 4794 -1238 4802
rect -1255 -4802 -1238 -4794
rect -1198 4794 -1181 4802
rect -1198 -4802 -1181 -4794
rect -1139 4794 -1122 4802
rect -1139 -4802 -1122 -4794
rect -1082 4794 -1065 4802
rect -1082 -4802 -1065 -4794
rect -1023 4794 -1006 4802
rect -1023 -4802 -1006 -4794
rect -966 4794 -949 4802
rect -966 -4802 -949 -4794
rect -907 4794 -890 4802
rect -907 -4802 -890 -4794
rect -850 4794 -833 4802
rect -850 -4802 -833 -4794
rect -791 4794 -774 4802
rect -791 -4802 -774 -4794
rect -734 4794 -717 4802
rect -734 -4802 -717 -4794
rect -675 4794 -658 4802
rect -675 -4802 -658 -4794
rect -618 4794 -601 4802
rect -618 -4802 -601 -4794
rect -559 4794 -542 4802
rect -559 -4802 -542 -4794
rect -502 4794 -485 4802
rect -502 -4802 -485 -4794
rect -443 4794 -426 4802
rect -443 -4802 -426 -4794
rect -386 4794 -369 4802
rect -386 -4802 -369 -4794
rect -327 4794 -310 4802
rect -327 -4802 -310 -4794
rect -270 4794 -253 4802
rect -270 -4802 -253 -4794
rect -211 4794 -194 4802
rect -211 -4802 -194 -4794
rect -154 4794 -137 4802
rect -154 -4802 -137 -4794
rect -95 4794 -78 4802
rect -95 -4802 -78 -4794
rect -38 4794 -21 4802
rect -38 -4802 -21 -4794
rect 21 4794 38 4802
rect 21 -4802 38 -4794
rect 78 4794 95 4802
rect 78 -4802 95 -4794
rect 137 4794 154 4802
rect 137 -4802 154 -4794
rect 194 4794 211 4802
rect 194 -4802 211 -4794
rect 253 4794 270 4802
rect 253 -4802 270 -4794
rect 310 4794 327 4802
rect 310 -4802 327 -4794
rect 369 4794 386 4802
rect 369 -4802 386 -4794
rect 426 4794 443 4802
rect 426 -4802 443 -4794
rect 485 4794 502 4802
rect 485 -4802 502 -4794
rect 542 4794 559 4802
rect 542 -4802 559 -4794
rect 601 4794 618 4802
rect 601 -4802 618 -4794
rect 658 4794 675 4802
rect 658 -4802 675 -4794
rect 717 4794 734 4802
rect 717 -4802 734 -4794
rect 774 4794 791 4802
rect 774 -4802 791 -4794
rect 833 4794 850 4802
rect 833 -4802 850 -4794
rect 890 4794 907 4802
rect 890 -4802 907 -4794
rect 949 4794 966 4802
rect 949 -4802 966 -4794
rect 1006 4794 1023 4802
rect 1006 -4802 1023 -4794
rect 1065 4794 1082 4802
rect 1065 -4802 1082 -4794
rect 1122 4794 1139 4802
rect 1122 -4802 1139 -4794
rect 1181 4794 1198 4802
rect 1181 -4802 1198 -4794
rect 1238 4794 1255 4802
rect 1238 -4802 1255 -4794
rect 1297 4794 1314 4802
rect 1297 -4802 1314 -4794
rect 1354 4794 1371 4802
rect 1354 -4802 1371 -4794
rect 1413 4794 1430 4802
rect 1413 -4802 1430 -4794
<< viali >>
rect -1430 -4794 -1413 4794
rect -1371 -4794 -1354 4794
rect -1314 -4794 -1297 4794
rect -1255 -4794 -1238 4794
rect -1198 -4794 -1181 4794
rect -1139 -4794 -1122 4794
rect -1082 -4794 -1065 4794
rect -1023 -4794 -1006 4794
rect -966 -4794 -949 4794
rect -907 -4794 -890 4794
rect -850 -4794 -833 4794
rect -791 -4794 -774 4794
rect -734 -4794 -717 4794
rect -675 -4794 -658 4794
rect -618 -4794 -601 4794
rect -559 -4794 -542 4794
rect -502 -4794 -485 4794
rect -443 -4794 -426 4794
rect -386 -4794 -369 4794
rect -327 -4794 -310 4794
rect -270 -4794 -253 4794
rect -211 -4794 -194 4794
rect -154 -4794 -137 4794
rect -95 -4794 -78 4794
rect -38 -4794 -21 4794
rect 21 -4794 38 4794
rect 78 -4794 95 4794
rect 137 -4794 154 4794
rect 194 -4794 211 4794
rect 253 -4794 270 4794
rect 310 -4794 327 4794
rect 369 -4794 386 4794
rect 426 -4794 443 4794
rect 485 -4794 502 4794
rect 542 -4794 559 4794
rect 601 -4794 618 4794
rect 658 -4794 675 4794
rect 717 -4794 734 4794
rect 774 -4794 791 4794
rect 833 -4794 850 4794
rect 890 -4794 907 4794
rect 949 -4794 966 4794
rect 1006 -4794 1023 4794
rect 1065 -4794 1082 4794
rect 1122 -4794 1139 4794
rect 1181 -4794 1198 4794
rect 1238 -4794 1255 4794
rect 1297 -4794 1314 4794
rect 1354 -4794 1371 4794
rect 1413 -4794 1430 4794
<< metal1 >>
rect -1433 4794 -1410 4800
rect -1433 -4794 -1430 4794
rect -1413 -4794 -1410 4794
rect -1433 -4800 -1410 -4794
rect -1374 4794 -1351 4800
rect -1374 -4794 -1371 4794
rect -1354 -4794 -1351 4794
rect -1374 -4800 -1351 -4794
rect -1317 4794 -1294 4800
rect -1317 -4794 -1314 4794
rect -1297 -4794 -1294 4794
rect -1317 -4800 -1294 -4794
rect -1258 4794 -1235 4800
rect -1258 -4794 -1255 4794
rect -1238 -4794 -1235 4794
rect -1258 -4800 -1235 -4794
rect -1201 4794 -1178 4800
rect -1201 -4794 -1198 4794
rect -1181 -4794 -1178 4794
rect -1201 -4800 -1178 -4794
rect -1142 4794 -1119 4800
rect -1142 -4794 -1139 4794
rect -1122 -4794 -1119 4794
rect -1142 -4800 -1119 -4794
rect -1085 4794 -1062 4800
rect -1085 -4794 -1082 4794
rect -1065 -4794 -1062 4794
rect -1085 -4800 -1062 -4794
rect -1026 4794 -1003 4800
rect -1026 -4794 -1023 4794
rect -1006 -4794 -1003 4794
rect -1026 -4800 -1003 -4794
rect -969 4794 -946 4800
rect -969 -4794 -966 4794
rect -949 -4794 -946 4794
rect -969 -4800 -946 -4794
rect -910 4794 -887 4800
rect -910 -4794 -907 4794
rect -890 -4794 -887 4794
rect -910 -4800 -887 -4794
rect -853 4794 -830 4800
rect -853 -4794 -850 4794
rect -833 -4794 -830 4794
rect -853 -4800 -830 -4794
rect -794 4794 -771 4800
rect -794 -4794 -791 4794
rect -774 -4794 -771 4794
rect -794 -4800 -771 -4794
rect -737 4794 -714 4800
rect -737 -4794 -734 4794
rect -717 -4794 -714 4794
rect -737 -4800 -714 -4794
rect -678 4794 -655 4800
rect -678 -4794 -675 4794
rect -658 -4794 -655 4794
rect -678 -4800 -655 -4794
rect -621 4794 -598 4800
rect -621 -4794 -618 4794
rect -601 -4794 -598 4794
rect -621 -4800 -598 -4794
rect -562 4794 -539 4800
rect -562 -4794 -559 4794
rect -542 -4794 -539 4794
rect -562 -4800 -539 -4794
rect -505 4794 -482 4800
rect -505 -4794 -502 4794
rect -485 -4794 -482 4794
rect -505 -4800 -482 -4794
rect -446 4794 -423 4800
rect -446 -4794 -443 4794
rect -426 -4794 -423 4794
rect -446 -4800 -423 -4794
rect -389 4794 -366 4800
rect -389 -4794 -386 4794
rect -369 -4794 -366 4794
rect -389 -4800 -366 -4794
rect -330 4794 -307 4800
rect -330 -4794 -327 4794
rect -310 -4794 -307 4794
rect -330 -4800 -307 -4794
rect -273 4794 -250 4800
rect -273 -4794 -270 4794
rect -253 -4794 -250 4794
rect -273 -4800 -250 -4794
rect -214 4794 -191 4800
rect -214 -4794 -211 4794
rect -194 -4794 -191 4794
rect -214 -4800 -191 -4794
rect -157 4794 -134 4800
rect -157 -4794 -154 4794
rect -137 -4794 -134 4794
rect -157 -4800 -134 -4794
rect -98 4794 -75 4800
rect -98 -4794 -95 4794
rect -78 -4794 -75 4794
rect -98 -4800 -75 -4794
rect -41 4794 -18 4800
rect -41 -4794 -38 4794
rect -21 -4794 -18 4794
rect -41 -4800 -18 -4794
rect 18 4794 41 4800
rect 18 -4794 21 4794
rect 38 -4794 41 4794
rect 18 -4800 41 -4794
rect 75 4794 98 4800
rect 75 -4794 78 4794
rect 95 -4794 98 4794
rect 75 -4800 98 -4794
rect 134 4794 157 4800
rect 134 -4794 137 4794
rect 154 -4794 157 4794
rect 134 -4800 157 -4794
rect 191 4794 214 4800
rect 191 -4794 194 4794
rect 211 -4794 214 4794
rect 191 -4800 214 -4794
rect 250 4794 273 4800
rect 250 -4794 253 4794
rect 270 -4794 273 4794
rect 250 -4800 273 -4794
rect 307 4794 330 4800
rect 307 -4794 310 4794
rect 327 -4794 330 4794
rect 307 -4800 330 -4794
rect 366 4794 389 4800
rect 366 -4794 369 4794
rect 386 -4794 389 4794
rect 366 -4800 389 -4794
rect 423 4794 446 4800
rect 423 -4794 426 4794
rect 443 -4794 446 4794
rect 423 -4800 446 -4794
rect 482 4794 505 4800
rect 482 -4794 485 4794
rect 502 -4794 505 4794
rect 482 -4800 505 -4794
rect 539 4794 562 4800
rect 539 -4794 542 4794
rect 559 -4794 562 4794
rect 539 -4800 562 -4794
rect 598 4794 621 4800
rect 598 -4794 601 4794
rect 618 -4794 621 4794
rect 598 -4800 621 -4794
rect 655 4794 678 4800
rect 655 -4794 658 4794
rect 675 -4794 678 4794
rect 655 -4800 678 -4794
rect 714 4794 737 4800
rect 714 -4794 717 4794
rect 734 -4794 737 4794
rect 714 -4800 737 -4794
rect 771 4794 794 4800
rect 771 -4794 774 4794
rect 791 -4794 794 4794
rect 771 -4800 794 -4794
rect 830 4794 853 4800
rect 830 -4794 833 4794
rect 850 -4794 853 4794
rect 830 -4800 853 -4794
rect 887 4794 910 4800
rect 887 -4794 890 4794
rect 907 -4794 910 4794
rect 887 -4800 910 -4794
rect 946 4794 969 4800
rect 946 -4794 949 4794
rect 966 -4794 969 4794
rect 946 -4800 969 -4794
rect 1003 4794 1026 4800
rect 1003 -4794 1006 4794
rect 1023 -4794 1026 4794
rect 1003 -4800 1026 -4794
rect 1062 4794 1085 4800
rect 1062 -4794 1065 4794
rect 1082 -4794 1085 4794
rect 1062 -4800 1085 -4794
rect 1119 4794 1142 4800
rect 1119 -4794 1122 4794
rect 1139 -4794 1142 4794
rect 1119 -4800 1142 -4794
rect 1178 4794 1201 4800
rect 1178 -4794 1181 4794
rect 1198 -4794 1201 4794
rect 1178 -4800 1201 -4794
rect 1235 4794 1258 4800
rect 1235 -4794 1238 4794
rect 1255 -4794 1258 4794
rect 1235 -4800 1258 -4794
rect 1294 4794 1317 4800
rect 1294 -4794 1297 4794
rect 1314 -4794 1317 4794
rect 1294 -4800 1317 -4794
rect 1351 4794 1374 4800
rect 1351 -4794 1354 4794
rect 1371 -4794 1374 4794
rect 1351 -4800 1374 -4794
rect 1410 4794 1433 4800
rect 1410 -4794 1413 4794
rect 1430 -4794 1433 4794
rect 1410 -4800 1433 -4794
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 96 l 0.3 m 1 nf 25 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
