magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -284 -157 284 95
<< nmos >>
rect -200 -131 200 69
<< ndiff >>
rect -258 54 -200 69
rect -258 20 -246 54
rect -212 20 -200 54
rect -258 -14 -200 20
rect -258 -48 -246 -14
rect -212 -48 -200 -14
rect -258 -82 -200 -48
rect -258 -116 -246 -82
rect -212 -116 -200 -82
rect -258 -131 -200 -116
rect 200 54 258 69
rect 200 20 212 54
rect 246 20 258 54
rect 200 -14 258 20
rect 200 -48 212 -14
rect 246 -48 258 -14
rect 200 -82 258 -48
rect 200 -116 212 -82
rect 246 -116 258 -82
rect 200 -131 258 -116
<< ndiffc >>
rect -246 20 -212 54
rect -246 -48 -212 -14
rect -246 -116 -212 -82
rect 212 20 246 54
rect 212 -48 246 -14
rect 212 -116 246 -82
<< poly >>
rect -200 141 200 157
rect -200 107 -153 141
rect -119 107 -85 141
rect -51 107 -17 141
rect 17 107 51 141
rect 85 107 119 141
rect 153 107 200 141
rect -200 69 200 107
rect -200 -157 200 -131
<< polycont >>
rect -153 107 -119 141
rect -85 107 -51 141
rect -17 107 17 141
rect 51 107 85 141
rect 119 107 153 141
<< locali >>
rect -200 107 -161 141
rect -119 107 -89 141
rect -51 107 -17 141
rect 17 107 51 141
rect 89 107 119 141
rect 161 107 200 141
rect -246 54 -212 73
rect -246 -14 -212 -12
rect -246 -50 -212 -48
rect -246 -135 -212 -116
rect 212 54 246 73
rect 212 -14 246 -12
rect 212 -50 246 -48
rect 212 -135 246 -116
<< viali >>
rect -161 107 -153 141
rect -153 107 -127 141
rect -89 107 -85 141
rect -85 107 -55 141
rect -17 107 17 141
rect 55 107 85 141
rect 85 107 89 141
rect 127 107 153 141
rect 153 107 161 141
rect -246 20 -212 22
rect -246 -12 -212 20
rect -246 -82 -212 -50
rect -246 -84 -212 -82
rect 212 20 246 22
rect 212 -12 246 20
rect 212 -82 246 -50
rect 212 -84 246 -82
<< metal1 >>
rect -196 141 196 147
rect -196 107 -161 141
rect -127 107 -89 141
rect -55 107 -17 141
rect 17 107 55 141
rect 89 107 127 141
rect 161 107 196 141
rect -196 101 196 107
rect -252 22 -206 69
rect -252 -12 -246 22
rect -212 -12 -206 22
rect -252 -50 -206 -12
rect -252 -84 -246 -50
rect -212 -84 -206 -50
rect -252 -131 -206 -84
rect 206 22 252 69
rect 206 -12 212 22
rect 246 -12 252 22
rect 206 -50 252 -12
rect 206 -84 212 -50
rect 246 -84 252 -50
rect 206 -131 252 -84
<< end >>
