magic
tech sky130A
magscale 1 2
timestamp 1666625676
<< error_p >>
rect -1466 45524 -1396 45668
rect -1148 45524 -1078 45668
rect -830 45524 -760 45668
rect -512 45524 -442 45668
rect -194 45524 -124 45668
rect 124 45524 194 45668
rect 442 45524 512 45668
rect 760 45524 830 45668
rect 1078 45524 1148 45668
rect 1396 45524 1466 45668
rect -1466 34156 -1396 34300
rect -1148 34156 -1078 34300
rect -830 34156 -760 34300
rect -512 34156 -442 34300
rect -194 34156 -124 34300
rect 124 34156 194 34300
rect 442 34156 512 34300
rect 760 34156 830 34300
rect 1078 34156 1148 34300
rect 1396 34156 1466 34300
rect -1466 22788 -1396 22932
rect -1148 22788 -1078 22932
rect -830 22788 -760 22932
rect -512 22788 -442 22932
rect -194 22788 -124 22932
rect 124 22788 194 22932
rect 442 22788 512 22932
rect 760 22788 830 22932
rect 1078 22788 1148 22932
rect 1396 22788 1466 22932
rect -1466 11420 -1396 11564
rect -1148 11420 -1078 11564
rect -830 11420 -760 11564
rect -512 11420 -442 11564
rect -194 11420 -124 11564
rect 124 11420 194 11564
rect 442 11420 512 11564
rect 760 11420 830 11564
rect 1078 11420 1148 11564
rect 1396 11420 1466 11564
rect -1466 52 -1396 196
rect -1148 52 -1078 196
rect -830 52 -760 196
rect -512 52 -442 196
rect -194 52 -124 196
rect 124 52 194 196
rect 442 52 512 196
rect 760 52 830 196
rect 1078 52 1148 196
rect 1396 52 1466 196
rect -1466 -11316 -1396 -11172
rect -1148 -11316 -1078 -11172
rect -830 -11316 -760 -11172
rect -512 -11316 -442 -11172
rect -194 -11316 -124 -11172
rect 124 -11316 194 -11172
rect 442 -11316 512 -11172
rect 760 -11316 830 -11172
rect 1078 -11316 1148 -11172
rect 1396 -11316 1466 -11172
rect -1466 -22684 -1396 -22540
rect -1148 -22684 -1078 -22540
rect -830 -22684 -760 -22540
rect -512 -22684 -442 -22540
rect -194 -22684 -124 -22540
rect 124 -22684 194 -22540
rect 442 -22684 512 -22540
rect 760 -22684 830 -22540
rect 1078 -22684 1148 -22540
rect 1396 -22684 1466 -22540
rect -1466 -34052 -1396 -33908
rect -1148 -34052 -1078 -33908
rect -830 -34052 -760 -33908
rect -512 -34052 -442 -33908
rect -194 -34052 -124 -33908
rect 124 -34052 194 -33908
rect 442 -34052 512 -33908
rect 760 -34052 830 -33908
rect 1078 -34052 1148 -33908
rect 1396 -34052 1466 -33908
rect -1466 -45420 -1396 -45276
rect -1148 -45420 -1078 -45276
rect -830 -45420 -760 -45276
rect -512 -45420 -442 -45276
rect -194 -45420 -124 -45276
rect 124 -45420 194 -45276
rect 442 -45420 512 -45276
rect 760 -45420 830 -45276
rect 1078 -45420 1148 -45276
rect 1396 -45420 1466 -45276
<< xpolycontact >>
rect -1466 56356 -1396 56788
rect -1466 45524 -1396 45956
rect -1148 56356 -1078 56788
rect -1148 45524 -1078 45956
rect -830 56356 -760 56788
rect -830 45524 -760 45956
rect -512 56356 -442 56788
rect -512 45524 -442 45956
rect -194 56356 -124 56788
rect -194 45524 -124 45956
rect 124 56356 194 56788
rect 124 45524 194 45956
rect 442 56356 512 56788
rect 442 45524 512 45956
rect 760 56356 830 56788
rect 760 45524 830 45956
rect 1078 56356 1148 56788
rect 1078 45524 1148 45956
rect 1396 56356 1466 56788
rect 1396 45524 1466 45956
rect -1466 44988 -1396 45420
rect -1466 34156 -1396 34588
rect -1148 44988 -1078 45420
rect -1148 34156 -1078 34588
rect -830 44988 -760 45420
rect -830 34156 -760 34588
rect -512 44988 -442 45420
rect -512 34156 -442 34588
rect -194 44988 -124 45420
rect -194 34156 -124 34588
rect 124 44988 194 45420
rect 124 34156 194 34588
rect 442 44988 512 45420
rect 442 34156 512 34588
rect 760 44988 830 45420
rect 760 34156 830 34588
rect 1078 44988 1148 45420
rect 1078 34156 1148 34588
rect 1396 44988 1466 45420
rect 1396 34156 1466 34588
rect -1466 33620 -1396 34052
rect -1466 22788 -1396 23220
rect -1148 33620 -1078 34052
rect -1148 22788 -1078 23220
rect -830 33620 -760 34052
rect -830 22788 -760 23220
rect -512 33620 -442 34052
rect -512 22788 -442 23220
rect -194 33620 -124 34052
rect -194 22788 -124 23220
rect 124 33620 194 34052
rect 124 22788 194 23220
rect 442 33620 512 34052
rect 442 22788 512 23220
rect 760 33620 830 34052
rect 760 22788 830 23220
rect 1078 33620 1148 34052
rect 1078 22788 1148 23220
rect 1396 33620 1466 34052
rect 1396 22788 1466 23220
rect -1466 22252 -1396 22684
rect -1466 11420 -1396 11852
rect -1148 22252 -1078 22684
rect -1148 11420 -1078 11852
rect -830 22252 -760 22684
rect -830 11420 -760 11852
rect -512 22252 -442 22684
rect -512 11420 -442 11852
rect -194 22252 -124 22684
rect -194 11420 -124 11852
rect 124 22252 194 22684
rect 124 11420 194 11852
rect 442 22252 512 22684
rect 442 11420 512 11852
rect 760 22252 830 22684
rect 760 11420 830 11852
rect 1078 22252 1148 22684
rect 1078 11420 1148 11852
rect 1396 22252 1466 22684
rect 1396 11420 1466 11852
rect -1466 10884 -1396 11316
rect -1466 52 -1396 484
rect -1148 10884 -1078 11316
rect -1148 52 -1078 484
rect -830 10884 -760 11316
rect -830 52 -760 484
rect -512 10884 -442 11316
rect -512 52 -442 484
rect -194 10884 -124 11316
rect -194 52 -124 484
rect 124 10884 194 11316
rect 124 52 194 484
rect 442 10884 512 11316
rect 442 52 512 484
rect 760 10884 830 11316
rect 760 52 830 484
rect 1078 10884 1148 11316
rect 1078 52 1148 484
rect 1396 10884 1466 11316
rect 1396 52 1466 484
rect -1466 -484 -1396 -52
rect -1466 -11316 -1396 -10884
rect -1148 -484 -1078 -52
rect -1148 -11316 -1078 -10884
rect -830 -484 -760 -52
rect -830 -11316 -760 -10884
rect -512 -484 -442 -52
rect -512 -11316 -442 -10884
rect -194 -484 -124 -52
rect -194 -11316 -124 -10884
rect 124 -484 194 -52
rect 124 -11316 194 -10884
rect 442 -484 512 -52
rect 442 -11316 512 -10884
rect 760 -484 830 -52
rect 760 -11316 830 -10884
rect 1078 -484 1148 -52
rect 1078 -11316 1148 -10884
rect 1396 -484 1466 -52
rect 1396 -11316 1466 -10884
rect -1466 -11852 -1396 -11420
rect -1466 -22684 -1396 -22252
rect -1148 -11852 -1078 -11420
rect -1148 -22684 -1078 -22252
rect -830 -11852 -760 -11420
rect -830 -22684 -760 -22252
rect -512 -11852 -442 -11420
rect -512 -22684 -442 -22252
rect -194 -11852 -124 -11420
rect -194 -22684 -124 -22252
rect 124 -11852 194 -11420
rect 124 -22684 194 -22252
rect 442 -11852 512 -11420
rect 442 -22684 512 -22252
rect 760 -11852 830 -11420
rect 760 -22684 830 -22252
rect 1078 -11852 1148 -11420
rect 1078 -22684 1148 -22252
rect 1396 -11852 1466 -11420
rect 1396 -22684 1466 -22252
rect -1466 -23220 -1396 -22788
rect -1466 -34052 -1396 -33620
rect -1148 -23220 -1078 -22788
rect -1148 -34052 -1078 -33620
rect -830 -23220 -760 -22788
rect -830 -34052 -760 -33620
rect -512 -23220 -442 -22788
rect -512 -34052 -442 -33620
rect -194 -23220 -124 -22788
rect -194 -34052 -124 -33620
rect 124 -23220 194 -22788
rect 124 -34052 194 -33620
rect 442 -23220 512 -22788
rect 442 -34052 512 -33620
rect 760 -23220 830 -22788
rect 760 -34052 830 -33620
rect 1078 -23220 1148 -22788
rect 1078 -34052 1148 -33620
rect 1396 -23220 1466 -22788
rect 1396 -34052 1466 -33620
rect -1466 -34588 -1396 -34156
rect -1466 -45420 -1396 -44988
rect -1148 -34588 -1078 -34156
rect -1148 -45420 -1078 -44988
rect -830 -34588 -760 -34156
rect -830 -45420 -760 -44988
rect -512 -34588 -442 -34156
rect -512 -45420 -442 -44988
rect -194 -34588 -124 -34156
rect -194 -45420 -124 -44988
rect 124 -34588 194 -34156
rect 124 -45420 194 -44988
rect 442 -34588 512 -34156
rect 442 -45420 512 -44988
rect 760 -34588 830 -34156
rect 760 -45420 830 -44988
rect 1078 -34588 1148 -34156
rect 1078 -45420 1148 -44988
rect 1396 -34588 1466 -34156
rect 1396 -45420 1466 -44988
rect -1466 -45956 -1396 -45524
rect -1466 -56788 -1396 -56356
rect -1148 -45956 -1078 -45524
rect -1148 -56788 -1078 -56356
rect -830 -45956 -760 -45524
rect -830 -56788 -760 -56356
rect -512 -45956 -442 -45524
rect -512 -56788 -442 -56356
rect -194 -45956 -124 -45524
rect -194 -56788 -124 -56356
rect 124 -45956 194 -45524
rect 124 -56788 194 -56356
rect 442 -45956 512 -45524
rect 442 -56788 512 -56356
rect 760 -45956 830 -45524
rect 760 -56788 830 -56356
rect 1078 -45956 1148 -45524
rect 1078 -56788 1148 -56356
rect 1396 -45956 1466 -45524
rect 1396 -56788 1466 -56356
<< xpolyres >>
rect -1466 45956 -1396 56356
rect -1148 45956 -1078 56356
rect -830 45956 -760 56356
rect -512 45956 -442 56356
rect -194 45956 -124 56356
rect 124 45956 194 56356
rect 442 45956 512 56356
rect 760 45956 830 56356
rect 1078 45956 1148 56356
rect 1396 45956 1466 56356
rect -1466 34588 -1396 44988
rect -1148 34588 -1078 44988
rect -830 34588 -760 44988
rect -512 34588 -442 44988
rect -194 34588 -124 44988
rect 124 34588 194 44988
rect 442 34588 512 44988
rect 760 34588 830 44988
rect 1078 34588 1148 44988
rect 1396 34588 1466 44988
rect -1466 23220 -1396 33620
rect -1148 23220 -1078 33620
rect -830 23220 -760 33620
rect -512 23220 -442 33620
rect -194 23220 -124 33620
rect 124 23220 194 33620
rect 442 23220 512 33620
rect 760 23220 830 33620
rect 1078 23220 1148 33620
rect 1396 23220 1466 33620
rect -1466 11852 -1396 22252
rect -1148 11852 -1078 22252
rect -830 11852 -760 22252
rect -512 11852 -442 22252
rect -194 11852 -124 22252
rect 124 11852 194 22252
rect 442 11852 512 22252
rect 760 11852 830 22252
rect 1078 11852 1148 22252
rect 1396 11852 1466 22252
rect -1466 484 -1396 10884
rect -1148 484 -1078 10884
rect -830 484 -760 10884
rect -512 484 -442 10884
rect -194 484 -124 10884
rect 124 484 194 10884
rect 442 484 512 10884
rect 760 484 830 10884
rect 1078 484 1148 10884
rect 1396 484 1466 10884
rect -1466 -10884 -1396 -484
rect -1148 -10884 -1078 -484
rect -830 -10884 -760 -484
rect -512 -10884 -442 -484
rect -194 -10884 -124 -484
rect 124 -10884 194 -484
rect 442 -10884 512 -484
rect 760 -10884 830 -484
rect 1078 -10884 1148 -484
rect 1396 -10884 1466 -484
rect -1466 -22252 -1396 -11852
rect -1148 -22252 -1078 -11852
rect -830 -22252 -760 -11852
rect -512 -22252 -442 -11852
rect -194 -22252 -124 -11852
rect 124 -22252 194 -11852
rect 442 -22252 512 -11852
rect 760 -22252 830 -11852
rect 1078 -22252 1148 -11852
rect 1396 -22252 1466 -11852
rect -1466 -33620 -1396 -23220
rect -1148 -33620 -1078 -23220
rect -830 -33620 -760 -23220
rect -512 -33620 -442 -23220
rect -194 -33620 -124 -23220
rect 124 -33620 194 -23220
rect 442 -33620 512 -23220
rect 760 -33620 830 -23220
rect 1078 -33620 1148 -23220
rect 1396 -33620 1466 -23220
rect -1466 -44988 -1396 -34588
rect -1148 -44988 -1078 -34588
rect -830 -44988 -760 -34588
rect -512 -44988 -442 -34588
rect -194 -44988 -124 -34588
rect 124 -44988 194 -34588
rect 442 -44988 512 -34588
rect 760 -44988 830 -34588
rect 1078 -44988 1148 -34588
rect 1396 -44988 1466 -34588
rect -1466 -56356 -1396 -45956
rect -1148 -56356 -1078 -45956
rect -830 -56356 -760 -45956
rect -512 -56356 -442 -45956
rect -194 -56356 -124 -45956
rect 124 -56356 194 -45956
rect 442 -56356 512 -45956
rect 760 -56356 830 -45956
rect 1078 -56356 1148 -45956
rect 1396 -56356 1466 -45956
<< viali >>
rect -1450 56373 -1412 56770
rect -1132 56373 -1094 56770
rect -814 56373 -776 56770
rect -496 56373 -458 56770
rect -178 56373 -140 56770
rect 140 56373 178 56770
rect 458 56373 496 56770
rect 776 56373 814 56770
rect 1094 56373 1132 56770
rect 1412 56373 1450 56770
rect -1450 45542 -1412 45939
rect -1132 45542 -1094 45939
rect -814 45542 -776 45939
rect -496 45542 -458 45939
rect -178 45542 -140 45939
rect 140 45542 178 45939
rect 458 45542 496 45939
rect 776 45542 814 45939
rect 1094 45542 1132 45939
rect 1412 45542 1450 45939
rect -1450 45005 -1412 45402
rect -1132 45005 -1094 45402
rect -814 45005 -776 45402
rect -496 45005 -458 45402
rect -178 45005 -140 45402
rect 140 45005 178 45402
rect 458 45005 496 45402
rect 776 45005 814 45402
rect 1094 45005 1132 45402
rect 1412 45005 1450 45402
rect -1450 34174 -1412 34571
rect -1132 34174 -1094 34571
rect -814 34174 -776 34571
rect -496 34174 -458 34571
rect -178 34174 -140 34571
rect 140 34174 178 34571
rect 458 34174 496 34571
rect 776 34174 814 34571
rect 1094 34174 1132 34571
rect 1412 34174 1450 34571
rect -1450 33637 -1412 34034
rect -1132 33637 -1094 34034
rect -814 33637 -776 34034
rect -496 33637 -458 34034
rect -178 33637 -140 34034
rect 140 33637 178 34034
rect 458 33637 496 34034
rect 776 33637 814 34034
rect 1094 33637 1132 34034
rect 1412 33637 1450 34034
rect -1450 22806 -1412 23203
rect -1132 22806 -1094 23203
rect -814 22806 -776 23203
rect -496 22806 -458 23203
rect -178 22806 -140 23203
rect 140 22806 178 23203
rect 458 22806 496 23203
rect 776 22806 814 23203
rect 1094 22806 1132 23203
rect 1412 22806 1450 23203
rect -1450 22269 -1412 22666
rect -1132 22269 -1094 22666
rect -814 22269 -776 22666
rect -496 22269 -458 22666
rect -178 22269 -140 22666
rect 140 22269 178 22666
rect 458 22269 496 22666
rect 776 22269 814 22666
rect 1094 22269 1132 22666
rect 1412 22269 1450 22666
rect -1450 11438 -1412 11835
rect -1132 11438 -1094 11835
rect -814 11438 -776 11835
rect -496 11438 -458 11835
rect -178 11438 -140 11835
rect 140 11438 178 11835
rect 458 11438 496 11835
rect 776 11438 814 11835
rect 1094 11438 1132 11835
rect 1412 11438 1450 11835
rect -1450 10901 -1412 11298
rect -1132 10901 -1094 11298
rect -814 10901 -776 11298
rect -496 10901 -458 11298
rect -178 10901 -140 11298
rect 140 10901 178 11298
rect 458 10901 496 11298
rect 776 10901 814 11298
rect 1094 10901 1132 11298
rect 1412 10901 1450 11298
rect -1450 70 -1412 467
rect -1132 70 -1094 467
rect -814 70 -776 467
rect -496 70 -458 467
rect -178 70 -140 467
rect 140 70 178 467
rect 458 70 496 467
rect 776 70 814 467
rect 1094 70 1132 467
rect 1412 70 1450 467
rect -1450 -467 -1412 -70
rect -1132 -467 -1094 -70
rect -814 -467 -776 -70
rect -496 -467 -458 -70
rect -178 -467 -140 -70
rect 140 -467 178 -70
rect 458 -467 496 -70
rect 776 -467 814 -70
rect 1094 -467 1132 -70
rect 1412 -467 1450 -70
rect -1450 -11298 -1412 -10901
rect -1132 -11298 -1094 -10901
rect -814 -11298 -776 -10901
rect -496 -11298 -458 -10901
rect -178 -11298 -140 -10901
rect 140 -11298 178 -10901
rect 458 -11298 496 -10901
rect 776 -11298 814 -10901
rect 1094 -11298 1132 -10901
rect 1412 -11298 1450 -10901
rect -1450 -11835 -1412 -11438
rect -1132 -11835 -1094 -11438
rect -814 -11835 -776 -11438
rect -496 -11835 -458 -11438
rect -178 -11835 -140 -11438
rect 140 -11835 178 -11438
rect 458 -11835 496 -11438
rect 776 -11835 814 -11438
rect 1094 -11835 1132 -11438
rect 1412 -11835 1450 -11438
rect -1450 -22666 -1412 -22269
rect -1132 -22666 -1094 -22269
rect -814 -22666 -776 -22269
rect -496 -22666 -458 -22269
rect -178 -22666 -140 -22269
rect 140 -22666 178 -22269
rect 458 -22666 496 -22269
rect 776 -22666 814 -22269
rect 1094 -22666 1132 -22269
rect 1412 -22666 1450 -22269
rect -1450 -23203 -1412 -22806
rect -1132 -23203 -1094 -22806
rect -814 -23203 -776 -22806
rect -496 -23203 -458 -22806
rect -178 -23203 -140 -22806
rect 140 -23203 178 -22806
rect 458 -23203 496 -22806
rect 776 -23203 814 -22806
rect 1094 -23203 1132 -22806
rect 1412 -23203 1450 -22806
rect -1450 -34034 -1412 -33637
rect -1132 -34034 -1094 -33637
rect -814 -34034 -776 -33637
rect -496 -34034 -458 -33637
rect -178 -34034 -140 -33637
rect 140 -34034 178 -33637
rect 458 -34034 496 -33637
rect 776 -34034 814 -33637
rect 1094 -34034 1132 -33637
rect 1412 -34034 1450 -33637
rect -1450 -34571 -1412 -34174
rect -1132 -34571 -1094 -34174
rect -814 -34571 -776 -34174
rect -496 -34571 -458 -34174
rect -178 -34571 -140 -34174
rect 140 -34571 178 -34174
rect 458 -34571 496 -34174
rect 776 -34571 814 -34174
rect 1094 -34571 1132 -34174
rect 1412 -34571 1450 -34174
rect -1450 -45402 -1412 -45005
rect -1132 -45402 -1094 -45005
rect -814 -45402 -776 -45005
rect -496 -45402 -458 -45005
rect -178 -45402 -140 -45005
rect 140 -45402 178 -45005
rect 458 -45402 496 -45005
rect 776 -45402 814 -45005
rect 1094 -45402 1132 -45005
rect 1412 -45402 1450 -45005
rect -1450 -45939 -1412 -45542
rect -1132 -45939 -1094 -45542
rect -814 -45939 -776 -45542
rect -496 -45939 -458 -45542
rect -178 -45939 -140 -45542
rect 140 -45939 178 -45542
rect 458 -45939 496 -45542
rect 776 -45939 814 -45542
rect 1094 -45939 1132 -45542
rect 1412 -45939 1450 -45542
rect -1450 -56770 -1412 -56373
rect -1132 -56770 -1094 -56373
rect -814 -56770 -776 -56373
rect -496 -56770 -458 -56373
rect -178 -56770 -140 -56373
rect 140 -56770 178 -56373
rect 458 -56770 496 -56373
rect 776 -56770 814 -56373
rect 1094 -56770 1132 -56373
rect 1412 -56770 1450 -56373
<< metal1 >>
rect -1456 56770 -1406 56782
rect -1456 56373 -1450 56770
rect -1412 56373 -1406 56770
rect -1456 56361 -1406 56373
rect -1138 56770 -1088 56782
rect -1138 56373 -1132 56770
rect -1094 56373 -1088 56770
rect -1138 56361 -1088 56373
rect -820 56770 -770 56782
rect -820 56373 -814 56770
rect -776 56373 -770 56770
rect -820 56361 -770 56373
rect -502 56770 -452 56782
rect -502 56373 -496 56770
rect -458 56373 -452 56770
rect -502 56361 -452 56373
rect -184 56770 -134 56782
rect -184 56373 -178 56770
rect -140 56373 -134 56770
rect -184 56361 -134 56373
rect 134 56770 184 56782
rect 134 56373 140 56770
rect 178 56373 184 56770
rect 134 56361 184 56373
rect 452 56770 502 56782
rect 452 56373 458 56770
rect 496 56373 502 56770
rect 452 56361 502 56373
rect 770 56770 820 56782
rect 770 56373 776 56770
rect 814 56373 820 56770
rect 770 56361 820 56373
rect 1088 56770 1138 56782
rect 1088 56373 1094 56770
rect 1132 56373 1138 56770
rect 1088 56361 1138 56373
rect 1406 56770 1456 56782
rect 1406 56373 1412 56770
rect 1450 56373 1456 56770
rect 1406 56361 1456 56373
rect -1456 45939 -1406 45951
rect -1456 45542 -1450 45939
rect -1412 45542 -1406 45939
rect -1456 45530 -1406 45542
rect -1138 45939 -1088 45951
rect -1138 45542 -1132 45939
rect -1094 45542 -1088 45939
rect -1138 45530 -1088 45542
rect -820 45939 -770 45951
rect -820 45542 -814 45939
rect -776 45542 -770 45939
rect -820 45530 -770 45542
rect -502 45939 -452 45951
rect -502 45542 -496 45939
rect -458 45542 -452 45939
rect -502 45530 -452 45542
rect -184 45939 -134 45951
rect -184 45542 -178 45939
rect -140 45542 -134 45939
rect -184 45530 -134 45542
rect 134 45939 184 45951
rect 134 45542 140 45939
rect 178 45542 184 45939
rect 134 45530 184 45542
rect 452 45939 502 45951
rect 452 45542 458 45939
rect 496 45542 502 45939
rect 452 45530 502 45542
rect 770 45939 820 45951
rect 770 45542 776 45939
rect 814 45542 820 45939
rect 770 45530 820 45542
rect 1088 45939 1138 45951
rect 1088 45542 1094 45939
rect 1132 45542 1138 45939
rect 1088 45530 1138 45542
rect 1406 45939 1456 45951
rect 1406 45542 1412 45939
rect 1450 45542 1456 45939
rect 1406 45530 1456 45542
rect -1456 45402 -1406 45414
rect -1456 45005 -1450 45402
rect -1412 45005 -1406 45402
rect -1456 44993 -1406 45005
rect -1138 45402 -1088 45414
rect -1138 45005 -1132 45402
rect -1094 45005 -1088 45402
rect -1138 44993 -1088 45005
rect -820 45402 -770 45414
rect -820 45005 -814 45402
rect -776 45005 -770 45402
rect -820 44993 -770 45005
rect -502 45402 -452 45414
rect -502 45005 -496 45402
rect -458 45005 -452 45402
rect -502 44993 -452 45005
rect -184 45402 -134 45414
rect -184 45005 -178 45402
rect -140 45005 -134 45402
rect -184 44993 -134 45005
rect 134 45402 184 45414
rect 134 45005 140 45402
rect 178 45005 184 45402
rect 134 44993 184 45005
rect 452 45402 502 45414
rect 452 45005 458 45402
rect 496 45005 502 45402
rect 452 44993 502 45005
rect 770 45402 820 45414
rect 770 45005 776 45402
rect 814 45005 820 45402
rect 770 44993 820 45005
rect 1088 45402 1138 45414
rect 1088 45005 1094 45402
rect 1132 45005 1138 45402
rect 1088 44993 1138 45005
rect 1406 45402 1456 45414
rect 1406 45005 1412 45402
rect 1450 45005 1456 45402
rect 1406 44993 1456 45005
rect -1456 34571 -1406 34583
rect -1456 34174 -1450 34571
rect -1412 34174 -1406 34571
rect -1456 34162 -1406 34174
rect -1138 34571 -1088 34583
rect -1138 34174 -1132 34571
rect -1094 34174 -1088 34571
rect -1138 34162 -1088 34174
rect -820 34571 -770 34583
rect -820 34174 -814 34571
rect -776 34174 -770 34571
rect -820 34162 -770 34174
rect -502 34571 -452 34583
rect -502 34174 -496 34571
rect -458 34174 -452 34571
rect -502 34162 -452 34174
rect -184 34571 -134 34583
rect -184 34174 -178 34571
rect -140 34174 -134 34571
rect -184 34162 -134 34174
rect 134 34571 184 34583
rect 134 34174 140 34571
rect 178 34174 184 34571
rect 134 34162 184 34174
rect 452 34571 502 34583
rect 452 34174 458 34571
rect 496 34174 502 34571
rect 452 34162 502 34174
rect 770 34571 820 34583
rect 770 34174 776 34571
rect 814 34174 820 34571
rect 770 34162 820 34174
rect 1088 34571 1138 34583
rect 1088 34174 1094 34571
rect 1132 34174 1138 34571
rect 1088 34162 1138 34174
rect 1406 34571 1456 34583
rect 1406 34174 1412 34571
rect 1450 34174 1456 34571
rect 1406 34162 1456 34174
rect -1456 34034 -1406 34046
rect -1456 33637 -1450 34034
rect -1412 33637 -1406 34034
rect -1456 33625 -1406 33637
rect -1138 34034 -1088 34046
rect -1138 33637 -1132 34034
rect -1094 33637 -1088 34034
rect -1138 33625 -1088 33637
rect -820 34034 -770 34046
rect -820 33637 -814 34034
rect -776 33637 -770 34034
rect -820 33625 -770 33637
rect -502 34034 -452 34046
rect -502 33637 -496 34034
rect -458 33637 -452 34034
rect -502 33625 -452 33637
rect -184 34034 -134 34046
rect -184 33637 -178 34034
rect -140 33637 -134 34034
rect -184 33625 -134 33637
rect 134 34034 184 34046
rect 134 33637 140 34034
rect 178 33637 184 34034
rect 134 33625 184 33637
rect 452 34034 502 34046
rect 452 33637 458 34034
rect 496 33637 502 34034
rect 452 33625 502 33637
rect 770 34034 820 34046
rect 770 33637 776 34034
rect 814 33637 820 34034
rect 770 33625 820 33637
rect 1088 34034 1138 34046
rect 1088 33637 1094 34034
rect 1132 33637 1138 34034
rect 1088 33625 1138 33637
rect 1406 34034 1456 34046
rect 1406 33637 1412 34034
rect 1450 33637 1456 34034
rect 1406 33625 1456 33637
rect -1456 23203 -1406 23215
rect -1456 22806 -1450 23203
rect -1412 22806 -1406 23203
rect -1456 22794 -1406 22806
rect -1138 23203 -1088 23215
rect -1138 22806 -1132 23203
rect -1094 22806 -1088 23203
rect -1138 22794 -1088 22806
rect -820 23203 -770 23215
rect -820 22806 -814 23203
rect -776 22806 -770 23203
rect -820 22794 -770 22806
rect -502 23203 -452 23215
rect -502 22806 -496 23203
rect -458 22806 -452 23203
rect -502 22794 -452 22806
rect -184 23203 -134 23215
rect -184 22806 -178 23203
rect -140 22806 -134 23203
rect -184 22794 -134 22806
rect 134 23203 184 23215
rect 134 22806 140 23203
rect 178 22806 184 23203
rect 134 22794 184 22806
rect 452 23203 502 23215
rect 452 22806 458 23203
rect 496 22806 502 23203
rect 452 22794 502 22806
rect 770 23203 820 23215
rect 770 22806 776 23203
rect 814 22806 820 23203
rect 770 22794 820 22806
rect 1088 23203 1138 23215
rect 1088 22806 1094 23203
rect 1132 22806 1138 23203
rect 1088 22794 1138 22806
rect 1406 23203 1456 23215
rect 1406 22806 1412 23203
rect 1450 22806 1456 23203
rect 1406 22794 1456 22806
rect -1456 22666 -1406 22678
rect -1456 22269 -1450 22666
rect -1412 22269 -1406 22666
rect -1456 22257 -1406 22269
rect -1138 22666 -1088 22678
rect -1138 22269 -1132 22666
rect -1094 22269 -1088 22666
rect -1138 22257 -1088 22269
rect -820 22666 -770 22678
rect -820 22269 -814 22666
rect -776 22269 -770 22666
rect -820 22257 -770 22269
rect -502 22666 -452 22678
rect -502 22269 -496 22666
rect -458 22269 -452 22666
rect -502 22257 -452 22269
rect -184 22666 -134 22678
rect -184 22269 -178 22666
rect -140 22269 -134 22666
rect -184 22257 -134 22269
rect 134 22666 184 22678
rect 134 22269 140 22666
rect 178 22269 184 22666
rect 134 22257 184 22269
rect 452 22666 502 22678
rect 452 22269 458 22666
rect 496 22269 502 22666
rect 452 22257 502 22269
rect 770 22666 820 22678
rect 770 22269 776 22666
rect 814 22269 820 22666
rect 770 22257 820 22269
rect 1088 22666 1138 22678
rect 1088 22269 1094 22666
rect 1132 22269 1138 22666
rect 1088 22257 1138 22269
rect 1406 22666 1456 22678
rect 1406 22269 1412 22666
rect 1450 22269 1456 22666
rect 1406 22257 1456 22269
rect -1456 11835 -1406 11847
rect -1456 11438 -1450 11835
rect -1412 11438 -1406 11835
rect -1456 11426 -1406 11438
rect -1138 11835 -1088 11847
rect -1138 11438 -1132 11835
rect -1094 11438 -1088 11835
rect -1138 11426 -1088 11438
rect -820 11835 -770 11847
rect -820 11438 -814 11835
rect -776 11438 -770 11835
rect -820 11426 -770 11438
rect -502 11835 -452 11847
rect -502 11438 -496 11835
rect -458 11438 -452 11835
rect -502 11426 -452 11438
rect -184 11835 -134 11847
rect -184 11438 -178 11835
rect -140 11438 -134 11835
rect -184 11426 -134 11438
rect 134 11835 184 11847
rect 134 11438 140 11835
rect 178 11438 184 11835
rect 134 11426 184 11438
rect 452 11835 502 11847
rect 452 11438 458 11835
rect 496 11438 502 11835
rect 452 11426 502 11438
rect 770 11835 820 11847
rect 770 11438 776 11835
rect 814 11438 820 11835
rect 770 11426 820 11438
rect 1088 11835 1138 11847
rect 1088 11438 1094 11835
rect 1132 11438 1138 11835
rect 1088 11426 1138 11438
rect 1406 11835 1456 11847
rect 1406 11438 1412 11835
rect 1450 11438 1456 11835
rect 1406 11426 1456 11438
rect -1456 11298 -1406 11310
rect -1456 10901 -1450 11298
rect -1412 10901 -1406 11298
rect -1456 10889 -1406 10901
rect -1138 11298 -1088 11310
rect -1138 10901 -1132 11298
rect -1094 10901 -1088 11298
rect -1138 10889 -1088 10901
rect -820 11298 -770 11310
rect -820 10901 -814 11298
rect -776 10901 -770 11298
rect -820 10889 -770 10901
rect -502 11298 -452 11310
rect -502 10901 -496 11298
rect -458 10901 -452 11298
rect -502 10889 -452 10901
rect -184 11298 -134 11310
rect -184 10901 -178 11298
rect -140 10901 -134 11298
rect -184 10889 -134 10901
rect 134 11298 184 11310
rect 134 10901 140 11298
rect 178 10901 184 11298
rect 134 10889 184 10901
rect 452 11298 502 11310
rect 452 10901 458 11298
rect 496 10901 502 11298
rect 452 10889 502 10901
rect 770 11298 820 11310
rect 770 10901 776 11298
rect 814 10901 820 11298
rect 770 10889 820 10901
rect 1088 11298 1138 11310
rect 1088 10901 1094 11298
rect 1132 10901 1138 11298
rect 1088 10889 1138 10901
rect 1406 11298 1456 11310
rect 1406 10901 1412 11298
rect 1450 10901 1456 11298
rect 1406 10889 1456 10901
rect -1456 467 -1406 479
rect -1456 70 -1450 467
rect -1412 70 -1406 467
rect -1456 58 -1406 70
rect -1138 467 -1088 479
rect -1138 70 -1132 467
rect -1094 70 -1088 467
rect -1138 58 -1088 70
rect -820 467 -770 479
rect -820 70 -814 467
rect -776 70 -770 467
rect -820 58 -770 70
rect -502 467 -452 479
rect -502 70 -496 467
rect -458 70 -452 467
rect -502 58 -452 70
rect -184 467 -134 479
rect -184 70 -178 467
rect -140 70 -134 467
rect -184 58 -134 70
rect 134 467 184 479
rect 134 70 140 467
rect 178 70 184 467
rect 134 58 184 70
rect 452 467 502 479
rect 452 70 458 467
rect 496 70 502 467
rect 452 58 502 70
rect 770 467 820 479
rect 770 70 776 467
rect 814 70 820 467
rect 770 58 820 70
rect 1088 467 1138 479
rect 1088 70 1094 467
rect 1132 70 1138 467
rect 1088 58 1138 70
rect 1406 467 1456 479
rect 1406 70 1412 467
rect 1450 70 1456 467
rect 1406 58 1456 70
rect -1456 -70 -1406 -58
rect -1456 -467 -1450 -70
rect -1412 -467 -1406 -70
rect -1456 -479 -1406 -467
rect -1138 -70 -1088 -58
rect -1138 -467 -1132 -70
rect -1094 -467 -1088 -70
rect -1138 -479 -1088 -467
rect -820 -70 -770 -58
rect -820 -467 -814 -70
rect -776 -467 -770 -70
rect -820 -479 -770 -467
rect -502 -70 -452 -58
rect -502 -467 -496 -70
rect -458 -467 -452 -70
rect -502 -479 -452 -467
rect -184 -70 -134 -58
rect -184 -467 -178 -70
rect -140 -467 -134 -70
rect -184 -479 -134 -467
rect 134 -70 184 -58
rect 134 -467 140 -70
rect 178 -467 184 -70
rect 134 -479 184 -467
rect 452 -70 502 -58
rect 452 -467 458 -70
rect 496 -467 502 -70
rect 452 -479 502 -467
rect 770 -70 820 -58
rect 770 -467 776 -70
rect 814 -467 820 -70
rect 770 -479 820 -467
rect 1088 -70 1138 -58
rect 1088 -467 1094 -70
rect 1132 -467 1138 -70
rect 1088 -479 1138 -467
rect 1406 -70 1456 -58
rect 1406 -467 1412 -70
rect 1450 -467 1456 -70
rect 1406 -479 1456 -467
rect -1456 -10901 -1406 -10889
rect -1456 -11298 -1450 -10901
rect -1412 -11298 -1406 -10901
rect -1456 -11310 -1406 -11298
rect -1138 -10901 -1088 -10889
rect -1138 -11298 -1132 -10901
rect -1094 -11298 -1088 -10901
rect -1138 -11310 -1088 -11298
rect -820 -10901 -770 -10889
rect -820 -11298 -814 -10901
rect -776 -11298 -770 -10901
rect -820 -11310 -770 -11298
rect -502 -10901 -452 -10889
rect -502 -11298 -496 -10901
rect -458 -11298 -452 -10901
rect -502 -11310 -452 -11298
rect -184 -10901 -134 -10889
rect -184 -11298 -178 -10901
rect -140 -11298 -134 -10901
rect -184 -11310 -134 -11298
rect 134 -10901 184 -10889
rect 134 -11298 140 -10901
rect 178 -11298 184 -10901
rect 134 -11310 184 -11298
rect 452 -10901 502 -10889
rect 452 -11298 458 -10901
rect 496 -11298 502 -10901
rect 452 -11310 502 -11298
rect 770 -10901 820 -10889
rect 770 -11298 776 -10901
rect 814 -11298 820 -10901
rect 770 -11310 820 -11298
rect 1088 -10901 1138 -10889
rect 1088 -11298 1094 -10901
rect 1132 -11298 1138 -10901
rect 1088 -11310 1138 -11298
rect 1406 -10901 1456 -10889
rect 1406 -11298 1412 -10901
rect 1450 -11298 1456 -10901
rect 1406 -11310 1456 -11298
rect -1456 -11438 -1406 -11426
rect -1456 -11835 -1450 -11438
rect -1412 -11835 -1406 -11438
rect -1456 -11847 -1406 -11835
rect -1138 -11438 -1088 -11426
rect -1138 -11835 -1132 -11438
rect -1094 -11835 -1088 -11438
rect -1138 -11847 -1088 -11835
rect -820 -11438 -770 -11426
rect -820 -11835 -814 -11438
rect -776 -11835 -770 -11438
rect -820 -11847 -770 -11835
rect -502 -11438 -452 -11426
rect -502 -11835 -496 -11438
rect -458 -11835 -452 -11438
rect -502 -11847 -452 -11835
rect -184 -11438 -134 -11426
rect -184 -11835 -178 -11438
rect -140 -11835 -134 -11438
rect -184 -11847 -134 -11835
rect 134 -11438 184 -11426
rect 134 -11835 140 -11438
rect 178 -11835 184 -11438
rect 134 -11847 184 -11835
rect 452 -11438 502 -11426
rect 452 -11835 458 -11438
rect 496 -11835 502 -11438
rect 452 -11847 502 -11835
rect 770 -11438 820 -11426
rect 770 -11835 776 -11438
rect 814 -11835 820 -11438
rect 770 -11847 820 -11835
rect 1088 -11438 1138 -11426
rect 1088 -11835 1094 -11438
rect 1132 -11835 1138 -11438
rect 1088 -11847 1138 -11835
rect 1406 -11438 1456 -11426
rect 1406 -11835 1412 -11438
rect 1450 -11835 1456 -11438
rect 1406 -11847 1456 -11835
rect -1456 -22269 -1406 -22257
rect -1456 -22666 -1450 -22269
rect -1412 -22666 -1406 -22269
rect -1456 -22678 -1406 -22666
rect -1138 -22269 -1088 -22257
rect -1138 -22666 -1132 -22269
rect -1094 -22666 -1088 -22269
rect -1138 -22678 -1088 -22666
rect -820 -22269 -770 -22257
rect -820 -22666 -814 -22269
rect -776 -22666 -770 -22269
rect -820 -22678 -770 -22666
rect -502 -22269 -452 -22257
rect -502 -22666 -496 -22269
rect -458 -22666 -452 -22269
rect -502 -22678 -452 -22666
rect -184 -22269 -134 -22257
rect -184 -22666 -178 -22269
rect -140 -22666 -134 -22269
rect -184 -22678 -134 -22666
rect 134 -22269 184 -22257
rect 134 -22666 140 -22269
rect 178 -22666 184 -22269
rect 134 -22678 184 -22666
rect 452 -22269 502 -22257
rect 452 -22666 458 -22269
rect 496 -22666 502 -22269
rect 452 -22678 502 -22666
rect 770 -22269 820 -22257
rect 770 -22666 776 -22269
rect 814 -22666 820 -22269
rect 770 -22678 820 -22666
rect 1088 -22269 1138 -22257
rect 1088 -22666 1094 -22269
rect 1132 -22666 1138 -22269
rect 1088 -22678 1138 -22666
rect 1406 -22269 1456 -22257
rect 1406 -22666 1412 -22269
rect 1450 -22666 1456 -22269
rect 1406 -22678 1456 -22666
rect -1456 -22806 -1406 -22794
rect -1456 -23203 -1450 -22806
rect -1412 -23203 -1406 -22806
rect -1456 -23215 -1406 -23203
rect -1138 -22806 -1088 -22794
rect -1138 -23203 -1132 -22806
rect -1094 -23203 -1088 -22806
rect -1138 -23215 -1088 -23203
rect -820 -22806 -770 -22794
rect -820 -23203 -814 -22806
rect -776 -23203 -770 -22806
rect -820 -23215 -770 -23203
rect -502 -22806 -452 -22794
rect -502 -23203 -496 -22806
rect -458 -23203 -452 -22806
rect -502 -23215 -452 -23203
rect -184 -22806 -134 -22794
rect -184 -23203 -178 -22806
rect -140 -23203 -134 -22806
rect -184 -23215 -134 -23203
rect 134 -22806 184 -22794
rect 134 -23203 140 -22806
rect 178 -23203 184 -22806
rect 134 -23215 184 -23203
rect 452 -22806 502 -22794
rect 452 -23203 458 -22806
rect 496 -23203 502 -22806
rect 452 -23215 502 -23203
rect 770 -22806 820 -22794
rect 770 -23203 776 -22806
rect 814 -23203 820 -22806
rect 770 -23215 820 -23203
rect 1088 -22806 1138 -22794
rect 1088 -23203 1094 -22806
rect 1132 -23203 1138 -22806
rect 1088 -23215 1138 -23203
rect 1406 -22806 1456 -22794
rect 1406 -23203 1412 -22806
rect 1450 -23203 1456 -22806
rect 1406 -23215 1456 -23203
rect -1456 -33637 -1406 -33625
rect -1456 -34034 -1450 -33637
rect -1412 -34034 -1406 -33637
rect -1456 -34046 -1406 -34034
rect -1138 -33637 -1088 -33625
rect -1138 -34034 -1132 -33637
rect -1094 -34034 -1088 -33637
rect -1138 -34046 -1088 -34034
rect -820 -33637 -770 -33625
rect -820 -34034 -814 -33637
rect -776 -34034 -770 -33637
rect -820 -34046 -770 -34034
rect -502 -33637 -452 -33625
rect -502 -34034 -496 -33637
rect -458 -34034 -452 -33637
rect -502 -34046 -452 -34034
rect -184 -33637 -134 -33625
rect -184 -34034 -178 -33637
rect -140 -34034 -134 -33637
rect -184 -34046 -134 -34034
rect 134 -33637 184 -33625
rect 134 -34034 140 -33637
rect 178 -34034 184 -33637
rect 134 -34046 184 -34034
rect 452 -33637 502 -33625
rect 452 -34034 458 -33637
rect 496 -34034 502 -33637
rect 452 -34046 502 -34034
rect 770 -33637 820 -33625
rect 770 -34034 776 -33637
rect 814 -34034 820 -33637
rect 770 -34046 820 -34034
rect 1088 -33637 1138 -33625
rect 1088 -34034 1094 -33637
rect 1132 -34034 1138 -33637
rect 1088 -34046 1138 -34034
rect 1406 -33637 1456 -33625
rect 1406 -34034 1412 -33637
rect 1450 -34034 1456 -33637
rect 1406 -34046 1456 -34034
rect -1456 -34174 -1406 -34162
rect -1456 -34571 -1450 -34174
rect -1412 -34571 -1406 -34174
rect -1456 -34583 -1406 -34571
rect -1138 -34174 -1088 -34162
rect -1138 -34571 -1132 -34174
rect -1094 -34571 -1088 -34174
rect -1138 -34583 -1088 -34571
rect -820 -34174 -770 -34162
rect -820 -34571 -814 -34174
rect -776 -34571 -770 -34174
rect -820 -34583 -770 -34571
rect -502 -34174 -452 -34162
rect -502 -34571 -496 -34174
rect -458 -34571 -452 -34174
rect -502 -34583 -452 -34571
rect -184 -34174 -134 -34162
rect -184 -34571 -178 -34174
rect -140 -34571 -134 -34174
rect -184 -34583 -134 -34571
rect 134 -34174 184 -34162
rect 134 -34571 140 -34174
rect 178 -34571 184 -34174
rect 134 -34583 184 -34571
rect 452 -34174 502 -34162
rect 452 -34571 458 -34174
rect 496 -34571 502 -34174
rect 452 -34583 502 -34571
rect 770 -34174 820 -34162
rect 770 -34571 776 -34174
rect 814 -34571 820 -34174
rect 770 -34583 820 -34571
rect 1088 -34174 1138 -34162
rect 1088 -34571 1094 -34174
rect 1132 -34571 1138 -34174
rect 1088 -34583 1138 -34571
rect 1406 -34174 1456 -34162
rect 1406 -34571 1412 -34174
rect 1450 -34571 1456 -34174
rect 1406 -34583 1456 -34571
rect -1456 -45005 -1406 -44993
rect -1456 -45402 -1450 -45005
rect -1412 -45402 -1406 -45005
rect -1456 -45414 -1406 -45402
rect -1138 -45005 -1088 -44993
rect -1138 -45402 -1132 -45005
rect -1094 -45402 -1088 -45005
rect -1138 -45414 -1088 -45402
rect -820 -45005 -770 -44993
rect -820 -45402 -814 -45005
rect -776 -45402 -770 -45005
rect -820 -45414 -770 -45402
rect -502 -45005 -452 -44993
rect -502 -45402 -496 -45005
rect -458 -45402 -452 -45005
rect -502 -45414 -452 -45402
rect -184 -45005 -134 -44993
rect -184 -45402 -178 -45005
rect -140 -45402 -134 -45005
rect -184 -45414 -134 -45402
rect 134 -45005 184 -44993
rect 134 -45402 140 -45005
rect 178 -45402 184 -45005
rect 134 -45414 184 -45402
rect 452 -45005 502 -44993
rect 452 -45402 458 -45005
rect 496 -45402 502 -45005
rect 452 -45414 502 -45402
rect 770 -45005 820 -44993
rect 770 -45402 776 -45005
rect 814 -45402 820 -45005
rect 770 -45414 820 -45402
rect 1088 -45005 1138 -44993
rect 1088 -45402 1094 -45005
rect 1132 -45402 1138 -45005
rect 1088 -45414 1138 -45402
rect 1406 -45005 1456 -44993
rect 1406 -45402 1412 -45005
rect 1450 -45402 1456 -45005
rect 1406 -45414 1456 -45402
rect -1456 -45542 -1406 -45530
rect -1456 -45939 -1450 -45542
rect -1412 -45939 -1406 -45542
rect -1456 -45951 -1406 -45939
rect -1138 -45542 -1088 -45530
rect -1138 -45939 -1132 -45542
rect -1094 -45939 -1088 -45542
rect -1138 -45951 -1088 -45939
rect -820 -45542 -770 -45530
rect -820 -45939 -814 -45542
rect -776 -45939 -770 -45542
rect -820 -45951 -770 -45939
rect -502 -45542 -452 -45530
rect -502 -45939 -496 -45542
rect -458 -45939 -452 -45542
rect -502 -45951 -452 -45939
rect -184 -45542 -134 -45530
rect -184 -45939 -178 -45542
rect -140 -45939 -134 -45542
rect -184 -45951 -134 -45939
rect 134 -45542 184 -45530
rect 134 -45939 140 -45542
rect 178 -45939 184 -45542
rect 134 -45951 184 -45939
rect 452 -45542 502 -45530
rect 452 -45939 458 -45542
rect 496 -45939 502 -45542
rect 452 -45951 502 -45939
rect 770 -45542 820 -45530
rect 770 -45939 776 -45542
rect 814 -45939 820 -45542
rect 770 -45951 820 -45939
rect 1088 -45542 1138 -45530
rect 1088 -45939 1094 -45542
rect 1132 -45939 1138 -45542
rect 1088 -45951 1138 -45939
rect 1406 -45542 1456 -45530
rect 1406 -45939 1412 -45542
rect 1450 -45939 1456 -45542
rect 1406 -45951 1456 -45939
rect -1456 -56373 -1406 -56361
rect -1456 -56770 -1450 -56373
rect -1412 -56770 -1406 -56373
rect -1456 -56782 -1406 -56770
rect -1138 -56373 -1088 -56361
rect -1138 -56770 -1132 -56373
rect -1094 -56770 -1088 -56373
rect -1138 -56782 -1088 -56770
rect -820 -56373 -770 -56361
rect -820 -56770 -814 -56373
rect -776 -56770 -770 -56373
rect -820 -56782 -770 -56770
rect -502 -56373 -452 -56361
rect -502 -56770 -496 -56373
rect -458 -56770 -452 -56373
rect -502 -56782 -452 -56770
rect -184 -56373 -134 -56361
rect -184 -56770 -178 -56373
rect -140 -56770 -134 -56373
rect -184 -56782 -134 -56770
rect 134 -56373 184 -56361
rect 134 -56770 140 -56373
rect 178 -56770 184 -56373
rect 134 -56782 184 -56770
rect 452 -56373 502 -56361
rect 452 -56770 458 -56373
rect 496 -56770 502 -56373
rect 452 -56782 502 -56770
rect 770 -56373 820 -56361
rect 770 -56770 776 -56373
rect 814 -56770 820 -56373
rect 770 -56782 820 -56770
rect 1088 -56373 1138 -56361
rect 1088 -56770 1094 -56373
rect 1132 -56770 1138 -56373
rect 1088 -56782 1138 -56770
rect 1406 -56373 1456 -56361
rect 1406 -56770 1412 -56373
rect 1450 -56770 1456 -56373
rect 1406 -56782 1456 -56770
<< res0p35 >>
rect -1468 45954 -1394 56358
rect -1150 45954 -1076 56358
rect -832 45954 -758 56358
rect -514 45954 -440 56358
rect -196 45954 -122 56358
rect 122 45954 196 56358
rect 440 45954 514 56358
rect 758 45954 832 56358
rect 1076 45954 1150 56358
rect 1394 45954 1468 56358
rect -1468 34586 -1394 44990
rect -1150 34586 -1076 44990
rect -832 34586 -758 44990
rect -514 34586 -440 44990
rect -196 34586 -122 44990
rect 122 34586 196 44990
rect 440 34586 514 44990
rect 758 34586 832 44990
rect 1076 34586 1150 44990
rect 1394 34586 1468 44990
rect -1468 23218 -1394 33622
rect -1150 23218 -1076 33622
rect -832 23218 -758 33622
rect -514 23218 -440 33622
rect -196 23218 -122 33622
rect 122 23218 196 33622
rect 440 23218 514 33622
rect 758 23218 832 33622
rect 1076 23218 1150 33622
rect 1394 23218 1468 33622
rect -1468 11850 -1394 22254
rect -1150 11850 -1076 22254
rect -832 11850 -758 22254
rect -514 11850 -440 22254
rect -196 11850 -122 22254
rect 122 11850 196 22254
rect 440 11850 514 22254
rect 758 11850 832 22254
rect 1076 11850 1150 22254
rect 1394 11850 1468 22254
rect -1468 482 -1394 10886
rect -1150 482 -1076 10886
rect -832 482 -758 10886
rect -514 482 -440 10886
rect -196 482 -122 10886
rect 122 482 196 10886
rect 440 482 514 10886
rect 758 482 832 10886
rect 1076 482 1150 10886
rect 1394 482 1468 10886
rect -1468 -10886 -1394 -482
rect -1150 -10886 -1076 -482
rect -832 -10886 -758 -482
rect -514 -10886 -440 -482
rect -196 -10886 -122 -482
rect 122 -10886 196 -482
rect 440 -10886 514 -482
rect 758 -10886 832 -482
rect 1076 -10886 1150 -482
rect 1394 -10886 1468 -482
rect -1468 -22254 -1394 -11850
rect -1150 -22254 -1076 -11850
rect -832 -22254 -758 -11850
rect -514 -22254 -440 -11850
rect -196 -22254 -122 -11850
rect 122 -22254 196 -11850
rect 440 -22254 514 -11850
rect 758 -22254 832 -11850
rect 1076 -22254 1150 -11850
rect 1394 -22254 1468 -11850
rect -1468 -33622 -1394 -23218
rect -1150 -33622 -1076 -23218
rect -832 -33622 -758 -23218
rect -514 -33622 -440 -23218
rect -196 -33622 -122 -23218
rect 122 -33622 196 -23218
rect 440 -33622 514 -23218
rect 758 -33622 832 -23218
rect 1076 -33622 1150 -23218
rect 1394 -33622 1468 -23218
rect -1468 -44990 -1394 -34586
rect -1150 -44990 -1076 -34586
rect -832 -44990 -758 -34586
rect -514 -44990 -440 -34586
rect -196 -44990 -122 -34586
rect 122 -44990 196 -34586
rect 440 -44990 514 -34586
rect 758 -44990 832 -34586
rect 1076 -44990 1150 -34586
rect 1394 -44990 1468 -34586
rect -1468 -56358 -1394 -45954
rect -1150 -56358 -1076 -45954
rect -832 -56358 -758 -45954
rect -514 -56358 -440 -45954
rect -196 -56358 -122 -45954
rect 122 -56358 196 -45954
rect 440 -56358 514 -45954
rect 758 -56358 832 -45954
rect 1076 -56358 1150 -45954
rect 1394 -56358 1468 -45954
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 52 m 10 nx 10 wmin 0.350 lmin 0.50 rho 2000 val 298.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
