magic
tech sky130A
magscale 1 2
timestamp 1668374365
<< error_p >>
rect -29 60617 29 60623
rect -29 60583 -17 60617
rect -29 60577 29 60583
rect -29 40507 29 40513
rect -29 40473 -17 40507
rect -29 40467 29 40473
rect -29 40399 29 40405
rect -29 40365 -17 40399
rect -29 40359 29 40365
rect -29 20289 29 20295
rect -29 20255 -17 20289
rect -29 20249 29 20255
rect -29 20181 29 20187
rect -29 20147 -17 20181
rect -29 20141 29 20147
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -20147 29 -20141
rect -29 -20181 -17 -20147
rect -29 -20187 29 -20181
rect -29 -20255 29 -20249
rect -29 -20289 -17 -20255
rect -29 -20295 29 -20289
rect -29 -40365 29 -40359
rect -29 -40399 -17 -40365
rect -29 -40405 29 -40399
rect -29 -40473 29 -40467
rect -29 -40507 -17 -40473
rect -29 -40513 29 -40507
rect -29 -60583 29 -60577
rect -29 -60617 -17 -60583
rect -29 -60623 29 -60617
<< pwell >>
rect -226 -60755 226 60755
<< nmos >>
rect -30 40545 30 60545
rect -30 20327 30 40327
rect -30 109 30 20109
rect -30 -20109 30 -109
rect -30 -40327 30 -20327
rect -30 -60545 30 -40545
<< ndiff >>
rect -88 60533 -30 60545
rect -88 40557 -76 60533
rect -42 40557 -30 60533
rect -88 40545 -30 40557
rect 30 60533 88 60545
rect 30 40557 42 60533
rect 76 40557 88 60533
rect 30 40545 88 40557
rect -88 40315 -30 40327
rect -88 20339 -76 40315
rect -42 20339 -30 40315
rect -88 20327 -30 20339
rect 30 40315 88 40327
rect 30 20339 42 40315
rect 76 20339 88 40315
rect 30 20327 88 20339
rect -88 20097 -30 20109
rect -88 121 -76 20097
rect -42 121 -30 20097
rect -88 109 -30 121
rect 30 20097 88 20109
rect 30 121 42 20097
rect 76 121 88 20097
rect 30 109 88 121
rect -88 -121 -30 -109
rect -88 -20097 -76 -121
rect -42 -20097 -30 -121
rect -88 -20109 -30 -20097
rect 30 -121 88 -109
rect 30 -20097 42 -121
rect 76 -20097 88 -121
rect 30 -20109 88 -20097
rect -88 -20339 -30 -20327
rect -88 -40315 -76 -20339
rect -42 -40315 -30 -20339
rect -88 -40327 -30 -40315
rect 30 -20339 88 -20327
rect 30 -40315 42 -20339
rect 76 -40315 88 -20339
rect 30 -40327 88 -40315
rect -88 -40557 -30 -40545
rect -88 -60533 -76 -40557
rect -42 -60533 -30 -40557
rect -88 -60545 -30 -60533
rect 30 -40557 88 -40545
rect 30 -60533 42 -40557
rect 76 -60533 88 -40557
rect 30 -60545 88 -60533
<< ndiffc >>
rect -76 40557 -42 60533
rect 42 40557 76 60533
rect -76 20339 -42 40315
rect 42 20339 76 40315
rect -76 121 -42 20097
rect 42 121 76 20097
rect -76 -20097 -42 -121
rect 42 -20097 76 -121
rect -76 -40315 -42 -20339
rect 42 -40315 76 -20339
rect -76 -60533 -42 -40557
rect 42 -60533 76 -40557
<< psubdiff >>
rect -190 60685 -94 60719
rect 94 60685 190 60719
rect -190 60623 -156 60685
rect 156 60623 190 60685
rect -190 -60685 -156 -60623
rect 156 -60685 190 -60623
rect -190 -60719 -94 -60685
rect 94 -60719 190 -60685
<< psubdiffcont >>
rect -94 60685 94 60719
rect -190 -60623 -156 60623
rect 156 -60623 190 60623
rect -94 -60719 94 -60685
<< poly >>
rect -33 60617 33 60633
rect -33 60583 -17 60617
rect 17 60583 33 60617
rect -33 60567 33 60583
rect -30 60545 30 60567
rect -30 40523 30 40545
rect -33 40507 33 40523
rect -33 40473 -17 40507
rect 17 40473 33 40507
rect -33 40457 33 40473
rect -33 40399 33 40415
rect -33 40365 -17 40399
rect 17 40365 33 40399
rect -33 40349 33 40365
rect -30 40327 30 40349
rect -30 20305 30 20327
rect -33 20289 33 20305
rect -33 20255 -17 20289
rect 17 20255 33 20289
rect -33 20239 33 20255
rect -33 20181 33 20197
rect -33 20147 -17 20181
rect 17 20147 33 20181
rect -33 20131 33 20147
rect -30 20109 30 20131
rect -30 87 30 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -109 30 -87
rect -30 -20131 30 -20109
rect -33 -20147 33 -20131
rect -33 -20181 -17 -20147
rect 17 -20181 33 -20147
rect -33 -20197 33 -20181
rect -33 -20255 33 -20239
rect -33 -20289 -17 -20255
rect 17 -20289 33 -20255
rect -33 -20305 33 -20289
rect -30 -20327 30 -20305
rect -30 -40349 30 -40327
rect -33 -40365 33 -40349
rect -33 -40399 -17 -40365
rect 17 -40399 33 -40365
rect -33 -40415 33 -40399
rect -33 -40473 33 -40457
rect -33 -40507 -17 -40473
rect 17 -40507 33 -40473
rect -33 -40523 33 -40507
rect -30 -40545 30 -40523
rect -30 -60567 30 -60545
rect -33 -60583 33 -60567
rect -33 -60617 -17 -60583
rect 17 -60617 33 -60583
rect -33 -60633 33 -60617
<< polycont >>
rect -17 60583 17 60617
rect -17 40473 17 40507
rect -17 40365 17 40399
rect -17 20255 17 20289
rect -17 20147 17 20181
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -20181 17 -20147
rect -17 -20289 17 -20255
rect -17 -40399 17 -40365
rect -17 -40507 17 -40473
rect -17 -60617 17 -60583
<< locali >>
rect -190 60685 -94 60719
rect 94 60685 190 60719
rect -190 60623 -156 60685
rect 156 60623 190 60685
rect -33 60583 -17 60617
rect 17 60583 33 60617
rect -76 60533 -42 60549
rect -76 40541 -42 40557
rect 42 60533 76 60549
rect 42 40541 76 40557
rect -33 40473 -17 40507
rect 17 40473 33 40507
rect -33 40365 -17 40399
rect 17 40365 33 40399
rect -76 40315 -42 40331
rect -76 20323 -42 20339
rect 42 40315 76 40331
rect 42 20323 76 20339
rect -33 20255 -17 20289
rect 17 20255 33 20289
rect -33 20147 -17 20181
rect 17 20147 33 20181
rect -76 20097 -42 20113
rect -76 105 -42 121
rect 42 20097 76 20113
rect 42 105 76 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -121 -42 -105
rect -76 -20113 -42 -20097
rect 42 -121 76 -105
rect 42 -20113 76 -20097
rect -33 -20181 -17 -20147
rect 17 -20181 33 -20147
rect -33 -20289 -17 -20255
rect 17 -20289 33 -20255
rect -76 -20339 -42 -20323
rect -76 -40331 -42 -40315
rect 42 -20339 76 -20323
rect 42 -40331 76 -40315
rect -33 -40399 -17 -40365
rect 17 -40399 33 -40365
rect -33 -40507 -17 -40473
rect 17 -40507 33 -40473
rect -76 -40557 -42 -40541
rect -76 -60549 -42 -60533
rect 42 -40557 76 -40541
rect 42 -60549 76 -60533
rect -33 -60617 -17 -60583
rect 17 -60617 33 -60583
rect -190 -60685 -156 -60623
rect 156 -60685 190 -60623
rect -190 -60719 -94 -60685
rect 94 -60719 190 -60685
<< viali >>
rect -17 60583 17 60617
rect -76 40557 -42 60533
rect 42 40557 76 60533
rect -17 40473 17 40507
rect -17 40365 17 40399
rect -76 20339 -42 40315
rect 42 20339 76 40315
rect -17 20255 17 20289
rect -17 20147 17 20181
rect -76 121 -42 20097
rect 42 121 76 20097
rect -17 37 17 71
rect -17 -71 17 -37
rect -76 -20097 -42 -121
rect 42 -20097 76 -121
rect -17 -20181 17 -20147
rect -17 -20289 17 -20255
rect -76 -40315 -42 -20339
rect 42 -40315 76 -20339
rect -17 -40399 17 -40365
rect -17 -40507 17 -40473
rect -76 -60533 -42 -40557
rect 42 -60533 76 -40557
rect -17 -60617 17 -60583
<< metal1 >>
rect -29 60617 29 60623
rect -29 60583 -17 60617
rect 17 60583 29 60617
rect -29 60577 29 60583
rect -82 60533 -36 60545
rect -82 40557 -76 60533
rect -42 40557 -36 60533
rect -82 40545 -36 40557
rect 36 60533 82 60545
rect 36 40557 42 60533
rect 76 40557 82 60533
rect 36 40545 82 40557
rect -29 40507 29 40513
rect -29 40473 -17 40507
rect 17 40473 29 40507
rect -29 40467 29 40473
rect -29 40399 29 40405
rect -29 40365 -17 40399
rect 17 40365 29 40399
rect -29 40359 29 40365
rect -82 40315 -36 40327
rect -82 20339 -76 40315
rect -42 20339 -36 40315
rect -82 20327 -36 20339
rect 36 40315 82 40327
rect 36 20339 42 40315
rect 76 20339 82 40315
rect 36 20327 82 20339
rect -29 20289 29 20295
rect -29 20255 -17 20289
rect 17 20255 29 20289
rect -29 20249 29 20255
rect -29 20181 29 20187
rect -29 20147 -17 20181
rect 17 20147 29 20181
rect -29 20141 29 20147
rect -82 20097 -36 20109
rect -82 121 -76 20097
rect -42 121 -36 20097
rect -82 109 -36 121
rect 36 20097 82 20109
rect 36 121 42 20097
rect 76 121 82 20097
rect 36 109 82 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -121 -36 -109
rect -82 -20097 -76 -121
rect -42 -20097 -36 -121
rect -82 -20109 -36 -20097
rect 36 -121 82 -109
rect 36 -20097 42 -121
rect 76 -20097 82 -121
rect 36 -20109 82 -20097
rect -29 -20147 29 -20141
rect -29 -20181 -17 -20147
rect 17 -20181 29 -20147
rect -29 -20187 29 -20181
rect -29 -20255 29 -20249
rect -29 -20289 -17 -20255
rect 17 -20289 29 -20255
rect -29 -20295 29 -20289
rect -82 -20339 -36 -20327
rect -82 -40315 -76 -20339
rect -42 -40315 -36 -20339
rect -82 -40327 -36 -40315
rect 36 -20339 82 -20327
rect 36 -40315 42 -20339
rect 76 -40315 82 -20339
rect 36 -40327 82 -40315
rect -29 -40365 29 -40359
rect -29 -40399 -17 -40365
rect 17 -40399 29 -40365
rect -29 -40405 29 -40399
rect -29 -40473 29 -40467
rect -29 -40507 -17 -40473
rect 17 -40507 29 -40473
rect -29 -40513 29 -40507
rect -82 -40557 -36 -40545
rect -82 -60533 -76 -40557
rect -42 -60533 -36 -40557
rect -82 -60545 -36 -60533
rect 36 -40557 82 -40545
rect 36 -60533 42 -40557
rect 76 -60533 82 -40557
rect 36 -60545 82 -60533
rect -29 -60583 29 -60577
rect -29 -60617 -17 -60583
rect 17 -60617 29 -60583
rect -29 -60623 29 -60617
<< properties >>
string FIXED_BBOX -173 -60702 173 60702
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 100.0 l 0.3 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
