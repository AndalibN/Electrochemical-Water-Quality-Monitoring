magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 341 29 347
rect -29 307 -17 341
rect -29 301 29 307
<< pwell >>
rect -114 -357 114 295
<< nmos >>
rect -30 -331 30 269
<< ndiff >>
rect -88 224 -30 269
rect -88 190 -76 224
rect -42 190 -30 224
rect -88 156 -30 190
rect -88 122 -76 156
rect -42 122 -30 156
rect -88 88 -30 122
rect -88 54 -76 88
rect -42 54 -30 88
rect -88 20 -30 54
rect -88 -14 -76 20
rect -42 -14 -30 20
rect -88 -48 -30 -14
rect -88 -82 -76 -48
rect -42 -82 -30 -48
rect -88 -116 -30 -82
rect -88 -150 -76 -116
rect -42 -150 -30 -116
rect -88 -184 -30 -150
rect -88 -218 -76 -184
rect -42 -218 -30 -184
rect -88 -252 -30 -218
rect -88 -286 -76 -252
rect -42 -286 -30 -252
rect -88 -331 -30 -286
rect 30 224 88 269
rect 30 190 42 224
rect 76 190 88 224
rect 30 156 88 190
rect 30 122 42 156
rect 76 122 88 156
rect 30 88 88 122
rect 30 54 42 88
rect 76 54 88 88
rect 30 20 88 54
rect 30 -14 42 20
rect 76 -14 88 20
rect 30 -48 88 -14
rect 30 -82 42 -48
rect 76 -82 88 -48
rect 30 -116 88 -82
rect 30 -150 42 -116
rect 76 -150 88 -116
rect 30 -184 88 -150
rect 30 -218 42 -184
rect 76 -218 88 -184
rect 30 -252 88 -218
rect 30 -286 42 -252
rect 76 -286 88 -252
rect 30 -331 88 -286
<< ndiffc >>
rect -76 190 -42 224
rect -76 122 -42 156
rect -76 54 -42 88
rect -76 -14 -42 20
rect -76 -82 -42 -48
rect -76 -150 -42 -116
rect -76 -218 -42 -184
rect -76 -286 -42 -252
rect 42 190 76 224
rect 42 122 76 156
rect 42 54 76 88
rect 42 -14 76 20
rect 42 -82 76 -48
rect 42 -150 76 -116
rect 42 -218 76 -184
rect 42 -286 76 -252
<< poly >>
rect -33 341 33 357
rect -33 307 -17 341
rect 17 307 33 341
rect -33 291 33 307
rect -30 269 30 291
rect -30 -357 30 -331
<< polycont >>
rect -17 307 17 341
<< locali >>
rect -33 307 -17 341
rect 17 307 33 341
rect -76 238 -42 273
rect -76 166 -42 190
rect -76 94 -42 122
rect -76 22 -42 54
rect -76 -48 -42 -14
rect -76 -116 -42 -84
rect -76 -184 -42 -156
rect -76 -252 -42 -228
rect -76 -335 -42 -300
rect 42 238 76 273
rect 42 166 76 190
rect 42 94 76 122
rect 42 22 76 54
rect 42 -48 76 -14
rect 42 -116 76 -84
rect 42 -184 76 -156
rect 42 -252 76 -228
rect 42 -335 76 -300
<< viali >>
rect -17 307 17 341
rect -76 224 -42 238
rect -76 204 -42 224
rect -76 156 -42 166
rect -76 132 -42 156
rect -76 88 -42 94
rect -76 60 -42 88
rect -76 20 -42 22
rect -76 -12 -42 20
rect -76 -82 -42 -50
rect -76 -84 -42 -82
rect -76 -150 -42 -122
rect -76 -156 -42 -150
rect -76 -218 -42 -194
rect -76 -228 -42 -218
rect -76 -286 -42 -266
rect -76 -300 -42 -286
rect 42 224 76 238
rect 42 204 76 224
rect 42 156 76 166
rect 42 132 76 156
rect 42 88 76 94
rect 42 60 76 88
rect 42 20 76 22
rect 42 -12 76 20
rect 42 -82 76 -50
rect 42 -84 76 -82
rect 42 -150 76 -122
rect 42 -156 76 -150
rect 42 -218 76 -194
rect 42 -228 76 -218
rect 42 -286 76 -266
rect 42 -300 76 -286
<< metal1 >>
rect -29 341 29 347
rect -29 307 -17 341
rect 17 307 29 341
rect -29 301 29 307
rect -82 238 -36 269
rect -82 204 -76 238
rect -42 204 -36 238
rect -82 166 -36 204
rect -82 132 -76 166
rect -42 132 -36 166
rect -82 94 -36 132
rect -82 60 -76 94
rect -42 60 -36 94
rect -82 22 -36 60
rect -82 -12 -76 22
rect -42 -12 -36 22
rect -82 -50 -36 -12
rect -82 -84 -76 -50
rect -42 -84 -36 -50
rect -82 -122 -36 -84
rect -82 -156 -76 -122
rect -42 -156 -36 -122
rect -82 -194 -36 -156
rect -82 -228 -76 -194
rect -42 -228 -36 -194
rect -82 -266 -36 -228
rect -82 -300 -76 -266
rect -42 -300 -36 -266
rect -82 -331 -36 -300
rect 36 238 82 269
rect 36 204 42 238
rect 76 204 82 238
rect 36 166 82 204
rect 36 132 42 166
rect 76 132 82 166
rect 36 94 82 132
rect 36 60 42 94
rect 76 60 82 94
rect 36 22 82 60
rect 36 -12 42 22
rect 76 -12 82 22
rect 36 -50 82 -12
rect 36 -84 42 -50
rect 76 -84 82 -50
rect 36 -122 82 -84
rect 36 -156 42 -122
rect 76 -156 82 -122
rect 36 -194 82 -156
rect 36 -228 42 -194
rect 76 -228 82 -194
rect 36 -266 82 -228
rect 36 -300 42 -266
rect 76 -300 82 -266
rect 36 -331 82 -300
<< end >>
