magic
tech sky130A
magscale 1 2
timestamp 1667937831
<< error_p >>
rect -88 -311 -30 -305
rect 30 -311 88 -305
rect -88 -345 -76 -311
rect 30 -345 42 -311
rect -88 -351 -30 -345
rect 30 -351 88 -345
<< nwell >>
rect -183 -364 183 398
<< pmos >>
rect -89 -264 -29 336
rect 29 -264 89 336
<< pdiff >>
rect -147 324 -89 336
rect -147 -252 -135 324
rect -101 -252 -89 324
rect -147 -264 -89 -252
rect -29 324 29 336
rect -29 -252 -17 324
rect 17 -252 29 324
rect -29 -264 29 -252
rect 89 324 147 336
rect 89 -252 101 324
rect 135 -252 147 324
rect 89 -264 147 -252
<< pdiffc >>
rect -135 -252 -101 324
rect -17 -252 17 324
rect 101 -252 135 324
<< poly >>
rect -89 336 -29 362
rect 29 336 89 362
rect -89 -295 -29 -264
rect 29 -295 89 -264
rect -92 -311 -26 -295
rect -92 -345 -76 -311
rect -42 -345 -26 -311
rect -92 -361 -26 -345
rect 26 -311 92 -295
rect 26 -345 42 -311
rect 76 -345 92 -311
rect 26 -361 92 -345
<< polycont >>
rect -76 -345 -42 -311
rect 42 -345 76 -311
<< locali >>
rect -135 324 -101 340
rect -135 -268 -101 -252
rect -17 324 17 340
rect -17 -268 17 -252
rect 101 324 135 340
rect 101 -268 135 -252
rect -92 -345 -76 -311
rect -42 -345 -26 -311
rect 26 -345 42 -311
rect 76 -345 92 -311
<< viali >>
rect -135 -252 -101 324
rect -17 -252 17 324
rect 101 -252 135 324
rect -76 -345 -42 -311
rect 42 -345 76 -311
<< metal1 >>
rect -141 324 -95 336
rect -141 -252 -135 324
rect -101 -252 -95 324
rect -141 -264 -95 -252
rect -23 324 23 336
rect -23 -252 -17 324
rect 17 -252 23 324
rect -23 -264 23 -252
rect 95 324 141 336
rect 95 -252 101 324
rect 135 -252 141 324
rect 95 -264 141 -252
rect -88 -311 -30 -305
rect -88 -345 -76 -311
rect -42 -345 -30 -311
rect -88 -351 -30 -345
rect 30 -311 88 -305
rect 30 -345 42 -311
rect 76 -345 88 -311
rect 30 -351 88 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.30 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
