magic
tech sky130A
magscale 1 2
timestamp 1668206180
<< error_s >>
rect 3542 -8176 3558 -5356
<< psubdiff >>
rect 12434 11388 12564 11412
rect 12434 10328 12564 10352
rect -10835 6139 -10678 6144
rect -9376 6139 -9219 6144
rect -10841 6120 -10817 6139
rect -9220 6120 -9196 6139
rect -10841 5954 -10835 6120
rect -9219 5954 -9196 6120
rect -3616 5306 -3514 5330
rect -4802 5234 -4778 5300
rect -3514 5234 -3500 5300
rect -10859 -141 -10835 -21
rect -9200 -141 -9176 -21
rect -10835 -165 -10678 -141
rect -9376 -165 -9219 -141
rect 16371 409 16762 433
rect 12326 372 12438 396
rect -4818 -484 -4794 -418
rect -3500 -484 -3476 -418
rect -4770 -500 -4712 -484
rect -3616 -524 -3514 -500
rect 16371 -550 16762 -526
rect 12326 -746 12438 -722
rect 12205 -946 12257 -928
rect 64564 -934 65024 -910
rect 11584 -974 11608 -946
rect 12248 -952 12272 -946
rect 11584 -995 11602 -974
rect 12257 -995 12272 -952
rect 11584 -2788 11602 -2748
rect 12257 -2782 12272 -2748
rect 64564 -2760 65024 -2736
rect 11584 -2797 11608 -2788
rect 12248 -2797 12272 -2782
rect 11602 -2812 11640 -2797
rect 12205 -2806 12257 -2797
rect 10746 -5214 10770 -4560
rect 11494 -5214 11518 -4560
rect -2578 -5530 -2296 -5506
rect -2578 -6762 -2296 -6738
<< psubdiffcont >>
rect 12434 10352 12564 11388
rect -10817 6120 -9220 6139
rect -10835 5954 -9219 6120
rect -10835 -21 -10678 5954
rect -9376 -21 -9219 5954
rect -3616 5300 -3514 5306
rect -4778 5234 -3514 5300
rect -10835 -141 -9200 -21
rect -4770 -418 -4712 5234
rect -3616 -418 -3514 5234
rect -4794 -484 -3500 -418
rect -3616 -500 -3514 -484
rect 12326 -722 12438 372
rect 16371 -526 16762 409
rect 11608 -952 12248 -946
rect 11608 -974 12257 -952
rect 11602 -995 12257 -974
rect 11602 -2748 11640 -995
rect 12205 -2748 12257 -995
rect 64564 -2736 65024 -934
rect 11602 -2782 12257 -2748
rect 11602 -2788 12248 -2782
rect 11608 -2797 12248 -2788
rect 10770 -5214 11494 -4560
rect -2578 -6738 -2296 -5530
<< locali >>
rect 12434 11388 12564 11404
rect 12434 10336 12564 10352
rect -10833 6136 -10817 6139
rect -10835 6120 -10817 6136
rect -9220 6120 -9204 6139
rect -9219 5954 -9204 6120
rect -9380 5178 -9376 5240
rect -10128 352 -10094 668
rect -9900 382 -9866 676
rect -9901 352 -9866 382
rect -10129 348 -9866 352
rect -10129 306 -9867 348
rect -3616 5306 -3514 5322
rect -4794 5240 -4778 5300
rect -9219 5234 -4778 5240
rect -3514 5234 -3508 5300
rect -9219 5178 -4770 5234
rect -10851 -141 -10835 -21
rect -9200 -141 -9184 -21
rect -10835 -157 -10678 -141
rect -9376 -157 -9219 -141
rect -4286 -326 -4252 -88
rect -4058 -326 -4024 -80
rect -4286 -364 -4024 -326
rect 4920 5196 5102 5197
rect -3514 5074 5102 5196
rect -4810 -484 -4794 -418
rect -3500 -484 -3484 -418
rect -4770 -492 -4712 -484
rect -3616 -516 -3514 -500
rect 2318 -4938 2814 5074
rect 4920 -1358 5102 5074
rect 12366 1476 12436 1485
rect 16600 1476 16646 1546
rect 12366 1444 16646 1476
rect 64730 1444 64828 6030
rect 12366 1386 64828 1444
rect 10890 780 10944 792
rect 12366 780 12436 1386
rect 16598 1228 64828 1386
rect 10890 716 12436 780
rect 10890 -1358 10944 716
rect 12366 388 12436 716
rect 16600 534 16646 1228
rect 12326 372 12438 388
rect 15860 66 16249 499
rect 16600 425 16670 534
rect 16371 409 16762 425
rect 15542 -680 15931 -247
rect 16371 -542 16762 -526
rect 12326 -738 12438 -722
rect 64730 -918 64828 1228
rect 64564 -934 65024 -918
rect 12205 -946 12257 -936
rect 11592 -974 11608 -946
rect 12248 -952 12264 -946
rect 11592 -995 11602 -974
rect 12257 -995 12264 -952
rect 11562 -1358 11602 -1350
rect 4920 -1460 11602 -1358
rect 11562 -1466 11602 -1460
rect 11592 -2788 11602 -2748
rect 12257 -2782 12264 -2748
rect 64564 -2752 65024 -2736
rect 11592 -2797 11608 -2788
rect 12248 -2797 12264 -2782
rect 11602 -2804 11640 -2797
rect 11302 -3404 11376 -3388
rect 11302 -3446 11310 -3404
rect 11370 -3446 11376 -3404
rect 11302 -4560 11376 -3446
rect 11854 -4448 11996 -4436
rect -2452 -5038 2814 -4938
rect -2458 -5096 2814 -5038
rect -2458 -5112 2424 -5096
rect -2458 -5514 -2380 -5112
rect 10754 -5214 10770 -4560
rect 11494 -4632 11510 -4560
rect 11854 -4564 11866 -4448
rect 11980 -4564 11996 -4448
rect 11854 -4632 11996 -4564
rect 11494 -4696 11996 -4632
rect 11494 -5067 11510 -4696
rect 12088 -5067 12164 -2797
rect 12205 -2798 12257 -2797
rect 11494 -5108 12164 -5067
rect 11494 -5116 12098 -5108
rect 11494 -5214 11510 -5116
rect -2578 -5530 -2296 -5514
rect -2578 -6754 -2296 -6738
<< viali >>
rect 11310 -3446 11370 -3404
rect 11866 -4564 11980 -4448
<< metal1 >>
rect -1748 19058 280 19160
rect -1748 18086 -1320 19058
rect -26 18086 280 19058
rect -1748 15844 280 18086
rect 11960 15844 12210 16334
rect -1748 15080 12210 15844
rect -1748 15012 280 15080
rect -1772 14346 280 15012
rect 11960 14432 12210 15080
rect 11948 14390 12210 14432
rect 11948 14294 12204 14390
rect 4618 13200 5094 13234
rect 4618 12912 4738 13200
rect 5000 12912 5094 13200
rect 4618 11938 5094 12912
rect 11994 12484 12194 14294
rect 13030 12484 13166 12504
rect 11994 12446 13166 12484
rect 12002 12294 13166 12446
rect 4786 9450 4984 11938
rect 13030 11468 13166 12294
rect 12694 11008 14488 11468
rect 12700 10342 14494 10802
rect 12964 9572 13116 10342
rect 12006 9530 13116 9572
rect 11994 9450 13116 9530
rect 4786 9382 13078 9450
rect 4786 9250 12382 9382
rect 11994 8234 12194 9250
rect 11756 7654 12194 8234
rect 11994 7232 12194 7654
rect 20136 7232 23624 7236
rect -10172 6974 -10054 6990
rect -10172 6888 -10146 6974
rect -10070 6888 -10054 6974
rect -10172 6586 -10054 6888
rect 11994 6964 23624 7232
rect -10156 6500 -10070 6586
rect -10128 5716 -10094 6500
rect 11994 5860 12194 6964
rect 11994 5842 12190 5860
rect 11266 5836 12190 5842
rect 9442 5832 12190 5836
rect 5786 5828 12190 5832
rect 3948 5824 12190 5828
rect 318 5822 12190 5824
rect -3232 5820 12190 5822
rect -5082 5818 12190 5820
rect -8278 5814 -7116 5816
rect -6022 5814 12190 5818
rect -9428 5810 12190 5814
rect -9632 5808 12190 5810
rect -9840 5792 12190 5808
rect -9840 5786 11310 5792
rect -9840 5782 9472 5786
rect -9840 5778 5816 5782
rect -9840 5774 3996 5778
rect -9840 5772 454 5774
rect -9840 5770 -5996 5772
rect -5082 5770 -3214 5772
rect -9840 5768 -9628 5770
rect -9428 5768 -8266 5770
rect -7158 5768 -5996 5770
rect -10128 5594 -10082 5716
rect -9840 5706 -9810 5768
rect -9856 5678 -9798 5706
rect -9836 5598 -9806 5678
rect -10242 148 -10208 5424
rect -10128 488 -10094 5594
rect -9856 5470 -9798 5598
rect 19960 5486 23624 6964
rect -10014 148 -9980 5424
rect -9900 488 -9866 5424
rect -9786 148 -9752 5424
rect 18778 5419 23624 5486
rect -5242 5076 -4606 5078
rect -7498 5074 -6336 5076
rect -5242 5074 -4600 5076
rect -8648 5070 -4600 5074
rect -8852 5068 -4600 5070
rect -9060 5032 -4600 5068
rect -9060 5030 -5216 5032
rect -9060 5028 -8848 5030
rect -8648 5028 -7486 5030
rect -6378 5028 -5216 5030
rect -9060 2670 -9030 5028
rect -4636 4984 -4600 5032
rect -4288 4984 -4058 4986
rect -4636 4956 -4058 4984
rect -4636 4954 -4252 4956
rect -4636 4738 -4600 4954
rect -9060 2644 -9028 2670
rect -9058 148 -9028 2644
rect -10420 120 -9028 148
rect -10420 114 -9032 120
rect -10420 112 -9702 114
rect -4400 -242 -4366 4828
rect -4286 -108 -4252 4954
rect -4018 4876 -3678 4922
rect -3708 4830 -3680 4876
rect -2972 4832 -2706 4834
rect -2972 4830 -2518 4832
rect -3730 4828 -2518 4830
rect -4172 -242 -4138 4828
rect -4058 -108 -4024 4828
rect -3944 3240 -3910 4828
rect -3730 4780 -2498 4828
rect -3730 4776 -2962 4780
rect -2856 4778 -2590 4780
rect -3944 3168 -2642 3240
rect -3944 3160 -2636 3168
rect -3944 3054 -2736 3160
rect -2646 3054 -2636 3160
rect -3944 3052 -2636 3054
rect -3944 3038 -2642 3052
rect -3944 -242 -3910 3038
rect -2556 2962 -2498 4780
rect 19960 4184 23624 5419
rect 19960 3693 20376 4184
rect 12622 3413 20376 3693
rect 12585 3064 20376 3413
rect 12585 3027 20196 3064
rect -2556 2956 -2496 2962
rect -2554 810 -2496 2956
rect -3294 790 -2496 810
rect -3302 674 -2496 790
rect -3302 664 -2504 674
rect -3302 -150 -3240 664
rect 12585 383 12808 3027
rect 12541 322 12808 383
rect 15188 734 15379 739
rect 15544 734 15612 738
rect 15188 664 15612 734
rect 12541 318 12711 322
rect 12541 171 12612 318
rect -3328 -166 -3088 -150
rect -4408 -286 -3896 -242
rect -3328 -272 -3188 -166
rect -3098 -272 -3088 -166
rect -3328 -286 -3088 -272
rect -4408 -288 -4126 -286
rect 15188 -413 15379 664
rect 15542 437 15612 664
rect 13001 -509 15379 -413
rect 13001 -575 15306 -509
rect 12540 -744 12611 -637
rect 12971 -707 15306 -575
rect 12971 -744 13037 -707
rect 12540 -770 13037 -744
rect 12015 -780 13037 -770
rect 12015 -818 13008 -780
rect 11831 -822 13008 -818
rect 11831 -869 12089 -822
rect 12540 -824 13008 -822
rect 12540 -825 12611 -824
rect 11942 -1060 12008 -1059
rect 12044 -1060 12089 -869
rect 16178 -884 16248 -592
rect 16174 -895 16289 -884
rect 12778 -975 16289 -895
rect 11942 -1092 12121 -1060
rect 11942 -1093 12008 -1092
rect 11883 -2912 11917 -1127
rect 12001 -1176 12035 -1127
rect 12090 -1176 12121 -1092
rect 12001 -1214 12121 -1176
rect 12778 -1114 12894 -975
rect 12778 -1204 12780 -1114
rect 12886 -1204 12894 -1114
rect 16174 -1152 16289 -975
rect 66364 -890 66598 -876
rect 66364 -1028 66390 -890
rect 66564 -1028 66598 -890
rect 66364 -1088 66598 -1028
rect 16178 -1160 16248 -1152
rect 12778 -1214 12894 -1204
rect 12001 -2469 12035 -1214
rect 12090 -1215 12121 -1214
rect 65290 -1750 67452 -1088
rect 65280 -2712 67406 -2156
rect 11169 -3006 11380 -3004
rect 11169 -3112 11179 -3006
rect 11269 -3112 11380 -3006
rect 11169 -3120 11380 -3112
rect 11300 -3404 11380 -3120
rect 11300 -3446 11310 -3404
rect 11370 -3446 11380 -3404
rect 11300 -3466 11380 -3446
rect 11846 -4448 11998 -2912
rect 66596 -3066 66804 -2712
rect 66590 -3170 66824 -3066
rect 66590 -3308 66624 -3170
rect 66798 -3308 66824 -3170
rect 66590 -3322 66824 -3308
rect 11846 -4564 11866 -4448
rect 11980 -4564 11998 -4448
rect 11846 -4590 11998 -4564
rect -3624 -5226 -3390 -5212
rect -3624 -5364 -3598 -5226
rect -3424 -5364 -3390 -5226
rect -3624 -5542 -3390 -5364
rect -4602 -6002 -2808 -5542
rect -4622 -6702 -2828 -6242
rect -3810 -7236 -3576 -6702
rect -3810 -7374 -3776 -7236
rect -3602 -7374 -3576 -7236
rect -3810 -7388 -3576 -7374
<< via1 >>
rect -1320 18086 -26 19058
rect 4738 12912 5000 13200
rect -10146 6888 -10070 6974
rect -2736 3054 -2646 3160
rect -3188 -272 -3098 -166
rect 12780 -1204 12886 -1114
rect 66390 -1028 66564 -890
rect 11179 -3112 11269 -3006
rect 66624 -3308 66798 -3170
rect -3598 -5364 -3424 -5226
rect -3776 -7374 -3602 -7236
<< metal2 >>
rect -1548 22396 300 22466
rect -1548 21500 -1250 22396
rect 158 21500 300 22396
rect -1548 19058 300 21500
rect -1548 18086 -1320 19058
rect -26 18086 300 19058
rect -1548 17946 300 18086
rect 4680 13790 5054 13830
rect 4680 13564 4738 13790
rect 4994 13564 5054 13790
rect 4680 13200 5054 13564
rect 4680 12912 4738 13200
rect 5000 12912 5054 13200
rect 4680 12840 5054 12912
rect -10172 7430 -10054 7442
rect -10172 7370 -10150 7430
rect -10070 7370 -10054 7430
rect -10172 6974 -10054 7370
rect -10172 6888 -10146 6974
rect -10070 6888 -10054 6974
rect -10172 6866 -10054 6888
rect -2752 3160 -2080 3176
rect -2752 3054 -2736 3160
rect -2646 3156 -2080 3160
rect -2646 3056 -2172 3156
rect -2090 3056 -2080 3156
rect -2646 3054 -2080 3056
rect -2752 3042 -2080 3054
rect -3204 -166 -2532 -150
rect -3204 -272 -3188 -166
rect -3098 -170 -2532 -166
rect -3098 -270 -2624 -170
rect -2542 -270 -2532 -170
rect -3098 -272 -2532 -270
rect -3204 -284 -2532 -272
rect 66360 -346 66624 -314
rect 66360 -484 66420 -346
rect 66576 -484 66624 -346
rect 66360 -890 66624 -484
rect 66360 -1028 66390 -890
rect 66564 -1028 66624 -890
rect 66360 -1066 66624 -1028
rect 12768 -1114 12902 -1098
rect 12768 -1204 12780 -1114
rect 12886 -1204 12902 -1114
rect 12768 -1678 12902 -1204
rect 12768 -1760 12782 -1678
rect 12882 -1760 12902 -1678
rect 12768 -1770 12902 -1760
rect 10613 -3006 11285 -2994
rect 10613 -3008 11179 -3006
rect 10613 -3108 10623 -3008
rect 10705 -3108 11179 -3008
rect 10613 -3112 11179 -3108
rect 11269 -3112 11285 -3006
rect 10613 -3128 11285 -3112
rect 66564 -3170 66828 -3132
rect 66564 -3308 66624 -3170
rect 66798 -3308 66828 -3170
rect 66564 -3714 66828 -3308
rect 66564 -3852 66612 -3714
rect 66768 -3852 66828 -3714
rect 66564 -3884 66828 -3852
rect -3628 -4682 -3364 -4650
rect -3628 -4820 -3568 -4682
rect -3412 -4820 -3364 -4682
rect -3628 -5226 -3364 -4820
rect -3628 -5364 -3598 -5226
rect -3424 -5364 -3364 -5226
rect -3628 -5402 -3364 -5364
rect -3836 -7236 -3572 -7198
rect -3836 -7374 -3776 -7236
rect -3602 -7374 -3572 -7236
rect -3836 -7780 -3572 -7374
rect -3836 -7918 -3788 -7780
rect -3632 -7918 -3572 -7780
rect -3836 -7950 -3572 -7918
<< via2 >>
rect -1250 21500 158 22396
rect 4738 13564 4994 13790
rect -10150 7370 -10070 7430
rect -2172 3056 -2090 3156
rect -2624 -270 -2542 -170
rect 66420 -484 66576 -346
rect 12782 -1760 12882 -1678
rect 10623 -3108 10705 -3008
rect 66612 -3852 66768 -3714
rect -3568 -4820 -3412 -4682
rect -3788 -7918 -3632 -7780
<< metal3 >>
rect -1942 33954 924 34392
rect -1942 32098 -1572 33954
rect 588 32098 924 33954
rect -1942 29400 924 32098
rect -1942 29264 934 29400
rect -1932 26332 934 29264
rect -1936 24272 934 26332
rect -1936 22396 930 24272
rect -1936 21500 -1250 22396
rect 158 21500 930 22396
rect -1936 21204 930 21500
rect 4682 14332 5048 14370
rect 4682 14114 4748 14332
rect 4982 14114 5048 14332
rect 4682 13790 5048 14114
rect 4682 13564 4738 13790
rect 4994 13564 5048 13790
rect 4682 13500 5048 13564
rect -10168 7804 -10044 7816
rect -10168 7740 -10146 7804
rect -10066 7740 -10044 7804
rect -10168 7430 -10044 7740
rect -10168 7370 -10150 7430
rect -10070 7370 -10044 7430
rect -10168 7352 -10044 7370
rect -2188 3156 -1704 3170
rect -2188 3056 -2172 3156
rect -2090 3148 -1704 3156
rect -2090 3056 -1792 3148
rect -2188 3048 -1792 3056
rect -1710 3048 -1704 3148
rect -2188 3042 -1704 3048
rect 66390 58 66630 80
rect 66390 -62 66442 58
rect 66582 -62 66630 58
rect -2640 -170 -2156 -156
rect -2640 -270 -2624 -170
rect -2542 -178 -2156 -170
rect -2542 -270 -2244 -178
rect -2640 -278 -2244 -270
rect -2162 -278 -2156 -178
rect 66390 -246 66630 -62
rect -2640 -284 -2156 -278
rect 66386 -346 66632 -246
rect 66386 -484 66420 -346
rect 66576 -484 66632 -346
rect 66386 -528 66632 -484
rect 12768 -1678 12896 -1662
rect 12768 -1760 12782 -1678
rect 12882 -1760 12896 -1678
rect 12768 -2058 12896 -1760
rect 12768 -2140 12774 -2058
rect 12874 -2140 12896 -2058
rect 12768 -2146 12896 -2140
rect 10237 -3000 10721 -2994
rect 10237 -3100 10243 -3000
rect 10325 -3008 10721 -3000
rect 10325 -3100 10623 -3008
rect 10237 -3108 10623 -3100
rect 10705 -3108 10721 -3008
rect 10237 -3122 10721 -3108
rect 66556 -3714 66802 -3670
rect 66556 -3852 66612 -3714
rect 66768 -3852 66802 -3714
rect 66556 -3952 66802 -3852
rect 66558 -4136 66798 -3952
rect 66558 -4256 66606 -4136
rect 66746 -4256 66798 -4136
rect -3598 -4278 -3358 -4256
rect 66558 -4278 66798 -4256
rect -3598 -4398 -3546 -4278
rect -3406 -4398 -3358 -4278
rect -3598 -4582 -3358 -4398
rect -3602 -4682 -3356 -4582
rect -3602 -4820 -3568 -4682
rect -3412 -4820 -3356 -4682
rect -3602 -4864 -3356 -4820
rect -3844 -7780 -3598 -7736
rect -3844 -7918 -3788 -7780
rect -3632 -7918 -3598 -7780
rect -3844 -8234 -3598 -7918
rect -3848 -8286 -3598 -8234
rect -3848 -8542 -3602 -8286
rect -3848 -8752 -3840 -8542
rect -3610 -8752 -3602 -8542
rect -3848 -8784 -3602 -8752
<< via3 >>
rect -1572 32098 588 33954
rect 4748 14114 4982 14332
rect -10146 7740 -10066 7804
rect -1792 3048 -1710 3148
rect 66442 -62 66582 58
rect -2244 -278 -2162 -178
rect 12774 -2140 12874 -2058
rect 10243 -3100 10325 -3000
rect 66606 -4256 66746 -4136
rect -3546 -4398 -3406 -4278
rect -3840 -8752 -3610 -8542
<< metal4 >>
rect -13386 54436 -11282 54590
rect -13386 52230 -13232 54436
rect -11540 52230 -11282 54436
rect -13386 26930 -11282 52230
rect -2874 33954 1832 42862
rect -2874 32098 -1572 33954
rect 588 32098 1832 33954
rect -2874 31566 1832 32098
rect 9000 26950 9318 26958
rect 4024 26946 9318 26950
rect 1880 26930 9318 26946
rect -13386 26352 9318 26930
rect -13386 26286 4644 26352
rect -13386 25482 1978 26286
rect -13386 15040 -11282 25482
rect 9000 23118 9318 26352
rect 16060 23290 16738 23780
rect 16030 23286 16738 23290
rect 13764 23162 16738 23286
rect 13764 23160 16210 23162
rect 8958 23036 12366 23118
rect 8958 22928 9068 23036
rect 10130 22892 10234 23036
rect 11300 22920 11402 23036
rect 12192 23034 12366 23036
rect 4708 19556 5026 19562
rect 8448 19556 8558 19696
rect 4708 19482 8558 19556
rect 9622 19482 9732 19704
rect 10790 19482 10900 19698
rect 4708 19396 10900 19482
rect 12224 19462 12366 23034
rect 13764 22928 13868 23160
rect 14936 22928 15038 23160
rect 16106 22928 16210 23160
rect 13332 19718 13358 19722
rect 13252 19462 13362 19716
rect 14422 19462 14532 19704
rect 15596 19462 15700 19708
rect 12224 19458 15700 19462
rect 4708 19018 5026 19396
rect 8448 19392 10900 19396
rect 12222 19336 15700 19458
rect 12222 19334 13246 19336
rect 12222 19240 12376 19334
rect 4708 18678 11736 19018
rect 4708 15760 5026 18678
rect 123252 16322 124372 27360
rect 118390 15820 124874 16322
rect 113334 15818 124874 15820
rect 4708 15750 5036 15760
rect -13386 14642 -10034 15040
rect 4698 14658 5036 15750
rect -13386 14624 -11282 14642
rect -10164 7966 -10070 14642
rect 4688 14332 5036 14658
rect 112330 15472 124874 15818
rect 112330 14506 113602 15472
rect 118390 15434 124874 15472
rect 4688 14114 4748 14332
rect 4982 14114 5036 14332
rect 4688 14026 5036 14114
rect 4688 14004 5010 14026
rect 111288 13734 113602 14506
rect 110206 13272 113602 13734
rect 110206 12770 112560 13272
rect 109396 11960 112560 12770
rect 109396 11188 111478 11960
rect 109396 11034 110668 11188
rect 107892 10224 110668 11034
rect 107892 8448 109976 10224
rect -10164 7804 -10040 7966
rect -10164 7740 -10146 7804
rect -10066 7740 -10040 7804
rect -10164 7726 -10040 7740
rect 105806 7058 109976 8448
rect 105806 6018 109588 7058
rect -1804 3148 -1643 3158
rect -1804 3048 -1792 3148
rect -1710 3048 -1643 3148
rect -1804 3038 -1643 3048
rect -1803 2938 -1647 3038
rect 1404 2982 1685 3201
rect 598 2940 1685 2982
rect 596 2938 1685 2940
rect -2053 2911 1685 2938
rect -2053 2849 659 2911
rect -1482 2770 -1378 2849
rect -464 2771 -360 2849
rect 544 2771 659 2849
rect -1923 -168 -1813 -44
rect -2256 -172 -1813 -168
rect -903 -172 -799 -47
rect 116 -172 220 -47
rect -2256 -178 686 -172
rect -2256 -278 -2244 -178
rect -2162 -278 686 -178
rect -2256 -288 686 -278
rect -1840 -608 -1503 -288
rect -7700 -769 -1503 -608
rect -7700 -1431 -7640 -769
rect -6676 -1431 -1503 -769
rect -7700 -1552 -1503 -1431
rect -1840 -1553 -1503 -1552
rect 1404 -3215 1685 2911
rect 103144 2774 109588 6018
rect 103144 2428 106926 2774
rect 100364 884 106926 2428
rect 66410 344 106926 884
rect 66410 58 104418 344
rect 66410 -62 66442 58
rect 66582 -62 104418 58
rect 66410 -94 104418 -62
rect 66416 -96 66634 -94
rect 12764 -2058 12884 -2046
rect 12764 -2140 12774 -2058
rect 12874 -2140 12884 -2058
rect 12764 -2249 12884 -2140
rect 12752 -2519 12939 -2249
rect 12698 -2665 12939 -2519
rect 3171 -2978 5778 -2970
rect 3171 -2990 10134 -2978
rect 3171 -3000 10337 -2990
rect 3171 -3057 10243 -3000
rect -3094 -3954 1711 -3215
rect 3171 -3425 3243 -3057
rect 3561 -3100 10243 -3057
rect 10325 -3100 10337 -3000
rect 3561 -3110 10337 -3100
rect 3561 -3165 10134 -3110
rect 12698 -3127 12914 -2665
rect 3561 -3425 5778 -3165
rect 3171 -3483 5778 -3425
rect -3572 -4078 1711 -3954
rect -3572 -4278 -3354 -4078
rect -3094 -4109 1711 -4078
rect -3572 -4398 -3546 -4278
rect -3406 -4398 -3354 -4278
rect -3572 -4432 -3354 -4398
rect -3594 -9656 -3128 -8516
rect -4016 -11684 -3126 -9656
rect -3608 -11702 -3126 -11684
rect -3606 -11707 -3126 -11702
rect 12347 -11292 12982 -3127
rect 100364 -3516 104418 -94
rect 66554 -4136 66772 -4102
rect 66554 -4256 66606 -4136
rect 66746 -4256 66772 -4136
rect 66554 -4300 66772 -4256
rect 58578 -4906 66808 -4300
rect 12347 -11697 12401 -11292
rect 12941 -11697 12982 -11292
rect 12347 -11751 12982 -11697
rect 58551 -5072 66808 -4906
rect 3806 -12852 4130 -12825
rect 58551 -12852 59016 -5072
rect 3755 -13273 59016 -12852
rect 3755 -13290 58709 -13273
rect 3806 -14863 4130 -13290
rect 3806 -14876 9858 -14863
rect 3433 -14978 9858 -14876
rect 3433 -14990 9891 -14978
rect 4266 -15282 4369 -14990
rect 6109 -15281 6213 -14990
rect 7947 -15280 8051 -14990
rect 9787 -15281 9891 -14990
rect 3447 -22395 3538 -22151
rect 3440 -22399 3897 -22395
rect 5291 -22399 5382 -22151
rect 7127 -22399 7218 -22152
rect 8960 -22399 9051 -22152
rect 3440 -22533 9924 -22399
rect 5005 -23084 5301 -22533
rect 4768 -23822 5588 -23084
<< via4 >>
rect -13232 52230 -11540 54436
rect -7640 -1431 -6676 -769
rect 3243 -3425 3561 -3057
rect 12401 -11697 12941 -11292
<< metal5 >>
rect -13406 54436 -11402 71972
rect -13406 52230 -13232 54436
rect -11540 52230 -11402 54436
rect -13406 51910 -11402 52230
rect -39997 -769 -6516 -611
rect -39997 -1431 -7640 -769
rect -6676 -1431 -6516 -769
rect -39997 -1590 -6516 -1431
rect -39997 -28361 -38928 -1590
rect 3192 -3057 3605 -2971
rect 3192 -3425 3243 -3057
rect 3561 -3425 3605 -3057
rect 3192 -5356 3605 -3425
rect 3238 -8176 3542 -5356
rect 3192 -8829 3605 -8176
rect 973 -8830 3605 -8829
rect -54 -8860 3605 -8830
rect -76 -9405 3605 -8860
rect -76 -9696 1186 -9405
rect 3192 -9407 3605 -9405
rect -76 -13282 720 -9696
rect 1748 -11292 12999 -11213
rect 1748 -11383 12401 -11292
rect 1662 -11697 12401 -11383
rect 12941 -11697 12999 -11292
rect 1662 -11769 12999 -11697
rect 1662 -28336 2090 -11769
rect 116008 -27840 117384 -21302
rect 64578 -28336 117384 -27840
rect -34584 -28361 117384 -28336
rect -40004 -29554 117384 -28361
rect -40004 -29561 117136 -29554
rect -40004 -29567 -34519 -29561
rect 64578 -29788 117136 -29561
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC1
timestamp 1667951165
transform 1 0 9723 0 1 21290
box -1711 -1620 1710 1640
use sky130_fd_pr__cap_mim_m3_1_FLZ2GZ  XC3
timestamp 1667951165
transform 1 0 6250 0 1 -18718
box -3568 -3440 3668 3440
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC4
timestamp 1667951165
transform 1 0 14527 0 1 21308
box -1711 -1620 1710 1640
use sky130_fd_pr__nfet_01v8_TAQE79  XM2
timestamp 1668019001
transform 1 0 -9997 0 1 2956
box -257 -2568 257 2568
use sky130_fd_pr__nfet_01v8_PAV6Y8  XM3
timestamp 1668017392
transform 1 0 11959 0 1 -1798
box -88 -755 88 755
use lg  lg_0
timestamp 1668127436
transform -1 0 114306 0 1 61558
box -81282 -83494 47246 55400
use lm  lm_0
timestamp 1668127496
transform 1 0 -6766 0 1 63380
box -63884 -36962 58600 50000
use ls  ls_0
timestamp 1668200762
transform 1 0 -2482 0 1 302
box -34810 -19320 2606 -3320
use sky130_fd_pr__cap_mim_m3_1_LJH8TW  sky130_fd_pr__cap_mim_m3_1_LJH8TW_1
timestamp 1667951165
transform 1 0 -801 0 1 1362
box -1489 -1410 1488 1410
use sky130_fd_pr__nfet_01v8_TAQE79  sky130_fd_pr__nfet_01v8_TAQE79_0
timestamp 1668019001
transform 1 0 -4155 0 1 2360
box -257 -2568 257 2568
use sky130_fd_pr__res_xhigh_po_0p35_BZ5JJG  sky130_fd_pr__res_xhigh_po_0p35_BZ5JJG_0
timestamp 1667951165
transform -1 0 15895 0 -1 -91
box -355 -589 355 589
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_0
timestamp 1667951165
transform -1 0 12576 0 1 -217
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_1
timestamp 1667951165
transform -1 0 12769 0 1 10908
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_2
timestamp 1667951165
transform -1 0 13345 0 1 10906
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_3
timestamp 1667951165
transform -1 0 13869 0 1 10898
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_4
timestamp 1667951165
transform -1 0 14403 0 1 10888
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_5
timestamp 1667951165
transform -1 0 -3519 0 1 -6142
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_6
timestamp 1667951165
transform -1 0 -2969 0 1 -6140
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_7
timestamp 1667951165
transform -1 0 -4001 0 1 -6122
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_8
timestamp 1667951165
transform -1 0 -4565 0 1 -6130
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_9
timestamp 1667951165
transform -1 0 65353 0 1 -1958
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_10
timestamp 1667951165
transform -1 0 65859 0 1 -1984
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_11
timestamp 1667951165
transform -1 0 66575 0 1 -1964
box -37 -502 37 502
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_12
timestamp 1667951165
transform -1 0 67273 0 1 -1990
box -37 -502 37 502
<< labels >>
rlabel metal4 16310 23440 16548 23660 1 RFOUT
port 1 n
rlabel metal4 4768 -23822 5588 -23084 1 RFIN
port 2 n
rlabel metal1 20408 4420 23150 6956 1 VDD
port 4 n
rlabel psubdiffcont 10770 -5214 11494 -4560 1 GND
port 3 n
<< end >>
