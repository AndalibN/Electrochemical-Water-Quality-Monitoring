magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< error_p >>
rect -78 2581 -20 2587
rect 118 2581 176 2587
rect -78 2547 -66 2581
rect 118 2547 130 2581
rect -78 2541 -20 2547
rect 118 2541 176 2547
rect -176 -2547 -118 -2541
rect 20 -2547 78 -2541
rect -176 -2581 -164 -2547
rect 20 -2581 32 -2547
rect -176 -2587 -118 -2581
rect 20 -2587 78 -2581
<< nwell >>
rect -163 2562 261 2600
rect -261 -2562 261 2562
rect -261 -2600 163 -2562
<< pmos >>
rect -167 -2500 -127 2500
rect -69 -2500 -29 2500
rect 29 -2500 69 2500
rect 127 -2500 167 2500
<< pdiff >>
rect -225 2488 -167 2500
rect -225 -2488 -213 2488
rect -179 -2488 -167 2488
rect -225 -2500 -167 -2488
rect -127 2488 -69 2500
rect -127 -2488 -115 2488
rect -81 -2488 -69 2488
rect -127 -2500 -69 -2488
rect -29 2488 29 2500
rect -29 -2488 -17 2488
rect 17 -2488 29 2488
rect -29 -2500 29 -2488
rect 69 2488 127 2500
rect 69 -2488 81 2488
rect 115 -2488 127 2488
rect 69 -2500 127 -2488
rect 167 2488 225 2500
rect 167 -2488 179 2488
rect 213 -2488 225 2488
rect 167 -2500 225 -2488
<< pdiffc >>
rect -213 -2488 -179 2488
rect -115 -2488 -81 2488
rect -17 -2488 17 2488
rect 81 -2488 115 2488
rect 179 -2488 213 2488
<< poly >>
rect -82 2581 -16 2597
rect -82 2547 -66 2581
rect -32 2547 -16 2581
rect -82 2531 -16 2547
rect 114 2581 180 2597
rect 114 2547 130 2581
rect 164 2547 180 2581
rect 114 2531 180 2547
rect -167 2500 -127 2526
rect -69 2500 -29 2531
rect 29 2500 69 2526
rect 127 2500 167 2531
rect -167 -2531 -127 -2500
rect -69 -2526 -29 -2500
rect 29 -2531 69 -2500
rect 127 -2526 167 -2500
rect -180 -2547 -114 -2531
rect -180 -2581 -164 -2547
rect -130 -2581 -114 -2547
rect -180 -2597 -114 -2581
rect 16 -2547 82 -2531
rect 16 -2581 32 -2547
rect 66 -2581 82 -2547
rect 16 -2597 82 -2581
<< polycont >>
rect -66 2547 -32 2581
rect 130 2547 164 2581
rect -164 -2581 -130 -2547
rect 32 -2581 66 -2547
<< locali >>
rect -82 2547 -66 2581
rect -32 2547 -16 2581
rect 114 2547 130 2581
rect 164 2547 180 2581
rect -213 2488 -179 2504
rect -213 -2504 -179 -2488
rect -115 2488 -81 2504
rect -115 -2504 -81 -2488
rect -17 2488 17 2504
rect -17 -2504 17 -2488
rect 81 2488 115 2504
rect 81 -2504 115 -2488
rect 179 2488 213 2504
rect 179 -2504 213 -2488
rect -180 -2581 -164 -2547
rect -130 -2581 -114 -2547
rect 16 -2581 32 -2547
rect 66 -2581 82 -2547
<< viali >>
rect -66 2547 -32 2581
rect 130 2547 164 2581
rect -213 -2488 -179 2488
rect -115 -2488 -81 2488
rect -17 -2488 17 2488
rect 81 -2488 115 2488
rect 179 -2488 213 2488
rect -164 -2581 -130 -2547
rect 32 -2581 66 -2547
<< metal1 >>
rect -78 2581 -20 2587
rect -78 2547 -66 2581
rect -32 2547 -20 2581
rect -78 2541 -20 2547
rect 118 2581 176 2587
rect 118 2547 130 2581
rect 164 2547 176 2581
rect 118 2541 176 2547
rect -219 2488 -173 2500
rect -219 -2488 -213 2488
rect -179 -2488 -173 2488
rect -219 -2500 -173 -2488
rect -121 2488 -75 2500
rect -121 -2488 -115 2488
rect -81 -2488 -75 2488
rect -121 -2500 -75 -2488
rect -23 2488 23 2500
rect -23 -2488 -17 2488
rect 17 -2488 23 2488
rect -23 -2500 23 -2488
rect 75 2488 121 2500
rect 75 -2488 81 2488
rect 115 -2488 121 2488
rect 75 -2500 121 -2488
rect 173 2488 219 2500
rect 173 -2488 179 2488
rect 213 -2488 219 2488
rect 173 -2500 219 -2488
rect -176 -2547 -118 -2541
rect -176 -2581 -164 -2547
rect -130 -2581 -118 -2547
rect -176 -2587 -118 -2581
rect 20 -2547 78 -2541
rect 20 -2581 32 -2547
rect 66 -2581 78 -2547
rect 20 -2587 78 -2581
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 25 l 0.2 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
