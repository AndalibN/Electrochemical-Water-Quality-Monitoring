magic
tech sky130A
timestamp 1668702877
<< pwell >>
rect -128 -21073 128 21073
<< nmos >>
rect -30 12668 30 20968
rect -30 4259 30 12559
rect -30 -4150 30 4150
rect -30 -12559 30 -4259
rect -30 -20968 30 -12668
<< ndiff >>
rect -59 20962 -30 20968
rect -59 12674 -53 20962
rect -36 12674 -30 20962
rect -59 12668 -30 12674
rect 30 20962 59 20968
rect 30 12674 36 20962
rect 53 12674 59 20962
rect 30 12668 59 12674
rect -59 12553 -30 12559
rect -59 4265 -53 12553
rect -36 4265 -30 12553
rect -59 4259 -30 4265
rect 30 12553 59 12559
rect 30 4265 36 12553
rect 53 4265 59 12553
rect 30 4259 59 4265
rect -59 4144 -30 4150
rect -59 -4144 -53 4144
rect -36 -4144 -30 4144
rect -59 -4150 -30 -4144
rect 30 4144 59 4150
rect 30 -4144 36 4144
rect 53 -4144 59 4144
rect 30 -4150 59 -4144
rect -59 -4265 -30 -4259
rect -59 -12553 -53 -4265
rect -36 -12553 -30 -4265
rect -59 -12559 -30 -12553
rect 30 -4265 59 -4259
rect 30 -12553 36 -4265
rect 53 -12553 59 -4265
rect 30 -12559 59 -12553
rect -59 -12674 -30 -12668
rect -59 -20962 -53 -12674
rect -36 -20962 -30 -12674
rect -59 -20968 -30 -20962
rect 30 -12674 59 -12668
rect 30 -20962 36 -12674
rect 53 -20962 59 -12674
rect 30 -20968 59 -20962
<< ndiffc >>
rect -53 12674 -36 20962
rect 36 12674 53 20962
rect -53 4265 -36 12553
rect 36 4265 53 12553
rect -53 -4144 -36 4144
rect 36 -4144 53 4144
rect -53 -12553 -36 -4265
rect 36 -12553 53 -4265
rect -53 -20962 -36 -12674
rect 36 -20962 53 -12674
<< psubdiff >>
rect -110 21038 -62 21055
rect 62 21038 110 21055
rect -110 21007 -93 21038
rect 93 21007 110 21038
rect -110 -21038 -93 -21007
rect 93 -21038 110 -21007
rect -110 -21055 -62 -21038
rect 62 -21055 110 -21038
<< psubdiffcont >>
rect -62 21038 62 21055
rect -110 -21007 -93 21007
rect 93 -21007 110 21007
rect -62 -21055 62 -21038
<< poly >>
rect -30 21004 30 21012
rect -30 20987 -22 21004
rect 22 20987 30 21004
rect -30 20968 30 20987
rect -30 12649 30 12668
rect -30 12632 -22 12649
rect 22 12632 30 12649
rect -30 12624 30 12632
rect -30 12595 30 12603
rect -30 12578 -22 12595
rect 22 12578 30 12595
rect -30 12559 30 12578
rect -30 4240 30 4259
rect -30 4223 -22 4240
rect 22 4223 30 4240
rect -30 4215 30 4223
rect -30 4186 30 4194
rect -30 4169 -22 4186
rect 22 4169 30 4186
rect -30 4150 30 4169
rect -30 -4169 30 -4150
rect -30 -4186 -22 -4169
rect 22 -4186 30 -4169
rect -30 -4194 30 -4186
rect -30 -4223 30 -4215
rect -30 -4240 -22 -4223
rect 22 -4240 30 -4223
rect -30 -4259 30 -4240
rect -30 -12578 30 -12559
rect -30 -12595 -22 -12578
rect 22 -12595 30 -12578
rect -30 -12603 30 -12595
rect -30 -12632 30 -12624
rect -30 -12649 -22 -12632
rect 22 -12649 30 -12632
rect -30 -12668 30 -12649
rect -30 -20987 30 -20968
rect -30 -21004 -22 -20987
rect 22 -21004 30 -20987
rect -30 -21012 30 -21004
<< polycont >>
rect -22 20987 22 21004
rect -22 12632 22 12649
rect -22 12578 22 12595
rect -22 4223 22 4240
rect -22 4169 22 4186
rect -22 -4186 22 -4169
rect -22 -4240 22 -4223
rect -22 -12595 22 -12578
rect -22 -12649 22 -12632
rect -22 -21004 22 -20987
<< locali >>
rect -110 21038 -62 21055
rect 62 21038 110 21055
rect -110 21007 -93 21038
rect 93 21007 110 21038
rect -30 20987 -22 21004
rect 22 20987 30 21004
rect -53 20962 -36 20970
rect -53 12666 -36 12674
rect 36 20962 53 20970
rect 36 12666 53 12674
rect -30 12632 -22 12649
rect 22 12632 30 12649
rect -30 12578 -22 12595
rect 22 12578 30 12595
rect -53 12553 -36 12561
rect -53 4257 -36 4265
rect 36 12553 53 12561
rect 36 4257 53 4265
rect -30 4223 -22 4240
rect 22 4223 30 4240
rect -30 4169 -22 4186
rect 22 4169 30 4186
rect -53 4144 -36 4152
rect -53 -4152 -36 -4144
rect 36 4144 53 4152
rect 36 -4152 53 -4144
rect -30 -4186 -22 -4169
rect 22 -4186 30 -4169
rect -30 -4240 -22 -4223
rect 22 -4240 30 -4223
rect -53 -4265 -36 -4257
rect -53 -12561 -36 -12553
rect 36 -4265 53 -4257
rect 36 -12561 53 -12553
rect -30 -12595 -22 -12578
rect 22 -12595 30 -12578
rect -30 -12649 -22 -12632
rect 22 -12649 30 -12632
rect -53 -12674 -36 -12666
rect -53 -20970 -36 -20962
rect 36 -12674 53 -12666
rect 36 -20970 53 -20962
rect -30 -21004 -22 -20987
rect 22 -21004 30 -20987
rect -110 -21038 -93 -21007
rect 93 -21038 110 -21007
rect -110 -21055 -62 -21038
rect 62 -21055 110 -21038
<< viali >>
rect -22 20987 22 21004
rect -53 12674 -36 20962
rect 36 12674 53 20962
rect -22 12632 22 12649
rect -22 12578 22 12595
rect -53 4265 -36 12553
rect 36 4265 53 12553
rect -22 4223 22 4240
rect -22 4169 22 4186
rect -53 -4144 -36 4144
rect 36 -4144 53 4144
rect -22 -4186 22 -4169
rect -22 -4240 22 -4223
rect -53 -12553 -36 -4265
rect 36 -12553 53 -4265
rect -22 -12595 22 -12578
rect -22 -12649 22 -12632
rect -53 -20962 -36 -12674
rect 36 -20962 53 -12674
rect -22 -21004 22 -20987
<< metal1 >>
rect -28 21004 28 21007
rect -28 20987 -22 21004
rect 22 20987 28 21004
rect -28 20984 28 20987
rect -56 20962 -33 20968
rect -56 12674 -53 20962
rect -36 12674 -33 20962
rect -56 12668 -33 12674
rect 33 20962 56 20968
rect 33 12674 36 20962
rect 53 12674 56 20962
rect 33 12668 56 12674
rect -28 12649 28 12652
rect -28 12632 -22 12649
rect 22 12632 28 12649
rect -28 12629 28 12632
rect -28 12595 28 12598
rect -28 12578 -22 12595
rect 22 12578 28 12595
rect -28 12575 28 12578
rect -56 12553 -33 12559
rect -56 4265 -53 12553
rect -36 4265 -33 12553
rect -56 4259 -33 4265
rect 33 12553 56 12559
rect 33 4265 36 12553
rect 53 4265 56 12553
rect 33 4259 56 4265
rect -28 4240 28 4243
rect -28 4223 -22 4240
rect 22 4223 28 4240
rect -28 4220 28 4223
rect -28 4186 28 4189
rect -28 4169 -22 4186
rect 22 4169 28 4186
rect -28 4166 28 4169
rect -56 4144 -33 4150
rect -56 -4144 -53 4144
rect -36 -4144 -33 4144
rect -56 -4150 -33 -4144
rect 33 4144 56 4150
rect 33 -4144 36 4144
rect 53 -4144 56 4144
rect 33 -4150 56 -4144
rect -28 -4169 28 -4166
rect -28 -4186 -22 -4169
rect 22 -4186 28 -4169
rect -28 -4189 28 -4186
rect -28 -4223 28 -4220
rect -28 -4240 -22 -4223
rect 22 -4240 28 -4223
rect -28 -4243 28 -4240
rect -56 -4265 -33 -4259
rect -56 -12553 -53 -4265
rect -36 -12553 -33 -4265
rect -56 -12559 -33 -12553
rect 33 -4265 56 -4259
rect 33 -12553 36 -4265
rect 53 -12553 56 -4265
rect 33 -12559 56 -12553
rect -28 -12578 28 -12575
rect -28 -12595 -22 -12578
rect 22 -12595 28 -12578
rect -28 -12598 28 -12595
rect -28 -12632 28 -12629
rect -28 -12649 -22 -12632
rect 22 -12649 28 -12632
rect -28 -12652 28 -12649
rect -56 -12674 -33 -12668
rect -56 -20962 -53 -12674
rect -36 -20962 -33 -12674
rect -56 -20968 -33 -20962
rect 33 -12674 56 -12668
rect 33 -20962 36 -12674
rect 53 -20962 56 -12674
rect 33 -20968 56 -20962
rect -28 -20987 28 -20984
rect -28 -21004 -22 -20987
rect 22 -21004 28 -20987
rect -28 -21007 28 -21004
<< properties >>
string FIXED_BBOX -101 -21046 101 21046
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 83.0 l 0.6 m 5 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
