magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -144 -357 144 295
<< nmos >>
rect -60 -331 60 269
<< ndiff >>
rect -118 224 -60 269
rect -118 190 -106 224
rect -72 190 -60 224
rect -118 156 -60 190
rect -118 122 -106 156
rect -72 122 -60 156
rect -118 88 -60 122
rect -118 54 -106 88
rect -72 54 -60 88
rect -118 20 -60 54
rect -118 -14 -106 20
rect -72 -14 -60 20
rect -118 -48 -60 -14
rect -118 -82 -106 -48
rect -72 -82 -60 -48
rect -118 -116 -60 -82
rect -118 -150 -106 -116
rect -72 -150 -60 -116
rect -118 -184 -60 -150
rect -118 -218 -106 -184
rect -72 -218 -60 -184
rect -118 -252 -60 -218
rect -118 -286 -106 -252
rect -72 -286 -60 -252
rect -118 -331 -60 -286
rect 60 224 118 269
rect 60 190 72 224
rect 106 190 118 224
rect 60 156 118 190
rect 60 122 72 156
rect 106 122 118 156
rect 60 88 118 122
rect 60 54 72 88
rect 106 54 118 88
rect 60 20 118 54
rect 60 -14 72 20
rect 106 -14 118 20
rect 60 -48 118 -14
rect 60 -82 72 -48
rect 106 -82 118 -48
rect 60 -116 118 -82
rect 60 -150 72 -116
rect 106 -150 118 -116
rect 60 -184 118 -150
rect 60 -218 72 -184
rect 106 -218 118 -184
rect 60 -252 118 -218
rect 60 -286 72 -252
rect 106 -286 118 -252
rect 60 -331 118 -286
<< ndiffc >>
rect -106 190 -72 224
rect -106 122 -72 156
rect -106 54 -72 88
rect -106 -14 -72 20
rect -106 -82 -72 -48
rect -106 -150 -72 -116
rect -106 -218 -72 -184
rect -106 -286 -72 -252
rect 72 190 106 224
rect 72 122 106 156
rect 72 54 106 88
rect 72 -14 106 20
rect 72 -82 106 -48
rect 72 -150 106 -116
rect 72 -218 106 -184
rect 72 -286 106 -252
<< poly >>
rect -60 341 60 357
rect -60 307 -17 341
rect 17 307 60 341
rect -60 269 60 307
rect -60 -357 60 -331
<< polycont >>
rect -17 307 17 341
<< locali >>
rect -60 307 -17 341
rect 17 307 60 341
rect -106 238 -72 273
rect -106 166 -72 190
rect -106 94 -72 122
rect -106 22 -72 54
rect -106 -48 -72 -14
rect -106 -116 -72 -84
rect -106 -184 -72 -156
rect -106 -252 -72 -228
rect -106 -335 -72 -300
rect 72 238 106 273
rect 72 166 106 190
rect 72 94 106 122
rect 72 22 106 54
rect 72 -48 106 -14
rect 72 -116 106 -84
rect 72 -184 106 -156
rect 72 -252 106 -228
rect 72 -335 106 -300
<< viali >>
rect -17 307 17 341
rect -106 224 -72 238
rect -106 204 -72 224
rect -106 156 -72 166
rect -106 132 -72 156
rect -106 88 -72 94
rect -106 60 -72 88
rect -106 20 -72 22
rect -106 -12 -72 20
rect -106 -82 -72 -50
rect -106 -84 -72 -82
rect -106 -150 -72 -122
rect -106 -156 -72 -150
rect -106 -218 -72 -194
rect -106 -228 -72 -218
rect -106 -286 -72 -266
rect -106 -300 -72 -286
rect 72 224 106 238
rect 72 204 106 224
rect 72 156 106 166
rect 72 132 106 156
rect 72 88 106 94
rect 72 60 106 88
rect 72 20 106 22
rect 72 -12 106 20
rect 72 -82 106 -50
rect 72 -84 106 -82
rect 72 -150 106 -122
rect 72 -156 106 -150
rect 72 -218 106 -194
rect 72 -228 106 -218
rect 72 -286 106 -266
rect 72 -300 106 -286
<< metal1 >>
rect -56 341 56 347
rect -56 307 -17 341
rect 17 307 56 341
rect -56 301 56 307
rect -112 238 -66 269
rect -112 204 -106 238
rect -72 204 -66 238
rect -112 166 -66 204
rect -112 132 -106 166
rect -72 132 -66 166
rect -112 94 -66 132
rect -112 60 -106 94
rect -72 60 -66 94
rect -112 22 -66 60
rect -112 -12 -106 22
rect -72 -12 -66 22
rect -112 -50 -66 -12
rect -112 -84 -106 -50
rect -72 -84 -66 -50
rect -112 -122 -66 -84
rect -112 -156 -106 -122
rect -72 -156 -66 -122
rect -112 -194 -66 -156
rect -112 -228 -106 -194
rect -72 -228 -66 -194
rect -112 -266 -66 -228
rect -112 -300 -106 -266
rect -72 -300 -66 -266
rect -112 -331 -66 -300
rect 66 238 112 269
rect 66 204 72 238
rect 106 204 112 238
rect 66 166 112 204
rect 66 132 72 166
rect 106 132 112 166
rect 66 94 112 132
rect 66 60 72 94
rect 106 60 112 94
rect 66 22 112 60
rect 66 -12 72 22
rect 106 -12 112 22
rect 66 -50 112 -12
rect 66 -84 72 -50
rect 106 -84 112 -50
rect 66 -122 112 -84
rect 66 -156 72 -122
rect 106 -156 112 -122
rect 66 -194 112 -156
rect 66 -228 72 -194
rect 106 -228 112 -194
rect 66 -266 112 -228
rect 66 -300 72 -266
rect 106 -300 112 -266
rect 66 -331 112 -300
<< end >>
