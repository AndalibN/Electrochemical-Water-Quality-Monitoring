magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -2346 6834 12460 7860
<< pwell >>
rect 3104 154 3411 557
rect -2278 -924 12580 154
<< psubdiff >>
rect 3130 316 3385 531
rect 3178 128 3347 316
rect -2252 -254 12554 128
rect -2252 -560 -1842 -254
rect 12200 -560 12554 -254
rect -2252 -898 12554 -560
<< nsubdiff >>
rect -2296 7814 -1974 7818
rect 12092 7814 12414 7818
rect -2296 7477 12414 7814
rect -2296 7171 -1964 7477
rect 12078 7171 12414 7477
rect -2296 6878 12414 7171
rect -1980 6876 12094 6878
<< psubdiffcont >>
rect -1842 -560 12200 -254
<< nsubdiffcont >>
rect -1964 7171 12078 7477
<< locali >>
rect -1980 7477 12094 7656
rect -1980 7171 -1964 7477
rect 12078 7171 12094 7477
rect -1980 7036 12094 7171
rect 3130 485 3385 531
rect 3130 316 3210 485
rect 3178 -46 3210 316
rect -2064 -254 3210 -46
rect 3316 316 3385 485
rect 6658 441 6922 504
rect 3316 -46 3347 316
rect 6658 276 6736 441
rect 6703 -46 6736 276
rect 3316 -241 6736 -46
rect 3316 -254 6021 -241
rect 6055 -254 6736 -241
rect 6842 276 6922 441
rect 6842 -46 6874 276
rect 6842 -254 12402 -46
rect -2064 -560 -1842 -254
rect 12200 -560 12402 -254
rect -2064 -563 6021 -560
rect 6055 -563 12402 -560
rect -2064 -738 12402 -563
<< viali >>
rect 4203 7218 4237 7252
rect 4275 7218 4309 7252
rect 4347 7218 4381 7252
rect 4540 7218 4574 7252
rect 4612 7218 4646 7252
rect 4684 7218 4718 7252
rect 3210 -254 3316 485
rect 6021 -254 6055 -241
rect 6736 -254 6842 441
rect 3210 -557 3316 -254
rect 6021 -275 6055 -254
rect 6021 -347 6055 -313
rect 6021 -419 6055 -385
rect 6021 -491 6055 -457
rect 6736 -529 6842 -254
rect 6021 -560 6055 -529
rect 6021 -563 6055 -560
<< metal1 >>
rect 4147 7252 4429 7304
rect 4147 7218 4203 7252
rect 4237 7218 4275 7252
rect 4309 7218 4347 7252
rect 4381 7218 4429 7252
rect 4147 7166 4429 7218
rect 4497 7252 4784 7304
rect 4497 7218 4540 7252
rect 4574 7218 4612 7252
rect 4646 7218 4684 7252
rect 4718 7218 4784 7252
rect 4497 7166 4784 7218
rect -2632 6718 -2404 6818
rect 3046 6733 3212 6756
rect 3046 6718 3071 6733
rect -2632 6636 3071 6718
rect -2632 6608 -2404 6636
rect 3046 6617 3071 6636
rect 3187 6617 3212 6733
rect 3046 6598 3212 6617
rect -2632 6498 -2406 6566
rect 3046 6515 3212 6538
rect 3046 6498 3071 6515
rect -2632 6424 3071 6498
rect -2632 6356 -2406 6424
rect 3046 6399 3071 6424
rect 3187 6399 3212 6515
rect 3046 6380 3212 6399
rect -2632 6246 -2408 6320
rect -2632 6172 3870 6246
rect -2632 6116 -2408 6172
rect 3798 4700 3870 6172
rect 4147 5705 4217 7166
rect 4272 6553 4438 6576
rect 4272 6437 4297 6553
rect 4413 6437 4438 6553
rect 4272 6418 4438 6437
rect 3898 5124 3984 5135
rect 3898 5072 3915 5124
rect 3967 5072 3984 5124
rect 3898 5036 3984 5072
rect 4147 5036 4217 5443
rect 3898 4986 4217 5036
rect 3898 4672 3941 4986
rect 4350 4692 4424 6418
rect 4713 5705 4783 7166
rect 13276 6728 13394 6758
rect 13448 6728 13604 6757
rect 13276 6726 13604 6728
rect 13276 6674 13303 6726
rect 13355 6674 13604 6726
rect 13276 6666 13604 6674
rect 13276 6642 13394 6666
rect 13448 6615 13604 6666
rect 13292 6387 13410 6412
rect 13491 6387 13715 6425
rect 13292 6380 13715 6387
rect 13292 6328 13319 6380
rect 13371 6328 13715 6380
rect 13292 6321 13715 6328
rect 13292 6296 13410 6321
rect 13491 6283 13715 6321
rect 5456 5781 5622 5804
rect 5456 5665 5481 5781
rect 5597 5665 5622 5781
rect 5456 5654 5622 5665
rect 5452 5646 5622 5654
rect 4452 5146 4549 5157
rect 4452 5094 4480 5146
rect 4532 5094 4549 5146
rect 4452 5043 4549 5094
rect 4713 5043 4783 5443
rect 4452 4993 4783 5043
rect 3752 890 3786 4659
rect 3882 1071 3941 4672
rect 4037 890 4071 4659
rect 4452 4647 4494 4993
rect 5452 4658 5524 5646
rect 5700 5085 5781 5095
rect 5700 5033 5715 5085
rect 5767 5033 5781 5085
rect 5700 4839 5781 5033
rect 5586 4802 5880 4839
rect 4305 890 4339 4647
rect 4435 1059 4494 4647
rect 4590 891 4624 4647
rect 5246 909 5318 912
rect 5246 891 5255 909
rect 4590 890 5255 891
rect 3752 857 5255 890
rect 5307 857 5318 909
rect 3752 850 5318 857
rect 5406 863 5440 4615
rect 5586 1027 5620 4802
rect 5716 863 5750 4615
rect 5846 1028 5880 4802
rect 5976 863 6010 4615
rect 5406 814 6071 863
rect 3130 487 3390 536
rect 3130 371 3172 487
rect 3352 371 3390 487
rect 3130 316 3210 371
rect 3178 -557 3210 316
rect 3316 320 3390 371
rect 3316 316 3385 320
rect 3316 -557 3347 316
rect 3178 -582 3347 -557
rect 6005 -241 6071 814
rect 6658 491 6922 504
rect 6655 442 6922 491
rect 6655 326 6697 442
rect 6877 326 6922 442
rect 6655 275 6736 326
rect 6005 -275 6021 -241
rect 6055 -275 6071 -241
rect 6005 -313 6071 -275
rect 6005 -347 6021 -313
rect 6055 -347 6071 -313
rect 6005 -385 6071 -347
rect 6005 -419 6021 -385
rect 6055 -419 6071 -385
rect 6005 -457 6071 -419
rect 6005 -491 6021 -457
rect 6055 -491 6071 -457
rect 6005 -529 6071 -491
rect 6005 -563 6021 -529
rect 6055 -563 6071 -529
rect 6005 -582 6071 -563
rect 6703 -529 6736 275
rect 6842 276 6922 326
rect 6842 275 6915 276
rect 6842 -529 6874 275
rect 6703 -574 6874 -529
<< via1 >>
rect 3071 6617 3187 6733
rect 3071 6399 3187 6515
rect 4297 6437 4413 6553
rect 3915 5072 3967 5124
rect 13303 6674 13355 6726
rect 13319 6328 13371 6380
rect 5481 5665 5597 5781
rect 4480 5094 4532 5146
rect 5715 5033 5767 5085
rect 5255 857 5307 909
rect 3172 485 3352 487
rect 3172 371 3210 485
rect 3210 371 3316 485
rect 3316 371 3352 485
rect 6697 441 6877 442
rect 6697 326 6736 441
rect 6736 326 6842 441
rect 6842 326 6877 441
<< metal2 >>
rect 3046 6733 3212 6756
rect 3046 6617 3071 6733
rect 3187 6617 3212 6733
rect 3046 6598 3212 6617
rect 3372 6726 13374 6735
rect 3372 6674 13303 6726
rect 13355 6674 13374 6726
rect 3372 6605 13374 6674
rect 3046 6515 3212 6538
rect 3046 6399 3071 6515
rect 3187 6399 3212 6515
rect 3046 6380 3212 6399
rect 3372 6021 3984 6605
rect 4272 6553 4438 6576
rect 4272 6437 4297 6553
rect 4413 6437 4438 6553
rect 4272 6418 4438 6437
rect 4462 6380 13390 6402
rect 4462 6328 13319 6380
rect 13371 6328 13390 6380
rect 4462 6260 13390 6328
rect 3111 5124 3984 6021
rect 3111 5072 3915 5124
rect 3967 5072 3984 5124
rect 4463 5146 4549 6260
rect 5456 5781 5622 5804
rect 5456 5665 5481 5781
rect 5597 5665 5622 5781
rect 5456 5646 5622 5665
rect 4463 5094 4480 5146
rect 4532 5094 4549 5146
rect 4463 5078 4549 5094
rect 5249 5085 5781 5095
rect 3111 5055 3984 5072
rect 5249 5033 5715 5085
rect 5767 5033 5781 5085
rect 5249 5024 5781 5033
rect 5249 909 5315 5024
rect 5249 857 5255 909
rect 5307 857 5315 909
rect 5249 850 5315 857
rect 3124 496 3398 546
rect 3124 487 3192 496
rect 3328 487 3398 496
rect 3124 371 3172 487
rect 3352 371 3398 487
rect 3124 360 3192 371
rect 3328 360 3398 371
rect 3124 312 3398 360
rect 6649 451 6923 501
rect 6649 442 6717 451
rect 6853 442 6923 451
rect 6649 326 6697 442
rect 6877 326 6923 442
rect 6649 315 6717 326
rect 6853 315 6923 326
rect 6649 267 6923 315
<< via2 >>
rect 3101 6647 3157 6703
rect 3101 6429 3157 6485
rect 4327 6467 4383 6523
rect 5511 5695 5567 5751
rect 3192 487 3328 496
rect 3192 371 3328 487
rect 3192 360 3328 371
rect 6717 442 6853 451
rect 6717 326 6853 442
rect 6717 315 6853 326
<< metal3 >>
rect 3046 6703 3212 6756
rect 3046 6647 3101 6703
rect 3157 6696 3212 6703
rect 3157 6647 5574 6696
rect 3046 6636 5574 6647
rect 3046 6598 3212 6636
rect 3046 6518 3212 6538
rect 4272 6523 4438 6576
rect 4272 6518 4327 6523
rect 3046 6485 4327 6518
rect 3046 6429 3101 6485
rect 3157 6467 4327 6485
rect 4383 6467 4438 6523
rect 3157 6452 4438 6467
rect 3157 6429 3212 6452
rect 3046 6380 3212 6429
rect 4272 6418 4438 6452
rect 3112 5055 3376 6023
rect 5512 5804 5574 6636
rect 8041 6300 8938 6411
rect 5456 5751 5622 5804
rect 5456 5695 5511 5751
rect 5567 5695 5622 5751
rect 5456 5646 5622 5695
rect 3118 500 3404 556
rect 3118 356 3188 500
rect 3332 356 3404 500
rect 3118 304 3404 356
rect 6643 455 6929 511
rect 6643 311 6713 455
rect 6857 311 6929 455
rect 6643 259 6929 311
<< via3 >>
rect 3188 496 3332 500
rect 3188 360 3192 496
rect 3192 360 3328 496
rect 3328 360 3332 496
rect 3188 356 3332 360
rect 6713 451 6857 455
rect 6713 315 6717 451
rect 6717 315 6853 451
rect 6853 315 6857 451
rect 6713 311 6857 315
<< metal4 >>
rect 2674 5055 3377 6022
rect 8041 6005 8938 6413
rect 3110 500 3416 566
rect 3110 480 3188 500
rect 2882 415 3188 480
rect 3110 356 3188 415
rect 3332 356 3416 500
rect 3110 294 3416 356
rect 6635 455 7108 539
rect 6635 311 6713 455
rect 6857 443 7108 455
rect 6857 311 6941 443
rect 6635 249 6941 311
use sky130_fd_pr__cap_mim_m3_1_NXL3SG  XC1
timestamp 1669522153
transform 0 1 9852 -1 0 3330
box -2890 -2840 2889 2840
use sky130_fd_pr__cap_mim_m3_1_NXL3SG  XC2
timestamp 1669522153
transform 0 1 94 -1 0 3285
box -2890 -2840 2889 2840
use sky130_fd_pr__nfet_01v8_FKEGQS  sky130_fd_pr__nfet_01v8_FKEGQS_0
timestamp 1669522153
transform -1 0 3924 0 -1 2865
box -185 -1894 210 1894
use sky130_fd_pr__nfet_01v8_FKEGQS  sky130_fd_pr__nfet_01v8_FKEGQS_1
timestamp 1669522153
transform -1 0 4477 0 -1 2853
box -185 -1894 210 1894
use sky130_fd_pr__nfet_01v8_S6EGL7  sky130_fd_pr__nfet_01v8_S6EGL7_0
timestamp 1669522153
transform 1 0 5733 0 1 2821
box -365 -1893 315 1894
use sky130_fd_pr__res_high_po_0p35_FJ8ACL  sky130_fd_pr__res_high_po_0p35_FJ8ACL_0
timestamp 1669522153
transform 1 0 4748 0 1 5645
box -35 -492 35 492
use sky130_fd_pr__res_high_po_0p35_FJ8ACL  sky130_fd_pr__res_high_po_0p35_FJ8ACL_1
timestamp 1669522153
transform 1 0 4182 0 1 5645
box -35 -492 35 492
<< labels >>
rlabel mvpsubdiff s 5174 -397 5174 -397 4 GND
rlabel metal1 s 13448 6615 13604 6757 4 IF_P
port 1 nsew
rlabel metal1 s -2630 6610 -2406 6816 4 RF
port 2 nsew
rlabel metal1 s 13491 6283 13715 6425 4 IF_N
port 3 nsew
rlabel metal1 s -2630 6358 -2408 6562 4 LO_N
port 4 nsew
rlabel metal1 s -2630 6116 -2410 6318 4 LO_P
port 5 nsew
rlabel metal2 s 5259 1052 5301 1198 4 mid
port 6 nsew
rlabel nwell s -1982 7162 12088 7506 4 VDD
port 7 nsew
<< end >>
