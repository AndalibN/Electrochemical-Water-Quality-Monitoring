magic
tech sky130A
magscale 1 2
timestamp 1669755697
<< error_p >>
rect -442 5260 -384 5266
rect -442 5226 -430 5260
rect -442 5220 -384 5226
<< nmos >>
rect -443 -5188 -383 5188
rect -325 -5188 -265 5188
rect -207 -5188 -147 5188
rect -89 -5188 -29 5188
rect 29 -5188 89 5188
rect 147 -5188 207 5188
rect 265 -5188 325 5188
rect 383 -5188 443 5188
<< ndiff >>
rect -501 5176 -443 5188
rect -501 -5176 -489 5176
rect -455 -5176 -443 5176
rect -501 -5188 -443 -5176
rect -383 5176 -325 5188
rect -383 -5176 -371 5176
rect -337 -5176 -325 5176
rect -383 -5188 -325 -5176
rect -265 5176 -207 5188
rect -265 -5176 -253 5176
rect -219 -5176 -207 5176
rect -265 -5188 -207 -5176
rect -147 5176 -89 5188
rect -147 -5176 -135 5176
rect -101 -5176 -89 5176
rect -147 -5188 -89 -5176
rect -29 5176 29 5188
rect -29 -5176 -17 5176
rect 17 -5176 29 5176
rect -29 -5188 29 -5176
rect 89 5176 147 5188
rect 89 -5176 101 5176
rect 135 -5176 147 5176
rect 89 -5188 147 -5176
rect 207 5176 265 5188
rect 207 -5176 219 5176
rect 253 -5176 265 5176
rect 207 -5188 265 -5176
rect 325 5176 383 5188
rect 325 -5176 337 5176
rect 371 -5176 383 5176
rect 325 -5188 383 -5176
rect 443 5176 501 5188
rect 443 -5176 455 5176
rect 489 -5176 501 5176
rect 443 -5188 501 -5176
<< ndiffc >>
rect -489 -5176 -455 5176
rect -371 -5176 -337 5176
rect -253 -5176 -219 5176
rect -135 -5176 -101 5176
rect -17 -5176 17 5176
rect 101 -5176 135 5176
rect 219 -5176 253 5176
rect 337 -5176 371 5176
rect 455 -5176 489 5176
<< poly >>
rect -446 5260 -380 5276
rect -446 5226 -430 5260
rect -396 5226 -380 5260
rect -446 5210 -380 5226
rect -328 5266 -262 5276
rect -210 5266 -144 5276
rect -328 5220 -144 5266
rect -328 5210 -262 5220
rect -210 5210 -144 5220
rect -92 5266 -26 5276
rect 26 5266 92 5276
rect -92 5220 92 5266
rect -92 5210 -26 5220
rect 26 5210 92 5220
rect 144 5266 210 5276
rect 262 5266 328 5276
rect 144 5220 328 5266
rect 144 5210 210 5220
rect 262 5210 328 5220
rect 380 5210 446 5276
rect -443 5188 -383 5210
rect -325 5188 -265 5210
rect -207 5188 -147 5210
rect -89 5188 -29 5210
rect 29 5188 89 5210
rect 147 5188 207 5210
rect 265 5188 325 5210
rect 383 5188 443 5210
rect -443 -5210 -383 -5188
rect -325 -5210 -265 -5188
rect -207 -5210 -147 -5188
rect -89 -5210 -29 -5188
rect 29 -5210 89 -5188
rect 147 -5210 207 -5188
rect 265 -5210 325 -5188
rect 383 -5210 443 -5188
rect -446 -5220 -380 -5210
rect -328 -5220 -262 -5210
rect -446 -5266 -262 -5220
rect -446 -5276 -380 -5266
rect -328 -5276 -262 -5266
rect -210 -5220 -144 -5210
rect -92 -5220 -26 -5210
rect -210 -5266 -26 -5220
rect -210 -5276 -144 -5266
rect -92 -5276 -26 -5266
rect 26 -5220 92 -5210
rect 144 -5220 210 -5210
rect 26 -5266 210 -5220
rect 26 -5276 92 -5266
rect 144 -5276 210 -5266
rect 262 -5220 328 -5210
rect 380 -5220 446 -5210
rect 262 -5266 446 -5220
rect 262 -5276 328 -5266
rect 380 -5276 446 -5266
<< polycont >>
rect -430 5226 -396 5260
<< locali >>
rect -446 5226 -430 5260
rect -396 5226 -380 5260
rect -489 5176 -455 5192
rect -489 -5192 -455 -5176
rect -371 5176 -337 5192
rect -371 -5192 -337 -5176
rect -253 5176 -219 5192
rect -253 -5192 -219 -5176
rect -135 5176 -101 5192
rect -135 -5192 -101 -5176
rect -17 5176 17 5192
rect -17 -5192 17 -5176
rect 101 5176 135 5192
rect 101 -5192 135 -5176
rect 219 5176 253 5192
rect 219 -5192 253 -5176
rect 337 5176 371 5192
rect 337 -5192 371 -5176
rect 455 5176 489 5192
rect 455 -5192 489 -5176
<< viali >>
rect -430 5226 -396 5260
rect -489 -5176 -455 5176
rect -371 -5176 -337 5176
rect -253 -5176 -219 5176
rect -135 -5176 -101 5176
rect -17 -5176 17 5176
rect 101 -5176 135 5176
rect 219 -5176 253 5176
rect 337 -5176 371 5176
rect 455 -5176 489 5176
<< metal1 >>
rect -442 5260 -384 5266
rect -442 5226 -430 5260
rect -396 5226 -384 5260
rect -442 5220 -384 5226
rect -495 5176 -449 5188
rect -495 -5176 -489 5176
rect -455 -5176 -449 5176
rect -495 -5188 -449 -5176
rect -377 5176 -331 5188
rect -377 -5176 -371 5176
rect -337 -5176 -331 5176
rect -377 -5188 -331 -5176
rect -259 5176 -213 5188
rect -259 -5176 -253 5176
rect -219 -5176 -213 5176
rect -259 -5188 -213 -5176
rect -141 5176 -95 5188
rect -141 -5176 -135 5176
rect -101 -5176 -95 5176
rect -141 -5188 -95 -5176
rect -23 5176 23 5188
rect -23 -5176 -17 5176
rect 17 -5176 23 5176
rect -23 -5188 23 -5176
rect 95 5176 141 5188
rect 95 -5176 101 5176
rect 135 -5176 141 5176
rect 95 -5188 141 -5176
rect 213 5176 259 5188
rect 213 -5176 219 5176
rect 253 -5176 259 5176
rect 213 -5188 259 -5176
rect 331 5176 377 5188
rect 331 -5176 337 5176
rect 371 -5176 377 5176
rect 331 -5188 377 -5176
rect 449 5176 495 5188
rect 449 -5176 455 5176
rect 489 -5176 495 5176
rect 449 -5188 495 -5176
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 51.875 l 0.3 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
