magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 1200 35 1632
rect -35 -1632 35 -1200
<< xpolyres >>
rect -35 -1200 35 1200
<< viali >>
rect -17 1578 17 1612
rect -17 1506 17 1540
rect -17 1434 17 1468
rect -17 1362 17 1396
rect -17 1290 17 1324
rect -17 1218 17 1252
rect -17 -1253 17 -1219
rect -17 -1325 17 -1291
rect -17 -1397 17 -1363
rect -17 -1469 17 -1435
rect -17 -1541 17 -1507
rect -17 -1613 17 -1579
<< metal1 >>
rect -25 1612 25 1626
rect -25 1578 -17 1612
rect 17 1578 25 1612
rect -25 1540 25 1578
rect -25 1506 -17 1540
rect 17 1506 25 1540
rect -25 1468 25 1506
rect -25 1434 -17 1468
rect 17 1434 25 1468
rect -25 1396 25 1434
rect -25 1362 -17 1396
rect 17 1362 25 1396
rect -25 1324 25 1362
rect -25 1290 -17 1324
rect 17 1290 25 1324
rect -25 1252 25 1290
rect -25 1218 -17 1252
rect 17 1218 25 1252
rect -25 1205 25 1218
rect -25 -1219 25 -1205
rect -25 -1253 -17 -1219
rect 17 -1253 25 -1219
rect -25 -1291 25 -1253
rect -25 -1325 -17 -1291
rect 17 -1325 25 -1291
rect -25 -1363 25 -1325
rect -25 -1397 -17 -1363
rect 17 -1397 25 -1363
rect -25 -1435 25 -1397
rect -25 -1469 -17 -1435
rect 17 -1469 25 -1435
rect -25 -1507 25 -1469
rect -25 -1541 -17 -1507
rect 17 -1541 25 -1507
rect -25 -1579 25 -1541
rect -25 -1613 -17 -1579
rect 17 -1613 25 -1579
rect -25 -1626 25 -1613
<< end >>
