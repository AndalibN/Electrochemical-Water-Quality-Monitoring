magic
tech sky130A
timestamp 1667443905
<< nmos >>
rect -50 -1400 50 1400
<< ndiff >>
rect -79 1394 -50 1400
rect -79 -1394 -73 1394
rect -56 -1394 -50 1394
rect -79 -1400 -50 -1394
rect 50 1394 79 1400
rect 50 -1394 56 1394
rect 73 -1394 79 1394
rect 50 -1400 79 -1394
<< ndiffc >>
rect -73 -1394 -56 1394
rect 56 -1394 73 1394
<< poly >>
rect -50 1436 50 1444
rect -50 1419 -42 1436
rect 42 1419 50 1436
rect -50 1400 50 1419
rect -50 -1419 50 -1400
rect -50 -1436 -42 -1419
rect 42 -1436 50 -1419
rect -50 -1444 50 -1436
<< polycont >>
rect -42 1419 42 1436
rect -42 -1436 42 -1419
<< locali >>
rect -50 1419 -42 1436
rect 42 1419 50 1436
rect -73 1394 -56 1402
rect -73 -1402 -56 -1394
rect 56 1394 73 1402
rect 56 -1402 73 -1394
rect -50 -1436 -42 -1419
rect 42 -1436 50 -1419
<< viali >>
rect -42 1419 42 1436
rect -73 -1394 -56 1394
rect 56 -1394 73 1394
rect -42 -1436 42 -1419
<< metal1 >>
rect -48 1436 48 1439
rect -48 1419 -42 1436
rect 42 1419 48 1436
rect -48 1416 48 1419
rect -76 1394 -53 1400
rect -76 -1394 -73 1394
rect -56 -1394 -53 1394
rect -76 -1400 -53 -1394
rect 53 1394 76 1400
rect 53 -1394 56 1394
rect 73 -1394 76 1394
rect 53 -1400 76 -1394
rect -48 -1419 48 -1416
rect -48 -1436 -42 -1419
rect 42 -1436 48 -1419
rect -48 -1439 48 -1436
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 28.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
