magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 -1031 29 -1025
rect -29 -1065 -17 -1031
rect -29 -1071 29 -1065
<< nwell >>
rect -124 -1084 124 1118
<< pmos >>
rect -30 -984 30 1056
<< pdiff >>
rect -88 1039 -30 1056
rect -88 1005 -76 1039
rect -42 1005 -30 1039
rect -88 971 -30 1005
rect -88 937 -76 971
rect -42 937 -30 971
rect -88 903 -30 937
rect -88 869 -76 903
rect -42 869 -30 903
rect -88 835 -30 869
rect -88 801 -76 835
rect -42 801 -30 835
rect -88 767 -30 801
rect -88 733 -76 767
rect -42 733 -30 767
rect -88 699 -30 733
rect -88 665 -76 699
rect -42 665 -30 699
rect -88 631 -30 665
rect -88 597 -76 631
rect -42 597 -30 631
rect -88 563 -30 597
rect -88 529 -76 563
rect -42 529 -30 563
rect -88 495 -30 529
rect -88 461 -76 495
rect -42 461 -30 495
rect -88 427 -30 461
rect -88 393 -76 427
rect -42 393 -30 427
rect -88 359 -30 393
rect -88 325 -76 359
rect -42 325 -30 359
rect -88 291 -30 325
rect -88 257 -76 291
rect -42 257 -30 291
rect -88 223 -30 257
rect -88 189 -76 223
rect -42 189 -30 223
rect -88 155 -30 189
rect -88 121 -76 155
rect -42 121 -30 155
rect -88 87 -30 121
rect -88 53 -76 87
rect -42 53 -30 87
rect -88 19 -30 53
rect -88 -15 -76 19
rect -42 -15 -30 19
rect -88 -49 -30 -15
rect -88 -83 -76 -49
rect -42 -83 -30 -49
rect -88 -117 -30 -83
rect -88 -151 -76 -117
rect -42 -151 -30 -117
rect -88 -185 -30 -151
rect -88 -219 -76 -185
rect -42 -219 -30 -185
rect -88 -253 -30 -219
rect -88 -287 -76 -253
rect -42 -287 -30 -253
rect -88 -321 -30 -287
rect -88 -355 -76 -321
rect -42 -355 -30 -321
rect -88 -389 -30 -355
rect -88 -423 -76 -389
rect -42 -423 -30 -389
rect -88 -457 -30 -423
rect -88 -491 -76 -457
rect -42 -491 -30 -457
rect -88 -525 -30 -491
rect -88 -559 -76 -525
rect -42 -559 -30 -525
rect -88 -593 -30 -559
rect -88 -627 -76 -593
rect -42 -627 -30 -593
rect -88 -661 -30 -627
rect -88 -695 -76 -661
rect -42 -695 -30 -661
rect -88 -729 -30 -695
rect -88 -763 -76 -729
rect -42 -763 -30 -729
rect -88 -797 -30 -763
rect -88 -831 -76 -797
rect -42 -831 -30 -797
rect -88 -865 -30 -831
rect -88 -899 -76 -865
rect -42 -899 -30 -865
rect -88 -933 -30 -899
rect -88 -967 -76 -933
rect -42 -967 -30 -933
rect -88 -984 -30 -967
rect 30 1039 88 1056
rect 30 1005 42 1039
rect 76 1005 88 1039
rect 30 971 88 1005
rect 30 937 42 971
rect 76 937 88 971
rect 30 903 88 937
rect 30 869 42 903
rect 76 869 88 903
rect 30 835 88 869
rect 30 801 42 835
rect 76 801 88 835
rect 30 767 88 801
rect 30 733 42 767
rect 76 733 88 767
rect 30 699 88 733
rect 30 665 42 699
rect 76 665 88 699
rect 30 631 88 665
rect 30 597 42 631
rect 76 597 88 631
rect 30 563 88 597
rect 30 529 42 563
rect 76 529 88 563
rect 30 495 88 529
rect 30 461 42 495
rect 76 461 88 495
rect 30 427 88 461
rect 30 393 42 427
rect 76 393 88 427
rect 30 359 88 393
rect 30 325 42 359
rect 76 325 88 359
rect 30 291 88 325
rect 30 257 42 291
rect 76 257 88 291
rect 30 223 88 257
rect 30 189 42 223
rect 76 189 88 223
rect 30 155 88 189
rect 30 121 42 155
rect 76 121 88 155
rect 30 87 88 121
rect 30 53 42 87
rect 76 53 88 87
rect 30 19 88 53
rect 30 -15 42 19
rect 76 -15 88 19
rect 30 -49 88 -15
rect 30 -83 42 -49
rect 76 -83 88 -49
rect 30 -117 88 -83
rect 30 -151 42 -117
rect 76 -151 88 -117
rect 30 -185 88 -151
rect 30 -219 42 -185
rect 76 -219 88 -185
rect 30 -253 88 -219
rect 30 -287 42 -253
rect 76 -287 88 -253
rect 30 -321 88 -287
rect 30 -355 42 -321
rect 76 -355 88 -321
rect 30 -389 88 -355
rect 30 -423 42 -389
rect 76 -423 88 -389
rect 30 -457 88 -423
rect 30 -491 42 -457
rect 76 -491 88 -457
rect 30 -525 88 -491
rect 30 -559 42 -525
rect 76 -559 88 -525
rect 30 -593 88 -559
rect 30 -627 42 -593
rect 76 -627 88 -593
rect 30 -661 88 -627
rect 30 -695 42 -661
rect 76 -695 88 -661
rect 30 -729 88 -695
rect 30 -763 42 -729
rect 76 -763 88 -729
rect 30 -797 88 -763
rect 30 -831 42 -797
rect 76 -831 88 -797
rect 30 -865 88 -831
rect 30 -899 42 -865
rect 76 -899 88 -865
rect 30 -933 88 -899
rect 30 -967 42 -933
rect 76 -967 88 -933
rect 30 -984 88 -967
<< pdiffc >>
rect -76 1005 -42 1039
rect -76 937 -42 971
rect -76 869 -42 903
rect -76 801 -42 835
rect -76 733 -42 767
rect -76 665 -42 699
rect -76 597 -42 631
rect -76 529 -42 563
rect -76 461 -42 495
rect -76 393 -42 427
rect -76 325 -42 359
rect -76 257 -42 291
rect -76 189 -42 223
rect -76 121 -42 155
rect -76 53 -42 87
rect -76 -15 -42 19
rect -76 -83 -42 -49
rect -76 -151 -42 -117
rect -76 -219 -42 -185
rect -76 -287 -42 -253
rect -76 -355 -42 -321
rect -76 -423 -42 -389
rect -76 -491 -42 -457
rect -76 -559 -42 -525
rect -76 -627 -42 -593
rect -76 -695 -42 -661
rect -76 -763 -42 -729
rect -76 -831 -42 -797
rect -76 -899 -42 -865
rect -76 -967 -42 -933
rect 42 1005 76 1039
rect 42 937 76 971
rect 42 869 76 903
rect 42 801 76 835
rect 42 733 76 767
rect 42 665 76 699
rect 42 597 76 631
rect 42 529 76 563
rect 42 461 76 495
rect 42 393 76 427
rect 42 325 76 359
rect 42 257 76 291
rect 42 189 76 223
rect 42 121 76 155
rect 42 53 76 87
rect 42 -15 76 19
rect 42 -83 76 -49
rect 42 -151 76 -117
rect 42 -219 76 -185
rect 42 -287 76 -253
rect 42 -355 76 -321
rect 42 -423 76 -389
rect 42 -491 76 -457
rect 42 -559 76 -525
rect 42 -627 76 -593
rect 42 -695 76 -661
rect 42 -763 76 -729
rect 42 -831 76 -797
rect 42 -899 76 -865
rect 42 -967 76 -933
<< poly >>
rect -30 1056 30 1082
rect -30 -1015 30 -984
rect -33 -1031 33 -1015
rect -33 -1065 -17 -1031
rect 17 -1065 33 -1031
rect -33 -1081 33 -1065
<< polycont >>
rect -17 -1065 17 -1031
<< locali >>
rect -76 1039 -42 1060
rect -76 971 -42 991
rect -76 903 -42 919
rect -76 835 -42 847
rect -76 767 -42 775
rect -76 699 -42 703
rect -76 593 -42 597
rect -76 521 -42 529
rect -76 449 -42 461
rect -76 377 -42 393
rect -76 305 -42 325
rect -76 233 -42 257
rect -76 161 -42 189
rect -76 89 -42 121
rect -76 19 -42 53
rect -76 -49 -42 -17
rect -76 -117 -42 -89
rect -76 -185 -42 -161
rect -76 -253 -42 -233
rect -76 -321 -42 -305
rect -76 -389 -42 -377
rect -76 -457 -42 -449
rect -76 -525 -42 -521
rect -76 -631 -42 -627
rect -76 -703 -42 -695
rect -76 -775 -42 -763
rect -76 -847 -42 -831
rect -76 -919 -42 -899
rect -76 -988 -42 -967
rect 42 1039 76 1060
rect 42 971 76 991
rect 42 903 76 919
rect 42 835 76 847
rect 42 767 76 775
rect 42 699 76 703
rect 42 593 76 597
rect 42 521 76 529
rect 42 449 76 461
rect 42 377 76 393
rect 42 305 76 325
rect 42 233 76 257
rect 42 161 76 189
rect 42 89 76 121
rect 42 19 76 53
rect 42 -49 76 -17
rect 42 -117 76 -89
rect 42 -185 76 -161
rect 42 -253 76 -233
rect 42 -321 76 -305
rect 42 -389 76 -377
rect 42 -457 76 -449
rect 42 -525 76 -521
rect 42 -631 76 -627
rect 42 -703 76 -695
rect 42 -775 76 -763
rect 42 -847 76 -831
rect 42 -919 76 -899
rect 42 -988 76 -967
rect -33 -1065 -17 -1031
rect 17 -1065 33 -1031
<< viali >>
rect -76 1005 -42 1025
rect -76 991 -42 1005
rect -76 937 -42 953
rect -76 919 -42 937
rect -76 869 -42 881
rect -76 847 -42 869
rect -76 801 -42 809
rect -76 775 -42 801
rect -76 733 -42 737
rect -76 703 -42 733
rect -76 631 -42 665
rect -76 563 -42 593
rect -76 559 -42 563
rect -76 495 -42 521
rect -76 487 -42 495
rect -76 427 -42 449
rect -76 415 -42 427
rect -76 359 -42 377
rect -76 343 -42 359
rect -76 291 -42 305
rect -76 271 -42 291
rect -76 223 -42 233
rect -76 199 -42 223
rect -76 155 -42 161
rect -76 127 -42 155
rect -76 87 -42 89
rect -76 55 -42 87
rect -76 -15 -42 17
rect -76 -17 -42 -15
rect -76 -83 -42 -55
rect -76 -89 -42 -83
rect -76 -151 -42 -127
rect -76 -161 -42 -151
rect -76 -219 -42 -199
rect -76 -233 -42 -219
rect -76 -287 -42 -271
rect -76 -305 -42 -287
rect -76 -355 -42 -343
rect -76 -377 -42 -355
rect -76 -423 -42 -415
rect -76 -449 -42 -423
rect -76 -491 -42 -487
rect -76 -521 -42 -491
rect -76 -593 -42 -559
rect -76 -661 -42 -631
rect -76 -665 -42 -661
rect -76 -729 -42 -703
rect -76 -737 -42 -729
rect -76 -797 -42 -775
rect -76 -809 -42 -797
rect -76 -865 -42 -847
rect -76 -881 -42 -865
rect -76 -933 -42 -919
rect -76 -953 -42 -933
rect 42 1005 76 1025
rect 42 991 76 1005
rect 42 937 76 953
rect 42 919 76 937
rect 42 869 76 881
rect 42 847 76 869
rect 42 801 76 809
rect 42 775 76 801
rect 42 733 76 737
rect 42 703 76 733
rect 42 631 76 665
rect 42 563 76 593
rect 42 559 76 563
rect 42 495 76 521
rect 42 487 76 495
rect 42 427 76 449
rect 42 415 76 427
rect 42 359 76 377
rect 42 343 76 359
rect 42 291 76 305
rect 42 271 76 291
rect 42 223 76 233
rect 42 199 76 223
rect 42 155 76 161
rect 42 127 76 155
rect 42 87 76 89
rect 42 55 76 87
rect 42 -15 76 17
rect 42 -17 76 -15
rect 42 -83 76 -55
rect 42 -89 76 -83
rect 42 -151 76 -127
rect 42 -161 76 -151
rect 42 -219 76 -199
rect 42 -233 76 -219
rect 42 -287 76 -271
rect 42 -305 76 -287
rect 42 -355 76 -343
rect 42 -377 76 -355
rect 42 -423 76 -415
rect 42 -449 76 -423
rect 42 -491 76 -487
rect 42 -521 76 -491
rect 42 -593 76 -559
rect 42 -661 76 -631
rect 42 -665 76 -661
rect 42 -729 76 -703
rect 42 -737 76 -729
rect 42 -797 76 -775
rect 42 -809 76 -797
rect 42 -865 76 -847
rect 42 -881 76 -865
rect 42 -933 76 -919
rect 42 -953 76 -933
rect -17 -1065 17 -1031
<< metal1 >>
rect -82 1025 -36 1056
rect -82 991 -76 1025
rect -42 991 -36 1025
rect -82 953 -36 991
rect -82 919 -76 953
rect -42 919 -36 953
rect -82 881 -36 919
rect -82 847 -76 881
rect -42 847 -36 881
rect -82 809 -36 847
rect -82 775 -76 809
rect -42 775 -36 809
rect -82 737 -36 775
rect -82 703 -76 737
rect -42 703 -36 737
rect -82 665 -36 703
rect -82 631 -76 665
rect -42 631 -36 665
rect -82 593 -36 631
rect -82 559 -76 593
rect -42 559 -36 593
rect -82 521 -36 559
rect -82 487 -76 521
rect -42 487 -36 521
rect -82 449 -36 487
rect -82 415 -76 449
rect -42 415 -36 449
rect -82 377 -36 415
rect -82 343 -76 377
rect -42 343 -36 377
rect -82 305 -36 343
rect -82 271 -76 305
rect -42 271 -36 305
rect -82 233 -36 271
rect -82 199 -76 233
rect -42 199 -36 233
rect -82 161 -36 199
rect -82 127 -76 161
rect -42 127 -36 161
rect -82 89 -36 127
rect -82 55 -76 89
rect -42 55 -36 89
rect -82 17 -36 55
rect -82 -17 -76 17
rect -42 -17 -36 17
rect -82 -55 -36 -17
rect -82 -89 -76 -55
rect -42 -89 -36 -55
rect -82 -127 -36 -89
rect -82 -161 -76 -127
rect -42 -161 -36 -127
rect -82 -199 -36 -161
rect -82 -233 -76 -199
rect -42 -233 -36 -199
rect -82 -271 -36 -233
rect -82 -305 -76 -271
rect -42 -305 -36 -271
rect -82 -343 -36 -305
rect -82 -377 -76 -343
rect -42 -377 -36 -343
rect -82 -415 -36 -377
rect -82 -449 -76 -415
rect -42 -449 -36 -415
rect -82 -487 -36 -449
rect -82 -521 -76 -487
rect -42 -521 -36 -487
rect -82 -559 -36 -521
rect -82 -593 -76 -559
rect -42 -593 -36 -559
rect -82 -631 -36 -593
rect -82 -665 -76 -631
rect -42 -665 -36 -631
rect -82 -703 -36 -665
rect -82 -737 -76 -703
rect -42 -737 -36 -703
rect -82 -775 -36 -737
rect -82 -809 -76 -775
rect -42 -809 -36 -775
rect -82 -847 -36 -809
rect -82 -881 -76 -847
rect -42 -881 -36 -847
rect -82 -919 -36 -881
rect -82 -953 -76 -919
rect -42 -953 -36 -919
rect -82 -984 -36 -953
rect 36 1025 82 1056
rect 36 991 42 1025
rect 76 991 82 1025
rect 36 953 82 991
rect 36 919 42 953
rect 76 919 82 953
rect 36 881 82 919
rect 36 847 42 881
rect 76 847 82 881
rect 36 809 82 847
rect 36 775 42 809
rect 76 775 82 809
rect 36 737 82 775
rect 36 703 42 737
rect 76 703 82 737
rect 36 665 82 703
rect 36 631 42 665
rect 76 631 82 665
rect 36 593 82 631
rect 36 559 42 593
rect 76 559 82 593
rect 36 521 82 559
rect 36 487 42 521
rect 76 487 82 521
rect 36 449 82 487
rect 36 415 42 449
rect 76 415 82 449
rect 36 377 82 415
rect 36 343 42 377
rect 76 343 82 377
rect 36 305 82 343
rect 36 271 42 305
rect 76 271 82 305
rect 36 233 82 271
rect 36 199 42 233
rect 76 199 82 233
rect 36 161 82 199
rect 36 127 42 161
rect 76 127 82 161
rect 36 89 82 127
rect 36 55 42 89
rect 76 55 82 89
rect 36 17 82 55
rect 36 -17 42 17
rect 76 -17 82 17
rect 36 -55 82 -17
rect 36 -89 42 -55
rect 76 -89 82 -55
rect 36 -127 82 -89
rect 36 -161 42 -127
rect 76 -161 82 -127
rect 36 -199 82 -161
rect 36 -233 42 -199
rect 76 -233 82 -199
rect 36 -271 82 -233
rect 36 -305 42 -271
rect 76 -305 82 -271
rect 36 -343 82 -305
rect 36 -377 42 -343
rect 76 -377 82 -343
rect 36 -415 82 -377
rect 36 -449 42 -415
rect 76 -449 82 -415
rect 36 -487 82 -449
rect 36 -521 42 -487
rect 76 -521 82 -487
rect 36 -559 82 -521
rect 36 -593 42 -559
rect 76 -593 82 -559
rect 36 -631 82 -593
rect 36 -665 42 -631
rect 76 -665 82 -631
rect 36 -703 82 -665
rect 36 -737 42 -703
rect 76 -737 82 -703
rect 36 -775 82 -737
rect 36 -809 42 -775
rect 76 -809 82 -775
rect 36 -847 82 -809
rect 36 -881 42 -847
rect 76 -881 82 -847
rect 36 -919 82 -881
rect 36 -953 42 -919
rect 76 -953 82 -919
rect 36 -984 82 -953
rect -29 -1031 29 -1025
rect -29 -1065 -17 -1031
rect 17 -1065 29 -1031
rect -29 -1071 29 -1065
<< end >>
