magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -1530 -9626 1530 9626
<< nmos >>
rect -1446 -9600 -1386 9600
rect -1328 -9600 -1268 9600
rect -1210 -9600 -1150 9600
rect -1092 -9600 -1032 9600
rect -974 -9600 -914 9600
rect -856 -9600 -796 9600
rect -738 -9600 -678 9600
rect -620 -9600 -560 9600
rect -502 -9600 -442 9600
rect -384 -9600 -324 9600
rect -266 -9600 -206 9600
rect -148 -9600 -88 9600
rect -30 -9600 30 9600
rect 88 -9600 148 9600
rect 206 -9600 266 9600
rect 324 -9600 384 9600
rect 442 -9600 502 9600
rect 560 -9600 620 9600
rect 678 -9600 738 9600
rect 796 -9600 856 9600
rect 914 -9600 974 9600
rect 1032 -9600 1092 9600
rect 1150 -9600 1210 9600
rect 1268 -9600 1328 9600
rect 1386 -9600 1446 9600
<< ndiff >>
rect -1504 9571 -1446 9600
rect -1504 9537 -1492 9571
rect -1458 9537 -1446 9571
rect -1504 9503 -1446 9537
rect -1504 9469 -1492 9503
rect -1458 9469 -1446 9503
rect -1504 9435 -1446 9469
rect -1504 9401 -1492 9435
rect -1458 9401 -1446 9435
rect -1504 9367 -1446 9401
rect -1504 9333 -1492 9367
rect -1458 9333 -1446 9367
rect -1504 9299 -1446 9333
rect -1504 9265 -1492 9299
rect -1458 9265 -1446 9299
rect -1504 9231 -1446 9265
rect -1504 9197 -1492 9231
rect -1458 9197 -1446 9231
rect -1504 9163 -1446 9197
rect -1504 9129 -1492 9163
rect -1458 9129 -1446 9163
rect -1504 9095 -1446 9129
rect -1504 9061 -1492 9095
rect -1458 9061 -1446 9095
rect -1504 9027 -1446 9061
rect -1504 8993 -1492 9027
rect -1458 8993 -1446 9027
rect -1504 8959 -1446 8993
rect -1504 8925 -1492 8959
rect -1458 8925 -1446 8959
rect -1504 8891 -1446 8925
rect -1504 8857 -1492 8891
rect -1458 8857 -1446 8891
rect -1504 8823 -1446 8857
rect -1504 8789 -1492 8823
rect -1458 8789 -1446 8823
rect -1504 8755 -1446 8789
rect -1504 8721 -1492 8755
rect -1458 8721 -1446 8755
rect -1504 8687 -1446 8721
rect -1504 8653 -1492 8687
rect -1458 8653 -1446 8687
rect -1504 8619 -1446 8653
rect -1504 8585 -1492 8619
rect -1458 8585 -1446 8619
rect -1504 8551 -1446 8585
rect -1504 8517 -1492 8551
rect -1458 8517 -1446 8551
rect -1504 8483 -1446 8517
rect -1504 8449 -1492 8483
rect -1458 8449 -1446 8483
rect -1504 8415 -1446 8449
rect -1504 8381 -1492 8415
rect -1458 8381 -1446 8415
rect -1504 8347 -1446 8381
rect -1504 8313 -1492 8347
rect -1458 8313 -1446 8347
rect -1504 8279 -1446 8313
rect -1504 8245 -1492 8279
rect -1458 8245 -1446 8279
rect -1504 8211 -1446 8245
rect -1504 8177 -1492 8211
rect -1458 8177 -1446 8211
rect -1504 8143 -1446 8177
rect -1504 8109 -1492 8143
rect -1458 8109 -1446 8143
rect -1504 8075 -1446 8109
rect -1504 8041 -1492 8075
rect -1458 8041 -1446 8075
rect -1504 8007 -1446 8041
rect -1504 7973 -1492 8007
rect -1458 7973 -1446 8007
rect -1504 7939 -1446 7973
rect -1504 7905 -1492 7939
rect -1458 7905 -1446 7939
rect -1504 7871 -1446 7905
rect -1504 7837 -1492 7871
rect -1458 7837 -1446 7871
rect -1504 7803 -1446 7837
rect -1504 7769 -1492 7803
rect -1458 7769 -1446 7803
rect -1504 7735 -1446 7769
rect -1504 7701 -1492 7735
rect -1458 7701 -1446 7735
rect -1504 7667 -1446 7701
rect -1504 7633 -1492 7667
rect -1458 7633 -1446 7667
rect -1504 7599 -1446 7633
rect -1504 7565 -1492 7599
rect -1458 7565 -1446 7599
rect -1504 7531 -1446 7565
rect -1504 7497 -1492 7531
rect -1458 7497 -1446 7531
rect -1504 7463 -1446 7497
rect -1504 7429 -1492 7463
rect -1458 7429 -1446 7463
rect -1504 7395 -1446 7429
rect -1504 7361 -1492 7395
rect -1458 7361 -1446 7395
rect -1504 7327 -1446 7361
rect -1504 7293 -1492 7327
rect -1458 7293 -1446 7327
rect -1504 7259 -1446 7293
rect -1504 7225 -1492 7259
rect -1458 7225 -1446 7259
rect -1504 7191 -1446 7225
rect -1504 7157 -1492 7191
rect -1458 7157 -1446 7191
rect -1504 7123 -1446 7157
rect -1504 7089 -1492 7123
rect -1458 7089 -1446 7123
rect -1504 7055 -1446 7089
rect -1504 7021 -1492 7055
rect -1458 7021 -1446 7055
rect -1504 6987 -1446 7021
rect -1504 6953 -1492 6987
rect -1458 6953 -1446 6987
rect -1504 6919 -1446 6953
rect -1504 6885 -1492 6919
rect -1458 6885 -1446 6919
rect -1504 6851 -1446 6885
rect -1504 6817 -1492 6851
rect -1458 6817 -1446 6851
rect -1504 6783 -1446 6817
rect -1504 6749 -1492 6783
rect -1458 6749 -1446 6783
rect -1504 6715 -1446 6749
rect -1504 6681 -1492 6715
rect -1458 6681 -1446 6715
rect -1504 6647 -1446 6681
rect -1504 6613 -1492 6647
rect -1458 6613 -1446 6647
rect -1504 6579 -1446 6613
rect -1504 6545 -1492 6579
rect -1458 6545 -1446 6579
rect -1504 6511 -1446 6545
rect -1504 6477 -1492 6511
rect -1458 6477 -1446 6511
rect -1504 6443 -1446 6477
rect -1504 6409 -1492 6443
rect -1458 6409 -1446 6443
rect -1504 6375 -1446 6409
rect -1504 6341 -1492 6375
rect -1458 6341 -1446 6375
rect -1504 6307 -1446 6341
rect -1504 6273 -1492 6307
rect -1458 6273 -1446 6307
rect -1504 6239 -1446 6273
rect -1504 6205 -1492 6239
rect -1458 6205 -1446 6239
rect -1504 6171 -1446 6205
rect -1504 6137 -1492 6171
rect -1458 6137 -1446 6171
rect -1504 6103 -1446 6137
rect -1504 6069 -1492 6103
rect -1458 6069 -1446 6103
rect -1504 6035 -1446 6069
rect -1504 6001 -1492 6035
rect -1458 6001 -1446 6035
rect -1504 5967 -1446 6001
rect -1504 5933 -1492 5967
rect -1458 5933 -1446 5967
rect -1504 5899 -1446 5933
rect -1504 5865 -1492 5899
rect -1458 5865 -1446 5899
rect -1504 5831 -1446 5865
rect -1504 5797 -1492 5831
rect -1458 5797 -1446 5831
rect -1504 5763 -1446 5797
rect -1504 5729 -1492 5763
rect -1458 5729 -1446 5763
rect -1504 5695 -1446 5729
rect -1504 5661 -1492 5695
rect -1458 5661 -1446 5695
rect -1504 5627 -1446 5661
rect -1504 5593 -1492 5627
rect -1458 5593 -1446 5627
rect -1504 5559 -1446 5593
rect -1504 5525 -1492 5559
rect -1458 5525 -1446 5559
rect -1504 5491 -1446 5525
rect -1504 5457 -1492 5491
rect -1458 5457 -1446 5491
rect -1504 5423 -1446 5457
rect -1504 5389 -1492 5423
rect -1458 5389 -1446 5423
rect -1504 5355 -1446 5389
rect -1504 5321 -1492 5355
rect -1458 5321 -1446 5355
rect -1504 5287 -1446 5321
rect -1504 5253 -1492 5287
rect -1458 5253 -1446 5287
rect -1504 5219 -1446 5253
rect -1504 5185 -1492 5219
rect -1458 5185 -1446 5219
rect -1504 5151 -1446 5185
rect -1504 5117 -1492 5151
rect -1458 5117 -1446 5151
rect -1504 5083 -1446 5117
rect -1504 5049 -1492 5083
rect -1458 5049 -1446 5083
rect -1504 5015 -1446 5049
rect -1504 4981 -1492 5015
rect -1458 4981 -1446 5015
rect -1504 4947 -1446 4981
rect -1504 4913 -1492 4947
rect -1458 4913 -1446 4947
rect -1504 4879 -1446 4913
rect -1504 4845 -1492 4879
rect -1458 4845 -1446 4879
rect -1504 4811 -1446 4845
rect -1504 4777 -1492 4811
rect -1458 4777 -1446 4811
rect -1504 4743 -1446 4777
rect -1504 4709 -1492 4743
rect -1458 4709 -1446 4743
rect -1504 4675 -1446 4709
rect -1504 4641 -1492 4675
rect -1458 4641 -1446 4675
rect -1504 4607 -1446 4641
rect -1504 4573 -1492 4607
rect -1458 4573 -1446 4607
rect -1504 4539 -1446 4573
rect -1504 4505 -1492 4539
rect -1458 4505 -1446 4539
rect -1504 4471 -1446 4505
rect -1504 4437 -1492 4471
rect -1458 4437 -1446 4471
rect -1504 4403 -1446 4437
rect -1504 4369 -1492 4403
rect -1458 4369 -1446 4403
rect -1504 4335 -1446 4369
rect -1504 4301 -1492 4335
rect -1458 4301 -1446 4335
rect -1504 4267 -1446 4301
rect -1504 4233 -1492 4267
rect -1458 4233 -1446 4267
rect -1504 4199 -1446 4233
rect -1504 4165 -1492 4199
rect -1458 4165 -1446 4199
rect -1504 4131 -1446 4165
rect -1504 4097 -1492 4131
rect -1458 4097 -1446 4131
rect -1504 4063 -1446 4097
rect -1504 4029 -1492 4063
rect -1458 4029 -1446 4063
rect -1504 3995 -1446 4029
rect -1504 3961 -1492 3995
rect -1458 3961 -1446 3995
rect -1504 3927 -1446 3961
rect -1504 3893 -1492 3927
rect -1458 3893 -1446 3927
rect -1504 3859 -1446 3893
rect -1504 3825 -1492 3859
rect -1458 3825 -1446 3859
rect -1504 3791 -1446 3825
rect -1504 3757 -1492 3791
rect -1458 3757 -1446 3791
rect -1504 3723 -1446 3757
rect -1504 3689 -1492 3723
rect -1458 3689 -1446 3723
rect -1504 3655 -1446 3689
rect -1504 3621 -1492 3655
rect -1458 3621 -1446 3655
rect -1504 3587 -1446 3621
rect -1504 3553 -1492 3587
rect -1458 3553 -1446 3587
rect -1504 3519 -1446 3553
rect -1504 3485 -1492 3519
rect -1458 3485 -1446 3519
rect -1504 3451 -1446 3485
rect -1504 3417 -1492 3451
rect -1458 3417 -1446 3451
rect -1504 3383 -1446 3417
rect -1504 3349 -1492 3383
rect -1458 3349 -1446 3383
rect -1504 3315 -1446 3349
rect -1504 3281 -1492 3315
rect -1458 3281 -1446 3315
rect -1504 3247 -1446 3281
rect -1504 3213 -1492 3247
rect -1458 3213 -1446 3247
rect -1504 3179 -1446 3213
rect -1504 3145 -1492 3179
rect -1458 3145 -1446 3179
rect -1504 3111 -1446 3145
rect -1504 3077 -1492 3111
rect -1458 3077 -1446 3111
rect -1504 3043 -1446 3077
rect -1504 3009 -1492 3043
rect -1458 3009 -1446 3043
rect -1504 2975 -1446 3009
rect -1504 2941 -1492 2975
rect -1458 2941 -1446 2975
rect -1504 2907 -1446 2941
rect -1504 2873 -1492 2907
rect -1458 2873 -1446 2907
rect -1504 2839 -1446 2873
rect -1504 2805 -1492 2839
rect -1458 2805 -1446 2839
rect -1504 2771 -1446 2805
rect -1504 2737 -1492 2771
rect -1458 2737 -1446 2771
rect -1504 2703 -1446 2737
rect -1504 2669 -1492 2703
rect -1458 2669 -1446 2703
rect -1504 2635 -1446 2669
rect -1504 2601 -1492 2635
rect -1458 2601 -1446 2635
rect -1504 2567 -1446 2601
rect -1504 2533 -1492 2567
rect -1458 2533 -1446 2567
rect -1504 2499 -1446 2533
rect -1504 2465 -1492 2499
rect -1458 2465 -1446 2499
rect -1504 2431 -1446 2465
rect -1504 2397 -1492 2431
rect -1458 2397 -1446 2431
rect -1504 2363 -1446 2397
rect -1504 2329 -1492 2363
rect -1458 2329 -1446 2363
rect -1504 2295 -1446 2329
rect -1504 2261 -1492 2295
rect -1458 2261 -1446 2295
rect -1504 2227 -1446 2261
rect -1504 2193 -1492 2227
rect -1458 2193 -1446 2227
rect -1504 2159 -1446 2193
rect -1504 2125 -1492 2159
rect -1458 2125 -1446 2159
rect -1504 2091 -1446 2125
rect -1504 2057 -1492 2091
rect -1458 2057 -1446 2091
rect -1504 2023 -1446 2057
rect -1504 1989 -1492 2023
rect -1458 1989 -1446 2023
rect -1504 1955 -1446 1989
rect -1504 1921 -1492 1955
rect -1458 1921 -1446 1955
rect -1504 1887 -1446 1921
rect -1504 1853 -1492 1887
rect -1458 1853 -1446 1887
rect -1504 1819 -1446 1853
rect -1504 1785 -1492 1819
rect -1458 1785 -1446 1819
rect -1504 1751 -1446 1785
rect -1504 1717 -1492 1751
rect -1458 1717 -1446 1751
rect -1504 1683 -1446 1717
rect -1504 1649 -1492 1683
rect -1458 1649 -1446 1683
rect -1504 1615 -1446 1649
rect -1504 1581 -1492 1615
rect -1458 1581 -1446 1615
rect -1504 1547 -1446 1581
rect -1504 1513 -1492 1547
rect -1458 1513 -1446 1547
rect -1504 1479 -1446 1513
rect -1504 1445 -1492 1479
rect -1458 1445 -1446 1479
rect -1504 1411 -1446 1445
rect -1504 1377 -1492 1411
rect -1458 1377 -1446 1411
rect -1504 1343 -1446 1377
rect -1504 1309 -1492 1343
rect -1458 1309 -1446 1343
rect -1504 1275 -1446 1309
rect -1504 1241 -1492 1275
rect -1458 1241 -1446 1275
rect -1504 1207 -1446 1241
rect -1504 1173 -1492 1207
rect -1458 1173 -1446 1207
rect -1504 1139 -1446 1173
rect -1504 1105 -1492 1139
rect -1458 1105 -1446 1139
rect -1504 1071 -1446 1105
rect -1504 1037 -1492 1071
rect -1458 1037 -1446 1071
rect -1504 1003 -1446 1037
rect -1504 969 -1492 1003
rect -1458 969 -1446 1003
rect -1504 935 -1446 969
rect -1504 901 -1492 935
rect -1458 901 -1446 935
rect -1504 867 -1446 901
rect -1504 833 -1492 867
rect -1458 833 -1446 867
rect -1504 799 -1446 833
rect -1504 765 -1492 799
rect -1458 765 -1446 799
rect -1504 731 -1446 765
rect -1504 697 -1492 731
rect -1458 697 -1446 731
rect -1504 663 -1446 697
rect -1504 629 -1492 663
rect -1458 629 -1446 663
rect -1504 595 -1446 629
rect -1504 561 -1492 595
rect -1458 561 -1446 595
rect -1504 527 -1446 561
rect -1504 493 -1492 527
rect -1458 493 -1446 527
rect -1504 459 -1446 493
rect -1504 425 -1492 459
rect -1458 425 -1446 459
rect -1504 391 -1446 425
rect -1504 357 -1492 391
rect -1458 357 -1446 391
rect -1504 323 -1446 357
rect -1504 289 -1492 323
rect -1458 289 -1446 323
rect -1504 255 -1446 289
rect -1504 221 -1492 255
rect -1458 221 -1446 255
rect -1504 187 -1446 221
rect -1504 153 -1492 187
rect -1458 153 -1446 187
rect -1504 119 -1446 153
rect -1504 85 -1492 119
rect -1458 85 -1446 119
rect -1504 51 -1446 85
rect -1504 17 -1492 51
rect -1458 17 -1446 51
rect -1504 -17 -1446 17
rect -1504 -51 -1492 -17
rect -1458 -51 -1446 -17
rect -1504 -85 -1446 -51
rect -1504 -119 -1492 -85
rect -1458 -119 -1446 -85
rect -1504 -153 -1446 -119
rect -1504 -187 -1492 -153
rect -1458 -187 -1446 -153
rect -1504 -221 -1446 -187
rect -1504 -255 -1492 -221
rect -1458 -255 -1446 -221
rect -1504 -289 -1446 -255
rect -1504 -323 -1492 -289
rect -1458 -323 -1446 -289
rect -1504 -357 -1446 -323
rect -1504 -391 -1492 -357
rect -1458 -391 -1446 -357
rect -1504 -425 -1446 -391
rect -1504 -459 -1492 -425
rect -1458 -459 -1446 -425
rect -1504 -493 -1446 -459
rect -1504 -527 -1492 -493
rect -1458 -527 -1446 -493
rect -1504 -561 -1446 -527
rect -1504 -595 -1492 -561
rect -1458 -595 -1446 -561
rect -1504 -629 -1446 -595
rect -1504 -663 -1492 -629
rect -1458 -663 -1446 -629
rect -1504 -697 -1446 -663
rect -1504 -731 -1492 -697
rect -1458 -731 -1446 -697
rect -1504 -765 -1446 -731
rect -1504 -799 -1492 -765
rect -1458 -799 -1446 -765
rect -1504 -833 -1446 -799
rect -1504 -867 -1492 -833
rect -1458 -867 -1446 -833
rect -1504 -901 -1446 -867
rect -1504 -935 -1492 -901
rect -1458 -935 -1446 -901
rect -1504 -969 -1446 -935
rect -1504 -1003 -1492 -969
rect -1458 -1003 -1446 -969
rect -1504 -1037 -1446 -1003
rect -1504 -1071 -1492 -1037
rect -1458 -1071 -1446 -1037
rect -1504 -1105 -1446 -1071
rect -1504 -1139 -1492 -1105
rect -1458 -1139 -1446 -1105
rect -1504 -1173 -1446 -1139
rect -1504 -1207 -1492 -1173
rect -1458 -1207 -1446 -1173
rect -1504 -1241 -1446 -1207
rect -1504 -1275 -1492 -1241
rect -1458 -1275 -1446 -1241
rect -1504 -1309 -1446 -1275
rect -1504 -1343 -1492 -1309
rect -1458 -1343 -1446 -1309
rect -1504 -1377 -1446 -1343
rect -1504 -1411 -1492 -1377
rect -1458 -1411 -1446 -1377
rect -1504 -1445 -1446 -1411
rect -1504 -1479 -1492 -1445
rect -1458 -1479 -1446 -1445
rect -1504 -1513 -1446 -1479
rect -1504 -1547 -1492 -1513
rect -1458 -1547 -1446 -1513
rect -1504 -1581 -1446 -1547
rect -1504 -1615 -1492 -1581
rect -1458 -1615 -1446 -1581
rect -1504 -1649 -1446 -1615
rect -1504 -1683 -1492 -1649
rect -1458 -1683 -1446 -1649
rect -1504 -1717 -1446 -1683
rect -1504 -1751 -1492 -1717
rect -1458 -1751 -1446 -1717
rect -1504 -1785 -1446 -1751
rect -1504 -1819 -1492 -1785
rect -1458 -1819 -1446 -1785
rect -1504 -1853 -1446 -1819
rect -1504 -1887 -1492 -1853
rect -1458 -1887 -1446 -1853
rect -1504 -1921 -1446 -1887
rect -1504 -1955 -1492 -1921
rect -1458 -1955 -1446 -1921
rect -1504 -1989 -1446 -1955
rect -1504 -2023 -1492 -1989
rect -1458 -2023 -1446 -1989
rect -1504 -2057 -1446 -2023
rect -1504 -2091 -1492 -2057
rect -1458 -2091 -1446 -2057
rect -1504 -2125 -1446 -2091
rect -1504 -2159 -1492 -2125
rect -1458 -2159 -1446 -2125
rect -1504 -2193 -1446 -2159
rect -1504 -2227 -1492 -2193
rect -1458 -2227 -1446 -2193
rect -1504 -2261 -1446 -2227
rect -1504 -2295 -1492 -2261
rect -1458 -2295 -1446 -2261
rect -1504 -2329 -1446 -2295
rect -1504 -2363 -1492 -2329
rect -1458 -2363 -1446 -2329
rect -1504 -2397 -1446 -2363
rect -1504 -2431 -1492 -2397
rect -1458 -2431 -1446 -2397
rect -1504 -2465 -1446 -2431
rect -1504 -2499 -1492 -2465
rect -1458 -2499 -1446 -2465
rect -1504 -2533 -1446 -2499
rect -1504 -2567 -1492 -2533
rect -1458 -2567 -1446 -2533
rect -1504 -2601 -1446 -2567
rect -1504 -2635 -1492 -2601
rect -1458 -2635 -1446 -2601
rect -1504 -2669 -1446 -2635
rect -1504 -2703 -1492 -2669
rect -1458 -2703 -1446 -2669
rect -1504 -2737 -1446 -2703
rect -1504 -2771 -1492 -2737
rect -1458 -2771 -1446 -2737
rect -1504 -2805 -1446 -2771
rect -1504 -2839 -1492 -2805
rect -1458 -2839 -1446 -2805
rect -1504 -2873 -1446 -2839
rect -1504 -2907 -1492 -2873
rect -1458 -2907 -1446 -2873
rect -1504 -2941 -1446 -2907
rect -1504 -2975 -1492 -2941
rect -1458 -2975 -1446 -2941
rect -1504 -3009 -1446 -2975
rect -1504 -3043 -1492 -3009
rect -1458 -3043 -1446 -3009
rect -1504 -3077 -1446 -3043
rect -1504 -3111 -1492 -3077
rect -1458 -3111 -1446 -3077
rect -1504 -3145 -1446 -3111
rect -1504 -3179 -1492 -3145
rect -1458 -3179 -1446 -3145
rect -1504 -3213 -1446 -3179
rect -1504 -3247 -1492 -3213
rect -1458 -3247 -1446 -3213
rect -1504 -3281 -1446 -3247
rect -1504 -3315 -1492 -3281
rect -1458 -3315 -1446 -3281
rect -1504 -3349 -1446 -3315
rect -1504 -3383 -1492 -3349
rect -1458 -3383 -1446 -3349
rect -1504 -3417 -1446 -3383
rect -1504 -3451 -1492 -3417
rect -1458 -3451 -1446 -3417
rect -1504 -3485 -1446 -3451
rect -1504 -3519 -1492 -3485
rect -1458 -3519 -1446 -3485
rect -1504 -3553 -1446 -3519
rect -1504 -3587 -1492 -3553
rect -1458 -3587 -1446 -3553
rect -1504 -3621 -1446 -3587
rect -1504 -3655 -1492 -3621
rect -1458 -3655 -1446 -3621
rect -1504 -3689 -1446 -3655
rect -1504 -3723 -1492 -3689
rect -1458 -3723 -1446 -3689
rect -1504 -3757 -1446 -3723
rect -1504 -3791 -1492 -3757
rect -1458 -3791 -1446 -3757
rect -1504 -3825 -1446 -3791
rect -1504 -3859 -1492 -3825
rect -1458 -3859 -1446 -3825
rect -1504 -3893 -1446 -3859
rect -1504 -3927 -1492 -3893
rect -1458 -3927 -1446 -3893
rect -1504 -3961 -1446 -3927
rect -1504 -3995 -1492 -3961
rect -1458 -3995 -1446 -3961
rect -1504 -4029 -1446 -3995
rect -1504 -4063 -1492 -4029
rect -1458 -4063 -1446 -4029
rect -1504 -4097 -1446 -4063
rect -1504 -4131 -1492 -4097
rect -1458 -4131 -1446 -4097
rect -1504 -4165 -1446 -4131
rect -1504 -4199 -1492 -4165
rect -1458 -4199 -1446 -4165
rect -1504 -4233 -1446 -4199
rect -1504 -4267 -1492 -4233
rect -1458 -4267 -1446 -4233
rect -1504 -4301 -1446 -4267
rect -1504 -4335 -1492 -4301
rect -1458 -4335 -1446 -4301
rect -1504 -4369 -1446 -4335
rect -1504 -4403 -1492 -4369
rect -1458 -4403 -1446 -4369
rect -1504 -4437 -1446 -4403
rect -1504 -4471 -1492 -4437
rect -1458 -4471 -1446 -4437
rect -1504 -4505 -1446 -4471
rect -1504 -4539 -1492 -4505
rect -1458 -4539 -1446 -4505
rect -1504 -4573 -1446 -4539
rect -1504 -4607 -1492 -4573
rect -1458 -4607 -1446 -4573
rect -1504 -4641 -1446 -4607
rect -1504 -4675 -1492 -4641
rect -1458 -4675 -1446 -4641
rect -1504 -4709 -1446 -4675
rect -1504 -4743 -1492 -4709
rect -1458 -4743 -1446 -4709
rect -1504 -4777 -1446 -4743
rect -1504 -4811 -1492 -4777
rect -1458 -4811 -1446 -4777
rect -1504 -4845 -1446 -4811
rect -1504 -4879 -1492 -4845
rect -1458 -4879 -1446 -4845
rect -1504 -4913 -1446 -4879
rect -1504 -4947 -1492 -4913
rect -1458 -4947 -1446 -4913
rect -1504 -4981 -1446 -4947
rect -1504 -5015 -1492 -4981
rect -1458 -5015 -1446 -4981
rect -1504 -5049 -1446 -5015
rect -1504 -5083 -1492 -5049
rect -1458 -5083 -1446 -5049
rect -1504 -5117 -1446 -5083
rect -1504 -5151 -1492 -5117
rect -1458 -5151 -1446 -5117
rect -1504 -5185 -1446 -5151
rect -1504 -5219 -1492 -5185
rect -1458 -5219 -1446 -5185
rect -1504 -5253 -1446 -5219
rect -1504 -5287 -1492 -5253
rect -1458 -5287 -1446 -5253
rect -1504 -5321 -1446 -5287
rect -1504 -5355 -1492 -5321
rect -1458 -5355 -1446 -5321
rect -1504 -5389 -1446 -5355
rect -1504 -5423 -1492 -5389
rect -1458 -5423 -1446 -5389
rect -1504 -5457 -1446 -5423
rect -1504 -5491 -1492 -5457
rect -1458 -5491 -1446 -5457
rect -1504 -5525 -1446 -5491
rect -1504 -5559 -1492 -5525
rect -1458 -5559 -1446 -5525
rect -1504 -5593 -1446 -5559
rect -1504 -5627 -1492 -5593
rect -1458 -5627 -1446 -5593
rect -1504 -5661 -1446 -5627
rect -1504 -5695 -1492 -5661
rect -1458 -5695 -1446 -5661
rect -1504 -5729 -1446 -5695
rect -1504 -5763 -1492 -5729
rect -1458 -5763 -1446 -5729
rect -1504 -5797 -1446 -5763
rect -1504 -5831 -1492 -5797
rect -1458 -5831 -1446 -5797
rect -1504 -5865 -1446 -5831
rect -1504 -5899 -1492 -5865
rect -1458 -5899 -1446 -5865
rect -1504 -5933 -1446 -5899
rect -1504 -5967 -1492 -5933
rect -1458 -5967 -1446 -5933
rect -1504 -6001 -1446 -5967
rect -1504 -6035 -1492 -6001
rect -1458 -6035 -1446 -6001
rect -1504 -6069 -1446 -6035
rect -1504 -6103 -1492 -6069
rect -1458 -6103 -1446 -6069
rect -1504 -6137 -1446 -6103
rect -1504 -6171 -1492 -6137
rect -1458 -6171 -1446 -6137
rect -1504 -6205 -1446 -6171
rect -1504 -6239 -1492 -6205
rect -1458 -6239 -1446 -6205
rect -1504 -6273 -1446 -6239
rect -1504 -6307 -1492 -6273
rect -1458 -6307 -1446 -6273
rect -1504 -6341 -1446 -6307
rect -1504 -6375 -1492 -6341
rect -1458 -6375 -1446 -6341
rect -1504 -6409 -1446 -6375
rect -1504 -6443 -1492 -6409
rect -1458 -6443 -1446 -6409
rect -1504 -6477 -1446 -6443
rect -1504 -6511 -1492 -6477
rect -1458 -6511 -1446 -6477
rect -1504 -6545 -1446 -6511
rect -1504 -6579 -1492 -6545
rect -1458 -6579 -1446 -6545
rect -1504 -6613 -1446 -6579
rect -1504 -6647 -1492 -6613
rect -1458 -6647 -1446 -6613
rect -1504 -6681 -1446 -6647
rect -1504 -6715 -1492 -6681
rect -1458 -6715 -1446 -6681
rect -1504 -6749 -1446 -6715
rect -1504 -6783 -1492 -6749
rect -1458 -6783 -1446 -6749
rect -1504 -6817 -1446 -6783
rect -1504 -6851 -1492 -6817
rect -1458 -6851 -1446 -6817
rect -1504 -6885 -1446 -6851
rect -1504 -6919 -1492 -6885
rect -1458 -6919 -1446 -6885
rect -1504 -6953 -1446 -6919
rect -1504 -6987 -1492 -6953
rect -1458 -6987 -1446 -6953
rect -1504 -7021 -1446 -6987
rect -1504 -7055 -1492 -7021
rect -1458 -7055 -1446 -7021
rect -1504 -7089 -1446 -7055
rect -1504 -7123 -1492 -7089
rect -1458 -7123 -1446 -7089
rect -1504 -7157 -1446 -7123
rect -1504 -7191 -1492 -7157
rect -1458 -7191 -1446 -7157
rect -1504 -7225 -1446 -7191
rect -1504 -7259 -1492 -7225
rect -1458 -7259 -1446 -7225
rect -1504 -7293 -1446 -7259
rect -1504 -7327 -1492 -7293
rect -1458 -7327 -1446 -7293
rect -1504 -7361 -1446 -7327
rect -1504 -7395 -1492 -7361
rect -1458 -7395 -1446 -7361
rect -1504 -7429 -1446 -7395
rect -1504 -7463 -1492 -7429
rect -1458 -7463 -1446 -7429
rect -1504 -7497 -1446 -7463
rect -1504 -7531 -1492 -7497
rect -1458 -7531 -1446 -7497
rect -1504 -7565 -1446 -7531
rect -1504 -7599 -1492 -7565
rect -1458 -7599 -1446 -7565
rect -1504 -7633 -1446 -7599
rect -1504 -7667 -1492 -7633
rect -1458 -7667 -1446 -7633
rect -1504 -7701 -1446 -7667
rect -1504 -7735 -1492 -7701
rect -1458 -7735 -1446 -7701
rect -1504 -7769 -1446 -7735
rect -1504 -7803 -1492 -7769
rect -1458 -7803 -1446 -7769
rect -1504 -7837 -1446 -7803
rect -1504 -7871 -1492 -7837
rect -1458 -7871 -1446 -7837
rect -1504 -7905 -1446 -7871
rect -1504 -7939 -1492 -7905
rect -1458 -7939 -1446 -7905
rect -1504 -7973 -1446 -7939
rect -1504 -8007 -1492 -7973
rect -1458 -8007 -1446 -7973
rect -1504 -8041 -1446 -8007
rect -1504 -8075 -1492 -8041
rect -1458 -8075 -1446 -8041
rect -1504 -8109 -1446 -8075
rect -1504 -8143 -1492 -8109
rect -1458 -8143 -1446 -8109
rect -1504 -8177 -1446 -8143
rect -1504 -8211 -1492 -8177
rect -1458 -8211 -1446 -8177
rect -1504 -8245 -1446 -8211
rect -1504 -8279 -1492 -8245
rect -1458 -8279 -1446 -8245
rect -1504 -8313 -1446 -8279
rect -1504 -8347 -1492 -8313
rect -1458 -8347 -1446 -8313
rect -1504 -8381 -1446 -8347
rect -1504 -8415 -1492 -8381
rect -1458 -8415 -1446 -8381
rect -1504 -8449 -1446 -8415
rect -1504 -8483 -1492 -8449
rect -1458 -8483 -1446 -8449
rect -1504 -8517 -1446 -8483
rect -1504 -8551 -1492 -8517
rect -1458 -8551 -1446 -8517
rect -1504 -8585 -1446 -8551
rect -1504 -8619 -1492 -8585
rect -1458 -8619 -1446 -8585
rect -1504 -8653 -1446 -8619
rect -1504 -8687 -1492 -8653
rect -1458 -8687 -1446 -8653
rect -1504 -8721 -1446 -8687
rect -1504 -8755 -1492 -8721
rect -1458 -8755 -1446 -8721
rect -1504 -8789 -1446 -8755
rect -1504 -8823 -1492 -8789
rect -1458 -8823 -1446 -8789
rect -1504 -8857 -1446 -8823
rect -1504 -8891 -1492 -8857
rect -1458 -8891 -1446 -8857
rect -1504 -8925 -1446 -8891
rect -1504 -8959 -1492 -8925
rect -1458 -8959 -1446 -8925
rect -1504 -8993 -1446 -8959
rect -1504 -9027 -1492 -8993
rect -1458 -9027 -1446 -8993
rect -1504 -9061 -1446 -9027
rect -1504 -9095 -1492 -9061
rect -1458 -9095 -1446 -9061
rect -1504 -9129 -1446 -9095
rect -1504 -9163 -1492 -9129
rect -1458 -9163 -1446 -9129
rect -1504 -9197 -1446 -9163
rect -1504 -9231 -1492 -9197
rect -1458 -9231 -1446 -9197
rect -1504 -9265 -1446 -9231
rect -1504 -9299 -1492 -9265
rect -1458 -9299 -1446 -9265
rect -1504 -9333 -1446 -9299
rect -1504 -9367 -1492 -9333
rect -1458 -9367 -1446 -9333
rect -1504 -9401 -1446 -9367
rect -1504 -9435 -1492 -9401
rect -1458 -9435 -1446 -9401
rect -1504 -9469 -1446 -9435
rect -1504 -9503 -1492 -9469
rect -1458 -9503 -1446 -9469
rect -1504 -9537 -1446 -9503
rect -1504 -9571 -1492 -9537
rect -1458 -9571 -1446 -9537
rect -1504 -9600 -1446 -9571
rect -1386 9571 -1328 9600
rect -1386 9537 -1374 9571
rect -1340 9537 -1328 9571
rect -1386 9503 -1328 9537
rect -1386 9469 -1374 9503
rect -1340 9469 -1328 9503
rect -1386 9435 -1328 9469
rect -1386 9401 -1374 9435
rect -1340 9401 -1328 9435
rect -1386 9367 -1328 9401
rect -1386 9333 -1374 9367
rect -1340 9333 -1328 9367
rect -1386 9299 -1328 9333
rect -1386 9265 -1374 9299
rect -1340 9265 -1328 9299
rect -1386 9231 -1328 9265
rect -1386 9197 -1374 9231
rect -1340 9197 -1328 9231
rect -1386 9163 -1328 9197
rect -1386 9129 -1374 9163
rect -1340 9129 -1328 9163
rect -1386 9095 -1328 9129
rect -1386 9061 -1374 9095
rect -1340 9061 -1328 9095
rect -1386 9027 -1328 9061
rect -1386 8993 -1374 9027
rect -1340 8993 -1328 9027
rect -1386 8959 -1328 8993
rect -1386 8925 -1374 8959
rect -1340 8925 -1328 8959
rect -1386 8891 -1328 8925
rect -1386 8857 -1374 8891
rect -1340 8857 -1328 8891
rect -1386 8823 -1328 8857
rect -1386 8789 -1374 8823
rect -1340 8789 -1328 8823
rect -1386 8755 -1328 8789
rect -1386 8721 -1374 8755
rect -1340 8721 -1328 8755
rect -1386 8687 -1328 8721
rect -1386 8653 -1374 8687
rect -1340 8653 -1328 8687
rect -1386 8619 -1328 8653
rect -1386 8585 -1374 8619
rect -1340 8585 -1328 8619
rect -1386 8551 -1328 8585
rect -1386 8517 -1374 8551
rect -1340 8517 -1328 8551
rect -1386 8483 -1328 8517
rect -1386 8449 -1374 8483
rect -1340 8449 -1328 8483
rect -1386 8415 -1328 8449
rect -1386 8381 -1374 8415
rect -1340 8381 -1328 8415
rect -1386 8347 -1328 8381
rect -1386 8313 -1374 8347
rect -1340 8313 -1328 8347
rect -1386 8279 -1328 8313
rect -1386 8245 -1374 8279
rect -1340 8245 -1328 8279
rect -1386 8211 -1328 8245
rect -1386 8177 -1374 8211
rect -1340 8177 -1328 8211
rect -1386 8143 -1328 8177
rect -1386 8109 -1374 8143
rect -1340 8109 -1328 8143
rect -1386 8075 -1328 8109
rect -1386 8041 -1374 8075
rect -1340 8041 -1328 8075
rect -1386 8007 -1328 8041
rect -1386 7973 -1374 8007
rect -1340 7973 -1328 8007
rect -1386 7939 -1328 7973
rect -1386 7905 -1374 7939
rect -1340 7905 -1328 7939
rect -1386 7871 -1328 7905
rect -1386 7837 -1374 7871
rect -1340 7837 -1328 7871
rect -1386 7803 -1328 7837
rect -1386 7769 -1374 7803
rect -1340 7769 -1328 7803
rect -1386 7735 -1328 7769
rect -1386 7701 -1374 7735
rect -1340 7701 -1328 7735
rect -1386 7667 -1328 7701
rect -1386 7633 -1374 7667
rect -1340 7633 -1328 7667
rect -1386 7599 -1328 7633
rect -1386 7565 -1374 7599
rect -1340 7565 -1328 7599
rect -1386 7531 -1328 7565
rect -1386 7497 -1374 7531
rect -1340 7497 -1328 7531
rect -1386 7463 -1328 7497
rect -1386 7429 -1374 7463
rect -1340 7429 -1328 7463
rect -1386 7395 -1328 7429
rect -1386 7361 -1374 7395
rect -1340 7361 -1328 7395
rect -1386 7327 -1328 7361
rect -1386 7293 -1374 7327
rect -1340 7293 -1328 7327
rect -1386 7259 -1328 7293
rect -1386 7225 -1374 7259
rect -1340 7225 -1328 7259
rect -1386 7191 -1328 7225
rect -1386 7157 -1374 7191
rect -1340 7157 -1328 7191
rect -1386 7123 -1328 7157
rect -1386 7089 -1374 7123
rect -1340 7089 -1328 7123
rect -1386 7055 -1328 7089
rect -1386 7021 -1374 7055
rect -1340 7021 -1328 7055
rect -1386 6987 -1328 7021
rect -1386 6953 -1374 6987
rect -1340 6953 -1328 6987
rect -1386 6919 -1328 6953
rect -1386 6885 -1374 6919
rect -1340 6885 -1328 6919
rect -1386 6851 -1328 6885
rect -1386 6817 -1374 6851
rect -1340 6817 -1328 6851
rect -1386 6783 -1328 6817
rect -1386 6749 -1374 6783
rect -1340 6749 -1328 6783
rect -1386 6715 -1328 6749
rect -1386 6681 -1374 6715
rect -1340 6681 -1328 6715
rect -1386 6647 -1328 6681
rect -1386 6613 -1374 6647
rect -1340 6613 -1328 6647
rect -1386 6579 -1328 6613
rect -1386 6545 -1374 6579
rect -1340 6545 -1328 6579
rect -1386 6511 -1328 6545
rect -1386 6477 -1374 6511
rect -1340 6477 -1328 6511
rect -1386 6443 -1328 6477
rect -1386 6409 -1374 6443
rect -1340 6409 -1328 6443
rect -1386 6375 -1328 6409
rect -1386 6341 -1374 6375
rect -1340 6341 -1328 6375
rect -1386 6307 -1328 6341
rect -1386 6273 -1374 6307
rect -1340 6273 -1328 6307
rect -1386 6239 -1328 6273
rect -1386 6205 -1374 6239
rect -1340 6205 -1328 6239
rect -1386 6171 -1328 6205
rect -1386 6137 -1374 6171
rect -1340 6137 -1328 6171
rect -1386 6103 -1328 6137
rect -1386 6069 -1374 6103
rect -1340 6069 -1328 6103
rect -1386 6035 -1328 6069
rect -1386 6001 -1374 6035
rect -1340 6001 -1328 6035
rect -1386 5967 -1328 6001
rect -1386 5933 -1374 5967
rect -1340 5933 -1328 5967
rect -1386 5899 -1328 5933
rect -1386 5865 -1374 5899
rect -1340 5865 -1328 5899
rect -1386 5831 -1328 5865
rect -1386 5797 -1374 5831
rect -1340 5797 -1328 5831
rect -1386 5763 -1328 5797
rect -1386 5729 -1374 5763
rect -1340 5729 -1328 5763
rect -1386 5695 -1328 5729
rect -1386 5661 -1374 5695
rect -1340 5661 -1328 5695
rect -1386 5627 -1328 5661
rect -1386 5593 -1374 5627
rect -1340 5593 -1328 5627
rect -1386 5559 -1328 5593
rect -1386 5525 -1374 5559
rect -1340 5525 -1328 5559
rect -1386 5491 -1328 5525
rect -1386 5457 -1374 5491
rect -1340 5457 -1328 5491
rect -1386 5423 -1328 5457
rect -1386 5389 -1374 5423
rect -1340 5389 -1328 5423
rect -1386 5355 -1328 5389
rect -1386 5321 -1374 5355
rect -1340 5321 -1328 5355
rect -1386 5287 -1328 5321
rect -1386 5253 -1374 5287
rect -1340 5253 -1328 5287
rect -1386 5219 -1328 5253
rect -1386 5185 -1374 5219
rect -1340 5185 -1328 5219
rect -1386 5151 -1328 5185
rect -1386 5117 -1374 5151
rect -1340 5117 -1328 5151
rect -1386 5083 -1328 5117
rect -1386 5049 -1374 5083
rect -1340 5049 -1328 5083
rect -1386 5015 -1328 5049
rect -1386 4981 -1374 5015
rect -1340 4981 -1328 5015
rect -1386 4947 -1328 4981
rect -1386 4913 -1374 4947
rect -1340 4913 -1328 4947
rect -1386 4879 -1328 4913
rect -1386 4845 -1374 4879
rect -1340 4845 -1328 4879
rect -1386 4811 -1328 4845
rect -1386 4777 -1374 4811
rect -1340 4777 -1328 4811
rect -1386 4743 -1328 4777
rect -1386 4709 -1374 4743
rect -1340 4709 -1328 4743
rect -1386 4675 -1328 4709
rect -1386 4641 -1374 4675
rect -1340 4641 -1328 4675
rect -1386 4607 -1328 4641
rect -1386 4573 -1374 4607
rect -1340 4573 -1328 4607
rect -1386 4539 -1328 4573
rect -1386 4505 -1374 4539
rect -1340 4505 -1328 4539
rect -1386 4471 -1328 4505
rect -1386 4437 -1374 4471
rect -1340 4437 -1328 4471
rect -1386 4403 -1328 4437
rect -1386 4369 -1374 4403
rect -1340 4369 -1328 4403
rect -1386 4335 -1328 4369
rect -1386 4301 -1374 4335
rect -1340 4301 -1328 4335
rect -1386 4267 -1328 4301
rect -1386 4233 -1374 4267
rect -1340 4233 -1328 4267
rect -1386 4199 -1328 4233
rect -1386 4165 -1374 4199
rect -1340 4165 -1328 4199
rect -1386 4131 -1328 4165
rect -1386 4097 -1374 4131
rect -1340 4097 -1328 4131
rect -1386 4063 -1328 4097
rect -1386 4029 -1374 4063
rect -1340 4029 -1328 4063
rect -1386 3995 -1328 4029
rect -1386 3961 -1374 3995
rect -1340 3961 -1328 3995
rect -1386 3927 -1328 3961
rect -1386 3893 -1374 3927
rect -1340 3893 -1328 3927
rect -1386 3859 -1328 3893
rect -1386 3825 -1374 3859
rect -1340 3825 -1328 3859
rect -1386 3791 -1328 3825
rect -1386 3757 -1374 3791
rect -1340 3757 -1328 3791
rect -1386 3723 -1328 3757
rect -1386 3689 -1374 3723
rect -1340 3689 -1328 3723
rect -1386 3655 -1328 3689
rect -1386 3621 -1374 3655
rect -1340 3621 -1328 3655
rect -1386 3587 -1328 3621
rect -1386 3553 -1374 3587
rect -1340 3553 -1328 3587
rect -1386 3519 -1328 3553
rect -1386 3485 -1374 3519
rect -1340 3485 -1328 3519
rect -1386 3451 -1328 3485
rect -1386 3417 -1374 3451
rect -1340 3417 -1328 3451
rect -1386 3383 -1328 3417
rect -1386 3349 -1374 3383
rect -1340 3349 -1328 3383
rect -1386 3315 -1328 3349
rect -1386 3281 -1374 3315
rect -1340 3281 -1328 3315
rect -1386 3247 -1328 3281
rect -1386 3213 -1374 3247
rect -1340 3213 -1328 3247
rect -1386 3179 -1328 3213
rect -1386 3145 -1374 3179
rect -1340 3145 -1328 3179
rect -1386 3111 -1328 3145
rect -1386 3077 -1374 3111
rect -1340 3077 -1328 3111
rect -1386 3043 -1328 3077
rect -1386 3009 -1374 3043
rect -1340 3009 -1328 3043
rect -1386 2975 -1328 3009
rect -1386 2941 -1374 2975
rect -1340 2941 -1328 2975
rect -1386 2907 -1328 2941
rect -1386 2873 -1374 2907
rect -1340 2873 -1328 2907
rect -1386 2839 -1328 2873
rect -1386 2805 -1374 2839
rect -1340 2805 -1328 2839
rect -1386 2771 -1328 2805
rect -1386 2737 -1374 2771
rect -1340 2737 -1328 2771
rect -1386 2703 -1328 2737
rect -1386 2669 -1374 2703
rect -1340 2669 -1328 2703
rect -1386 2635 -1328 2669
rect -1386 2601 -1374 2635
rect -1340 2601 -1328 2635
rect -1386 2567 -1328 2601
rect -1386 2533 -1374 2567
rect -1340 2533 -1328 2567
rect -1386 2499 -1328 2533
rect -1386 2465 -1374 2499
rect -1340 2465 -1328 2499
rect -1386 2431 -1328 2465
rect -1386 2397 -1374 2431
rect -1340 2397 -1328 2431
rect -1386 2363 -1328 2397
rect -1386 2329 -1374 2363
rect -1340 2329 -1328 2363
rect -1386 2295 -1328 2329
rect -1386 2261 -1374 2295
rect -1340 2261 -1328 2295
rect -1386 2227 -1328 2261
rect -1386 2193 -1374 2227
rect -1340 2193 -1328 2227
rect -1386 2159 -1328 2193
rect -1386 2125 -1374 2159
rect -1340 2125 -1328 2159
rect -1386 2091 -1328 2125
rect -1386 2057 -1374 2091
rect -1340 2057 -1328 2091
rect -1386 2023 -1328 2057
rect -1386 1989 -1374 2023
rect -1340 1989 -1328 2023
rect -1386 1955 -1328 1989
rect -1386 1921 -1374 1955
rect -1340 1921 -1328 1955
rect -1386 1887 -1328 1921
rect -1386 1853 -1374 1887
rect -1340 1853 -1328 1887
rect -1386 1819 -1328 1853
rect -1386 1785 -1374 1819
rect -1340 1785 -1328 1819
rect -1386 1751 -1328 1785
rect -1386 1717 -1374 1751
rect -1340 1717 -1328 1751
rect -1386 1683 -1328 1717
rect -1386 1649 -1374 1683
rect -1340 1649 -1328 1683
rect -1386 1615 -1328 1649
rect -1386 1581 -1374 1615
rect -1340 1581 -1328 1615
rect -1386 1547 -1328 1581
rect -1386 1513 -1374 1547
rect -1340 1513 -1328 1547
rect -1386 1479 -1328 1513
rect -1386 1445 -1374 1479
rect -1340 1445 -1328 1479
rect -1386 1411 -1328 1445
rect -1386 1377 -1374 1411
rect -1340 1377 -1328 1411
rect -1386 1343 -1328 1377
rect -1386 1309 -1374 1343
rect -1340 1309 -1328 1343
rect -1386 1275 -1328 1309
rect -1386 1241 -1374 1275
rect -1340 1241 -1328 1275
rect -1386 1207 -1328 1241
rect -1386 1173 -1374 1207
rect -1340 1173 -1328 1207
rect -1386 1139 -1328 1173
rect -1386 1105 -1374 1139
rect -1340 1105 -1328 1139
rect -1386 1071 -1328 1105
rect -1386 1037 -1374 1071
rect -1340 1037 -1328 1071
rect -1386 1003 -1328 1037
rect -1386 969 -1374 1003
rect -1340 969 -1328 1003
rect -1386 935 -1328 969
rect -1386 901 -1374 935
rect -1340 901 -1328 935
rect -1386 867 -1328 901
rect -1386 833 -1374 867
rect -1340 833 -1328 867
rect -1386 799 -1328 833
rect -1386 765 -1374 799
rect -1340 765 -1328 799
rect -1386 731 -1328 765
rect -1386 697 -1374 731
rect -1340 697 -1328 731
rect -1386 663 -1328 697
rect -1386 629 -1374 663
rect -1340 629 -1328 663
rect -1386 595 -1328 629
rect -1386 561 -1374 595
rect -1340 561 -1328 595
rect -1386 527 -1328 561
rect -1386 493 -1374 527
rect -1340 493 -1328 527
rect -1386 459 -1328 493
rect -1386 425 -1374 459
rect -1340 425 -1328 459
rect -1386 391 -1328 425
rect -1386 357 -1374 391
rect -1340 357 -1328 391
rect -1386 323 -1328 357
rect -1386 289 -1374 323
rect -1340 289 -1328 323
rect -1386 255 -1328 289
rect -1386 221 -1374 255
rect -1340 221 -1328 255
rect -1386 187 -1328 221
rect -1386 153 -1374 187
rect -1340 153 -1328 187
rect -1386 119 -1328 153
rect -1386 85 -1374 119
rect -1340 85 -1328 119
rect -1386 51 -1328 85
rect -1386 17 -1374 51
rect -1340 17 -1328 51
rect -1386 -17 -1328 17
rect -1386 -51 -1374 -17
rect -1340 -51 -1328 -17
rect -1386 -85 -1328 -51
rect -1386 -119 -1374 -85
rect -1340 -119 -1328 -85
rect -1386 -153 -1328 -119
rect -1386 -187 -1374 -153
rect -1340 -187 -1328 -153
rect -1386 -221 -1328 -187
rect -1386 -255 -1374 -221
rect -1340 -255 -1328 -221
rect -1386 -289 -1328 -255
rect -1386 -323 -1374 -289
rect -1340 -323 -1328 -289
rect -1386 -357 -1328 -323
rect -1386 -391 -1374 -357
rect -1340 -391 -1328 -357
rect -1386 -425 -1328 -391
rect -1386 -459 -1374 -425
rect -1340 -459 -1328 -425
rect -1386 -493 -1328 -459
rect -1386 -527 -1374 -493
rect -1340 -527 -1328 -493
rect -1386 -561 -1328 -527
rect -1386 -595 -1374 -561
rect -1340 -595 -1328 -561
rect -1386 -629 -1328 -595
rect -1386 -663 -1374 -629
rect -1340 -663 -1328 -629
rect -1386 -697 -1328 -663
rect -1386 -731 -1374 -697
rect -1340 -731 -1328 -697
rect -1386 -765 -1328 -731
rect -1386 -799 -1374 -765
rect -1340 -799 -1328 -765
rect -1386 -833 -1328 -799
rect -1386 -867 -1374 -833
rect -1340 -867 -1328 -833
rect -1386 -901 -1328 -867
rect -1386 -935 -1374 -901
rect -1340 -935 -1328 -901
rect -1386 -969 -1328 -935
rect -1386 -1003 -1374 -969
rect -1340 -1003 -1328 -969
rect -1386 -1037 -1328 -1003
rect -1386 -1071 -1374 -1037
rect -1340 -1071 -1328 -1037
rect -1386 -1105 -1328 -1071
rect -1386 -1139 -1374 -1105
rect -1340 -1139 -1328 -1105
rect -1386 -1173 -1328 -1139
rect -1386 -1207 -1374 -1173
rect -1340 -1207 -1328 -1173
rect -1386 -1241 -1328 -1207
rect -1386 -1275 -1374 -1241
rect -1340 -1275 -1328 -1241
rect -1386 -1309 -1328 -1275
rect -1386 -1343 -1374 -1309
rect -1340 -1343 -1328 -1309
rect -1386 -1377 -1328 -1343
rect -1386 -1411 -1374 -1377
rect -1340 -1411 -1328 -1377
rect -1386 -1445 -1328 -1411
rect -1386 -1479 -1374 -1445
rect -1340 -1479 -1328 -1445
rect -1386 -1513 -1328 -1479
rect -1386 -1547 -1374 -1513
rect -1340 -1547 -1328 -1513
rect -1386 -1581 -1328 -1547
rect -1386 -1615 -1374 -1581
rect -1340 -1615 -1328 -1581
rect -1386 -1649 -1328 -1615
rect -1386 -1683 -1374 -1649
rect -1340 -1683 -1328 -1649
rect -1386 -1717 -1328 -1683
rect -1386 -1751 -1374 -1717
rect -1340 -1751 -1328 -1717
rect -1386 -1785 -1328 -1751
rect -1386 -1819 -1374 -1785
rect -1340 -1819 -1328 -1785
rect -1386 -1853 -1328 -1819
rect -1386 -1887 -1374 -1853
rect -1340 -1887 -1328 -1853
rect -1386 -1921 -1328 -1887
rect -1386 -1955 -1374 -1921
rect -1340 -1955 -1328 -1921
rect -1386 -1989 -1328 -1955
rect -1386 -2023 -1374 -1989
rect -1340 -2023 -1328 -1989
rect -1386 -2057 -1328 -2023
rect -1386 -2091 -1374 -2057
rect -1340 -2091 -1328 -2057
rect -1386 -2125 -1328 -2091
rect -1386 -2159 -1374 -2125
rect -1340 -2159 -1328 -2125
rect -1386 -2193 -1328 -2159
rect -1386 -2227 -1374 -2193
rect -1340 -2227 -1328 -2193
rect -1386 -2261 -1328 -2227
rect -1386 -2295 -1374 -2261
rect -1340 -2295 -1328 -2261
rect -1386 -2329 -1328 -2295
rect -1386 -2363 -1374 -2329
rect -1340 -2363 -1328 -2329
rect -1386 -2397 -1328 -2363
rect -1386 -2431 -1374 -2397
rect -1340 -2431 -1328 -2397
rect -1386 -2465 -1328 -2431
rect -1386 -2499 -1374 -2465
rect -1340 -2499 -1328 -2465
rect -1386 -2533 -1328 -2499
rect -1386 -2567 -1374 -2533
rect -1340 -2567 -1328 -2533
rect -1386 -2601 -1328 -2567
rect -1386 -2635 -1374 -2601
rect -1340 -2635 -1328 -2601
rect -1386 -2669 -1328 -2635
rect -1386 -2703 -1374 -2669
rect -1340 -2703 -1328 -2669
rect -1386 -2737 -1328 -2703
rect -1386 -2771 -1374 -2737
rect -1340 -2771 -1328 -2737
rect -1386 -2805 -1328 -2771
rect -1386 -2839 -1374 -2805
rect -1340 -2839 -1328 -2805
rect -1386 -2873 -1328 -2839
rect -1386 -2907 -1374 -2873
rect -1340 -2907 -1328 -2873
rect -1386 -2941 -1328 -2907
rect -1386 -2975 -1374 -2941
rect -1340 -2975 -1328 -2941
rect -1386 -3009 -1328 -2975
rect -1386 -3043 -1374 -3009
rect -1340 -3043 -1328 -3009
rect -1386 -3077 -1328 -3043
rect -1386 -3111 -1374 -3077
rect -1340 -3111 -1328 -3077
rect -1386 -3145 -1328 -3111
rect -1386 -3179 -1374 -3145
rect -1340 -3179 -1328 -3145
rect -1386 -3213 -1328 -3179
rect -1386 -3247 -1374 -3213
rect -1340 -3247 -1328 -3213
rect -1386 -3281 -1328 -3247
rect -1386 -3315 -1374 -3281
rect -1340 -3315 -1328 -3281
rect -1386 -3349 -1328 -3315
rect -1386 -3383 -1374 -3349
rect -1340 -3383 -1328 -3349
rect -1386 -3417 -1328 -3383
rect -1386 -3451 -1374 -3417
rect -1340 -3451 -1328 -3417
rect -1386 -3485 -1328 -3451
rect -1386 -3519 -1374 -3485
rect -1340 -3519 -1328 -3485
rect -1386 -3553 -1328 -3519
rect -1386 -3587 -1374 -3553
rect -1340 -3587 -1328 -3553
rect -1386 -3621 -1328 -3587
rect -1386 -3655 -1374 -3621
rect -1340 -3655 -1328 -3621
rect -1386 -3689 -1328 -3655
rect -1386 -3723 -1374 -3689
rect -1340 -3723 -1328 -3689
rect -1386 -3757 -1328 -3723
rect -1386 -3791 -1374 -3757
rect -1340 -3791 -1328 -3757
rect -1386 -3825 -1328 -3791
rect -1386 -3859 -1374 -3825
rect -1340 -3859 -1328 -3825
rect -1386 -3893 -1328 -3859
rect -1386 -3927 -1374 -3893
rect -1340 -3927 -1328 -3893
rect -1386 -3961 -1328 -3927
rect -1386 -3995 -1374 -3961
rect -1340 -3995 -1328 -3961
rect -1386 -4029 -1328 -3995
rect -1386 -4063 -1374 -4029
rect -1340 -4063 -1328 -4029
rect -1386 -4097 -1328 -4063
rect -1386 -4131 -1374 -4097
rect -1340 -4131 -1328 -4097
rect -1386 -4165 -1328 -4131
rect -1386 -4199 -1374 -4165
rect -1340 -4199 -1328 -4165
rect -1386 -4233 -1328 -4199
rect -1386 -4267 -1374 -4233
rect -1340 -4267 -1328 -4233
rect -1386 -4301 -1328 -4267
rect -1386 -4335 -1374 -4301
rect -1340 -4335 -1328 -4301
rect -1386 -4369 -1328 -4335
rect -1386 -4403 -1374 -4369
rect -1340 -4403 -1328 -4369
rect -1386 -4437 -1328 -4403
rect -1386 -4471 -1374 -4437
rect -1340 -4471 -1328 -4437
rect -1386 -4505 -1328 -4471
rect -1386 -4539 -1374 -4505
rect -1340 -4539 -1328 -4505
rect -1386 -4573 -1328 -4539
rect -1386 -4607 -1374 -4573
rect -1340 -4607 -1328 -4573
rect -1386 -4641 -1328 -4607
rect -1386 -4675 -1374 -4641
rect -1340 -4675 -1328 -4641
rect -1386 -4709 -1328 -4675
rect -1386 -4743 -1374 -4709
rect -1340 -4743 -1328 -4709
rect -1386 -4777 -1328 -4743
rect -1386 -4811 -1374 -4777
rect -1340 -4811 -1328 -4777
rect -1386 -4845 -1328 -4811
rect -1386 -4879 -1374 -4845
rect -1340 -4879 -1328 -4845
rect -1386 -4913 -1328 -4879
rect -1386 -4947 -1374 -4913
rect -1340 -4947 -1328 -4913
rect -1386 -4981 -1328 -4947
rect -1386 -5015 -1374 -4981
rect -1340 -5015 -1328 -4981
rect -1386 -5049 -1328 -5015
rect -1386 -5083 -1374 -5049
rect -1340 -5083 -1328 -5049
rect -1386 -5117 -1328 -5083
rect -1386 -5151 -1374 -5117
rect -1340 -5151 -1328 -5117
rect -1386 -5185 -1328 -5151
rect -1386 -5219 -1374 -5185
rect -1340 -5219 -1328 -5185
rect -1386 -5253 -1328 -5219
rect -1386 -5287 -1374 -5253
rect -1340 -5287 -1328 -5253
rect -1386 -5321 -1328 -5287
rect -1386 -5355 -1374 -5321
rect -1340 -5355 -1328 -5321
rect -1386 -5389 -1328 -5355
rect -1386 -5423 -1374 -5389
rect -1340 -5423 -1328 -5389
rect -1386 -5457 -1328 -5423
rect -1386 -5491 -1374 -5457
rect -1340 -5491 -1328 -5457
rect -1386 -5525 -1328 -5491
rect -1386 -5559 -1374 -5525
rect -1340 -5559 -1328 -5525
rect -1386 -5593 -1328 -5559
rect -1386 -5627 -1374 -5593
rect -1340 -5627 -1328 -5593
rect -1386 -5661 -1328 -5627
rect -1386 -5695 -1374 -5661
rect -1340 -5695 -1328 -5661
rect -1386 -5729 -1328 -5695
rect -1386 -5763 -1374 -5729
rect -1340 -5763 -1328 -5729
rect -1386 -5797 -1328 -5763
rect -1386 -5831 -1374 -5797
rect -1340 -5831 -1328 -5797
rect -1386 -5865 -1328 -5831
rect -1386 -5899 -1374 -5865
rect -1340 -5899 -1328 -5865
rect -1386 -5933 -1328 -5899
rect -1386 -5967 -1374 -5933
rect -1340 -5967 -1328 -5933
rect -1386 -6001 -1328 -5967
rect -1386 -6035 -1374 -6001
rect -1340 -6035 -1328 -6001
rect -1386 -6069 -1328 -6035
rect -1386 -6103 -1374 -6069
rect -1340 -6103 -1328 -6069
rect -1386 -6137 -1328 -6103
rect -1386 -6171 -1374 -6137
rect -1340 -6171 -1328 -6137
rect -1386 -6205 -1328 -6171
rect -1386 -6239 -1374 -6205
rect -1340 -6239 -1328 -6205
rect -1386 -6273 -1328 -6239
rect -1386 -6307 -1374 -6273
rect -1340 -6307 -1328 -6273
rect -1386 -6341 -1328 -6307
rect -1386 -6375 -1374 -6341
rect -1340 -6375 -1328 -6341
rect -1386 -6409 -1328 -6375
rect -1386 -6443 -1374 -6409
rect -1340 -6443 -1328 -6409
rect -1386 -6477 -1328 -6443
rect -1386 -6511 -1374 -6477
rect -1340 -6511 -1328 -6477
rect -1386 -6545 -1328 -6511
rect -1386 -6579 -1374 -6545
rect -1340 -6579 -1328 -6545
rect -1386 -6613 -1328 -6579
rect -1386 -6647 -1374 -6613
rect -1340 -6647 -1328 -6613
rect -1386 -6681 -1328 -6647
rect -1386 -6715 -1374 -6681
rect -1340 -6715 -1328 -6681
rect -1386 -6749 -1328 -6715
rect -1386 -6783 -1374 -6749
rect -1340 -6783 -1328 -6749
rect -1386 -6817 -1328 -6783
rect -1386 -6851 -1374 -6817
rect -1340 -6851 -1328 -6817
rect -1386 -6885 -1328 -6851
rect -1386 -6919 -1374 -6885
rect -1340 -6919 -1328 -6885
rect -1386 -6953 -1328 -6919
rect -1386 -6987 -1374 -6953
rect -1340 -6987 -1328 -6953
rect -1386 -7021 -1328 -6987
rect -1386 -7055 -1374 -7021
rect -1340 -7055 -1328 -7021
rect -1386 -7089 -1328 -7055
rect -1386 -7123 -1374 -7089
rect -1340 -7123 -1328 -7089
rect -1386 -7157 -1328 -7123
rect -1386 -7191 -1374 -7157
rect -1340 -7191 -1328 -7157
rect -1386 -7225 -1328 -7191
rect -1386 -7259 -1374 -7225
rect -1340 -7259 -1328 -7225
rect -1386 -7293 -1328 -7259
rect -1386 -7327 -1374 -7293
rect -1340 -7327 -1328 -7293
rect -1386 -7361 -1328 -7327
rect -1386 -7395 -1374 -7361
rect -1340 -7395 -1328 -7361
rect -1386 -7429 -1328 -7395
rect -1386 -7463 -1374 -7429
rect -1340 -7463 -1328 -7429
rect -1386 -7497 -1328 -7463
rect -1386 -7531 -1374 -7497
rect -1340 -7531 -1328 -7497
rect -1386 -7565 -1328 -7531
rect -1386 -7599 -1374 -7565
rect -1340 -7599 -1328 -7565
rect -1386 -7633 -1328 -7599
rect -1386 -7667 -1374 -7633
rect -1340 -7667 -1328 -7633
rect -1386 -7701 -1328 -7667
rect -1386 -7735 -1374 -7701
rect -1340 -7735 -1328 -7701
rect -1386 -7769 -1328 -7735
rect -1386 -7803 -1374 -7769
rect -1340 -7803 -1328 -7769
rect -1386 -7837 -1328 -7803
rect -1386 -7871 -1374 -7837
rect -1340 -7871 -1328 -7837
rect -1386 -7905 -1328 -7871
rect -1386 -7939 -1374 -7905
rect -1340 -7939 -1328 -7905
rect -1386 -7973 -1328 -7939
rect -1386 -8007 -1374 -7973
rect -1340 -8007 -1328 -7973
rect -1386 -8041 -1328 -8007
rect -1386 -8075 -1374 -8041
rect -1340 -8075 -1328 -8041
rect -1386 -8109 -1328 -8075
rect -1386 -8143 -1374 -8109
rect -1340 -8143 -1328 -8109
rect -1386 -8177 -1328 -8143
rect -1386 -8211 -1374 -8177
rect -1340 -8211 -1328 -8177
rect -1386 -8245 -1328 -8211
rect -1386 -8279 -1374 -8245
rect -1340 -8279 -1328 -8245
rect -1386 -8313 -1328 -8279
rect -1386 -8347 -1374 -8313
rect -1340 -8347 -1328 -8313
rect -1386 -8381 -1328 -8347
rect -1386 -8415 -1374 -8381
rect -1340 -8415 -1328 -8381
rect -1386 -8449 -1328 -8415
rect -1386 -8483 -1374 -8449
rect -1340 -8483 -1328 -8449
rect -1386 -8517 -1328 -8483
rect -1386 -8551 -1374 -8517
rect -1340 -8551 -1328 -8517
rect -1386 -8585 -1328 -8551
rect -1386 -8619 -1374 -8585
rect -1340 -8619 -1328 -8585
rect -1386 -8653 -1328 -8619
rect -1386 -8687 -1374 -8653
rect -1340 -8687 -1328 -8653
rect -1386 -8721 -1328 -8687
rect -1386 -8755 -1374 -8721
rect -1340 -8755 -1328 -8721
rect -1386 -8789 -1328 -8755
rect -1386 -8823 -1374 -8789
rect -1340 -8823 -1328 -8789
rect -1386 -8857 -1328 -8823
rect -1386 -8891 -1374 -8857
rect -1340 -8891 -1328 -8857
rect -1386 -8925 -1328 -8891
rect -1386 -8959 -1374 -8925
rect -1340 -8959 -1328 -8925
rect -1386 -8993 -1328 -8959
rect -1386 -9027 -1374 -8993
rect -1340 -9027 -1328 -8993
rect -1386 -9061 -1328 -9027
rect -1386 -9095 -1374 -9061
rect -1340 -9095 -1328 -9061
rect -1386 -9129 -1328 -9095
rect -1386 -9163 -1374 -9129
rect -1340 -9163 -1328 -9129
rect -1386 -9197 -1328 -9163
rect -1386 -9231 -1374 -9197
rect -1340 -9231 -1328 -9197
rect -1386 -9265 -1328 -9231
rect -1386 -9299 -1374 -9265
rect -1340 -9299 -1328 -9265
rect -1386 -9333 -1328 -9299
rect -1386 -9367 -1374 -9333
rect -1340 -9367 -1328 -9333
rect -1386 -9401 -1328 -9367
rect -1386 -9435 -1374 -9401
rect -1340 -9435 -1328 -9401
rect -1386 -9469 -1328 -9435
rect -1386 -9503 -1374 -9469
rect -1340 -9503 -1328 -9469
rect -1386 -9537 -1328 -9503
rect -1386 -9571 -1374 -9537
rect -1340 -9571 -1328 -9537
rect -1386 -9600 -1328 -9571
rect -1268 9571 -1210 9600
rect -1268 9537 -1256 9571
rect -1222 9537 -1210 9571
rect -1268 9503 -1210 9537
rect -1268 9469 -1256 9503
rect -1222 9469 -1210 9503
rect -1268 9435 -1210 9469
rect -1268 9401 -1256 9435
rect -1222 9401 -1210 9435
rect -1268 9367 -1210 9401
rect -1268 9333 -1256 9367
rect -1222 9333 -1210 9367
rect -1268 9299 -1210 9333
rect -1268 9265 -1256 9299
rect -1222 9265 -1210 9299
rect -1268 9231 -1210 9265
rect -1268 9197 -1256 9231
rect -1222 9197 -1210 9231
rect -1268 9163 -1210 9197
rect -1268 9129 -1256 9163
rect -1222 9129 -1210 9163
rect -1268 9095 -1210 9129
rect -1268 9061 -1256 9095
rect -1222 9061 -1210 9095
rect -1268 9027 -1210 9061
rect -1268 8993 -1256 9027
rect -1222 8993 -1210 9027
rect -1268 8959 -1210 8993
rect -1268 8925 -1256 8959
rect -1222 8925 -1210 8959
rect -1268 8891 -1210 8925
rect -1268 8857 -1256 8891
rect -1222 8857 -1210 8891
rect -1268 8823 -1210 8857
rect -1268 8789 -1256 8823
rect -1222 8789 -1210 8823
rect -1268 8755 -1210 8789
rect -1268 8721 -1256 8755
rect -1222 8721 -1210 8755
rect -1268 8687 -1210 8721
rect -1268 8653 -1256 8687
rect -1222 8653 -1210 8687
rect -1268 8619 -1210 8653
rect -1268 8585 -1256 8619
rect -1222 8585 -1210 8619
rect -1268 8551 -1210 8585
rect -1268 8517 -1256 8551
rect -1222 8517 -1210 8551
rect -1268 8483 -1210 8517
rect -1268 8449 -1256 8483
rect -1222 8449 -1210 8483
rect -1268 8415 -1210 8449
rect -1268 8381 -1256 8415
rect -1222 8381 -1210 8415
rect -1268 8347 -1210 8381
rect -1268 8313 -1256 8347
rect -1222 8313 -1210 8347
rect -1268 8279 -1210 8313
rect -1268 8245 -1256 8279
rect -1222 8245 -1210 8279
rect -1268 8211 -1210 8245
rect -1268 8177 -1256 8211
rect -1222 8177 -1210 8211
rect -1268 8143 -1210 8177
rect -1268 8109 -1256 8143
rect -1222 8109 -1210 8143
rect -1268 8075 -1210 8109
rect -1268 8041 -1256 8075
rect -1222 8041 -1210 8075
rect -1268 8007 -1210 8041
rect -1268 7973 -1256 8007
rect -1222 7973 -1210 8007
rect -1268 7939 -1210 7973
rect -1268 7905 -1256 7939
rect -1222 7905 -1210 7939
rect -1268 7871 -1210 7905
rect -1268 7837 -1256 7871
rect -1222 7837 -1210 7871
rect -1268 7803 -1210 7837
rect -1268 7769 -1256 7803
rect -1222 7769 -1210 7803
rect -1268 7735 -1210 7769
rect -1268 7701 -1256 7735
rect -1222 7701 -1210 7735
rect -1268 7667 -1210 7701
rect -1268 7633 -1256 7667
rect -1222 7633 -1210 7667
rect -1268 7599 -1210 7633
rect -1268 7565 -1256 7599
rect -1222 7565 -1210 7599
rect -1268 7531 -1210 7565
rect -1268 7497 -1256 7531
rect -1222 7497 -1210 7531
rect -1268 7463 -1210 7497
rect -1268 7429 -1256 7463
rect -1222 7429 -1210 7463
rect -1268 7395 -1210 7429
rect -1268 7361 -1256 7395
rect -1222 7361 -1210 7395
rect -1268 7327 -1210 7361
rect -1268 7293 -1256 7327
rect -1222 7293 -1210 7327
rect -1268 7259 -1210 7293
rect -1268 7225 -1256 7259
rect -1222 7225 -1210 7259
rect -1268 7191 -1210 7225
rect -1268 7157 -1256 7191
rect -1222 7157 -1210 7191
rect -1268 7123 -1210 7157
rect -1268 7089 -1256 7123
rect -1222 7089 -1210 7123
rect -1268 7055 -1210 7089
rect -1268 7021 -1256 7055
rect -1222 7021 -1210 7055
rect -1268 6987 -1210 7021
rect -1268 6953 -1256 6987
rect -1222 6953 -1210 6987
rect -1268 6919 -1210 6953
rect -1268 6885 -1256 6919
rect -1222 6885 -1210 6919
rect -1268 6851 -1210 6885
rect -1268 6817 -1256 6851
rect -1222 6817 -1210 6851
rect -1268 6783 -1210 6817
rect -1268 6749 -1256 6783
rect -1222 6749 -1210 6783
rect -1268 6715 -1210 6749
rect -1268 6681 -1256 6715
rect -1222 6681 -1210 6715
rect -1268 6647 -1210 6681
rect -1268 6613 -1256 6647
rect -1222 6613 -1210 6647
rect -1268 6579 -1210 6613
rect -1268 6545 -1256 6579
rect -1222 6545 -1210 6579
rect -1268 6511 -1210 6545
rect -1268 6477 -1256 6511
rect -1222 6477 -1210 6511
rect -1268 6443 -1210 6477
rect -1268 6409 -1256 6443
rect -1222 6409 -1210 6443
rect -1268 6375 -1210 6409
rect -1268 6341 -1256 6375
rect -1222 6341 -1210 6375
rect -1268 6307 -1210 6341
rect -1268 6273 -1256 6307
rect -1222 6273 -1210 6307
rect -1268 6239 -1210 6273
rect -1268 6205 -1256 6239
rect -1222 6205 -1210 6239
rect -1268 6171 -1210 6205
rect -1268 6137 -1256 6171
rect -1222 6137 -1210 6171
rect -1268 6103 -1210 6137
rect -1268 6069 -1256 6103
rect -1222 6069 -1210 6103
rect -1268 6035 -1210 6069
rect -1268 6001 -1256 6035
rect -1222 6001 -1210 6035
rect -1268 5967 -1210 6001
rect -1268 5933 -1256 5967
rect -1222 5933 -1210 5967
rect -1268 5899 -1210 5933
rect -1268 5865 -1256 5899
rect -1222 5865 -1210 5899
rect -1268 5831 -1210 5865
rect -1268 5797 -1256 5831
rect -1222 5797 -1210 5831
rect -1268 5763 -1210 5797
rect -1268 5729 -1256 5763
rect -1222 5729 -1210 5763
rect -1268 5695 -1210 5729
rect -1268 5661 -1256 5695
rect -1222 5661 -1210 5695
rect -1268 5627 -1210 5661
rect -1268 5593 -1256 5627
rect -1222 5593 -1210 5627
rect -1268 5559 -1210 5593
rect -1268 5525 -1256 5559
rect -1222 5525 -1210 5559
rect -1268 5491 -1210 5525
rect -1268 5457 -1256 5491
rect -1222 5457 -1210 5491
rect -1268 5423 -1210 5457
rect -1268 5389 -1256 5423
rect -1222 5389 -1210 5423
rect -1268 5355 -1210 5389
rect -1268 5321 -1256 5355
rect -1222 5321 -1210 5355
rect -1268 5287 -1210 5321
rect -1268 5253 -1256 5287
rect -1222 5253 -1210 5287
rect -1268 5219 -1210 5253
rect -1268 5185 -1256 5219
rect -1222 5185 -1210 5219
rect -1268 5151 -1210 5185
rect -1268 5117 -1256 5151
rect -1222 5117 -1210 5151
rect -1268 5083 -1210 5117
rect -1268 5049 -1256 5083
rect -1222 5049 -1210 5083
rect -1268 5015 -1210 5049
rect -1268 4981 -1256 5015
rect -1222 4981 -1210 5015
rect -1268 4947 -1210 4981
rect -1268 4913 -1256 4947
rect -1222 4913 -1210 4947
rect -1268 4879 -1210 4913
rect -1268 4845 -1256 4879
rect -1222 4845 -1210 4879
rect -1268 4811 -1210 4845
rect -1268 4777 -1256 4811
rect -1222 4777 -1210 4811
rect -1268 4743 -1210 4777
rect -1268 4709 -1256 4743
rect -1222 4709 -1210 4743
rect -1268 4675 -1210 4709
rect -1268 4641 -1256 4675
rect -1222 4641 -1210 4675
rect -1268 4607 -1210 4641
rect -1268 4573 -1256 4607
rect -1222 4573 -1210 4607
rect -1268 4539 -1210 4573
rect -1268 4505 -1256 4539
rect -1222 4505 -1210 4539
rect -1268 4471 -1210 4505
rect -1268 4437 -1256 4471
rect -1222 4437 -1210 4471
rect -1268 4403 -1210 4437
rect -1268 4369 -1256 4403
rect -1222 4369 -1210 4403
rect -1268 4335 -1210 4369
rect -1268 4301 -1256 4335
rect -1222 4301 -1210 4335
rect -1268 4267 -1210 4301
rect -1268 4233 -1256 4267
rect -1222 4233 -1210 4267
rect -1268 4199 -1210 4233
rect -1268 4165 -1256 4199
rect -1222 4165 -1210 4199
rect -1268 4131 -1210 4165
rect -1268 4097 -1256 4131
rect -1222 4097 -1210 4131
rect -1268 4063 -1210 4097
rect -1268 4029 -1256 4063
rect -1222 4029 -1210 4063
rect -1268 3995 -1210 4029
rect -1268 3961 -1256 3995
rect -1222 3961 -1210 3995
rect -1268 3927 -1210 3961
rect -1268 3893 -1256 3927
rect -1222 3893 -1210 3927
rect -1268 3859 -1210 3893
rect -1268 3825 -1256 3859
rect -1222 3825 -1210 3859
rect -1268 3791 -1210 3825
rect -1268 3757 -1256 3791
rect -1222 3757 -1210 3791
rect -1268 3723 -1210 3757
rect -1268 3689 -1256 3723
rect -1222 3689 -1210 3723
rect -1268 3655 -1210 3689
rect -1268 3621 -1256 3655
rect -1222 3621 -1210 3655
rect -1268 3587 -1210 3621
rect -1268 3553 -1256 3587
rect -1222 3553 -1210 3587
rect -1268 3519 -1210 3553
rect -1268 3485 -1256 3519
rect -1222 3485 -1210 3519
rect -1268 3451 -1210 3485
rect -1268 3417 -1256 3451
rect -1222 3417 -1210 3451
rect -1268 3383 -1210 3417
rect -1268 3349 -1256 3383
rect -1222 3349 -1210 3383
rect -1268 3315 -1210 3349
rect -1268 3281 -1256 3315
rect -1222 3281 -1210 3315
rect -1268 3247 -1210 3281
rect -1268 3213 -1256 3247
rect -1222 3213 -1210 3247
rect -1268 3179 -1210 3213
rect -1268 3145 -1256 3179
rect -1222 3145 -1210 3179
rect -1268 3111 -1210 3145
rect -1268 3077 -1256 3111
rect -1222 3077 -1210 3111
rect -1268 3043 -1210 3077
rect -1268 3009 -1256 3043
rect -1222 3009 -1210 3043
rect -1268 2975 -1210 3009
rect -1268 2941 -1256 2975
rect -1222 2941 -1210 2975
rect -1268 2907 -1210 2941
rect -1268 2873 -1256 2907
rect -1222 2873 -1210 2907
rect -1268 2839 -1210 2873
rect -1268 2805 -1256 2839
rect -1222 2805 -1210 2839
rect -1268 2771 -1210 2805
rect -1268 2737 -1256 2771
rect -1222 2737 -1210 2771
rect -1268 2703 -1210 2737
rect -1268 2669 -1256 2703
rect -1222 2669 -1210 2703
rect -1268 2635 -1210 2669
rect -1268 2601 -1256 2635
rect -1222 2601 -1210 2635
rect -1268 2567 -1210 2601
rect -1268 2533 -1256 2567
rect -1222 2533 -1210 2567
rect -1268 2499 -1210 2533
rect -1268 2465 -1256 2499
rect -1222 2465 -1210 2499
rect -1268 2431 -1210 2465
rect -1268 2397 -1256 2431
rect -1222 2397 -1210 2431
rect -1268 2363 -1210 2397
rect -1268 2329 -1256 2363
rect -1222 2329 -1210 2363
rect -1268 2295 -1210 2329
rect -1268 2261 -1256 2295
rect -1222 2261 -1210 2295
rect -1268 2227 -1210 2261
rect -1268 2193 -1256 2227
rect -1222 2193 -1210 2227
rect -1268 2159 -1210 2193
rect -1268 2125 -1256 2159
rect -1222 2125 -1210 2159
rect -1268 2091 -1210 2125
rect -1268 2057 -1256 2091
rect -1222 2057 -1210 2091
rect -1268 2023 -1210 2057
rect -1268 1989 -1256 2023
rect -1222 1989 -1210 2023
rect -1268 1955 -1210 1989
rect -1268 1921 -1256 1955
rect -1222 1921 -1210 1955
rect -1268 1887 -1210 1921
rect -1268 1853 -1256 1887
rect -1222 1853 -1210 1887
rect -1268 1819 -1210 1853
rect -1268 1785 -1256 1819
rect -1222 1785 -1210 1819
rect -1268 1751 -1210 1785
rect -1268 1717 -1256 1751
rect -1222 1717 -1210 1751
rect -1268 1683 -1210 1717
rect -1268 1649 -1256 1683
rect -1222 1649 -1210 1683
rect -1268 1615 -1210 1649
rect -1268 1581 -1256 1615
rect -1222 1581 -1210 1615
rect -1268 1547 -1210 1581
rect -1268 1513 -1256 1547
rect -1222 1513 -1210 1547
rect -1268 1479 -1210 1513
rect -1268 1445 -1256 1479
rect -1222 1445 -1210 1479
rect -1268 1411 -1210 1445
rect -1268 1377 -1256 1411
rect -1222 1377 -1210 1411
rect -1268 1343 -1210 1377
rect -1268 1309 -1256 1343
rect -1222 1309 -1210 1343
rect -1268 1275 -1210 1309
rect -1268 1241 -1256 1275
rect -1222 1241 -1210 1275
rect -1268 1207 -1210 1241
rect -1268 1173 -1256 1207
rect -1222 1173 -1210 1207
rect -1268 1139 -1210 1173
rect -1268 1105 -1256 1139
rect -1222 1105 -1210 1139
rect -1268 1071 -1210 1105
rect -1268 1037 -1256 1071
rect -1222 1037 -1210 1071
rect -1268 1003 -1210 1037
rect -1268 969 -1256 1003
rect -1222 969 -1210 1003
rect -1268 935 -1210 969
rect -1268 901 -1256 935
rect -1222 901 -1210 935
rect -1268 867 -1210 901
rect -1268 833 -1256 867
rect -1222 833 -1210 867
rect -1268 799 -1210 833
rect -1268 765 -1256 799
rect -1222 765 -1210 799
rect -1268 731 -1210 765
rect -1268 697 -1256 731
rect -1222 697 -1210 731
rect -1268 663 -1210 697
rect -1268 629 -1256 663
rect -1222 629 -1210 663
rect -1268 595 -1210 629
rect -1268 561 -1256 595
rect -1222 561 -1210 595
rect -1268 527 -1210 561
rect -1268 493 -1256 527
rect -1222 493 -1210 527
rect -1268 459 -1210 493
rect -1268 425 -1256 459
rect -1222 425 -1210 459
rect -1268 391 -1210 425
rect -1268 357 -1256 391
rect -1222 357 -1210 391
rect -1268 323 -1210 357
rect -1268 289 -1256 323
rect -1222 289 -1210 323
rect -1268 255 -1210 289
rect -1268 221 -1256 255
rect -1222 221 -1210 255
rect -1268 187 -1210 221
rect -1268 153 -1256 187
rect -1222 153 -1210 187
rect -1268 119 -1210 153
rect -1268 85 -1256 119
rect -1222 85 -1210 119
rect -1268 51 -1210 85
rect -1268 17 -1256 51
rect -1222 17 -1210 51
rect -1268 -17 -1210 17
rect -1268 -51 -1256 -17
rect -1222 -51 -1210 -17
rect -1268 -85 -1210 -51
rect -1268 -119 -1256 -85
rect -1222 -119 -1210 -85
rect -1268 -153 -1210 -119
rect -1268 -187 -1256 -153
rect -1222 -187 -1210 -153
rect -1268 -221 -1210 -187
rect -1268 -255 -1256 -221
rect -1222 -255 -1210 -221
rect -1268 -289 -1210 -255
rect -1268 -323 -1256 -289
rect -1222 -323 -1210 -289
rect -1268 -357 -1210 -323
rect -1268 -391 -1256 -357
rect -1222 -391 -1210 -357
rect -1268 -425 -1210 -391
rect -1268 -459 -1256 -425
rect -1222 -459 -1210 -425
rect -1268 -493 -1210 -459
rect -1268 -527 -1256 -493
rect -1222 -527 -1210 -493
rect -1268 -561 -1210 -527
rect -1268 -595 -1256 -561
rect -1222 -595 -1210 -561
rect -1268 -629 -1210 -595
rect -1268 -663 -1256 -629
rect -1222 -663 -1210 -629
rect -1268 -697 -1210 -663
rect -1268 -731 -1256 -697
rect -1222 -731 -1210 -697
rect -1268 -765 -1210 -731
rect -1268 -799 -1256 -765
rect -1222 -799 -1210 -765
rect -1268 -833 -1210 -799
rect -1268 -867 -1256 -833
rect -1222 -867 -1210 -833
rect -1268 -901 -1210 -867
rect -1268 -935 -1256 -901
rect -1222 -935 -1210 -901
rect -1268 -969 -1210 -935
rect -1268 -1003 -1256 -969
rect -1222 -1003 -1210 -969
rect -1268 -1037 -1210 -1003
rect -1268 -1071 -1256 -1037
rect -1222 -1071 -1210 -1037
rect -1268 -1105 -1210 -1071
rect -1268 -1139 -1256 -1105
rect -1222 -1139 -1210 -1105
rect -1268 -1173 -1210 -1139
rect -1268 -1207 -1256 -1173
rect -1222 -1207 -1210 -1173
rect -1268 -1241 -1210 -1207
rect -1268 -1275 -1256 -1241
rect -1222 -1275 -1210 -1241
rect -1268 -1309 -1210 -1275
rect -1268 -1343 -1256 -1309
rect -1222 -1343 -1210 -1309
rect -1268 -1377 -1210 -1343
rect -1268 -1411 -1256 -1377
rect -1222 -1411 -1210 -1377
rect -1268 -1445 -1210 -1411
rect -1268 -1479 -1256 -1445
rect -1222 -1479 -1210 -1445
rect -1268 -1513 -1210 -1479
rect -1268 -1547 -1256 -1513
rect -1222 -1547 -1210 -1513
rect -1268 -1581 -1210 -1547
rect -1268 -1615 -1256 -1581
rect -1222 -1615 -1210 -1581
rect -1268 -1649 -1210 -1615
rect -1268 -1683 -1256 -1649
rect -1222 -1683 -1210 -1649
rect -1268 -1717 -1210 -1683
rect -1268 -1751 -1256 -1717
rect -1222 -1751 -1210 -1717
rect -1268 -1785 -1210 -1751
rect -1268 -1819 -1256 -1785
rect -1222 -1819 -1210 -1785
rect -1268 -1853 -1210 -1819
rect -1268 -1887 -1256 -1853
rect -1222 -1887 -1210 -1853
rect -1268 -1921 -1210 -1887
rect -1268 -1955 -1256 -1921
rect -1222 -1955 -1210 -1921
rect -1268 -1989 -1210 -1955
rect -1268 -2023 -1256 -1989
rect -1222 -2023 -1210 -1989
rect -1268 -2057 -1210 -2023
rect -1268 -2091 -1256 -2057
rect -1222 -2091 -1210 -2057
rect -1268 -2125 -1210 -2091
rect -1268 -2159 -1256 -2125
rect -1222 -2159 -1210 -2125
rect -1268 -2193 -1210 -2159
rect -1268 -2227 -1256 -2193
rect -1222 -2227 -1210 -2193
rect -1268 -2261 -1210 -2227
rect -1268 -2295 -1256 -2261
rect -1222 -2295 -1210 -2261
rect -1268 -2329 -1210 -2295
rect -1268 -2363 -1256 -2329
rect -1222 -2363 -1210 -2329
rect -1268 -2397 -1210 -2363
rect -1268 -2431 -1256 -2397
rect -1222 -2431 -1210 -2397
rect -1268 -2465 -1210 -2431
rect -1268 -2499 -1256 -2465
rect -1222 -2499 -1210 -2465
rect -1268 -2533 -1210 -2499
rect -1268 -2567 -1256 -2533
rect -1222 -2567 -1210 -2533
rect -1268 -2601 -1210 -2567
rect -1268 -2635 -1256 -2601
rect -1222 -2635 -1210 -2601
rect -1268 -2669 -1210 -2635
rect -1268 -2703 -1256 -2669
rect -1222 -2703 -1210 -2669
rect -1268 -2737 -1210 -2703
rect -1268 -2771 -1256 -2737
rect -1222 -2771 -1210 -2737
rect -1268 -2805 -1210 -2771
rect -1268 -2839 -1256 -2805
rect -1222 -2839 -1210 -2805
rect -1268 -2873 -1210 -2839
rect -1268 -2907 -1256 -2873
rect -1222 -2907 -1210 -2873
rect -1268 -2941 -1210 -2907
rect -1268 -2975 -1256 -2941
rect -1222 -2975 -1210 -2941
rect -1268 -3009 -1210 -2975
rect -1268 -3043 -1256 -3009
rect -1222 -3043 -1210 -3009
rect -1268 -3077 -1210 -3043
rect -1268 -3111 -1256 -3077
rect -1222 -3111 -1210 -3077
rect -1268 -3145 -1210 -3111
rect -1268 -3179 -1256 -3145
rect -1222 -3179 -1210 -3145
rect -1268 -3213 -1210 -3179
rect -1268 -3247 -1256 -3213
rect -1222 -3247 -1210 -3213
rect -1268 -3281 -1210 -3247
rect -1268 -3315 -1256 -3281
rect -1222 -3315 -1210 -3281
rect -1268 -3349 -1210 -3315
rect -1268 -3383 -1256 -3349
rect -1222 -3383 -1210 -3349
rect -1268 -3417 -1210 -3383
rect -1268 -3451 -1256 -3417
rect -1222 -3451 -1210 -3417
rect -1268 -3485 -1210 -3451
rect -1268 -3519 -1256 -3485
rect -1222 -3519 -1210 -3485
rect -1268 -3553 -1210 -3519
rect -1268 -3587 -1256 -3553
rect -1222 -3587 -1210 -3553
rect -1268 -3621 -1210 -3587
rect -1268 -3655 -1256 -3621
rect -1222 -3655 -1210 -3621
rect -1268 -3689 -1210 -3655
rect -1268 -3723 -1256 -3689
rect -1222 -3723 -1210 -3689
rect -1268 -3757 -1210 -3723
rect -1268 -3791 -1256 -3757
rect -1222 -3791 -1210 -3757
rect -1268 -3825 -1210 -3791
rect -1268 -3859 -1256 -3825
rect -1222 -3859 -1210 -3825
rect -1268 -3893 -1210 -3859
rect -1268 -3927 -1256 -3893
rect -1222 -3927 -1210 -3893
rect -1268 -3961 -1210 -3927
rect -1268 -3995 -1256 -3961
rect -1222 -3995 -1210 -3961
rect -1268 -4029 -1210 -3995
rect -1268 -4063 -1256 -4029
rect -1222 -4063 -1210 -4029
rect -1268 -4097 -1210 -4063
rect -1268 -4131 -1256 -4097
rect -1222 -4131 -1210 -4097
rect -1268 -4165 -1210 -4131
rect -1268 -4199 -1256 -4165
rect -1222 -4199 -1210 -4165
rect -1268 -4233 -1210 -4199
rect -1268 -4267 -1256 -4233
rect -1222 -4267 -1210 -4233
rect -1268 -4301 -1210 -4267
rect -1268 -4335 -1256 -4301
rect -1222 -4335 -1210 -4301
rect -1268 -4369 -1210 -4335
rect -1268 -4403 -1256 -4369
rect -1222 -4403 -1210 -4369
rect -1268 -4437 -1210 -4403
rect -1268 -4471 -1256 -4437
rect -1222 -4471 -1210 -4437
rect -1268 -4505 -1210 -4471
rect -1268 -4539 -1256 -4505
rect -1222 -4539 -1210 -4505
rect -1268 -4573 -1210 -4539
rect -1268 -4607 -1256 -4573
rect -1222 -4607 -1210 -4573
rect -1268 -4641 -1210 -4607
rect -1268 -4675 -1256 -4641
rect -1222 -4675 -1210 -4641
rect -1268 -4709 -1210 -4675
rect -1268 -4743 -1256 -4709
rect -1222 -4743 -1210 -4709
rect -1268 -4777 -1210 -4743
rect -1268 -4811 -1256 -4777
rect -1222 -4811 -1210 -4777
rect -1268 -4845 -1210 -4811
rect -1268 -4879 -1256 -4845
rect -1222 -4879 -1210 -4845
rect -1268 -4913 -1210 -4879
rect -1268 -4947 -1256 -4913
rect -1222 -4947 -1210 -4913
rect -1268 -4981 -1210 -4947
rect -1268 -5015 -1256 -4981
rect -1222 -5015 -1210 -4981
rect -1268 -5049 -1210 -5015
rect -1268 -5083 -1256 -5049
rect -1222 -5083 -1210 -5049
rect -1268 -5117 -1210 -5083
rect -1268 -5151 -1256 -5117
rect -1222 -5151 -1210 -5117
rect -1268 -5185 -1210 -5151
rect -1268 -5219 -1256 -5185
rect -1222 -5219 -1210 -5185
rect -1268 -5253 -1210 -5219
rect -1268 -5287 -1256 -5253
rect -1222 -5287 -1210 -5253
rect -1268 -5321 -1210 -5287
rect -1268 -5355 -1256 -5321
rect -1222 -5355 -1210 -5321
rect -1268 -5389 -1210 -5355
rect -1268 -5423 -1256 -5389
rect -1222 -5423 -1210 -5389
rect -1268 -5457 -1210 -5423
rect -1268 -5491 -1256 -5457
rect -1222 -5491 -1210 -5457
rect -1268 -5525 -1210 -5491
rect -1268 -5559 -1256 -5525
rect -1222 -5559 -1210 -5525
rect -1268 -5593 -1210 -5559
rect -1268 -5627 -1256 -5593
rect -1222 -5627 -1210 -5593
rect -1268 -5661 -1210 -5627
rect -1268 -5695 -1256 -5661
rect -1222 -5695 -1210 -5661
rect -1268 -5729 -1210 -5695
rect -1268 -5763 -1256 -5729
rect -1222 -5763 -1210 -5729
rect -1268 -5797 -1210 -5763
rect -1268 -5831 -1256 -5797
rect -1222 -5831 -1210 -5797
rect -1268 -5865 -1210 -5831
rect -1268 -5899 -1256 -5865
rect -1222 -5899 -1210 -5865
rect -1268 -5933 -1210 -5899
rect -1268 -5967 -1256 -5933
rect -1222 -5967 -1210 -5933
rect -1268 -6001 -1210 -5967
rect -1268 -6035 -1256 -6001
rect -1222 -6035 -1210 -6001
rect -1268 -6069 -1210 -6035
rect -1268 -6103 -1256 -6069
rect -1222 -6103 -1210 -6069
rect -1268 -6137 -1210 -6103
rect -1268 -6171 -1256 -6137
rect -1222 -6171 -1210 -6137
rect -1268 -6205 -1210 -6171
rect -1268 -6239 -1256 -6205
rect -1222 -6239 -1210 -6205
rect -1268 -6273 -1210 -6239
rect -1268 -6307 -1256 -6273
rect -1222 -6307 -1210 -6273
rect -1268 -6341 -1210 -6307
rect -1268 -6375 -1256 -6341
rect -1222 -6375 -1210 -6341
rect -1268 -6409 -1210 -6375
rect -1268 -6443 -1256 -6409
rect -1222 -6443 -1210 -6409
rect -1268 -6477 -1210 -6443
rect -1268 -6511 -1256 -6477
rect -1222 -6511 -1210 -6477
rect -1268 -6545 -1210 -6511
rect -1268 -6579 -1256 -6545
rect -1222 -6579 -1210 -6545
rect -1268 -6613 -1210 -6579
rect -1268 -6647 -1256 -6613
rect -1222 -6647 -1210 -6613
rect -1268 -6681 -1210 -6647
rect -1268 -6715 -1256 -6681
rect -1222 -6715 -1210 -6681
rect -1268 -6749 -1210 -6715
rect -1268 -6783 -1256 -6749
rect -1222 -6783 -1210 -6749
rect -1268 -6817 -1210 -6783
rect -1268 -6851 -1256 -6817
rect -1222 -6851 -1210 -6817
rect -1268 -6885 -1210 -6851
rect -1268 -6919 -1256 -6885
rect -1222 -6919 -1210 -6885
rect -1268 -6953 -1210 -6919
rect -1268 -6987 -1256 -6953
rect -1222 -6987 -1210 -6953
rect -1268 -7021 -1210 -6987
rect -1268 -7055 -1256 -7021
rect -1222 -7055 -1210 -7021
rect -1268 -7089 -1210 -7055
rect -1268 -7123 -1256 -7089
rect -1222 -7123 -1210 -7089
rect -1268 -7157 -1210 -7123
rect -1268 -7191 -1256 -7157
rect -1222 -7191 -1210 -7157
rect -1268 -7225 -1210 -7191
rect -1268 -7259 -1256 -7225
rect -1222 -7259 -1210 -7225
rect -1268 -7293 -1210 -7259
rect -1268 -7327 -1256 -7293
rect -1222 -7327 -1210 -7293
rect -1268 -7361 -1210 -7327
rect -1268 -7395 -1256 -7361
rect -1222 -7395 -1210 -7361
rect -1268 -7429 -1210 -7395
rect -1268 -7463 -1256 -7429
rect -1222 -7463 -1210 -7429
rect -1268 -7497 -1210 -7463
rect -1268 -7531 -1256 -7497
rect -1222 -7531 -1210 -7497
rect -1268 -7565 -1210 -7531
rect -1268 -7599 -1256 -7565
rect -1222 -7599 -1210 -7565
rect -1268 -7633 -1210 -7599
rect -1268 -7667 -1256 -7633
rect -1222 -7667 -1210 -7633
rect -1268 -7701 -1210 -7667
rect -1268 -7735 -1256 -7701
rect -1222 -7735 -1210 -7701
rect -1268 -7769 -1210 -7735
rect -1268 -7803 -1256 -7769
rect -1222 -7803 -1210 -7769
rect -1268 -7837 -1210 -7803
rect -1268 -7871 -1256 -7837
rect -1222 -7871 -1210 -7837
rect -1268 -7905 -1210 -7871
rect -1268 -7939 -1256 -7905
rect -1222 -7939 -1210 -7905
rect -1268 -7973 -1210 -7939
rect -1268 -8007 -1256 -7973
rect -1222 -8007 -1210 -7973
rect -1268 -8041 -1210 -8007
rect -1268 -8075 -1256 -8041
rect -1222 -8075 -1210 -8041
rect -1268 -8109 -1210 -8075
rect -1268 -8143 -1256 -8109
rect -1222 -8143 -1210 -8109
rect -1268 -8177 -1210 -8143
rect -1268 -8211 -1256 -8177
rect -1222 -8211 -1210 -8177
rect -1268 -8245 -1210 -8211
rect -1268 -8279 -1256 -8245
rect -1222 -8279 -1210 -8245
rect -1268 -8313 -1210 -8279
rect -1268 -8347 -1256 -8313
rect -1222 -8347 -1210 -8313
rect -1268 -8381 -1210 -8347
rect -1268 -8415 -1256 -8381
rect -1222 -8415 -1210 -8381
rect -1268 -8449 -1210 -8415
rect -1268 -8483 -1256 -8449
rect -1222 -8483 -1210 -8449
rect -1268 -8517 -1210 -8483
rect -1268 -8551 -1256 -8517
rect -1222 -8551 -1210 -8517
rect -1268 -8585 -1210 -8551
rect -1268 -8619 -1256 -8585
rect -1222 -8619 -1210 -8585
rect -1268 -8653 -1210 -8619
rect -1268 -8687 -1256 -8653
rect -1222 -8687 -1210 -8653
rect -1268 -8721 -1210 -8687
rect -1268 -8755 -1256 -8721
rect -1222 -8755 -1210 -8721
rect -1268 -8789 -1210 -8755
rect -1268 -8823 -1256 -8789
rect -1222 -8823 -1210 -8789
rect -1268 -8857 -1210 -8823
rect -1268 -8891 -1256 -8857
rect -1222 -8891 -1210 -8857
rect -1268 -8925 -1210 -8891
rect -1268 -8959 -1256 -8925
rect -1222 -8959 -1210 -8925
rect -1268 -8993 -1210 -8959
rect -1268 -9027 -1256 -8993
rect -1222 -9027 -1210 -8993
rect -1268 -9061 -1210 -9027
rect -1268 -9095 -1256 -9061
rect -1222 -9095 -1210 -9061
rect -1268 -9129 -1210 -9095
rect -1268 -9163 -1256 -9129
rect -1222 -9163 -1210 -9129
rect -1268 -9197 -1210 -9163
rect -1268 -9231 -1256 -9197
rect -1222 -9231 -1210 -9197
rect -1268 -9265 -1210 -9231
rect -1268 -9299 -1256 -9265
rect -1222 -9299 -1210 -9265
rect -1268 -9333 -1210 -9299
rect -1268 -9367 -1256 -9333
rect -1222 -9367 -1210 -9333
rect -1268 -9401 -1210 -9367
rect -1268 -9435 -1256 -9401
rect -1222 -9435 -1210 -9401
rect -1268 -9469 -1210 -9435
rect -1268 -9503 -1256 -9469
rect -1222 -9503 -1210 -9469
rect -1268 -9537 -1210 -9503
rect -1268 -9571 -1256 -9537
rect -1222 -9571 -1210 -9537
rect -1268 -9600 -1210 -9571
rect -1150 9571 -1092 9600
rect -1150 9537 -1138 9571
rect -1104 9537 -1092 9571
rect -1150 9503 -1092 9537
rect -1150 9469 -1138 9503
rect -1104 9469 -1092 9503
rect -1150 9435 -1092 9469
rect -1150 9401 -1138 9435
rect -1104 9401 -1092 9435
rect -1150 9367 -1092 9401
rect -1150 9333 -1138 9367
rect -1104 9333 -1092 9367
rect -1150 9299 -1092 9333
rect -1150 9265 -1138 9299
rect -1104 9265 -1092 9299
rect -1150 9231 -1092 9265
rect -1150 9197 -1138 9231
rect -1104 9197 -1092 9231
rect -1150 9163 -1092 9197
rect -1150 9129 -1138 9163
rect -1104 9129 -1092 9163
rect -1150 9095 -1092 9129
rect -1150 9061 -1138 9095
rect -1104 9061 -1092 9095
rect -1150 9027 -1092 9061
rect -1150 8993 -1138 9027
rect -1104 8993 -1092 9027
rect -1150 8959 -1092 8993
rect -1150 8925 -1138 8959
rect -1104 8925 -1092 8959
rect -1150 8891 -1092 8925
rect -1150 8857 -1138 8891
rect -1104 8857 -1092 8891
rect -1150 8823 -1092 8857
rect -1150 8789 -1138 8823
rect -1104 8789 -1092 8823
rect -1150 8755 -1092 8789
rect -1150 8721 -1138 8755
rect -1104 8721 -1092 8755
rect -1150 8687 -1092 8721
rect -1150 8653 -1138 8687
rect -1104 8653 -1092 8687
rect -1150 8619 -1092 8653
rect -1150 8585 -1138 8619
rect -1104 8585 -1092 8619
rect -1150 8551 -1092 8585
rect -1150 8517 -1138 8551
rect -1104 8517 -1092 8551
rect -1150 8483 -1092 8517
rect -1150 8449 -1138 8483
rect -1104 8449 -1092 8483
rect -1150 8415 -1092 8449
rect -1150 8381 -1138 8415
rect -1104 8381 -1092 8415
rect -1150 8347 -1092 8381
rect -1150 8313 -1138 8347
rect -1104 8313 -1092 8347
rect -1150 8279 -1092 8313
rect -1150 8245 -1138 8279
rect -1104 8245 -1092 8279
rect -1150 8211 -1092 8245
rect -1150 8177 -1138 8211
rect -1104 8177 -1092 8211
rect -1150 8143 -1092 8177
rect -1150 8109 -1138 8143
rect -1104 8109 -1092 8143
rect -1150 8075 -1092 8109
rect -1150 8041 -1138 8075
rect -1104 8041 -1092 8075
rect -1150 8007 -1092 8041
rect -1150 7973 -1138 8007
rect -1104 7973 -1092 8007
rect -1150 7939 -1092 7973
rect -1150 7905 -1138 7939
rect -1104 7905 -1092 7939
rect -1150 7871 -1092 7905
rect -1150 7837 -1138 7871
rect -1104 7837 -1092 7871
rect -1150 7803 -1092 7837
rect -1150 7769 -1138 7803
rect -1104 7769 -1092 7803
rect -1150 7735 -1092 7769
rect -1150 7701 -1138 7735
rect -1104 7701 -1092 7735
rect -1150 7667 -1092 7701
rect -1150 7633 -1138 7667
rect -1104 7633 -1092 7667
rect -1150 7599 -1092 7633
rect -1150 7565 -1138 7599
rect -1104 7565 -1092 7599
rect -1150 7531 -1092 7565
rect -1150 7497 -1138 7531
rect -1104 7497 -1092 7531
rect -1150 7463 -1092 7497
rect -1150 7429 -1138 7463
rect -1104 7429 -1092 7463
rect -1150 7395 -1092 7429
rect -1150 7361 -1138 7395
rect -1104 7361 -1092 7395
rect -1150 7327 -1092 7361
rect -1150 7293 -1138 7327
rect -1104 7293 -1092 7327
rect -1150 7259 -1092 7293
rect -1150 7225 -1138 7259
rect -1104 7225 -1092 7259
rect -1150 7191 -1092 7225
rect -1150 7157 -1138 7191
rect -1104 7157 -1092 7191
rect -1150 7123 -1092 7157
rect -1150 7089 -1138 7123
rect -1104 7089 -1092 7123
rect -1150 7055 -1092 7089
rect -1150 7021 -1138 7055
rect -1104 7021 -1092 7055
rect -1150 6987 -1092 7021
rect -1150 6953 -1138 6987
rect -1104 6953 -1092 6987
rect -1150 6919 -1092 6953
rect -1150 6885 -1138 6919
rect -1104 6885 -1092 6919
rect -1150 6851 -1092 6885
rect -1150 6817 -1138 6851
rect -1104 6817 -1092 6851
rect -1150 6783 -1092 6817
rect -1150 6749 -1138 6783
rect -1104 6749 -1092 6783
rect -1150 6715 -1092 6749
rect -1150 6681 -1138 6715
rect -1104 6681 -1092 6715
rect -1150 6647 -1092 6681
rect -1150 6613 -1138 6647
rect -1104 6613 -1092 6647
rect -1150 6579 -1092 6613
rect -1150 6545 -1138 6579
rect -1104 6545 -1092 6579
rect -1150 6511 -1092 6545
rect -1150 6477 -1138 6511
rect -1104 6477 -1092 6511
rect -1150 6443 -1092 6477
rect -1150 6409 -1138 6443
rect -1104 6409 -1092 6443
rect -1150 6375 -1092 6409
rect -1150 6341 -1138 6375
rect -1104 6341 -1092 6375
rect -1150 6307 -1092 6341
rect -1150 6273 -1138 6307
rect -1104 6273 -1092 6307
rect -1150 6239 -1092 6273
rect -1150 6205 -1138 6239
rect -1104 6205 -1092 6239
rect -1150 6171 -1092 6205
rect -1150 6137 -1138 6171
rect -1104 6137 -1092 6171
rect -1150 6103 -1092 6137
rect -1150 6069 -1138 6103
rect -1104 6069 -1092 6103
rect -1150 6035 -1092 6069
rect -1150 6001 -1138 6035
rect -1104 6001 -1092 6035
rect -1150 5967 -1092 6001
rect -1150 5933 -1138 5967
rect -1104 5933 -1092 5967
rect -1150 5899 -1092 5933
rect -1150 5865 -1138 5899
rect -1104 5865 -1092 5899
rect -1150 5831 -1092 5865
rect -1150 5797 -1138 5831
rect -1104 5797 -1092 5831
rect -1150 5763 -1092 5797
rect -1150 5729 -1138 5763
rect -1104 5729 -1092 5763
rect -1150 5695 -1092 5729
rect -1150 5661 -1138 5695
rect -1104 5661 -1092 5695
rect -1150 5627 -1092 5661
rect -1150 5593 -1138 5627
rect -1104 5593 -1092 5627
rect -1150 5559 -1092 5593
rect -1150 5525 -1138 5559
rect -1104 5525 -1092 5559
rect -1150 5491 -1092 5525
rect -1150 5457 -1138 5491
rect -1104 5457 -1092 5491
rect -1150 5423 -1092 5457
rect -1150 5389 -1138 5423
rect -1104 5389 -1092 5423
rect -1150 5355 -1092 5389
rect -1150 5321 -1138 5355
rect -1104 5321 -1092 5355
rect -1150 5287 -1092 5321
rect -1150 5253 -1138 5287
rect -1104 5253 -1092 5287
rect -1150 5219 -1092 5253
rect -1150 5185 -1138 5219
rect -1104 5185 -1092 5219
rect -1150 5151 -1092 5185
rect -1150 5117 -1138 5151
rect -1104 5117 -1092 5151
rect -1150 5083 -1092 5117
rect -1150 5049 -1138 5083
rect -1104 5049 -1092 5083
rect -1150 5015 -1092 5049
rect -1150 4981 -1138 5015
rect -1104 4981 -1092 5015
rect -1150 4947 -1092 4981
rect -1150 4913 -1138 4947
rect -1104 4913 -1092 4947
rect -1150 4879 -1092 4913
rect -1150 4845 -1138 4879
rect -1104 4845 -1092 4879
rect -1150 4811 -1092 4845
rect -1150 4777 -1138 4811
rect -1104 4777 -1092 4811
rect -1150 4743 -1092 4777
rect -1150 4709 -1138 4743
rect -1104 4709 -1092 4743
rect -1150 4675 -1092 4709
rect -1150 4641 -1138 4675
rect -1104 4641 -1092 4675
rect -1150 4607 -1092 4641
rect -1150 4573 -1138 4607
rect -1104 4573 -1092 4607
rect -1150 4539 -1092 4573
rect -1150 4505 -1138 4539
rect -1104 4505 -1092 4539
rect -1150 4471 -1092 4505
rect -1150 4437 -1138 4471
rect -1104 4437 -1092 4471
rect -1150 4403 -1092 4437
rect -1150 4369 -1138 4403
rect -1104 4369 -1092 4403
rect -1150 4335 -1092 4369
rect -1150 4301 -1138 4335
rect -1104 4301 -1092 4335
rect -1150 4267 -1092 4301
rect -1150 4233 -1138 4267
rect -1104 4233 -1092 4267
rect -1150 4199 -1092 4233
rect -1150 4165 -1138 4199
rect -1104 4165 -1092 4199
rect -1150 4131 -1092 4165
rect -1150 4097 -1138 4131
rect -1104 4097 -1092 4131
rect -1150 4063 -1092 4097
rect -1150 4029 -1138 4063
rect -1104 4029 -1092 4063
rect -1150 3995 -1092 4029
rect -1150 3961 -1138 3995
rect -1104 3961 -1092 3995
rect -1150 3927 -1092 3961
rect -1150 3893 -1138 3927
rect -1104 3893 -1092 3927
rect -1150 3859 -1092 3893
rect -1150 3825 -1138 3859
rect -1104 3825 -1092 3859
rect -1150 3791 -1092 3825
rect -1150 3757 -1138 3791
rect -1104 3757 -1092 3791
rect -1150 3723 -1092 3757
rect -1150 3689 -1138 3723
rect -1104 3689 -1092 3723
rect -1150 3655 -1092 3689
rect -1150 3621 -1138 3655
rect -1104 3621 -1092 3655
rect -1150 3587 -1092 3621
rect -1150 3553 -1138 3587
rect -1104 3553 -1092 3587
rect -1150 3519 -1092 3553
rect -1150 3485 -1138 3519
rect -1104 3485 -1092 3519
rect -1150 3451 -1092 3485
rect -1150 3417 -1138 3451
rect -1104 3417 -1092 3451
rect -1150 3383 -1092 3417
rect -1150 3349 -1138 3383
rect -1104 3349 -1092 3383
rect -1150 3315 -1092 3349
rect -1150 3281 -1138 3315
rect -1104 3281 -1092 3315
rect -1150 3247 -1092 3281
rect -1150 3213 -1138 3247
rect -1104 3213 -1092 3247
rect -1150 3179 -1092 3213
rect -1150 3145 -1138 3179
rect -1104 3145 -1092 3179
rect -1150 3111 -1092 3145
rect -1150 3077 -1138 3111
rect -1104 3077 -1092 3111
rect -1150 3043 -1092 3077
rect -1150 3009 -1138 3043
rect -1104 3009 -1092 3043
rect -1150 2975 -1092 3009
rect -1150 2941 -1138 2975
rect -1104 2941 -1092 2975
rect -1150 2907 -1092 2941
rect -1150 2873 -1138 2907
rect -1104 2873 -1092 2907
rect -1150 2839 -1092 2873
rect -1150 2805 -1138 2839
rect -1104 2805 -1092 2839
rect -1150 2771 -1092 2805
rect -1150 2737 -1138 2771
rect -1104 2737 -1092 2771
rect -1150 2703 -1092 2737
rect -1150 2669 -1138 2703
rect -1104 2669 -1092 2703
rect -1150 2635 -1092 2669
rect -1150 2601 -1138 2635
rect -1104 2601 -1092 2635
rect -1150 2567 -1092 2601
rect -1150 2533 -1138 2567
rect -1104 2533 -1092 2567
rect -1150 2499 -1092 2533
rect -1150 2465 -1138 2499
rect -1104 2465 -1092 2499
rect -1150 2431 -1092 2465
rect -1150 2397 -1138 2431
rect -1104 2397 -1092 2431
rect -1150 2363 -1092 2397
rect -1150 2329 -1138 2363
rect -1104 2329 -1092 2363
rect -1150 2295 -1092 2329
rect -1150 2261 -1138 2295
rect -1104 2261 -1092 2295
rect -1150 2227 -1092 2261
rect -1150 2193 -1138 2227
rect -1104 2193 -1092 2227
rect -1150 2159 -1092 2193
rect -1150 2125 -1138 2159
rect -1104 2125 -1092 2159
rect -1150 2091 -1092 2125
rect -1150 2057 -1138 2091
rect -1104 2057 -1092 2091
rect -1150 2023 -1092 2057
rect -1150 1989 -1138 2023
rect -1104 1989 -1092 2023
rect -1150 1955 -1092 1989
rect -1150 1921 -1138 1955
rect -1104 1921 -1092 1955
rect -1150 1887 -1092 1921
rect -1150 1853 -1138 1887
rect -1104 1853 -1092 1887
rect -1150 1819 -1092 1853
rect -1150 1785 -1138 1819
rect -1104 1785 -1092 1819
rect -1150 1751 -1092 1785
rect -1150 1717 -1138 1751
rect -1104 1717 -1092 1751
rect -1150 1683 -1092 1717
rect -1150 1649 -1138 1683
rect -1104 1649 -1092 1683
rect -1150 1615 -1092 1649
rect -1150 1581 -1138 1615
rect -1104 1581 -1092 1615
rect -1150 1547 -1092 1581
rect -1150 1513 -1138 1547
rect -1104 1513 -1092 1547
rect -1150 1479 -1092 1513
rect -1150 1445 -1138 1479
rect -1104 1445 -1092 1479
rect -1150 1411 -1092 1445
rect -1150 1377 -1138 1411
rect -1104 1377 -1092 1411
rect -1150 1343 -1092 1377
rect -1150 1309 -1138 1343
rect -1104 1309 -1092 1343
rect -1150 1275 -1092 1309
rect -1150 1241 -1138 1275
rect -1104 1241 -1092 1275
rect -1150 1207 -1092 1241
rect -1150 1173 -1138 1207
rect -1104 1173 -1092 1207
rect -1150 1139 -1092 1173
rect -1150 1105 -1138 1139
rect -1104 1105 -1092 1139
rect -1150 1071 -1092 1105
rect -1150 1037 -1138 1071
rect -1104 1037 -1092 1071
rect -1150 1003 -1092 1037
rect -1150 969 -1138 1003
rect -1104 969 -1092 1003
rect -1150 935 -1092 969
rect -1150 901 -1138 935
rect -1104 901 -1092 935
rect -1150 867 -1092 901
rect -1150 833 -1138 867
rect -1104 833 -1092 867
rect -1150 799 -1092 833
rect -1150 765 -1138 799
rect -1104 765 -1092 799
rect -1150 731 -1092 765
rect -1150 697 -1138 731
rect -1104 697 -1092 731
rect -1150 663 -1092 697
rect -1150 629 -1138 663
rect -1104 629 -1092 663
rect -1150 595 -1092 629
rect -1150 561 -1138 595
rect -1104 561 -1092 595
rect -1150 527 -1092 561
rect -1150 493 -1138 527
rect -1104 493 -1092 527
rect -1150 459 -1092 493
rect -1150 425 -1138 459
rect -1104 425 -1092 459
rect -1150 391 -1092 425
rect -1150 357 -1138 391
rect -1104 357 -1092 391
rect -1150 323 -1092 357
rect -1150 289 -1138 323
rect -1104 289 -1092 323
rect -1150 255 -1092 289
rect -1150 221 -1138 255
rect -1104 221 -1092 255
rect -1150 187 -1092 221
rect -1150 153 -1138 187
rect -1104 153 -1092 187
rect -1150 119 -1092 153
rect -1150 85 -1138 119
rect -1104 85 -1092 119
rect -1150 51 -1092 85
rect -1150 17 -1138 51
rect -1104 17 -1092 51
rect -1150 -17 -1092 17
rect -1150 -51 -1138 -17
rect -1104 -51 -1092 -17
rect -1150 -85 -1092 -51
rect -1150 -119 -1138 -85
rect -1104 -119 -1092 -85
rect -1150 -153 -1092 -119
rect -1150 -187 -1138 -153
rect -1104 -187 -1092 -153
rect -1150 -221 -1092 -187
rect -1150 -255 -1138 -221
rect -1104 -255 -1092 -221
rect -1150 -289 -1092 -255
rect -1150 -323 -1138 -289
rect -1104 -323 -1092 -289
rect -1150 -357 -1092 -323
rect -1150 -391 -1138 -357
rect -1104 -391 -1092 -357
rect -1150 -425 -1092 -391
rect -1150 -459 -1138 -425
rect -1104 -459 -1092 -425
rect -1150 -493 -1092 -459
rect -1150 -527 -1138 -493
rect -1104 -527 -1092 -493
rect -1150 -561 -1092 -527
rect -1150 -595 -1138 -561
rect -1104 -595 -1092 -561
rect -1150 -629 -1092 -595
rect -1150 -663 -1138 -629
rect -1104 -663 -1092 -629
rect -1150 -697 -1092 -663
rect -1150 -731 -1138 -697
rect -1104 -731 -1092 -697
rect -1150 -765 -1092 -731
rect -1150 -799 -1138 -765
rect -1104 -799 -1092 -765
rect -1150 -833 -1092 -799
rect -1150 -867 -1138 -833
rect -1104 -867 -1092 -833
rect -1150 -901 -1092 -867
rect -1150 -935 -1138 -901
rect -1104 -935 -1092 -901
rect -1150 -969 -1092 -935
rect -1150 -1003 -1138 -969
rect -1104 -1003 -1092 -969
rect -1150 -1037 -1092 -1003
rect -1150 -1071 -1138 -1037
rect -1104 -1071 -1092 -1037
rect -1150 -1105 -1092 -1071
rect -1150 -1139 -1138 -1105
rect -1104 -1139 -1092 -1105
rect -1150 -1173 -1092 -1139
rect -1150 -1207 -1138 -1173
rect -1104 -1207 -1092 -1173
rect -1150 -1241 -1092 -1207
rect -1150 -1275 -1138 -1241
rect -1104 -1275 -1092 -1241
rect -1150 -1309 -1092 -1275
rect -1150 -1343 -1138 -1309
rect -1104 -1343 -1092 -1309
rect -1150 -1377 -1092 -1343
rect -1150 -1411 -1138 -1377
rect -1104 -1411 -1092 -1377
rect -1150 -1445 -1092 -1411
rect -1150 -1479 -1138 -1445
rect -1104 -1479 -1092 -1445
rect -1150 -1513 -1092 -1479
rect -1150 -1547 -1138 -1513
rect -1104 -1547 -1092 -1513
rect -1150 -1581 -1092 -1547
rect -1150 -1615 -1138 -1581
rect -1104 -1615 -1092 -1581
rect -1150 -1649 -1092 -1615
rect -1150 -1683 -1138 -1649
rect -1104 -1683 -1092 -1649
rect -1150 -1717 -1092 -1683
rect -1150 -1751 -1138 -1717
rect -1104 -1751 -1092 -1717
rect -1150 -1785 -1092 -1751
rect -1150 -1819 -1138 -1785
rect -1104 -1819 -1092 -1785
rect -1150 -1853 -1092 -1819
rect -1150 -1887 -1138 -1853
rect -1104 -1887 -1092 -1853
rect -1150 -1921 -1092 -1887
rect -1150 -1955 -1138 -1921
rect -1104 -1955 -1092 -1921
rect -1150 -1989 -1092 -1955
rect -1150 -2023 -1138 -1989
rect -1104 -2023 -1092 -1989
rect -1150 -2057 -1092 -2023
rect -1150 -2091 -1138 -2057
rect -1104 -2091 -1092 -2057
rect -1150 -2125 -1092 -2091
rect -1150 -2159 -1138 -2125
rect -1104 -2159 -1092 -2125
rect -1150 -2193 -1092 -2159
rect -1150 -2227 -1138 -2193
rect -1104 -2227 -1092 -2193
rect -1150 -2261 -1092 -2227
rect -1150 -2295 -1138 -2261
rect -1104 -2295 -1092 -2261
rect -1150 -2329 -1092 -2295
rect -1150 -2363 -1138 -2329
rect -1104 -2363 -1092 -2329
rect -1150 -2397 -1092 -2363
rect -1150 -2431 -1138 -2397
rect -1104 -2431 -1092 -2397
rect -1150 -2465 -1092 -2431
rect -1150 -2499 -1138 -2465
rect -1104 -2499 -1092 -2465
rect -1150 -2533 -1092 -2499
rect -1150 -2567 -1138 -2533
rect -1104 -2567 -1092 -2533
rect -1150 -2601 -1092 -2567
rect -1150 -2635 -1138 -2601
rect -1104 -2635 -1092 -2601
rect -1150 -2669 -1092 -2635
rect -1150 -2703 -1138 -2669
rect -1104 -2703 -1092 -2669
rect -1150 -2737 -1092 -2703
rect -1150 -2771 -1138 -2737
rect -1104 -2771 -1092 -2737
rect -1150 -2805 -1092 -2771
rect -1150 -2839 -1138 -2805
rect -1104 -2839 -1092 -2805
rect -1150 -2873 -1092 -2839
rect -1150 -2907 -1138 -2873
rect -1104 -2907 -1092 -2873
rect -1150 -2941 -1092 -2907
rect -1150 -2975 -1138 -2941
rect -1104 -2975 -1092 -2941
rect -1150 -3009 -1092 -2975
rect -1150 -3043 -1138 -3009
rect -1104 -3043 -1092 -3009
rect -1150 -3077 -1092 -3043
rect -1150 -3111 -1138 -3077
rect -1104 -3111 -1092 -3077
rect -1150 -3145 -1092 -3111
rect -1150 -3179 -1138 -3145
rect -1104 -3179 -1092 -3145
rect -1150 -3213 -1092 -3179
rect -1150 -3247 -1138 -3213
rect -1104 -3247 -1092 -3213
rect -1150 -3281 -1092 -3247
rect -1150 -3315 -1138 -3281
rect -1104 -3315 -1092 -3281
rect -1150 -3349 -1092 -3315
rect -1150 -3383 -1138 -3349
rect -1104 -3383 -1092 -3349
rect -1150 -3417 -1092 -3383
rect -1150 -3451 -1138 -3417
rect -1104 -3451 -1092 -3417
rect -1150 -3485 -1092 -3451
rect -1150 -3519 -1138 -3485
rect -1104 -3519 -1092 -3485
rect -1150 -3553 -1092 -3519
rect -1150 -3587 -1138 -3553
rect -1104 -3587 -1092 -3553
rect -1150 -3621 -1092 -3587
rect -1150 -3655 -1138 -3621
rect -1104 -3655 -1092 -3621
rect -1150 -3689 -1092 -3655
rect -1150 -3723 -1138 -3689
rect -1104 -3723 -1092 -3689
rect -1150 -3757 -1092 -3723
rect -1150 -3791 -1138 -3757
rect -1104 -3791 -1092 -3757
rect -1150 -3825 -1092 -3791
rect -1150 -3859 -1138 -3825
rect -1104 -3859 -1092 -3825
rect -1150 -3893 -1092 -3859
rect -1150 -3927 -1138 -3893
rect -1104 -3927 -1092 -3893
rect -1150 -3961 -1092 -3927
rect -1150 -3995 -1138 -3961
rect -1104 -3995 -1092 -3961
rect -1150 -4029 -1092 -3995
rect -1150 -4063 -1138 -4029
rect -1104 -4063 -1092 -4029
rect -1150 -4097 -1092 -4063
rect -1150 -4131 -1138 -4097
rect -1104 -4131 -1092 -4097
rect -1150 -4165 -1092 -4131
rect -1150 -4199 -1138 -4165
rect -1104 -4199 -1092 -4165
rect -1150 -4233 -1092 -4199
rect -1150 -4267 -1138 -4233
rect -1104 -4267 -1092 -4233
rect -1150 -4301 -1092 -4267
rect -1150 -4335 -1138 -4301
rect -1104 -4335 -1092 -4301
rect -1150 -4369 -1092 -4335
rect -1150 -4403 -1138 -4369
rect -1104 -4403 -1092 -4369
rect -1150 -4437 -1092 -4403
rect -1150 -4471 -1138 -4437
rect -1104 -4471 -1092 -4437
rect -1150 -4505 -1092 -4471
rect -1150 -4539 -1138 -4505
rect -1104 -4539 -1092 -4505
rect -1150 -4573 -1092 -4539
rect -1150 -4607 -1138 -4573
rect -1104 -4607 -1092 -4573
rect -1150 -4641 -1092 -4607
rect -1150 -4675 -1138 -4641
rect -1104 -4675 -1092 -4641
rect -1150 -4709 -1092 -4675
rect -1150 -4743 -1138 -4709
rect -1104 -4743 -1092 -4709
rect -1150 -4777 -1092 -4743
rect -1150 -4811 -1138 -4777
rect -1104 -4811 -1092 -4777
rect -1150 -4845 -1092 -4811
rect -1150 -4879 -1138 -4845
rect -1104 -4879 -1092 -4845
rect -1150 -4913 -1092 -4879
rect -1150 -4947 -1138 -4913
rect -1104 -4947 -1092 -4913
rect -1150 -4981 -1092 -4947
rect -1150 -5015 -1138 -4981
rect -1104 -5015 -1092 -4981
rect -1150 -5049 -1092 -5015
rect -1150 -5083 -1138 -5049
rect -1104 -5083 -1092 -5049
rect -1150 -5117 -1092 -5083
rect -1150 -5151 -1138 -5117
rect -1104 -5151 -1092 -5117
rect -1150 -5185 -1092 -5151
rect -1150 -5219 -1138 -5185
rect -1104 -5219 -1092 -5185
rect -1150 -5253 -1092 -5219
rect -1150 -5287 -1138 -5253
rect -1104 -5287 -1092 -5253
rect -1150 -5321 -1092 -5287
rect -1150 -5355 -1138 -5321
rect -1104 -5355 -1092 -5321
rect -1150 -5389 -1092 -5355
rect -1150 -5423 -1138 -5389
rect -1104 -5423 -1092 -5389
rect -1150 -5457 -1092 -5423
rect -1150 -5491 -1138 -5457
rect -1104 -5491 -1092 -5457
rect -1150 -5525 -1092 -5491
rect -1150 -5559 -1138 -5525
rect -1104 -5559 -1092 -5525
rect -1150 -5593 -1092 -5559
rect -1150 -5627 -1138 -5593
rect -1104 -5627 -1092 -5593
rect -1150 -5661 -1092 -5627
rect -1150 -5695 -1138 -5661
rect -1104 -5695 -1092 -5661
rect -1150 -5729 -1092 -5695
rect -1150 -5763 -1138 -5729
rect -1104 -5763 -1092 -5729
rect -1150 -5797 -1092 -5763
rect -1150 -5831 -1138 -5797
rect -1104 -5831 -1092 -5797
rect -1150 -5865 -1092 -5831
rect -1150 -5899 -1138 -5865
rect -1104 -5899 -1092 -5865
rect -1150 -5933 -1092 -5899
rect -1150 -5967 -1138 -5933
rect -1104 -5967 -1092 -5933
rect -1150 -6001 -1092 -5967
rect -1150 -6035 -1138 -6001
rect -1104 -6035 -1092 -6001
rect -1150 -6069 -1092 -6035
rect -1150 -6103 -1138 -6069
rect -1104 -6103 -1092 -6069
rect -1150 -6137 -1092 -6103
rect -1150 -6171 -1138 -6137
rect -1104 -6171 -1092 -6137
rect -1150 -6205 -1092 -6171
rect -1150 -6239 -1138 -6205
rect -1104 -6239 -1092 -6205
rect -1150 -6273 -1092 -6239
rect -1150 -6307 -1138 -6273
rect -1104 -6307 -1092 -6273
rect -1150 -6341 -1092 -6307
rect -1150 -6375 -1138 -6341
rect -1104 -6375 -1092 -6341
rect -1150 -6409 -1092 -6375
rect -1150 -6443 -1138 -6409
rect -1104 -6443 -1092 -6409
rect -1150 -6477 -1092 -6443
rect -1150 -6511 -1138 -6477
rect -1104 -6511 -1092 -6477
rect -1150 -6545 -1092 -6511
rect -1150 -6579 -1138 -6545
rect -1104 -6579 -1092 -6545
rect -1150 -6613 -1092 -6579
rect -1150 -6647 -1138 -6613
rect -1104 -6647 -1092 -6613
rect -1150 -6681 -1092 -6647
rect -1150 -6715 -1138 -6681
rect -1104 -6715 -1092 -6681
rect -1150 -6749 -1092 -6715
rect -1150 -6783 -1138 -6749
rect -1104 -6783 -1092 -6749
rect -1150 -6817 -1092 -6783
rect -1150 -6851 -1138 -6817
rect -1104 -6851 -1092 -6817
rect -1150 -6885 -1092 -6851
rect -1150 -6919 -1138 -6885
rect -1104 -6919 -1092 -6885
rect -1150 -6953 -1092 -6919
rect -1150 -6987 -1138 -6953
rect -1104 -6987 -1092 -6953
rect -1150 -7021 -1092 -6987
rect -1150 -7055 -1138 -7021
rect -1104 -7055 -1092 -7021
rect -1150 -7089 -1092 -7055
rect -1150 -7123 -1138 -7089
rect -1104 -7123 -1092 -7089
rect -1150 -7157 -1092 -7123
rect -1150 -7191 -1138 -7157
rect -1104 -7191 -1092 -7157
rect -1150 -7225 -1092 -7191
rect -1150 -7259 -1138 -7225
rect -1104 -7259 -1092 -7225
rect -1150 -7293 -1092 -7259
rect -1150 -7327 -1138 -7293
rect -1104 -7327 -1092 -7293
rect -1150 -7361 -1092 -7327
rect -1150 -7395 -1138 -7361
rect -1104 -7395 -1092 -7361
rect -1150 -7429 -1092 -7395
rect -1150 -7463 -1138 -7429
rect -1104 -7463 -1092 -7429
rect -1150 -7497 -1092 -7463
rect -1150 -7531 -1138 -7497
rect -1104 -7531 -1092 -7497
rect -1150 -7565 -1092 -7531
rect -1150 -7599 -1138 -7565
rect -1104 -7599 -1092 -7565
rect -1150 -7633 -1092 -7599
rect -1150 -7667 -1138 -7633
rect -1104 -7667 -1092 -7633
rect -1150 -7701 -1092 -7667
rect -1150 -7735 -1138 -7701
rect -1104 -7735 -1092 -7701
rect -1150 -7769 -1092 -7735
rect -1150 -7803 -1138 -7769
rect -1104 -7803 -1092 -7769
rect -1150 -7837 -1092 -7803
rect -1150 -7871 -1138 -7837
rect -1104 -7871 -1092 -7837
rect -1150 -7905 -1092 -7871
rect -1150 -7939 -1138 -7905
rect -1104 -7939 -1092 -7905
rect -1150 -7973 -1092 -7939
rect -1150 -8007 -1138 -7973
rect -1104 -8007 -1092 -7973
rect -1150 -8041 -1092 -8007
rect -1150 -8075 -1138 -8041
rect -1104 -8075 -1092 -8041
rect -1150 -8109 -1092 -8075
rect -1150 -8143 -1138 -8109
rect -1104 -8143 -1092 -8109
rect -1150 -8177 -1092 -8143
rect -1150 -8211 -1138 -8177
rect -1104 -8211 -1092 -8177
rect -1150 -8245 -1092 -8211
rect -1150 -8279 -1138 -8245
rect -1104 -8279 -1092 -8245
rect -1150 -8313 -1092 -8279
rect -1150 -8347 -1138 -8313
rect -1104 -8347 -1092 -8313
rect -1150 -8381 -1092 -8347
rect -1150 -8415 -1138 -8381
rect -1104 -8415 -1092 -8381
rect -1150 -8449 -1092 -8415
rect -1150 -8483 -1138 -8449
rect -1104 -8483 -1092 -8449
rect -1150 -8517 -1092 -8483
rect -1150 -8551 -1138 -8517
rect -1104 -8551 -1092 -8517
rect -1150 -8585 -1092 -8551
rect -1150 -8619 -1138 -8585
rect -1104 -8619 -1092 -8585
rect -1150 -8653 -1092 -8619
rect -1150 -8687 -1138 -8653
rect -1104 -8687 -1092 -8653
rect -1150 -8721 -1092 -8687
rect -1150 -8755 -1138 -8721
rect -1104 -8755 -1092 -8721
rect -1150 -8789 -1092 -8755
rect -1150 -8823 -1138 -8789
rect -1104 -8823 -1092 -8789
rect -1150 -8857 -1092 -8823
rect -1150 -8891 -1138 -8857
rect -1104 -8891 -1092 -8857
rect -1150 -8925 -1092 -8891
rect -1150 -8959 -1138 -8925
rect -1104 -8959 -1092 -8925
rect -1150 -8993 -1092 -8959
rect -1150 -9027 -1138 -8993
rect -1104 -9027 -1092 -8993
rect -1150 -9061 -1092 -9027
rect -1150 -9095 -1138 -9061
rect -1104 -9095 -1092 -9061
rect -1150 -9129 -1092 -9095
rect -1150 -9163 -1138 -9129
rect -1104 -9163 -1092 -9129
rect -1150 -9197 -1092 -9163
rect -1150 -9231 -1138 -9197
rect -1104 -9231 -1092 -9197
rect -1150 -9265 -1092 -9231
rect -1150 -9299 -1138 -9265
rect -1104 -9299 -1092 -9265
rect -1150 -9333 -1092 -9299
rect -1150 -9367 -1138 -9333
rect -1104 -9367 -1092 -9333
rect -1150 -9401 -1092 -9367
rect -1150 -9435 -1138 -9401
rect -1104 -9435 -1092 -9401
rect -1150 -9469 -1092 -9435
rect -1150 -9503 -1138 -9469
rect -1104 -9503 -1092 -9469
rect -1150 -9537 -1092 -9503
rect -1150 -9571 -1138 -9537
rect -1104 -9571 -1092 -9537
rect -1150 -9600 -1092 -9571
rect -1032 9571 -974 9600
rect -1032 9537 -1020 9571
rect -986 9537 -974 9571
rect -1032 9503 -974 9537
rect -1032 9469 -1020 9503
rect -986 9469 -974 9503
rect -1032 9435 -974 9469
rect -1032 9401 -1020 9435
rect -986 9401 -974 9435
rect -1032 9367 -974 9401
rect -1032 9333 -1020 9367
rect -986 9333 -974 9367
rect -1032 9299 -974 9333
rect -1032 9265 -1020 9299
rect -986 9265 -974 9299
rect -1032 9231 -974 9265
rect -1032 9197 -1020 9231
rect -986 9197 -974 9231
rect -1032 9163 -974 9197
rect -1032 9129 -1020 9163
rect -986 9129 -974 9163
rect -1032 9095 -974 9129
rect -1032 9061 -1020 9095
rect -986 9061 -974 9095
rect -1032 9027 -974 9061
rect -1032 8993 -1020 9027
rect -986 8993 -974 9027
rect -1032 8959 -974 8993
rect -1032 8925 -1020 8959
rect -986 8925 -974 8959
rect -1032 8891 -974 8925
rect -1032 8857 -1020 8891
rect -986 8857 -974 8891
rect -1032 8823 -974 8857
rect -1032 8789 -1020 8823
rect -986 8789 -974 8823
rect -1032 8755 -974 8789
rect -1032 8721 -1020 8755
rect -986 8721 -974 8755
rect -1032 8687 -974 8721
rect -1032 8653 -1020 8687
rect -986 8653 -974 8687
rect -1032 8619 -974 8653
rect -1032 8585 -1020 8619
rect -986 8585 -974 8619
rect -1032 8551 -974 8585
rect -1032 8517 -1020 8551
rect -986 8517 -974 8551
rect -1032 8483 -974 8517
rect -1032 8449 -1020 8483
rect -986 8449 -974 8483
rect -1032 8415 -974 8449
rect -1032 8381 -1020 8415
rect -986 8381 -974 8415
rect -1032 8347 -974 8381
rect -1032 8313 -1020 8347
rect -986 8313 -974 8347
rect -1032 8279 -974 8313
rect -1032 8245 -1020 8279
rect -986 8245 -974 8279
rect -1032 8211 -974 8245
rect -1032 8177 -1020 8211
rect -986 8177 -974 8211
rect -1032 8143 -974 8177
rect -1032 8109 -1020 8143
rect -986 8109 -974 8143
rect -1032 8075 -974 8109
rect -1032 8041 -1020 8075
rect -986 8041 -974 8075
rect -1032 8007 -974 8041
rect -1032 7973 -1020 8007
rect -986 7973 -974 8007
rect -1032 7939 -974 7973
rect -1032 7905 -1020 7939
rect -986 7905 -974 7939
rect -1032 7871 -974 7905
rect -1032 7837 -1020 7871
rect -986 7837 -974 7871
rect -1032 7803 -974 7837
rect -1032 7769 -1020 7803
rect -986 7769 -974 7803
rect -1032 7735 -974 7769
rect -1032 7701 -1020 7735
rect -986 7701 -974 7735
rect -1032 7667 -974 7701
rect -1032 7633 -1020 7667
rect -986 7633 -974 7667
rect -1032 7599 -974 7633
rect -1032 7565 -1020 7599
rect -986 7565 -974 7599
rect -1032 7531 -974 7565
rect -1032 7497 -1020 7531
rect -986 7497 -974 7531
rect -1032 7463 -974 7497
rect -1032 7429 -1020 7463
rect -986 7429 -974 7463
rect -1032 7395 -974 7429
rect -1032 7361 -1020 7395
rect -986 7361 -974 7395
rect -1032 7327 -974 7361
rect -1032 7293 -1020 7327
rect -986 7293 -974 7327
rect -1032 7259 -974 7293
rect -1032 7225 -1020 7259
rect -986 7225 -974 7259
rect -1032 7191 -974 7225
rect -1032 7157 -1020 7191
rect -986 7157 -974 7191
rect -1032 7123 -974 7157
rect -1032 7089 -1020 7123
rect -986 7089 -974 7123
rect -1032 7055 -974 7089
rect -1032 7021 -1020 7055
rect -986 7021 -974 7055
rect -1032 6987 -974 7021
rect -1032 6953 -1020 6987
rect -986 6953 -974 6987
rect -1032 6919 -974 6953
rect -1032 6885 -1020 6919
rect -986 6885 -974 6919
rect -1032 6851 -974 6885
rect -1032 6817 -1020 6851
rect -986 6817 -974 6851
rect -1032 6783 -974 6817
rect -1032 6749 -1020 6783
rect -986 6749 -974 6783
rect -1032 6715 -974 6749
rect -1032 6681 -1020 6715
rect -986 6681 -974 6715
rect -1032 6647 -974 6681
rect -1032 6613 -1020 6647
rect -986 6613 -974 6647
rect -1032 6579 -974 6613
rect -1032 6545 -1020 6579
rect -986 6545 -974 6579
rect -1032 6511 -974 6545
rect -1032 6477 -1020 6511
rect -986 6477 -974 6511
rect -1032 6443 -974 6477
rect -1032 6409 -1020 6443
rect -986 6409 -974 6443
rect -1032 6375 -974 6409
rect -1032 6341 -1020 6375
rect -986 6341 -974 6375
rect -1032 6307 -974 6341
rect -1032 6273 -1020 6307
rect -986 6273 -974 6307
rect -1032 6239 -974 6273
rect -1032 6205 -1020 6239
rect -986 6205 -974 6239
rect -1032 6171 -974 6205
rect -1032 6137 -1020 6171
rect -986 6137 -974 6171
rect -1032 6103 -974 6137
rect -1032 6069 -1020 6103
rect -986 6069 -974 6103
rect -1032 6035 -974 6069
rect -1032 6001 -1020 6035
rect -986 6001 -974 6035
rect -1032 5967 -974 6001
rect -1032 5933 -1020 5967
rect -986 5933 -974 5967
rect -1032 5899 -974 5933
rect -1032 5865 -1020 5899
rect -986 5865 -974 5899
rect -1032 5831 -974 5865
rect -1032 5797 -1020 5831
rect -986 5797 -974 5831
rect -1032 5763 -974 5797
rect -1032 5729 -1020 5763
rect -986 5729 -974 5763
rect -1032 5695 -974 5729
rect -1032 5661 -1020 5695
rect -986 5661 -974 5695
rect -1032 5627 -974 5661
rect -1032 5593 -1020 5627
rect -986 5593 -974 5627
rect -1032 5559 -974 5593
rect -1032 5525 -1020 5559
rect -986 5525 -974 5559
rect -1032 5491 -974 5525
rect -1032 5457 -1020 5491
rect -986 5457 -974 5491
rect -1032 5423 -974 5457
rect -1032 5389 -1020 5423
rect -986 5389 -974 5423
rect -1032 5355 -974 5389
rect -1032 5321 -1020 5355
rect -986 5321 -974 5355
rect -1032 5287 -974 5321
rect -1032 5253 -1020 5287
rect -986 5253 -974 5287
rect -1032 5219 -974 5253
rect -1032 5185 -1020 5219
rect -986 5185 -974 5219
rect -1032 5151 -974 5185
rect -1032 5117 -1020 5151
rect -986 5117 -974 5151
rect -1032 5083 -974 5117
rect -1032 5049 -1020 5083
rect -986 5049 -974 5083
rect -1032 5015 -974 5049
rect -1032 4981 -1020 5015
rect -986 4981 -974 5015
rect -1032 4947 -974 4981
rect -1032 4913 -1020 4947
rect -986 4913 -974 4947
rect -1032 4879 -974 4913
rect -1032 4845 -1020 4879
rect -986 4845 -974 4879
rect -1032 4811 -974 4845
rect -1032 4777 -1020 4811
rect -986 4777 -974 4811
rect -1032 4743 -974 4777
rect -1032 4709 -1020 4743
rect -986 4709 -974 4743
rect -1032 4675 -974 4709
rect -1032 4641 -1020 4675
rect -986 4641 -974 4675
rect -1032 4607 -974 4641
rect -1032 4573 -1020 4607
rect -986 4573 -974 4607
rect -1032 4539 -974 4573
rect -1032 4505 -1020 4539
rect -986 4505 -974 4539
rect -1032 4471 -974 4505
rect -1032 4437 -1020 4471
rect -986 4437 -974 4471
rect -1032 4403 -974 4437
rect -1032 4369 -1020 4403
rect -986 4369 -974 4403
rect -1032 4335 -974 4369
rect -1032 4301 -1020 4335
rect -986 4301 -974 4335
rect -1032 4267 -974 4301
rect -1032 4233 -1020 4267
rect -986 4233 -974 4267
rect -1032 4199 -974 4233
rect -1032 4165 -1020 4199
rect -986 4165 -974 4199
rect -1032 4131 -974 4165
rect -1032 4097 -1020 4131
rect -986 4097 -974 4131
rect -1032 4063 -974 4097
rect -1032 4029 -1020 4063
rect -986 4029 -974 4063
rect -1032 3995 -974 4029
rect -1032 3961 -1020 3995
rect -986 3961 -974 3995
rect -1032 3927 -974 3961
rect -1032 3893 -1020 3927
rect -986 3893 -974 3927
rect -1032 3859 -974 3893
rect -1032 3825 -1020 3859
rect -986 3825 -974 3859
rect -1032 3791 -974 3825
rect -1032 3757 -1020 3791
rect -986 3757 -974 3791
rect -1032 3723 -974 3757
rect -1032 3689 -1020 3723
rect -986 3689 -974 3723
rect -1032 3655 -974 3689
rect -1032 3621 -1020 3655
rect -986 3621 -974 3655
rect -1032 3587 -974 3621
rect -1032 3553 -1020 3587
rect -986 3553 -974 3587
rect -1032 3519 -974 3553
rect -1032 3485 -1020 3519
rect -986 3485 -974 3519
rect -1032 3451 -974 3485
rect -1032 3417 -1020 3451
rect -986 3417 -974 3451
rect -1032 3383 -974 3417
rect -1032 3349 -1020 3383
rect -986 3349 -974 3383
rect -1032 3315 -974 3349
rect -1032 3281 -1020 3315
rect -986 3281 -974 3315
rect -1032 3247 -974 3281
rect -1032 3213 -1020 3247
rect -986 3213 -974 3247
rect -1032 3179 -974 3213
rect -1032 3145 -1020 3179
rect -986 3145 -974 3179
rect -1032 3111 -974 3145
rect -1032 3077 -1020 3111
rect -986 3077 -974 3111
rect -1032 3043 -974 3077
rect -1032 3009 -1020 3043
rect -986 3009 -974 3043
rect -1032 2975 -974 3009
rect -1032 2941 -1020 2975
rect -986 2941 -974 2975
rect -1032 2907 -974 2941
rect -1032 2873 -1020 2907
rect -986 2873 -974 2907
rect -1032 2839 -974 2873
rect -1032 2805 -1020 2839
rect -986 2805 -974 2839
rect -1032 2771 -974 2805
rect -1032 2737 -1020 2771
rect -986 2737 -974 2771
rect -1032 2703 -974 2737
rect -1032 2669 -1020 2703
rect -986 2669 -974 2703
rect -1032 2635 -974 2669
rect -1032 2601 -1020 2635
rect -986 2601 -974 2635
rect -1032 2567 -974 2601
rect -1032 2533 -1020 2567
rect -986 2533 -974 2567
rect -1032 2499 -974 2533
rect -1032 2465 -1020 2499
rect -986 2465 -974 2499
rect -1032 2431 -974 2465
rect -1032 2397 -1020 2431
rect -986 2397 -974 2431
rect -1032 2363 -974 2397
rect -1032 2329 -1020 2363
rect -986 2329 -974 2363
rect -1032 2295 -974 2329
rect -1032 2261 -1020 2295
rect -986 2261 -974 2295
rect -1032 2227 -974 2261
rect -1032 2193 -1020 2227
rect -986 2193 -974 2227
rect -1032 2159 -974 2193
rect -1032 2125 -1020 2159
rect -986 2125 -974 2159
rect -1032 2091 -974 2125
rect -1032 2057 -1020 2091
rect -986 2057 -974 2091
rect -1032 2023 -974 2057
rect -1032 1989 -1020 2023
rect -986 1989 -974 2023
rect -1032 1955 -974 1989
rect -1032 1921 -1020 1955
rect -986 1921 -974 1955
rect -1032 1887 -974 1921
rect -1032 1853 -1020 1887
rect -986 1853 -974 1887
rect -1032 1819 -974 1853
rect -1032 1785 -1020 1819
rect -986 1785 -974 1819
rect -1032 1751 -974 1785
rect -1032 1717 -1020 1751
rect -986 1717 -974 1751
rect -1032 1683 -974 1717
rect -1032 1649 -1020 1683
rect -986 1649 -974 1683
rect -1032 1615 -974 1649
rect -1032 1581 -1020 1615
rect -986 1581 -974 1615
rect -1032 1547 -974 1581
rect -1032 1513 -1020 1547
rect -986 1513 -974 1547
rect -1032 1479 -974 1513
rect -1032 1445 -1020 1479
rect -986 1445 -974 1479
rect -1032 1411 -974 1445
rect -1032 1377 -1020 1411
rect -986 1377 -974 1411
rect -1032 1343 -974 1377
rect -1032 1309 -1020 1343
rect -986 1309 -974 1343
rect -1032 1275 -974 1309
rect -1032 1241 -1020 1275
rect -986 1241 -974 1275
rect -1032 1207 -974 1241
rect -1032 1173 -1020 1207
rect -986 1173 -974 1207
rect -1032 1139 -974 1173
rect -1032 1105 -1020 1139
rect -986 1105 -974 1139
rect -1032 1071 -974 1105
rect -1032 1037 -1020 1071
rect -986 1037 -974 1071
rect -1032 1003 -974 1037
rect -1032 969 -1020 1003
rect -986 969 -974 1003
rect -1032 935 -974 969
rect -1032 901 -1020 935
rect -986 901 -974 935
rect -1032 867 -974 901
rect -1032 833 -1020 867
rect -986 833 -974 867
rect -1032 799 -974 833
rect -1032 765 -1020 799
rect -986 765 -974 799
rect -1032 731 -974 765
rect -1032 697 -1020 731
rect -986 697 -974 731
rect -1032 663 -974 697
rect -1032 629 -1020 663
rect -986 629 -974 663
rect -1032 595 -974 629
rect -1032 561 -1020 595
rect -986 561 -974 595
rect -1032 527 -974 561
rect -1032 493 -1020 527
rect -986 493 -974 527
rect -1032 459 -974 493
rect -1032 425 -1020 459
rect -986 425 -974 459
rect -1032 391 -974 425
rect -1032 357 -1020 391
rect -986 357 -974 391
rect -1032 323 -974 357
rect -1032 289 -1020 323
rect -986 289 -974 323
rect -1032 255 -974 289
rect -1032 221 -1020 255
rect -986 221 -974 255
rect -1032 187 -974 221
rect -1032 153 -1020 187
rect -986 153 -974 187
rect -1032 119 -974 153
rect -1032 85 -1020 119
rect -986 85 -974 119
rect -1032 51 -974 85
rect -1032 17 -1020 51
rect -986 17 -974 51
rect -1032 -17 -974 17
rect -1032 -51 -1020 -17
rect -986 -51 -974 -17
rect -1032 -85 -974 -51
rect -1032 -119 -1020 -85
rect -986 -119 -974 -85
rect -1032 -153 -974 -119
rect -1032 -187 -1020 -153
rect -986 -187 -974 -153
rect -1032 -221 -974 -187
rect -1032 -255 -1020 -221
rect -986 -255 -974 -221
rect -1032 -289 -974 -255
rect -1032 -323 -1020 -289
rect -986 -323 -974 -289
rect -1032 -357 -974 -323
rect -1032 -391 -1020 -357
rect -986 -391 -974 -357
rect -1032 -425 -974 -391
rect -1032 -459 -1020 -425
rect -986 -459 -974 -425
rect -1032 -493 -974 -459
rect -1032 -527 -1020 -493
rect -986 -527 -974 -493
rect -1032 -561 -974 -527
rect -1032 -595 -1020 -561
rect -986 -595 -974 -561
rect -1032 -629 -974 -595
rect -1032 -663 -1020 -629
rect -986 -663 -974 -629
rect -1032 -697 -974 -663
rect -1032 -731 -1020 -697
rect -986 -731 -974 -697
rect -1032 -765 -974 -731
rect -1032 -799 -1020 -765
rect -986 -799 -974 -765
rect -1032 -833 -974 -799
rect -1032 -867 -1020 -833
rect -986 -867 -974 -833
rect -1032 -901 -974 -867
rect -1032 -935 -1020 -901
rect -986 -935 -974 -901
rect -1032 -969 -974 -935
rect -1032 -1003 -1020 -969
rect -986 -1003 -974 -969
rect -1032 -1037 -974 -1003
rect -1032 -1071 -1020 -1037
rect -986 -1071 -974 -1037
rect -1032 -1105 -974 -1071
rect -1032 -1139 -1020 -1105
rect -986 -1139 -974 -1105
rect -1032 -1173 -974 -1139
rect -1032 -1207 -1020 -1173
rect -986 -1207 -974 -1173
rect -1032 -1241 -974 -1207
rect -1032 -1275 -1020 -1241
rect -986 -1275 -974 -1241
rect -1032 -1309 -974 -1275
rect -1032 -1343 -1020 -1309
rect -986 -1343 -974 -1309
rect -1032 -1377 -974 -1343
rect -1032 -1411 -1020 -1377
rect -986 -1411 -974 -1377
rect -1032 -1445 -974 -1411
rect -1032 -1479 -1020 -1445
rect -986 -1479 -974 -1445
rect -1032 -1513 -974 -1479
rect -1032 -1547 -1020 -1513
rect -986 -1547 -974 -1513
rect -1032 -1581 -974 -1547
rect -1032 -1615 -1020 -1581
rect -986 -1615 -974 -1581
rect -1032 -1649 -974 -1615
rect -1032 -1683 -1020 -1649
rect -986 -1683 -974 -1649
rect -1032 -1717 -974 -1683
rect -1032 -1751 -1020 -1717
rect -986 -1751 -974 -1717
rect -1032 -1785 -974 -1751
rect -1032 -1819 -1020 -1785
rect -986 -1819 -974 -1785
rect -1032 -1853 -974 -1819
rect -1032 -1887 -1020 -1853
rect -986 -1887 -974 -1853
rect -1032 -1921 -974 -1887
rect -1032 -1955 -1020 -1921
rect -986 -1955 -974 -1921
rect -1032 -1989 -974 -1955
rect -1032 -2023 -1020 -1989
rect -986 -2023 -974 -1989
rect -1032 -2057 -974 -2023
rect -1032 -2091 -1020 -2057
rect -986 -2091 -974 -2057
rect -1032 -2125 -974 -2091
rect -1032 -2159 -1020 -2125
rect -986 -2159 -974 -2125
rect -1032 -2193 -974 -2159
rect -1032 -2227 -1020 -2193
rect -986 -2227 -974 -2193
rect -1032 -2261 -974 -2227
rect -1032 -2295 -1020 -2261
rect -986 -2295 -974 -2261
rect -1032 -2329 -974 -2295
rect -1032 -2363 -1020 -2329
rect -986 -2363 -974 -2329
rect -1032 -2397 -974 -2363
rect -1032 -2431 -1020 -2397
rect -986 -2431 -974 -2397
rect -1032 -2465 -974 -2431
rect -1032 -2499 -1020 -2465
rect -986 -2499 -974 -2465
rect -1032 -2533 -974 -2499
rect -1032 -2567 -1020 -2533
rect -986 -2567 -974 -2533
rect -1032 -2601 -974 -2567
rect -1032 -2635 -1020 -2601
rect -986 -2635 -974 -2601
rect -1032 -2669 -974 -2635
rect -1032 -2703 -1020 -2669
rect -986 -2703 -974 -2669
rect -1032 -2737 -974 -2703
rect -1032 -2771 -1020 -2737
rect -986 -2771 -974 -2737
rect -1032 -2805 -974 -2771
rect -1032 -2839 -1020 -2805
rect -986 -2839 -974 -2805
rect -1032 -2873 -974 -2839
rect -1032 -2907 -1020 -2873
rect -986 -2907 -974 -2873
rect -1032 -2941 -974 -2907
rect -1032 -2975 -1020 -2941
rect -986 -2975 -974 -2941
rect -1032 -3009 -974 -2975
rect -1032 -3043 -1020 -3009
rect -986 -3043 -974 -3009
rect -1032 -3077 -974 -3043
rect -1032 -3111 -1020 -3077
rect -986 -3111 -974 -3077
rect -1032 -3145 -974 -3111
rect -1032 -3179 -1020 -3145
rect -986 -3179 -974 -3145
rect -1032 -3213 -974 -3179
rect -1032 -3247 -1020 -3213
rect -986 -3247 -974 -3213
rect -1032 -3281 -974 -3247
rect -1032 -3315 -1020 -3281
rect -986 -3315 -974 -3281
rect -1032 -3349 -974 -3315
rect -1032 -3383 -1020 -3349
rect -986 -3383 -974 -3349
rect -1032 -3417 -974 -3383
rect -1032 -3451 -1020 -3417
rect -986 -3451 -974 -3417
rect -1032 -3485 -974 -3451
rect -1032 -3519 -1020 -3485
rect -986 -3519 -974 -3485
rect -1032 -3553 -974 -3519
rect -1032 -3587 -1020 -3553
rect -986 -3587 -974 -3553
rect -1032 -3621 -974 -3587
rect -1032 -3655 -1020 -3621
rect -986 -3655 -974 -3621
rect -1032 -3689 -974 -3655
rect -1032 -3723 -1020 -3689
rect -986 -3723 -974 -3689
rect -1032 -3757 -974 -3723
rect -1032 -3791 -1020 -3757
rect -986 -3791 -974 -3757
rect -1032 -3825 -974 -3791
rect -1032 -3859 -1020 -3825
rect -986 -3859 -974 -3825
rect -1032 -3893 -974 -3859
rect -1032 -3927 -1020 -3893
rect -986 -3927 -974 -3893
rect -1032 -3961 -974 -3927
rect -1032 -3995 -1020 -3961
rect -986 -3995 -974 -3961
rect -1032 -4029 -974 -3995
rect -1032 -4063 -1020 -4029
rect -986 -4063 -974 -4029
rect -1032 -4097 -974 -4063
rect -1032 -4131 -1020 -4097
rect -986 -4131 -974 -4097
rect -1032 -4165 -974 -4131
rect -1032 -4199 -1020 -4165
rect -986 -4199 -974 -4165
rect -1032 -4233 -974 -4199
rect -1032 -4267 -1020 -4233
rect -986 -4267 -974 -4233
rect -1032 -4301 -974 -4267
rect -1032 -4335 -1020 -4301
rect -986 -4335 -974 -4301
rect -1032 -4369 -974 -4335
rect -1032 -4403 -1020 -4369
rect -986 -4403 -974 -4369
rect -1032 -4437 -974 -4403
rect -1032 -4471 -1020 -4437
rect -986 -4471 -974 -4437
rect -1032 -4505 -974 -4471
rect -1032 -4539 -1020 -4505
rect -986 -4539 -974 -4505
rect -1032 -4573 -974 -4539
rect -1032 -4607 -1020 -4573
rect -986 -4607 -974 -4573
rect -1032 -4641 -974 -4607
rect -1032 -4675 -1020 -4641
rect -986 -4675 -974 -4641
rect -1032 -4709 -974 -4675
rect -1032 -4743 -1020 -4709
rect -986 -4743 -974 -4709
rect -1032 -4777 -974 -4743
rect -1032 -4811 -1020 -4777
rect -986 -4811 -974 -4777
rect -1032 -4845 -974 -4811
rect -1032 -4879 -1020 -4845
rect -986 -4879 -974 -4845
rect -1032 -4913 -974 -4879
rect -1032 -4947 -1020 -4913
rect -986 -4947 -974 -4913
rect -1032 -4981 -974 -4947
rect -1032 -5015 -1020 -4981
rect -986 -5015 -974 -4981
rect -1032 -5049 -974 -5015
rect -1032 -5083 -1020 -5049
rect -986 -5083 -974 -5049
rect -1032 -5117 -974 -5083
rect -1032 -5151 -1020 -5117
rect -986 -5151 -974 -5117
rect -1032 -5185 -974 -5151
rect -1032 -5219 -1020 -5185
rect -986 -5219 -974 -5185
rect -1032 -5253 -974 -5219
rect -1032 -5287 -1020 -5253
rect -986 -5287 -974 -5253
rect -1032 -5321 -974 -5287
rect -1032 -5355 -1020 -5321
rect -986 -5355 -974 -5321
rect -1032 -5389 -974 -5355
rect -1032 -5423 -1020 -5389
rect -986 -5423 -974 -5389
rect -1032 -5457 -974 -5423
rect -1032 -5491 -1020 -5457
rect -986 -5491 -974 -5457
rect -1032 -5525 -974 -5491
rect -1032 -5559 -1020 -5525
rect -986 -5559 -974 -5525
rect -1032 -5593 -974 -5559
rect -1032 -5627 -1020 -5593
rect -986 -5627 -974 -5593
rect -1032 -5661 -974 -5627
rect -1032 -5695 -1020 -5661
rect -986 -5695 -974 -5661
rect -1032 -5729 -974 -5695
rect -1032 -5763 -1020 -5729
rect -986 -5763 -974 -5729
rect -1032 -5797 -974 -5763
rect -1032 -5831 -1020 -5797
rect -986 -5831 -974 -5797
rect -1032 -5865 -974 -5831
rect -1032 -5899 -1020 -5865
rect -986 -5899 -974 -5865
rect -1032 -5933 -974 -5899
rect -1032 -5967 -1020 -5933
rect -986 -5967 -974 -5933
rect -1032 -6001 -974 -5967
rect -1032 -6035 -1020 -6001
rect -986 -6035 -974 -6001
rect -1032 -6069 -974 -6035
rect -1032 -6103 -1020 -6069
rect -986 -6103 -974 -6069
rect -1032 -6137 -974 -6103
rect -1032 -6171 -1020 -6137
rect -986 -6171 -974 -6137
rect -1032 -6205 -974 -6171
rect -1032 -6239 -1020 -6205
rect -986 -6239 -974 -6205
rect -1032 -6273 -974 -6239
rect -1032 -6307 -1020 -6273
rect -986 -6307 -974 -6273
rect -1032 -6341 -974 -6307
rect -1032 -6375 -1020 -6341
rect -986 -6375 -974 -6341
rect -1032 -6409 -974 -6375
rect -1032 -6443 -1020 -6409
rect -986 -6443 -974 -6409
rect -1032 -6477 -974 -6443
rect -1032 -6511 -1020 -6477
rect -986 -6511 -974 -6477
rect -1032 -6545 -974 -6511
rect -1032 -6579 -1020 -6545
rect -986 -6579 -974 -6545
rect -1032 -6613 -974 -6579
rect -1032 -6647 -1020 -6613
rect -986 -6647 -974 -6613
rect -1032 -6681 -974 -6647
rect -1032 -6715 -1020 -6681
rect -986 -6715 -974 -6681
rect -1032 -6749 -974 -6715
rect -1032 -6783 -1020 -6749
rect -986 -6783 -974 -6749
rect -1032 -6817 -974 -6783
rect -1032 -6851 -1020 -6817
rect -986 -6851 -974 -6817
rect -1032 -6885 -974 -6851
rect -1032 -6919 -1020 -6885
rect -986 -6919 -974 -6885
rect -1032 -6953 -974 -6919
rect -1032 -6987 -1020 -6953
rect -986 -6987 -974 -6953
rect -1032 -7021 -974 -6987
rect -1032 -7055 -1020 -7021
rect -986 -7055 -974 -7021
rect -1032 -7089 -974 -7055
rect -1032 -7123 -1020 -7089
rect -986 -7123 -974 -7089
rect -1032 -7157 -974 -7123
rect -1032 -7191 -1020 -7157
rect -986 -7191 -974 -7157
rect -1032 -7225 -974 -7191
rect -1032 -7259 -1020 -7225
rect -986 -7259 -974 -7225
rect -1032 -7293 -974 -7259
rect -1032 -7327 -1020 -7293
rect -986 -7327 -974 -7293
rect -1032 -7361 -974 -7327
rect -1032 -7395 -1020 -7361
rect -986 -7395 -974 -7361
rect -1032 -7429 -974 -7395
rect -1032 -7463 -1020 -7429
rect -986 -7463 -974 -7429
rect -1032 -7497 -974 -7463
rect -1032 -7531 -1020 -7497
rect -986 -7531 -974 -7497
rect -1032 -7565 -974 -7531
rect -1032 -7599 -1020 -7565
rect -986 -7599 -974 -7565
rect -1032 -7633 -974 -7599
rect -1032 -7667 -1020 -7633
rect -986 -7667 -974 -7633
rect -1032 -7701 -974 -7667
rect -1032 -7735 -1020 -7701
rect -986 -7735 -974 -7701
rect -1032 -7769 -974 -7735
rect -1032 -7803 -1020 -7769
rect -986 -7803 -974 -7769
rect -1032 -7837 -974 -7803
rect -1032 -7871 -1020 -7837
rect -986 -7871 -974 -7837
rect -1032 -7905 -974 -7871
rect -1032 -7939 -1020 -7905
rect -986 -7939 -974 -7905
rect -1032 -7973 -974 -7939
rect -1032 -8007 -1020 -7973
rect -986 -8007 -974 -7973
rect -1032 -8041 -974 -8007
rect -1032 -8075 -1020 -8041
rect -986 -8075 -974 -8041
rect -1032 -8109 -974 -8075
rect -1032 -8143 -1020 -8109
rect -986 -8143 -974 -8109
rect -1032 -8177 -974 -8143
rect -1032 -8211 -1020 -8177
rect -986 -8211 -974 -8177
rect -1032 -8245 -974 -8211
rect -1032 -8279 -1020 -8245
rect -986 -8279 -974 -8245
rect -1032 -8313 -974 -8279
rect -1032 -8347 -1020 -8313
rect -986 -8347 -974 -8313
rect -1032 -8381 -974 -8347
rect -1032 -8415 -1020 -8381
rect -986 -8415 -974 -8381
rect -1032 -8449 -974 -8415
rect -1032 -8483 -1020 -8449
rect -986 -8483 -974 -8449
rect -1032 -8517 -974 -8483
rect -1032 -8551 -1020 -8517
rect -986 -8551 -974 -8517
rect -1032 -8585 -974 -8551
rect -1032 -8619 -1020 -8585
rect -986 -8619 -974 -8585
rect -1032 -8653 -974 -8619
rect -1032 -8687 -1020 -8653
rect -986 -8687 -974 -8653
rect -1032 -8721 -974 -8687
rect -1032 -8755 -1020 -8721
rect -986 -8755 -974 -8721
rect -1032 -8789 -974 -8755
rect -1032 -8823 -1020 -8789
rect -986 -8823 -974 -8789
rect -1032 -8857 -974 -8823
rect -1032 -8891 -1020 -8857
rect -986 -8891 -974 -8857
rect -1032 -8925 -974 -8891
rect -1032 -8959 -1020 -8925
rect -986 -8959 -974 -8925
rect -1032 -8993 -974 -8959
rect -1032 -9027 -1020 -8993
rect -986 -9027 -974 -8993
rect -1032 -9061 -974 -9027
rect -1032 -9095 -1020 -9061
rect -986 -9095 -974 -9061
rect -1032 -9129 -974 -9095
rect -1032 -9163 -1020 -9129
rect -986 -9163 -974 -9129
rect -1032 -9197 -974 -9163
rect -1032 -9231 -1020 -9197
rect -986 -9231 -974 -9197
rect -1032 -9265 -974 -9231
rect -1032 -9299 -1020 -9265
rect -986 -9299 -974 -9265
rect -1032 -9333 -974 -9299
rect -1032 -9367 -1020 -9333
rect -986 -9367 -974 -9333
rect -1032 -9401 -974 -9367
rect -1032 -9435 -1020 -9401
rect -986 -9435 -974 -9401
rect -1032 -9469 -974 -9435
rect -1032 -9503 -1020 -9469
rect -986 -9503 -974 -9469
rect -1032 -9537 -974 -9503
rect -1032 -9571 -1020 -9537
rect -986 -9571 -974 -9537
rect -1032 -9600 -974 -9571
rect -914 9571 -856 9600
rect -914 9537 -902 9571
rect -868 9537 -856 9571
rect -914 9503 -856 9537
rect -914 9469 -902 9503
rect -868 9469 -856 9503
rect -914 9435 -856 9469
rect -914 9401 -902 9435
rect -868 9401 -856 9435
rect -914 9367 -856 9401
rect -914 9333 -902 9367
rect -868 9333 -856 9367
rect -914 9299 -856 9333
rect -914 9265 -902 9299
rect -868 9265 -856 9299
rect -914 9231 -856 9265
rect -914 9197 -902 9231
rect -868 9197 -856 9231
rect -914 9163 -856 9197
rect -914 9129 -902 9163
rect -868 9129 -856 9163
rect -914 9095 -856 9129
rect -914 9061 -902 9095
rect -868 9061 -856 9095
rect -914 9027 -856 9061
rect -914 8993 -902 9027
rect -868 8993 -856 9027
rect -914 8959 -856 8993
rect -914 8925 -902 8959
rect -868 8925 -856 8959
rect -914 8891 -856 8925
rect -914 8857 -902 8891
rect -868 8857 -856 8891
rect -914 8823 -856 8857
rect -914 8789 -902 8823
rect -868 8789 -856 8823
rect -914 8755 -856 8789
rect -914 8721 -902 8755
rect -868 8721 -856 8755
rect -914 8687 -856 8721
rect -914 8653 -902 8687
rect -868 8653 -856 8687
rect -914 8619 -856 8653
rect -914 8585 -902 8619
rect -868 8585 -856 8619
rect -914 8551 -856 8585
rect -914 8517 -902 8551
rect -868 8517 -856 8551
rect -914 8483 -856 8517
rect -914 8449 -902 8483
rect -868 8449 -856 8483
rect -914 8415 -856 8449
rect -914 8381 -902 8415
rect -868 8381 -856 8415
rect -914 8347 -856 8381
rect -914 8313 -902 8347
rect -868 8313 -856 8347
rect -914 8279 -856 8313
rect -914 8245 -902 8279
rect -868 8245 -856 8279
rect -914 8211 -856 8245
rect -914 8177 -902 8211
rect -868 8177 -856 8211
rect -914 8143 -856 8177
rect -914 8109 -902 8143
rect -868 8109 -856 8143
rect -914 8075 -856 8109
rect -914 8041 -902 8075
rect -868 8041 -856 8075
rect -914 8007 -856 8041
rect -914 7973 -902 8007
rect -868 7973 -856 8007
rect -914 7939 -856 7973
rect -914 7905 -902 7939
rect -868 7905 -856 7939
rect -914 7871 -856 7905
rect -914 7837 -902 7871
rect -868 7837 -856 7871
rect -914 7803 -856 7837
rect -914 7769 -902 7803
rect -868 7769 -856 7803
rect -914 7735 -856 7769
rect -914 7701 -902 7735
rect -868 7701 -856 7735
rect -914 7667 -856 7701
rect -914 7633 -902 7667
rect -868 7633 -856 7667
rect -914 7599 -856 7633
rect -914 7565 -902 7599
rect -868 7565 -856 7599
rect -914 7531 -856 7565
rect -914 7497 -902 7531
rect -868 7497 -856 7531
rect -914 7463 -856 7497
rect -914 7429 -902 7463
rect -868 7429 -856 7463
rect -914 7395 -856 7429
rect -914 7361 -902 7395
rect -868 7361 -856 7395
rect -914 7327 -856 7361
rect -914 7293 -902 7327
rect -868 7293 -856 7327
rect -914 7259 -856 7293
rect -914 7225 -902 7259
rect -868 7225 -856 7259
rect -914 7191 -856 7225
rect -914 7157 -902 7191
rect -868 7157 -856 7191
rect -914 7123 -856 7157
rect -914 7089 -902 7123
rect -868 7089 -856 7123
rect -914 7055 -856 7089
rect -914 7021 -902 7055
rect -868 7021 -856 7055
rect -914 6987 -856 7021
rect -914 6953 -902 6987
rect -868 6953 -856 6987
rect -914 6919 -856 6953
rect -914 6885 -902 6919
rect -868 6885 -856 6919
rect -914 6851 -856 6885
rect -914 6817 -902 6851
rect -868 6817 -856 6851
rect -914 6783 -856 6817
rect -914 6749 -902 6783
rect -868 6749 -856 6783
rect -914 6715 -856 6749
rect -914 6681 -902 6715
rect -868 6681 -856 6715
rect -914 6647 -856 6681
rect -914 6613 -902 6647
rect -868 6613 -856 6647
rect -914 6579 -856 6613
rect -914 6545 -902 6579
rect -868 6545 -856 6579
rect -914 6511 -856 6545
rect -914 6477 -902 6511
rect -868 6477 -856 6511
rect -914 6443 -856 6477
rect -914 6409 -902 6443
rect -868 6409 -856 6443
rect -914 6375 -856 6409
rect -914 6341 -902 6375
rect -868 6341 -856 6375
rect -914 6307 -856 6341
rect -914 6273 -902 6307
rect -868 6273 -856 6307
rect -914 6239 -856 6273
rect -914 6205 -902 6239
rect -868 6205 -856 6239
rect -914 6171 -856 6205
rect -914 6137 -902 6171
rect -868 6137 -856 6171
rect -914 6103 -856 6137
rect -914 6069 -902 6103
rect -868 6069 -856 6103
rect -914 6035 -856 6069
rect -914 6001 -902 6035
rect -868 6001 -856 6035
rect -914 5967 -856 6001
rect -914 5933 -902 5967
rect -868 5933 -856 5967
rect -914 5899 -856 5933
rect -914 5865 -902 5899
rect -868 5865 -856 5899
rect -914 5831 -856 5865
rect -914 5797 -902 5831
rect -868 5797 -856 5831
rect -914 5763 -856 5797
rect -914 5729 -902 5763
rect -868 5729 -856 5763
rect -914 5695 -856 5729
rect -914 5661 -902 5695
rect -868 5661 -856 5695
rect -914 5627 -856 5661
rect -914 5593 -902 5627
rect -868 5593 -856 5627
rect -914 5559 -856 5593
rect -914 5525 -902 5559
rect -868 5525 -856 5559
rect -914 5491 -856 5525
rect -914 5457 -902 5491
rect -868 5457 -856 5491
rect -914 5423 -856 5457
rect -914 5389 -902 5423
rect -868 5389 -856 5423
rect -914 5355 -856 5389
rect -914 5321 -902 5355
rect -868 5321 -856 5355
rect -914 5287 -856 5321
rect -914 5253 -902 5287
rect -868 5253 -856 5287
rect -914 5219 -856 5253
rect -914 5185 -902 5219
rect -868 5185 -856 5219
rect -914 5151 -856 5185
rect -914 5117 -902 5151
rect -868 5117 -856 5151
rect -914 5083 -856 5117
rect -914 5049 -902 5083
rect -868 5049 -856 5083
rect -914 5015 -856 5049
rect -914 4981 -902 5015
rect -868 4981 -856 5015
rect -914 4947 -856 4981
rect -914 4913 -902 4947
rect -868 4913 -856 4947
rect -914 4879 -856 4913
rect -914 4845 -902 4879
rect -868 4845 -856 4879
rect -914 4811 -856 4845
rect -914 4777 -902 4811
rect -868 4777 -856 4811
rect -914 4743 -856 4777
rect -914 4709 -902 4743
rect -868 4709 -856 4743
rect -914 4675 -856 4709
rect -914 4641 -902 4675
rect -868 4641 -856 4675
rect -914 4607 -856 4641
rect -914 4573 -902 4607
rect -868 4573 -856 4607
rect -914 4539 -856 4573
rect -914 4505 -902 4539
rect -868 4505 -856 4539
rect -914 4471 -856 4505
rect -914 4437 -902 4471
rect -868 4437 -856 4471
rect -914 4403 -856 4437
rect -914 4369 -902 4403
rect -868 4369 -856 4403
rect -914 4335 -856 4369
rect -914 4301 -902 4335
rect -868 4301 -856 4335
rect -914 4267 -856 4301
rect -914 4233 -902 4267
rect -868 4233 -856 4267
rect -914 4199 -856 4233
rect -914 4165 -902 4199
rect -868 4165 -856 4199
rect -914 4131 -856 4165
rect -914 4097 -902 4131
rect -868 4097 -856 4131
rect -914 4063 -856 4097
rect -914 4029 -902 4063
rect -868 4029 -856 4063
rect -914 3995 -856 4029
rect -914 3961 -902 3995
rect -868 3961 -856 3995
rect -914 3927 -856 3961
rect -914 3893 -902 3927
rect -868 3893 -856 3927
rect -914 3859 -856 3893
rect -914 3825 -902 3859
rect -868 3825 -856 3859
rect -914 3791 -856 3825
rect -914 3757 -902 3791
rect -868 3757 -856 3791
rect -914 3723 -856 3757
rect -914 3689 -902 3723
rect -868 3689 -856 3723
rect -914 3655 -856 3689
rect -914 3621 -902 3655
rect -868 3621 -856 3655
rect -914 3587 -856 3621
rect -914 3553 -902 3587
rect -868 3553 -856 3587
rect -914 3519 -856 3553
rect -914 3485 -902 3519
rect -868 3485 -856 3519
rect -914 3451 -856 3485
rect -914 3417 -902 3451
rect -868 3417 -856 3451
rect -914 3383 -856 3417
rect -914 3349 -902 3383
rect -868 3349 -856 3383
rect -914 3315 -856 3349
rect -914 3281 -902 3315
rect -868 3281 -856 3315
rect -914 3247 -856 3281
rect -914 3213 -902 3247
rect -868 3213 -856 3247
rect -914 3179 -856 3213
rect -914 3145 -902 3179
rect -868 3145 -856 3179
rect -914 3111 -856 3145
rect -914 3077 -902 3111
rect -868 3077 -856 3111
rect -914 3043 -856 3077
rect -914 3009 -902 3043
rect -868 3009 -856 3043
rect -914 2975 -856 3009
rect -914 2941 -902 2975
rect -868 2941 -856 2975
rect -914 2907 -856 2941
rect -914 2873 -902 2907
rect -868 2873 -856 2907
rect -914 2839 -856 2873
rect -914 2805 -902 2839
rect -868 2805 -856 2839
rect -914 2771 -856 2805
rect -914 2737 -902 2771
rect -868 2737 -856 2771
rect -914 2703 -856 2737
rect -914 2669 -902 2703
rect -868 2669 -856 2703
rect -914 2635 -856 2669
rect -914 2601 -902 2635
rect -868 2601 -856 2635
rect -914 2567 -856 2601
rect -914 2533 -902 2567
rect -868 2533 -856 2567
rect -914 2499 -856 2533
rect -914 2465 -902 2499
rect -868 2465 -856 2499
rect -914 2431 -856 2465
rect -914 2397 -902 2431
rect -868 2397 -856 2431
rect -914 2363 -856 2397
rect -914 2329 -902 2363
rect -868 2329 -856 2363
rect -914 2295 -856 2329
rect -914 2261 -902 2295
rect -868 2261 -856 2295
rect -914 2227 -856 2261
rect -914 2193 -902 2227
rect -868 2193 -856 2227
rect -914 2159 -856 2193
rect -914 2125 -902 2159
rect -868 2125 -856 2159
rect -914 2091 -856 2125
rect -914 2057 -902 2091
rect -868 2057 -856 2091
rect -914 2023 -856 2057
rect -914 1989 -902 2023
rect -868 1989 -856 2023
rect -914 1955 -856 1989
rect -914 1921 -902 1955
rect -868 1921 -856 1955
rect -914 1887 -856 1921
rect -914 1853 -902 1887
rect -868 1853 -856 1887
rect -914 1819 -856 1853
rect -914 1785 -902 1819
rect -868 1785 -856 1819
rect -914 1751 -856 1785
rect -914 1717 -902 1751
rect -868 1717 -856 1751
rect -914 1683 -856 1717
rect -914 1649 -902 1683
rect -868 1649 -856 1683
rect -914 1615 -856 1649
rect -914 1581 -902 1615
rect -868 1581 -856 1615
rect -914 1547 -856 1581
rect -914 1513 -902 1547
rect -868 1513 -856 1547
rect -914 1479 -856 1513
rect -914 1445 -902 1479
rect -868 1445 -856 1479
rect -914 1411 -856 1445
rect -914 1377 -902 1411
rect -868 1377 -856 1411
rect -914 1343 -856 1377
rect -914 1309 -902 1343
rect -868 1309 -856 1343
rect -914 1275 -856 1309
rect -914 1241 -902 1275
rect -868 1241 -856 1275
rect -914 1207 -856 1241
rect -914 1173 -902 1207
rect -868 1173 -856 1207
rect -914 1139 -856 1173
rect -914 1105 -902 1139
rect -868 1105 -856 1139
rect -914 1071 -856 1105
rect -914 1037 -902 1071
rect -868 1037 -856 1071
rect -914 1003 -856 1037
rect -914 969 -902 1003
rect -868 969 -856 1003
rect -914 935 -856 969
rect -914 901 -902 935
rect -868 901 -856 935
rect -914 867 -856 901
rect -914 833 -902 867
rect -868 833 -856 867
rect -914 799 -856 833
rect -914 765 -902 799
rect -868 765 -856 799
rect -914 731 -856 765
rect -914 697 -902 731
rect -868 697 -856 731
rect -914 663 -856 697
rect -914 629 -902 663
rect -868 629 -856 663
rect -914 595 -856 629
rect -914 561 -902 595
rect -868 561 -856 595
rect -914 527 -856 561
rect -914 493 -902 527
rect -868 493 -856 527
rect -914 459 -856 493
rect -914 425 -902 459
rect -868 425 -856 459
rect -914 391 -856 425
rect -914 357 -902 391
rect -868 357 -856 391
rect -914 323 -856 357
rect -914 289 -902 323
rect -868 289 -856 323
rect -914 255 -856 289
rect -914 221 -902 255
rect -868 221 -856 255
rect -914 187 -856 221
rect -914 153 -902 187
rect -868 153 -856 187
rect -914 119 -856 153
rect -914 85 -902 119
rect -868 85 -856 119
rect -914 51 -856 85
rect -914 17 -902 51
rect -868 17 -856 51
rect -914 -17 -856 17
rect -914 -51 -902 -17
rect -868 -51 -856 -17
rect -914 -85 -856 -51
rect -914 -119 -902 -85
rect -868 -119 -856 -85
rect -914 -153 -856 -119
rect -914 -187 -902 -153
rect -868 -187 -856 -153
rect -914 -221 -856 -187
rect -914 -255 -902 -221
rect -868 -255 -856 -221
rect -914 -289 -856 -255
rect -914 -323 -902 -289
rect -868 -323 -856 -289
rect -914 -357 -856 -323
rect -914 -391 -902 -357
rect -868 -391 -856 -357
rect -914 -425 -856 -391
rect -914 -459 -902 -425
rect -868 -459 -856 -425
rect -914 -493 -856 -459
rect -914 -527 -902 -493
rect -868 -527 -856 -493
rect -914 -561 -856 -527
rect -914 -595 -902 -561
rect -868 -595 -856 -561
rect -914 -629 -856 -595
rect -914 -663 -902 -629
rect -868 -663 -856 -629
rect -914 -697 -856 -663
rect -914 -731 -902 -697
rect -868 -731 -856 -697
rect -914 -765 -856 -731
rect -914 -799 -902 -765
rect -868 -799 -856 -765
rect -914 -833 -856 -799
rect -914 -867 -902 -833
rect -868 -867 -856 -833
rect -914 -901 -856 -867
rect -914 -935 -902 -901
rect -868 -935 -856 -901
rect -914 -969 -856 -935
rect -914 -1003 -902 -969
rect -868 -1003 -856 -969
rect -914 -1037 -856 -1003
rect -914 -1071 -902 -1037
rect -868 -1071 -856 -1037
rect -914 -1105 -856 -1071
rect -914 -1139 -902 -1105
rect -868 -1139 -856 -1105
rect -914 -1173 -856 -1139
rect -914 -1207 -902 -1173
rect -868 -1207 -856 -1173
rect -914 -1241 -856 -1207
rect -914 -1275 -902 -1241
rect -868 -1275 -856 -1241
rect -914 -1309 -856 -1275
rect -914 -1343 -902 -1309
rect -868 -1343 -856 -1309
rect -914 -1377 -856 -1343
rect -914 -1411 -902 -1377
rect -868 -1411 -856 -1377
rect -914 -1445 -856 -1411
rect -914 -1479 -902 -1445
rect -868 -1479 -856 -1445
rect -914 -1513 -856 -1479
rect -914 -1547 -902 -1513
rect -868 -1547 -856 -1513
rect -914 -1581 -856 -1547
rect -914 -1615 -902 -1581
rect -868 -1615 -856 -1581
rect -914 -1649 -856 -1615
rect -914 -1683 -902 -1649
rect -868 -1683 -856 -1649
rect -914 -1717 -856 -1683
rect -914 -1751 -902 -1717
rect -868 -1751 -856 -1717
rect -914 -1785 -856 -1751
rect -914 -1819 -902 -1785
rect -868 -1819 -856 -1785
rect -914 -1853 -856 -1819
rect -914 -1887 -902 -1853
rect -868 -1887 -856 -1853
rect -914 -1921 -856 -1887
rect -914 -1955 -902 -1921
rect -868 -1955 -856 -1921
rect -914 -1989 -856 -1955
rect -914 -2023 -902 -1989
rect -868 -2023 -856 -1989
rect -914 -2057 -856 -2023
rect -914 -2091 -902 -2057
rect -868 -2091 -856 -2057
rect -914 -2125 -856 -2091
rect -914 -2159 -902 -2125
rect -868 -2159 -856 -2125
rect -914 -2193 -856 -2159
rect -914 -2227 -902 -2193
rect -868 -2227 -856 -2193
rect -914 -2261 -856 -2227
rect -914 -2295 -902 -2261
rect -868 -2295 -856 -2261
rect -914 -2329 -856 -2295
rect -914 -2363 -902 -2329
rect -868 -2363 -856 -2329
rect -914 -2397 -856 -2363
rect -914 -2431 -902 -2397
rect -868 -2431 -856 -2397
rect -914 -2465 -856 -2431
rect -914 -2499 -902 -2465
rect -868 -2499 -856 -2465
rect -914 -2533 -856 -2499
rect -914 -2567 -902 -2533
rect -868 -2567 -856 -2533
rect -914 -2601 -856 -2567
rect -914 -2635 -902 -2601
rect -868 -2635 -856 -2601
rect -914 -2669 -856 -2635
rect -914 -2703 -902 -2669
rect -868 -2703 -856 -2669
rect -914 -2737 -856 -2703
rect -914 -2771 -902 -2737
rect -868 -2771 -856 -2737
rect -914 -2805 -856 -2771
rect -914 -2839 -902 -2805
rect -868 -2839 -856 -2805
rect -914 -2873 -856 -2839
rect -914 -2907 -902 -2873
rect -868 -2907 -856 -2873
rect -914 -2941 -856 -2907
rect -914 -2975 -902 -2941
rect -868 -2975 -856 -2941
rect -914 -3009 -856 -2975
rect -914 -3043 -902 -3009
rect -868 -3043 -856 -3009
rect -914 -3077 -856 -3043
rect -914 -3111 -902 -3077
rect -868 -3111 -856 -3077
rect -914 -3145 -856 -3111
rect -914 -3179 -902 -3145
rect -868 -3179 -856 -3145
rect -914 -3213 -856 -3179
rect -914 -3247 -902 -3213
rect -868 -3247 -856 -3213
rect -914 -3281 -856 -3247
rect -914 -3315 -902 -3281
rect -868 -3315 -856 -3281
rect -914 -3349 -856 -3315
rect -914 -3383 -902 -3349
rect -868 -3383 -856 -3349
rect -914 -3417 -856 -3383
rect -914 -3451 -902 -3417
rect -868 -3451 -856 -3417
rect -914 -3485 -856 -3451
rect -914 -3519 -902 -3485
rect -868 -3519 -856 -3485
rect -914 -3553 -856 -3519
rect -914 -3587 -902 -3553
rect -868 -3587 -856 -3553
rect -914 -3621 -856 -3587
rect -914 -3655 -902 -3621
rect -868 -3655 -856 -3621
rect -914 -3689 -856 -3655
rect -914 -3723 -902 -3689
rect -868 -3723 -856 -3689
rect -914 -3757 -856 -3723
rect -914 -3791 -902 -3757
rect -868 -3791 -856 -3757
rect -914 -3825 -856 -3791
rect -914 -3859 -902 -3825
rect -868 -3859 -856 -3825
rect -914 -3893 -856 -3859
rect -914 -3927 -902 -3893
rect -868 -3927 -856 -3893
rect -914 -3961 -856 -3927
rect -914 -3995 -902 -3961
rect -868 -3995 -856 -3961
rect -914 -4029 -856 -3995
rect -914 -4063 -902 -4029
rect -868 -4063 -856 -4029
rect -914 -4097 -856 -4063
rect -914 -4131 -902 -4097
rect -868 -4131 -856 -4097
rect -914 -4165 -856 -4131
rect -914 -4199 -902 -4165
rect -868 -4199 -856 -4165
rect -914 -4233 -856 -4199
rect -914 -4267 -902 -4233
rect -868 -4267 -856 -4233
rect -914 -4301 -856 -4267
rect -914 -4335 -902 -4301
rect -868 -4335 -856 -4301
rect -914 -4369 -856 -4335
rect -914 -4403 -902 -4369
rect -868 -4403 -856 -4369
rect -914 -4437 -856 -4403
rect -914 -4471 -902 -4437
rect -868 -4471 -856 -4437
rect -914 -4505 -856 -4471
rect -914 -4539 -902 -4505
rect -868 -4539 -856 -4505
rect -914 -4573 -856 -4539
rect -914 -4607 -902 -4573
rect -868 -4607 -856 -4573
rect -914 -4641 -856 -4607
rect -914 -4675 -902 -4641
rect -868 -4675 -856 -4641
rect -914 -4709 -856 -4675
rect -914 -4743 -902 -4709
rect -868 -4743 -856 -4709
rect -914 -4777 -856 -4743
rect -914 -4811 -902 -4777
rect -868 -4811 -856 -4777
rect -914 -4845 -856 -4811
rect -914 -4879 -902 -4845
rect -868 -4879 -856 -4845
rect -914 -4913 -856 -4879
rect -914 -4947 -902 -4913
rect -868 -4947 -856 -4913
rect -914 -4981 -856 -4947
rect -914 -5015 -902 -4981
rect -868 -5015 -856 -4981
rect -914 -5049 -856 -5015
rect -914 -5083 -902 -5049
rect -868 -5083 -856 -5049
rect -914 -5117 -856 -5083
rect -914 -5151 -902 -5117
rect -868 -5151 -856 -5117
rect -914 -5185 -856 -5151
rect -914 -5219 -902 -5185
rect -868 -5219 -856 -5185
rect -914 -5253 -856 -5219
rect -914 -5287 -902 -5253
rect -868 -5287 -856 -5253
rect -914 -5321 -856 -5287
rect -914 -5355 -902 -5321
rect -868 -5355 -856 -5321
rect -914 -5389 -856 -5355
rect -914 -5423 -902 -5389
rect -868 -5423 -856 -5389
rect -914 -5457 -856 -5423
rect -914 -5491 -902 -5457
rect -868 -5491 -856 -5457
rect -914 -5525 -856 -5491
rect -914 -5559 -902 -5525
rect -868 -5559 -856 -5525
rect -914 -5593 -856 -5559
rect -914 -5627 -902 -5593
rect -868 -5627 -856 -5593
rect -914 -5661 -856 -5627
rect -914 -5695 -902 -5661
rect -868 -5695 -856 -5661
rect -914 -5729 -856 -5695
rect -914 -5763 -902 -5729
rect -868 -5763 -856 -5729
rect -914 -5797 -856 -5763
rect -914 -5831 -902 -5797
rect -868 -5831 -856 -5797
rect -914 -5865 -856 -5831
rect -914 -5899 -902 -5865
rect -868 -5899 -856 -5865
rect -914 -5933 -856 -5899
rect -914 -5967 -902 -5933
rect -868 -5967 -856 -5933
rect -914 -6001 -856 -5967
rect -914 -6035 -902 -6001
rect -868 -6035 -856 -6001
rect -914 -6069 -856 -6035
rect -914 -6103 -902 -6069
rect -868 -6103 -856 -6069
rect -914 -6137 -856 -6103
rect -914 -6171 -902 -6137
rect -868 -6171 -856 -6137
rect -914 -6205 -856 -6171
rect -914 -6239 -902 -6205
rect -868 -6239 -856 -6205
rect -914 -6273 -856 -6239
rect -914 -6307 -902 -6273
rect -868 -6307 -856 -6273
rect -914 -6341 -856 -6307
rect -914 -6375 -902 -6341
rect -868 -6375 -856 -6341
rect -914 -6409 -856 -6375
rect -914 -6443 -902 -6409
rect -868 -6443 -856 -6409
rect -914 -6477 -856 -6443
rect -914 -6511 -902 -6477
rect -868 -6511 -856 -6477
rect -914 -6545 -856 -6511
rect -914 -6579 -902 -6545
rect -868 -6579 -856 -6545
rect -914 -6613 -856 -6579
rect -914 -6647 -902 -6613
rect -868 -6647 -856 -6613
rect -914 -6681 -856 -6647
rect -914 -6715 -902 -6681
rect -868 -6715 -856 -6681
rect -914 -6749 -856 -6715
rect -914 -6783 -902 -6749
rect -868 -6783 -856 -6749
rect -914 -6817 -856 -6783
rect -914 -6851 -902 -6817
rect -868 -6851 -856 -6817
rect -914 -6885 -856 -6851
rect -914 -6919 -902 -6885
rect -868 -6919 -856 -6885
rect -914 -6953 -856 -6919
rect -914 -6987 -902 -6953
rect -868 -6987 -856 -6953
rect -914 -7021 -856 -6987
rect -914 -7055 -902 -7021
rect -868 -7055 -856 -7021
rect -914 -7089 -856 -7055
rect -914 -7123 -902 -7089
rect -868 -7123 -856 -7089
rect -914 -7157 -856 -7123
rect -914 -7191 -902 -7157
rect -868 -7191 -856 -7157
rect -914 -7225 -856 -7191
rect -914 -7259 -902 -7225
rect -868 -7259 -856 -7225
rect -914 -7293 -856 -7259
rect -914 -7327 -902 -7293
rect -868 -7327 -856 -7293
rect -914 -7361 -856 -7327
rect -914 -7395 -902 -7361
rect -868 -7395 -856 -7361
rect -914 -7429 -856 -7395
rect -914 -7463 -902 -7429
rect -868 -7463 -856 -7429
rect -914 -7497 -856 -7463
rect -914 -7531 -902 -7497
rect -868 -7531 -856 -7497
rect -914 -7565 -856 -7531
rect -914 -7599 -902 -7565
rect -868 -7599 -856 -7565
rect -914 -7633 -856 -7599
rect -914 -7667 -902 -7633
rect -868 -7667 -856 -7633
rect -914 -7701 -856 -7667
rect -914 -7735 -902 -7701
rect -868 -7735 -856 -7701
rect -914 -7769 -856 -7735
rect -914 -7803 -902 -7769
rect -868 -7803 -856 -7769
rect -914 -7837 -856 -7803
rect -914 -7871 -902 -7837
rect -868 -7871 -856 -7837
rect -914 -7905 -856 -7871
rect -914 -7939 -902 -7905
rect -868 -7939 -856 -7905
rect -914 -7973 -856 -7939
rect -914 -8007 -902 -7973
rect -868 -8007 -856 -7973
rect -914 -8041 -856 -8007
rect -914 -8075 -902 -8041
rect -868 -8075 -856 -8041
rect -914 -8109 -856 -8075
rect -914 -8143 -902 -8109
rect -868 -8143 -856 -8109
rect -914 -8177 -856 -8143
rect -914 -8211 -902 -8177
rect -868 -8211 -856 -8177
rect -914 -8245 -856 -8211
rect -914 -8279 -902 -8245
rect -868 -8279 -856 -8245
rect -914 -8313 -856 -8279
rect -914 -8347 -902 -8313
rect -868 -8347 -856 -8313
rect -914 -8381 -856 -8347
rect -914 -8415 -902 -8381
rect -868 -8415 -856 -8381
rect -914 -8449 -856 -8415
rect -914 -8483 -902 -8449
rect -868 -8483 -856 -8449
rect -914 -8517 -856 -8483
rect -914 -8551 -902 -8517
rect -868 -8551 -856 -8517
rect -914 -8585 -856 -8551
rect -914 -8619 -902 -8585
rect -868 -8619 -856 -8585
rect -914 -8653 -856 -8619
rect -914 -8687 -902 -8653
rect -868 -8687 -856 -8653
rect -914 -8721 -856 -8687
rect -914 -8755 -902 -8721
rect -868 -8755 -856 -8721
rect -914 -8789 -856 -8755
rect -914 -8823 -902 -8789
rect -868 -8823 -856 -8789
rect -914 -8857 -856 -8823
rect -914 -8891 -902 -8857
rect -868 -8891 -856 -8857
rect -914 -8925 -856 -8891
rect -914 -8959 -902 -8925
rect -868 -8959 -856 -8925
rect -914 -8993 -856 -8959
rect -914 -9027 -902 -8993
rect -868 -9027 -856 -8993
rect -914 -9061 -856 -9027
rect -914 -9095 -902 -9061
rect -868 -9095 -856 -9061
rect -914 -9129 -856 -9095
rect -914 -9163 -902 -9129
rect -868 -9163 -856 -9129
rect -914 -9197 -856 -9163
rect -914 -9231 -902 -9197
rect -868 -9231 -856 -9197
rect -914 -9265 -856 -9231
rect -914 -9299 -902 -9265
rect -868 -9299 -856 -9265
rect -914 -9333 -856 -9299
rect -914 -9367 -902 -9333
rect -868 -9367 -856 -9333
rect -914 -9401 -856 -9367
rect -914 -9435 -902 -9401
rect -868 -9435 -856 -9401
rect -914 -9469 -856 -9435
rect -914 -9503 -902 -9469
rect -868 -9503 -856 -9469
rect -914 -9537 -856 -9503
rect -914 -9571 -902 -9537
rect -868 -9571 -856 -9537
rect -914 -9600 -856 -9571
rect -796 9571 -738 9600
rect -796 9537 -784 9571
rect -750 9537 -738 9571
rect -796 9503 -738 9537
rect -796 9469 -784 9503
rect -750 9469 -738 9503
rect -796 9435 -738 9469
rect -796 9401 -784 9435
rect -750 9401 -738 9435
rect -796 9367 -738 9401
rect -796 9333 -784 9367
rect -750 9333 -738 9367
rect -796 9299 -738 9333
rect -796 9265 -784 9299
rect -750 9265 -738 9299
rect -796 9231 -738 9265
rect -796 9197 -784 9231
rect -750 9197 -738 9231
rect -796 9163 -738 9197
rect -796 9129 -784 9163
rect -750 9129 -738 9163
rect -796 9095 -738 9129
rect -796 9061 -784 9095
rect -750 9061 -738 9095
rect -796 9027 -738 9061
rect -796 8993 -784 9027
rect -750 8993 -738 9027
rect -796 8959 -738 8993
rect -796 8925 -784 8959
rect -750 8925 -738 8959
rect -796 8891 -738 8925
rect -796 8857 -784 8891
rect -750 8857 -738 8891
rect -796 8823 -738 8857
rect -796 8789 -784 8823
rect -750 8789 -738 8823
rect -796 8755 -738 8789
rect -796 8721 -784 8755
rect -750 8721 -738 8755
rect -796 8687 -738 8721
rect -796 8653 -784 8687
rect -750 8653 -738 8687
rect -796 8619 -738 8653
rect -796 8585 -784 8619
rect -750 8585 -738 8619
rect -796 8551 -738 8585
rect -796 8517 -784 8551
rect -750 8517 -738 8551
rect -796 8483 -738 8517
rect -796 8449 -784 8483
rect -750 8449 -738 8483
rect -796 8415 -738 8449
rect -796 8381 -784 8415
rect -750 8381 -738 8415
rect -796 8347 -738 8381
rect -796 8313 -784 8347
rect -750 8313 -738 8347
rect -796 8279 -738 8313
rect -796 8245 -784 8279
rect -750 8245 -738 8279
rect -796 8211 -738 8245
rect -796 8177 -784 8211
rect -750 8177 -738 8211
rect -796 8143 -738 8177
rect -796 8109 -784 8143
rect -750 8109 -738 8143
rect -796 8075 -738 8109
rect -796 8041 -784 8075
rect -750 8041 -738 8075
rect -796 8007 -738 8041
rect -796 7973 -784 8007
rect -750 7973 -738 8007
rect -796 7939 -738 7973
rect -796 7905 -784 7939
rect -750 7905 -738 7939
rect -796 7871 -738 7905
rect -796 7837 -784 7871
rect -750 7837 -738 7871
rect -796 7803 -738 7837
rect -796 7769 -784 7803
rect -750 7769 -738 7803
rect -796 7735 -738 7769
rect -796 7701 -784 7735
rect -750 7701 -738 7735
rect -796 7667 -738 7701
rect -796 7633 -784 7667
rect -750 7633 -738 7667
rect -796 7599 -738 7633
rect -796 7565 -784 7599
rect -750 7565 -738 7599
rect -796 7531 -738 7565
rect -796 7497 -784 7531
rect -750 7497 -738 7531
rect -796 7463 -738 7497
rect -796 7429 -784 7463
rect -750 7429 -738 7463
rect -796 7395 -738 7429
rect -796 7361 -784 7395
rect -750 7361 -738 7395
rect -796 7327 -738 7361
rect -796 7293 -784 7327
rect -750 7293 -738 7327
rect -796 7259 -738 7293
rect -796 7225 -784 7259
rect -750 7225 -738 7259
rect -796 7191 -738 7225
rect -796 7157 -784 7191
rect -750 7157 -738 7191
rect -796 7123 -738 7157
rect -796 7089 -784 7123
rect -750 7089 -738 7123
rect -796 7055 -738 7089
rect -796 7021 -784 7055
rect -750 7021 -738 7055
rect -796 6987 -738 7021
rect -796 6953 -784 6987
rect -750 6953 -738 6987
rect -796 6919 -738 6953
rect -796 6885 -784 6919
rect -750 6885 -738 6919
rect -796 6851 -738 6885
rect -796 6817 -784 6851
rect -750 6817 -738 6851
rect -796 6783 -738 6817
rect -796 6749 -784 6783
rect -750 6749 -738 6783
rect -796 6715 -738 6749
rect -796 6681 -784 6715
rect -750 6681 -738 6715
rect -796 6647 -738 6681
rect -796 6613 -784 6647
rect -750 6613 -738 6647
rect -796 6579 -738 6613
rect -796 6545 -784 6579
rect -750 6545 -738 6579
rect -796 6511 -738 6545
rect -796 6477 -784 6511
rect -750 6477 -738 6511
rect -796 6443 -738 6477
rect -796 6409 -784 6443
rect -750 6409 -738 6443
rect -796 6375 -738 6409
rect -796 6341 -784 6375
rect -750 6341 -738 6375
rect -796 6307 -738 6341
rect -796 6273 -784 6307
rect -750 6273 -738 6307
rect -796 6239 -738 6273
rect -796 6205 -784 6239
rect -750 6205 -738 6239
rect -796 6171 -738 6205
rect -796 6137 -784 6171
rect -750 6137 -738 6171
rect -796 6103 -738 6137
rect -796 6069 -784 6103
rect -750 6069 -738 6103
rect -796 6035 -738 6069
rect -796 6001 -784 6035
rect -750 6001 -738 6035
rect -796 5967 -738 6001
rect -796 5933 -784 5967
rect -750 5933 -738 5967
rect -796 5899 -738 5933
rect -796 5865 -784 5899
rect -750 5865 -738 5899
rect -796 5831 -738 5865
rect -796 5797 -784 5831
rect -750 5797 -738 5831
rect -796 5763 -738 5797
rect -796 5729 -784 5763
rect -750 5729 -738 5763
rect -796 5695 -738 5729
rect -796 5661 -784 5695
rect -750 5661 -738 5695
rect -796 5627 -738 5661
rect -796 5593 -784 5627
rect -750 5593 -738 5627
rect -796 5559 -738 5593
rect -796 5525 -784 5559
rect -750 5525 -738 5559
rect -796 5491 -738 5525
rect -796 5457 -784 5491
rect -750 5457 -738 5491
rect -796 5423 -738 5457
rect -796 5389 -784 5423
rect -750 5389 -738 5423
rect -796 5355 -738 5389
rect -796 5321 -784 5355
rect -750 5321 -738 5355
rect -796 5287 -738 5321
rect -796 5253 -784 5287
rect -750 5253 -738 5287
rect -796 5219 -738 5253
rect -796 5185 -784 5219
rect -750 5185 -738 5219
rect -796 5151 -738 5185
rect -796 5117 -784 5151
rect -750 5117 -738 5151
rect -796 5083 -738 5117
rect -796 5049 -784 5083
rect -750 5049 -738 5083
rect -796 5015 -738 5049
rect -796 4981 -784 5015
rect -750 4981 -738 5015
rect -796 4947 -738 4981
rect -796 4913 -784 4947
rect -750 4913 -738 4947
rect -796 4879 -738 4913
rect -796 4845 -784 4879
rect -750 4845 -738 4879
rect -796 4811 -738 4845
rect -796 4777 -784 4811
rect -750 4777 -738 4811
rect -796 4743 -738 4777
rect -796 4709 -784 4743
rect -750 4709 -738 4743
rect -796 4675 -738 4709
rect -796 4641 -784 4675
rect -750 4641 -738 4675
rect -796 4607 -738 4641
rect -796 4573 -784 4607
rect -750 4573 -738 4607
rect -796 4539 -738 4573
rect -796 4505 -784 4539
rect -750 4505 -738 4539
rect -796 4471 -738 4505
rect -796 4437 -784 4471
rect -750 4437 -738 4471
rect -796 4403 -738 4437
rect -796 4369 -784 4403
rect -750 4369 -738 4403
rect -796 4335 -738 4369
rect -796 4301 -784 4335
rect -750 4301 -738 4335
rect -796 4267 -738 4301
rect -796 4233 -784 4267
rect -750 4233 -738 4267
rect -796 4199 -738 4233
rect -796 4165 -784 4199
rect -750 4165 -738 4199
rect -796 4131 -738 4165
rect -796 4097 -784 4131
rect -750 4097 -738 4131
rect -796 4063 -738 4097
rect -796 4029 -784 4063
rect -750 4029 -738 4063
rect -796 3995 -738 4029
rect -796 3961 -784 3995
rect -750 3961 -738 3995
rect -796 3927 -738 3961
rect -796 3893 -784 3927
rect -750 3893 -738 3927
rect -796 3859 -738 3893
rect -796 3825 -784 3859
rect -750 3825 -738 3859
rect -796 3791 -738 3825
rect -796 3757 -784 3791
rect -750 3757 -738 3791
rect -796 3723 -738 3757
rect -796 3689 -784 3723
rect -750 3689 -738 3723
rect -796 3655 -738 3689
rect -796 3621 -784 3655
rect -750 3621 -738 3655
rect -796 3587 -738 3621
rect -796 3553 -784 3587
rect -750 3553 -738 3587
rect -796 3519 -738 3553
rect -796 3485 -784 3519
rect -750 3485 -738 3519
rect -796 3451 -738 3485
rect -796 3417 -784 3451
rect -750 3417 -738 3451
rect -796 3383 -738 3417
rect -796 3349 -784 3383
rect -750 3349 -738 3383
rect -796 3315 -738 3349
rect -796 3281 -784 3315
rect -750 3281 -738 3315
rect -796 3247 -738 3281
rect -796 3213 -784 3247
rect -750 3213 -738 3247
rect -796 3179 -738 3213
rect -796 3145 -784 3179
rect -750 3145 -738 3179
rect -796 3111 -738 3145
rect -796 3077 -784 3111
rect -750 3077 -738 3111
rect -796 3043 -738 3077
rect -796 3009 -784 3043
rect -750 3009 -738 3043
rect -796 2975 -738 3009
rect -796 2941 -784 2975
rect -750 2941 -738 2975
rect -796 2907 -738 2941
rect -796 2873 -784 2907
rect -750 2873 -738 2907
rect -796 2839 -738 2873
rect -796 2805 -784 2839
rect -750 2805 -738 2839
rect -796 2771 -738 2805
rect -796 2737 -784 2771
rect -750 2737 -738 2771
rect -796 2703 -738 2737
rect -796 2669 -784 2703
rect -750 2669 -738 2703
rect -796 2635 -738 2669
rect -796 2601 -784 2635
rect -750 2601 -738 2635
rect -796 2567 -738 2601
rect -796 2533 -784 2567
rect -750 2533 -738 2567
rect -796 2499 -738 2533
rect -796 2465 -784 2499
rect -750 2465 -738 2499
rect -796 2431 -738 2465
rect -796 2397 -784 2431
rect -750 2397 -738 2431
rect -796 2363 -738 2397
rect -796 2329 -784 2363
rect -750 2329 -738 2363
rect -796 2295 -738 2329
rect -796 2261 -784 2295
rect -750 2261 -738 2295
rect -796 2227 -738 2261
rect -796 2193 -784 2227
rect -750 2193 -738 2227
rect -796 2159 -738 2193
rect -796 2125 -784 2159
rect -750 2125 -738 2159
rect -796 2091 -738 2125
rect -796 2057 -784 2091
rect -750 2057 -738 2091
rect -796 2023 -738 2057
rect -796 1989 -784 2023
rect -750 1989 -738 2023
rect -796 1955 -738 1989
rect -796 1921 -784 1955
rect -750 1921 -738 1955
rect -796 1887 -738 1921
rect -796 1853 -784 1887
rect -750 1853 -738 1887
rect -796 1819 -738 1853
rect -796 1785 -784 1819
rect -750 1785 -738 1819
rect -796 1751 -738 1785
rect -796 1717 -784 1751
rect -750 1717 -738 1751
rect -796 1683 -738 1717
rect -796 1649 -784 1683
rect -750 1649 -738 1683
rect -796 1615 -738 1649
rect -796 1581 -784 1615
rect -750 1581 -738 1615
rect -796 1547 -738 1581
rect -796 1513 -784 1547
rect -750 1513 -738 1547
rect -796 1479 -738 1513
rect -796 1445 -784 1479
rect -750 1445 -738 1479
rect -796 1411 -738 1445
rect -796 1377 -784 1411
rect -750 1377 -738 1411
rect -796 1343 -738 1377
rect -796 1309 -784 1343
rect -750 1309 -738 1343
rect -796 1275 -738 1309
rect -796 1241 -784 1275
rect -750 1241 -738 1275
rect -796 1207 -738 1241
rect -796 1173 -784 1207
rect -750 1173 -738 1207
rect -796 1139 -738 1173
rect -796 1105 -784 1139
rect -750 1105 -738 1139
rect -796 1071 -738 1105
rect -796 1037 -784 1071
rect -750 1037 -738 1071
rect -796 1003 -738 1037
rect -796 969 -784 1003
rect -750 969 -738 1003
rect -796 935 -738 969
rect -796 901 -784 935
rect -750 901 -738 935
rect -796 867 -738 901
rect -796 833 -784 867
rect -750 833 -738 867
rect -796 799 -738 833
rect -796 765 -784 799
rect -750 765 -738 799
rect -796 731 -738 765
rect -796 697 -784 731
rect -750 697 -738 731
rect -796 663 -738 697
rect -796 629 -784 663
rect -750 629 -738 663
rect -796 595 -738 629
rect -796 561 -784 595
rect -750 561 -738 595
rect -796 527 -738 561
rect -796 493 -784 527
rect -750 493 -738 527
rect -796 459 -738 493
rect -796 425 -784 459
rect -750 425 -738 459
rect -796 391 -738 425
rect -796 357 -784 391
rect -750 357 -738 391
rect -796 323 -738 357
rect -796 289 -784 323
rect -750 289 -738 323
rect -796 255 -738 289
rect -796 221 -784 255
rect -750 221 -738 255
rect -796 187 -738 221
rect -796 153 -784 187
rect -750 153 -738 187
rect -796 119 -738 153
rect -796 85 -784 119
rect -750 85 -738 119
rect -796 51 -738 85
rect -796 17 -784 51
rect -750 17 -738 51
rect -796 -17 -738 17
rect -796 -51 -784 -17
rect -750 -51 -738 -17
rect -796 -85 -738 -51
rect -796 -119 -784 -85
rect -750 -119 -738 -85
rect -796 -153 -738 -119
rect -796 -187 -784 -153
rect -750 -187 -738 -153
rect -796 -221 -738 -187
rect -796 -255 -784 -221
rect -750 -255 -738 -221
rect -796 -289 -738 -255
rect -796 -323 -784 -289
rect -750 -323 -738 -289
rect -796 -357 -738 -323
rect -796 -391 -784 -357
rect -750 -391 -738 -357
rect -796 -425 -738 -391
rect -796 -459 -784 -425
rect -750 -459 -738 -425
rect -796 -493 -738 -459
rect -796 -527 -784 -493
rect -750 -527 -738 -493
rect -796 -561 -738 -527
rect -796 -595 -784 -561
rect -750 -595 -738 -561
rect -796 -629 -738 -595
rect -796 -663 -784 -629
rect -750 -663 -738 -629
rect -796 -697 -738 -663
rect -796 -731 -784 -697
rect -750 -731 -738 -697
rect -796 -765 -738 -731
rect -796 -799 -784 -765
rect -750 -799 -738 -765
rect -796 -833 -738 -799
rect -796 -867 -784 -833
rect -750 -867 -738 -833
rect -796 -901 -738 -867
rect -796 -935 -784 -901
rect -750 -935 -738 -901
rect -796 -969 -738 -935
rect -796 -1003 -784 -969
rect -750 -1003 -738 -969
rect -796 -1037 -738 -1003
rect -796 -1071 -784 -1037
rect -750 -1071 -738 -1037
rect -796 -1105 -738 -1071
rect -796 -1139 -784 -1105
rect -750 -1139 -738 -1105
rect -796 -1173 -738 -1139
rect -796 -1207 -784 -1173
rect -750 -1207 -738 -1173
rect -796 -1241 -738 -1207
rect -796 -1275 -784 -1241
rect -750 -1275 -738 -1241
rect -796 -1309 -738 -1275
rect -796 -1343 -784 -1309
rect -750 -1343 -738 -1309
rect -796 -1377 -738 -1343
rect -796 -1411 -784 -1377
rect -750 -1411 -738 -1377
rect -796 -1445 -738 -1411
rect -796 -1479 -784 -1445
rect -750 -1479 -738 -1445
rect -796 -1513 -738 -1479
rect -796 -1547 -784 -1513
rect -750 -1547 -738 -1513
rect -796 -1581 -738 -1547
rect -796 -1615 -784 -1581
rect -750 -1615 -738 -1581
rect -796 -1649 -738 -1615
rect -796 -1683 -784 -1649
rect -750 -1683 -738 -1649
rect -796 -1717 -738 -1683
rect -796 -1751 -784 -1717
rect -750 -1751 -738 -1717
rect -796 -1785 -738 -1751
rect -796 -1819 -784 -1785
rect -750 -1819 -738 -1785
rect -796 -1853 -738 -1819
rect -796 -1887 -784 -1853
rect -750 -1887 -738 -1853
rect -796 -1921 -738 -1887
rect -796 -1955 -784 -1921
rect -750 -1955 -738 -1921
rect -796 -1989 -738 -1955
rect -796 -2023 -784 -1989
rect -750 -2023 -738 -1989
rect -796 -2057 -738 -2023
rect -796 -2091 -784 -2057
rect -750 -2091 -738 -2057
rect -796 -2125 -738 -2091
rect -796 -2159 -784 -2125
rect -750 -2159 -738 -2125
rect -796 -2193 -738 -2159
rect -796 -2227 -784 -2193
rect -750 -2227 -738 -2193
rect -796 -2261 -738 -2227
rect -796 -2295 -784 -2261
rect -750 -2295 -738 -2261
rect -796 -2329 -738 -2295
rect -796 -2363 -784 -2329
rect -750 -2363 -738 -2329
rect -796 -2397 -738 -2363
rect -796 -2431 -784 -2397
rect -750 -2431 -738 -2397
rect -796 -2465 -738 -2431
rect -796 -2499 -784 -2465
rect -750 -2499 -738 -2465
rect -796 -2533 -738 -2499
rect -796 -2567 -784 -2533
rect -750 -2567 -738 -2533
rect -796 -2601 -738 -2567
rect -796 -2635 -784 -2601
rect -750 -2635 -738 -2601
rect -796 -2669 -738 -2635
rect -796 -2703 -784 -2669
rect -750 -2703 -738 -2669
rect -796 -2737 -738 -2703
rect -796 -2771 -784 -2737
rect -750 -2771 -738 -2737
rect -796 -2805 -738 -2771
rect -796 -2839 -784 -2805
rect -750 -2839 -738 -2805
rect -796 -2873 -738 -2839
rect -796 -2907 -784 -2873
rect -750 -2907 -738 -2873
rect -796 -2941 -738 -2907
rect -796 -2975 -784 -2941
rect -750 -2975 -738 -2941
rect -796 -3009 -738 -2975
rect -796 -3043 -784 -3009
rect -750 -3043 -738 -3009
rect -796 -3077 -738 -3043
rect -796 -3111 -784 -3077
rect -750 -3111 -738 -3077
rect -796 -3145 -738 -3111
rect -796 -3179 -784 -3145
rect -750 -3179 -738 -3145
rect -796 -3213 -738 -3179
rect -796 -3247 -784 -3213
rect -750 -3247 -738 -3213
rect -796 -3281 -738 -3247
rect -796 -3315 -784 -3281
rect -750 -3315 -738 -3281
rect -796 -3349 -738 -3315
rect -796 -3383 -784 -3349
rect -750 -3383 -738 -3349
rect -796 -3417 -738 -3383
rect -796 -3451 -784 -3417
rect -750 -3451 -738 -3417
rect -796 -3485 -738 -3451
rect -796 -3519 -784 -3485
rect -750 -3519 -738 -3485
rect -796 -3553 -738 -3519
rect -796 -3587 -784 -3553
rect -750 -3587 -738 -3553
rect -796 -3621 -738 -3587
rect -796 -3655 -784 -3621
rect -750 -3655 -738 -3621
rect -796 -3689 -738 -3655
rect -796 -3723 -784 -3689
rect -750 -3723 -738 -3689
rect -796 -3757 -738 -3723
rect -796 -3791 -784 -3757
rect -750 -3791 -738 -3757
rect -796 -3825 -738 -3791
rect -796 -3859 -784 -3825
rect -750 -3859 -738 -3825
rect -796 -3893 -738 -3859
rect -796 -3927 -784 -3893
rect -750 -3927 -738 -3893
rect -796 -3961 -738 -3927
rect -796 -3995 -784 -3961
rect -750 -3995 -738 -3961
rect -796 -4029 -738 -3995
rect -796 -4063 -784 -4029
rect -750 -4063 -738 -4029
rect -796 -4097 -738 -4063
rect -796 -4131 -784 -4097
rect -750 -4131 -738 -4097
rect -796 -4165 -738 -4131
rect -796 -4199 -784 -4165
rect -750 -4199 -738 -4165
rect -796 -4233 -738 -4199
rect -796 -4267 -784 -4233
rect -750 -4267 -738 -4233
rect -796 -4301 -738 -4267
rect -796 -4335 -784 -4301
rect -750 -4335 -738 -4301
rect -796 -4369 -738 -4335
rect -796 -4403 -784 -4369
rect -750 -4403 -738 -4369
rect -796 -4437 -738 -4403
rect -796 -4471 -784 -4437
rect -750 -4471 -738 -4437
rect -796 -4505 -738 -4471
rect -796 -4539 -784 -4505
rect -750 -4539 -738 -4505
rect -796 -4573 -738 -4539
rect -796 -4607 -784 -4573
rect -750 -4607 -738 -4573
rect -796 -4641 -738 -4607
rect -796 -4675 -784 -4641
rect -750 -4675 -738 -4641
rect -796 -4709 -738 -4675
rect -796 -4743 -784 -4709
rect -750 -4743 -738 -4709
rect -796 -4777 -738 -4743
rect -796 -4811 -784 -4777
rect -750 -4811 -738 -4777
rect -796 -4845 -738 -4811
rect -796 -4879 -784 -4845
rect -750 -4879 -738 -4845
rect -796 -4913 -738 -4879
rect -796 -4947 -784 -4913
rect -750 -4947 -738 -4913
rect -796 -4981 -738 -4947
rect -796 -5015 -784 -4981
rect -750 -5015 -738 -4981
rect -796 -5049 -738 -5015
rect -796 -5083 -784 -5049
rect -750 -5083 -738 -5049
rect -796 -5117 -738 -5083
rect -796 -5151 -784 -5117
rect -750 -5151 -738 -5117
rect -796 -5185 -738 -5151
rect -796 -5219 -784 -5185
rect -750 -5219 -738 -5185
rect -796 -5253 -738 -5219
rect -796 -5287 -784 -5253
rect -750 -5287 -738 -5253
rect -796 -5321 -738 -5287
rect -796 -5355 -784 -5321
rect -750 -5355 -738 -5321
rect -796 -5389 -738 -5355
rect -796 -5423 -784 -5389
rect -750 -5423 -738 -5389
rect -796 -5457 -738 -5423
rect -796 -5491 -784 -5457
rect -750 -5491 -738 -5457
rect -796 -5525 -738 -5491
rect -796 -5559 -784 -5525
rect -750 -5559 -738 -5525
rect -796 -5593 -738 -5559
rect -796 -5627 -784 -5593
rect -750 -5627 -738 -5593
rect -796 -5661 -738 -5627
rect -796 -5695 -784 -5661
rect -750 -5695 -738 -5661
rect -796 -5729 -738 -5695
rect -796 -5763 -784 -5729
rect -750 -5763 -738 -5729
rect -796 -5797 -738 -5763
rect -796 -5831 -784 -5797
rect -750 -5831 -738 -5797
rect -796 -5865 -738 -5831
rect -796 -5899 -784 -5865
rect -750 -5899 -738 -5865
rect -796 -5933 -738 -5899
rect -796 -5967 -784 -5933
rect -750 -5967 -738 -5933
rect -796 -6001 -738 -5967
rect -796 -6035 -784 -6001
rect -750 -6035 -738 -6001
rect -796 -6069 -738 -6035
rect -796 -6103 -784 -6069
rect -750 -6103 -738 -6069
rect -796 -6137 -738 -6103
rect -796 -6171 -784 -6137
rect -750 -6171 -738 -6137
rect -796 -6205 -738 -6171
rect -796 -6239 -784 -6205
rect -750 -6239 -738 -6205
rect -796 -6273 -738 -6239
rect -796 -6307 -784 -6273
rect -750 -6307 -738 -6273
rect -796 -6341 -738 -6307
rect -796 -6375 -784 -6341
rect -750 -6375 -738 -6341
rect -796 -6409 -738 -6375
rect -796 -6443 -784 -6409
rect -750 -6443 -738 -6409
rect -796 -6477 -738 -6443
rect -796 -6511 -784 -6477
rect -750 -6511 -738 -6477
rect -796 -6545 -738 -6511
rect -796 -6579 -784 -6545
rect -750 -6579 -738 -6545
rect -796 -6613 -738 -6579
rect -796 -6647 -784 -6613
rect -750 -6647 -738 -6613
rect -796 -6681 -738 -6647
rect -796 -6715 -784 -6681
rect -750 -6715 -738 -6681
rect -796 -6749 -738 -6715
rect -796 -6783 -784 -6749
rect -750 -6783 -738 -6749
rect -796 -6817 -738 -6783
rect -796 -6851 -784 -6817
rect -750 -6851 -738 -6817
rect -796 -6885 -738 -6851
rect -796 -6919 -784 -6885
rect -750 -6919 -738 -6885
rect -796 -6953 -738 -6919
rect -796 -6987 -784 -6953
rect -750 -6987 -738 -6953
rect -796 -7021 -738 -6987
rect -796 -7055 -784 -7021
rect -750 -7055 -738 -7021
rect -796 -7089 -738 -7055
rect -796 -7123 -784 -7089
rect -750 -7123 -738 -7089
rect -796 -7157 -738 -7123
rect -796 -7191 -784 -7157
rect -750 -7191 -738 -7157
rect -796 -7225 -738 -7191
rect -796 -7259 -784 -7225
rect -750 -7259 -738 -7225
rect -796 -7293 -738 -7259
rect -796 -7327 -784 -7293
rect -750 -7327 -738 -7293
rect -796 -7361 -738 -7327
rect -796 -7395 -784 -7361
rect -750 -7395 -738 -7361
rect -796 -7429 -738 -7395
rect -796 -7463 -784 -7429
rect -750 -7463 -738 -7429
rect -796 -7497 -738 -7463
rect -796 -7531 -784 -7497
rect -750 -7531 -738 -7497
rect -796 -7565 -738 -7531
rect -796 -7599 -784 -7565
rect -750 -7599 -738 -7565
rect -796 -7633 -738 -7599
rect -796 -7667 -784 -7633
rect -750 -7667 -738 -7633
rect -796 -7701 -738 -7667
rect -796 -7735 -784 -7701
rect -750 -7735 -738 -7701
rect -796 -7769 -738 -7735
rect -796 -7803 -784 -7769
rect -750 -7803 -738 -7769
rect -796 -7837 -738 -7803
rect -796 -7871 -784 -7837
rect -750 -7871 -738 -7837
rect -796 -7905 -738 -7871
rect -796 -7939 -784 -7905
rect -750 -7939 -738 -7905
rect -796 -7973 -738 -7939
rect -796 -8007 -784 -7973
rect -750 -8007 -738 -7973
rect -796 -8041 -738 -8007
rect -796 -8075 -784 -8041
rect -750 -8075 -738 -8041
rect -796 -8109 -738 -8075
rect -796 -8143 -784 -8109
rect -750 -8143 -738 -8109
rect -796 -8177 -738 -8143
rect -796 -8211 -784 -8177
rect -750 -8211 -738 -8177
rect -796 -8245 -738 -8211
rect -796 -8279 -784 -8245
rect -750 -8279 -738 -8245
rect -796 -8313 -738 -8279
rect -796 -8347 -784 -8313
rect -750 -8347 -738 -8313
rect -796 -8381 -738 -8347
rect -796 -8415 -784 -8381
rect -750 -8415 -738 -8381
rect -796 -8449 -738 -8415
rect -796 -8483 -784 -8449
rect -750 -8483 -738 -8449
rect -796 -8517 -738 -8483
rect -796 -8551 -784 -8517
rect -750 -8551 -738 -8517
rect -796 -8585 -738 -8551
rect -796 -8619 -784 -8585
rect -750 -8619 -738 -8585
rect -796 -8653 -738 -8619
rect -796 -8687 -784 -8653
rect -750 -8687 -738 -8653
rect -796 -8721 -738 -8687
rect -796 -8755 -784 -8721
rect -750 -8755 -738 -8721
rect -796 -8789 -738 -8755
rect -796 -8823 -784 -8789
rect -750 -8823 -738 -8789
rect -796 -8857 -738 -8823
rect -796 -8891 -784 -8857
rect -750 -8891 -738 -8857
rect -796 -8925 -738 -8891
rect -796 -8959 -784 -8925
rect -750 -8959 -738 -8925
rect -796 -8993 -738 -8959
rect -796 -9027 -784 -8993
rect -750 -9027 -738 -8993
rect -796 -9061 -738 -9027
rect -796 -9095 -784 -9061
rect -750 -9095 -738 -9061
rect -796 -9129 -738 -9095
rect -796 -9163 -784 -9129
rect -750 -9163 -738 -9129
rect -796 -9197 -738 -9163
rect -796 -9231 -784 -9197
rect -750 -9231 -738 -9197
rect -796 -9265 -738 -9231
rect -796 -9299 -784 -9265
rect -750 -9299 -738 -9265
rect -796 -9333 -738 -9299
rect -796 -9367 -784 -9333
rect -750 -9367 -738 -9333
rect -796 -9401 -738 -9367
rect -796 -9435 -784 -9401
rect -750 -9435 -738 -9401
rect -796 -9469 -738 -9435
rect -796 -9503 -784 -9469
rect -750 -9503 -738 -9469
rect -796 -9537 -738 -9503
rect -796 -9571 -784 -9537
rect -750 -9571 -738 -9537
rect -796 -9600 -738 -9571
rect -678 9571 -620 9600
rect -678 9537 -666 9571
rect -632 9537 -620 9571
rect -678 9503 -620 9537
rect -678 9469 -666 9503
rect -632 9469 -620 9503
rect -678 9435 -620 9469
rect -678 9401 -666 9435
rect -632 9401 -620 9435
rect -678 9367 -620 9401
rect -678 9333 -666 9367
rect -632 9333 -620 9367
rect -678 9299 -620 9333
rect -678 9265 -666 9299
rect -632 9265 -620 9299
rect -678 9231 -620 9265
rect -678 9197 -666 9231
rect -632 9197 -620 9231
rect -678 9163 -620 9197
rect -678 9129 -666 9163
rect -632 9129 -620 9163
rect -678 9095 -620 9129
rect -678 9061 -666 9095
rect -632 9061 -620 9095
rect -678 9027 -620 9061
rect -678 8993 -666 9027
rect -632 8993 -620 9027
rect -678 8959 -620 8993
rect -678 8925 -666 8959
rect -632 8925 -620 8959
rect -678 8891 -620 8925
rect -678 8857 -666 8891
rect -632 8857 -620 8891
rect -678 8823 -620 8857
rect -678 8789 -666 8823
rect -632 8789 -620 8823
rect -678 8755 -620 8789
rect -678 8721 -666 8755
rect -632 8721 -620 8755
rect -678 8687 -620 8721
rect -678 8653 -666 8687
rect -632 8653 -620 8687
rect -678 8619 -620 8653
rect -678 8585 -666 8619
rect -632 8585 -620 8619
rect -678 8551 -620 8585
rect -678 8517 -666 8551
rect -632 8517 -620 8551
rect -678 8483 -620 8517
rect -678 8449 -666 8483
rect -632 8449 -620 8483
rect -678 8415 -620 8449
rect -678 8381 -666 8415
rect -632 8381 -620 8415
rect -678 8347 -620 8381
rect -678 8313 -666 8347
rect -632 8313 -620 8347
rect -678 8279 -620 8313
rect -678 8245 -666 8279
rect -632 8245 -620 8279
rect -678 8211 -620 8245
rect -678 8177 -666 8211
rect -632 8177 -620 8211
rect -678 8143 -620 8177
rect -678 8109 -666 8143
rect -632 8109 -620 8143
rect -678 8075 -620 8109
rect -678 8041 -666 8075
rect -632 8041 -620 8075
rect -678 8007 -620 8041
rect -678 7973 -666 8007
rect -632 7973 -620 8007
rect -678 7939 -620 7973
rect -678 7905 -666 7939
rect -632 7905 -620 7939
rect -678 7871 -620 7905
rect -678 7837 -666 7871
rect -632 7837 -620 7871
rect -678 7803 -620 7837
rect -678 7769 -666 7803
rect -632 7769 -620 7803
rect -678 7735 -620 7769
rect -678 7701 -666 7735
rect -632 7701 -620 7735
rect -678 7667 -620 7701
rect -678 7633 -666 7667
rect -632 7633 -620 7667
rect -678 7599 -620 7633
rect -678 7565 -666 7599
rect -632 7565 -620 7599
rect -678 7531 -620 7565
rect -678 7497 -666 7531
rect -632 7497 -620 7531
rect -678 7463 -620 7497
rect -678 7429 -666 7463
rect -632 7429 -620 7463
rect -678 7395 -620 7429
rect -678 7361 -666 7395
rect -632 7361 -620 7395
rect -678 7327 -620 7361
rect -678 7293 -666 7327
rect -632 7293 -620 7327
rect -678 7259 -620 7293
rect -678 7225 -666 7259
rect -632 7225 -620 7259
rect -678 7191 -620 7225
rect -678 7157 -666 7191
rect -632 7157 -620 7191
rect -678 7123 -620 7157
rect -678 7089 -666 7123
rect -632 7089 -620 7123
rect -678 7055 -620 7089
rect -678 7021 -666 7055
rect -632 7021 -620 7055
rect -678 6987 -620 7021
rect -678 6953 -666 6987
rect -632 6953 -620 6987
rect -678 6919 -620 6953
rect -678 6885 -666 6919
rect -632 6885 -620 6919
rect -678 6851 -620 6885
rect -678 6817 -666 6851
rect -632 6817 -620 6851
rect -678 6783 -620 6817
rect -678 6749 -666 6783
rect -632 6749 -620 6783
rect -678 6715 -620 6749
rect -678 6681 -666 6715
rect -632 6681 -620 6715
rect -678 6647 -620 6681
rect -678 6613 -666 6647
rect -632 6613 -620 6647
rect -678 6579 -620 6613
rect -678 6545 -666 6579
rect -632 6545 -620 6579
rect -678 6511 -620 6545
rect -678 6477 -666 6511
rect -632 6477 -620 6511
rect -678 6443 -620 6477
rect -678 6409 -666 6443
rect -632 6409 -620 6443
rect -678 6375 -620 6409
rect -678 6341 -666 6375
rect -632 6341 -620 6375
rect -678 6307 -620 6341
rect -678 6273 -666 6307
rect -632 6273 -620 6307
rect -678 6239 -620 6273
rect -678 6205 -666 6239
rect -632 6205 -620 6239
rect -678 6171 -620 6205
rect -678 6137 -666 6171
rect -632 6137 -620 6171
rect -678 6103 -620 6137
rect -678 6069 -666 6103
rect -632 6069 -620 6103
rect -678 6035 -620 6069
rect -678 6001 -666 6035
rect -632 6001 -620 6035
rect -678 5967 -620 6001
rect -678 5933 -666 5967
rect -632 5933 -620 5967
rect -678 5899 -620 5933
rect -678 5865 -666 5899
rect -632 5865 -620 5899
rect -678 5831 -620 5865
rect -678 5797 -666 5831
rect -632 5797 -620 5831
rect -678 5763 -620 5797
rect -678 5729 -666 5763
rect -632 5729 -620 5763
rect -678 5695 -620 5729
rect -678 5661 -666 5695
rect -632 5661 -620 5695
rect -678 5627 -620 5661
rect -678 5593 -666 5627
rect -632 5593 -620 5627
rect -678 5559 -620 5593
rect -678 5525 -666 5559
rect -632 5525 -620 5559
rect -678 5491 -620 5525
rect -678 5457 -666 5491
rect -632 5457 -620 5491
rect -678 5423 -620 5457
rect -678 5389 -666 5423
rect -632 5389 -620 5423
rect -678 5355 -620 5389
rect -678 5321 -666 5355
rect -632 5321 -620 5355
rect -678 5287 -620 5321
rect -678 5253 -666 5287
rect -632 5253 -620 5287
rect -678 5219 -620 5253
rect -678 5185 -666 5219
rect -632 5185 -620 5219
rect -678 5151 -620 5185
rect -678 5117 -666 5151
rect -632 5117 -620 5151
rect -678 5083 -620 5117
rect -678 5049 -666 5083
rect -632 5049 -620 5083
rect -678 5015 -620 5049
rect -678 4981 -666 5015
rect -632 4981 -620 5015
rect -678 4947 -620 4981
rect -678 4913 -666 4947
rect -632 4913 -620 4947
rect -678 4879 -620 4913
rect -678 4845 -666 4879
rect -632 4845 -620 4879
rect -678 4811 -620 4845
rect -678 4777 -666 4811
rect -632 4777 -620 4811
rect -678 4743 -620 4777
rect -678 4709 -666 4743
rect -632 4709 -620 4743
rect -678 4675 -620 4709
rect -678 4641 -666 4675
rect -632 4641 -620 4675
rect -678 4607 -620 4641
rect -678 4573 -666 4607
rect -632 4573 -620 4607
rect -678 4539 -620 4573
rect -678 4505 -666 4539
rect -632 4505 -620 4539
rect -678 4471 -620 4505
rect -678 4437 -666 4471
rect -632 4437 -620 4471
rect -678 4403 -620 4437
rect -678 4369 -666 4403
rect -632 4369 -620 4403
rect -678 4335 -620 4369
rect -678 4301 -666 4335
rect -632 4301 -620 4335
rect -678 4267 -620 4301
rect -678 4233 -666 4267
rect -632 4233 -620 4267
rect -678 4199 -620 4233
rect -678 4165 -666 4199
rect -632 4165 -620 4199
rect -678 4131 -620 4165
rect -678 4097 -666 4131
rect -632 4097 -620 4131
rect -678 4063 -620 4097
rect -678 4029 -666 4063
rect -632 4029 -620 4063
rect -678 3995 -620 4029
rect -678 3961 -666 3995
rect -632 3961 -620 3995
rect -678 3927 -620 3961
rect -678 3893 -666 3927
rect -632 3893 -620 3927
rect -678 3859 -620 3893
rect -678 3825 -666 3859
rect -632 3825 -620 3859
rect -678 3791 -620 3825
rect -678 3757 -666 3791
rect -632 3757 -620 3791
rect -678 3723 -620 3757
rect -678 3689 -666 3723
rect -632 3689 -620 3723
rect -678 3655 -620 3689
rect -678 3621 -666 3655
rect -632 3621 -620 3655
rect -678 3587 -620 3621
rect -678 3553 -666 3587
rect -632 3553 -620 3587
rect -678 3519 -620 3553
rect -678 3485 -666 3519
rect -632 3485 -620 3519
rect -678 3451 -620 3485
rect -678 3417 -666 3451
rect -632 3417 -620 3451
rect -678 3383 -620 3417
rect -678 3349 -666 3383
rect -632 3349 -620 3383
rect -678 3315 -620 3349
rect -678 3281 -666 3315
rect -632 3281 -620 3315
rect -678 3247 -620 3281
rect -678 3213 -666 3247
rect -632 3213 -620 3247
rect -678 3179 -620 3213
rect -678 3145 -666 3179
rect -632 3145 -620 3179
rect -678 3111 -620 3145
rect -678 3077 -666 3111
rect -632 3077 -620 3111
rect -678 3043 -620 3077
rect -678 3009 -666 3043
rect -632 3009 -620 3043
rect -678 2975 -620 3009
rect -678 2941 -666 2975
rect -632 2941 -620 2975
rect -678 2907 -620 2941
rect -678 2873 -666 2907
rect -632 2873 -620 2907
rect -678 2839 -620 2873
rect -678 2805 -666 2839
rect -632 2805 -620 2839
rect -678 2771 -620 2805
rect -678 2737 -666 2771
rect -632 2737 -620 2771
rect -678 2703 -620 2737
rect -678 2669 -666 2703
rect -632 2669 -620 2703
rect -678 2635 -620 2669
rect -678 2601 -666 2635
rect -632 2601 -620 2635
rect -678 2567 -620 2601
rect -678 2533 -666 2567
rect -632 2533 -620 2567
rect -678 2499 -620 2533
rect -678 2465 -666 2499
rect -632 2465 -620 2499
rect -678 2431 -620 2465
rect -678 2397 -666 2431
rect -632 2397 -620 2431
rect -678 2363 -620 2397
rect -678 2329 -666 2363
rect -632 2329 -620 2363
rect -678 2295 -620 2329
rect -678 2261 -666 2295
rect -632 2261 -620 2295
rect -678 2227 -620 2261
rect -678 2193 -666 2227
rect -632 2193 -620 2227
rect -678 2159 -620 2193
rect -678 2125 -666 2159
rect -632 2125 -620 2159
rect -678 2091 -620 2125
rect -678 2057 -666 2091
rect -632 2057 -620 2091
rect -678 2023 -620 2057
rect -678 1989 -666 2023
rect -632 1989 -620 2023
rect -678 1955 -620 1989
rect -678 1921 -666 1955
rect -632 1921 -620 1955
rect -678 1887 -620 1921
rect -678 1853 -666 1887
rect -632 1853 -620 1887
rect -678 1819 -620 1853
rect -678 1785 -666 1819
rect -632 1785 -620 1819
rect -678 1751 -620 1785
rect -678 1717 -666 1751
rect -632 1717 -620 1751
rect -678 1683 -620 1717
rect -678 1649 -666 1683
rect -632 1649 -620 1683
rect -678 1615 -620 1649
rect -678 1581 -666 1615
rect -632 1581 -620 1615
rect -678 1547 -620 1581
rect -678 1513 -666 1547
rect -632 1513 -620 1547
rect -678 1479 -620 1513
rect -678 1445 -666 1479
rect -632 1445 -620 1479
rect -678 1411 -620 1445
rect -678 1377 -666 1411
rect -632 1377 -620 1411
rect -678 1343 -620 1377
rect -678 1309 -666 1343
rect -632 1309 -620 1343
rect -678 1275 -620 1309
rect -678 1241 -666 1275
rect -632 1241 -620 1275
rect -678 1207 -620 1241
rect -678 1173 -666 1207
rect -632 1173 -620 1207
rect -678 1139 -620 1173
rect -678 1105 -666 1139
rect -632 1105 -620 1139
rect -678 1071 -620 1105
rect -678 1037 -666 1071
rect -632 1037 -620 1071
rect -678 1003 -620 1037
rect -678 969 -666 1003
rect -632 969 -620 1003
rect -678 935 -620 969
rect -678 901 -666 935
rect -632 901 -620 935
rect -678 867 -620 901
rect -678 833 -666 867
rect -632 833 -620 867
rect -678 799 -620 833
rect -678 765 -666 799
rect -632 765 -620 799
rect -678 731 -620 765
rect -678 697 -666 731
rect -632 697 -620 731
rect -678 663 -620 697
rect -678 629 -666 663
rect -632 629 -620 663
rect -678 595 -620 629
rect -678 561 -666 595
rect -632 561 -620 595
rect -678 527 -620 561
rect -678 493 -666 527
rect -632 493 -620 527
rect -678 459 -620 493
rect -678 425 -666 459
rect -632 425 -620 459
rect -678 391 -620 425
rect -678 357 -666 391
rect -632 357 -620 391
rect -678 323 -620 357
rect -678 289 -666 323
rect -632 289 -620 323
rect -678 255 -620 289
rect -678 221 -666 255
rect -632 221 -620 255
rect -678 187 -620 221
rect -678 153 -666 187
rect -632 153 -620 187
rect -678 119 -620 153
rect -678 85 -666 119
rect -632 85 -620 119
rect -678 51 -620 85
rect -678 17 -666 51
rect -632 17 -620 51
rect -678 -17 -620 17
rect -678 -51 -666 -17
rect -632 -51 -620 -17
rect -678 -85 -620 -51
rect -678 -119 -666 -85
rect -632 -119 -620 -85
rect -678 -153 -620 -119
rect -678 -187 -666 -153
rect -632 -187 -620 -153
rect -678 -221 -620 -187
rect -678 -255 -666 -221
rect -632 -255 -620 -221
rect -678 -289 -620 -255
rect -678 -323 -666 -289
rect -632 -323 -620 -289
rect -678 -357 -620 -323
rect -678 -391 -666 -357
rect -632 -391 -620 -357
rect -678 -425 -620 -391
rect -678 -459 -666 -425
rect -632 -459 -620 -425
rect -678 -493 -620 -459
rect -678 -527 -666 -493
rect -632 -527 -620 -493
rect -678 -561 -620 -527
rect -678 -595 -666 -561
rect -632 -595 -620 -561
rect -678 -629 -620 -595
rect -678 -663 -666 -629
rect -632 -663 -620 -629
rect -678 -697 -620 -663
rect -678 -731 -666 -697
rect -632 -731 -620 -697
rect -678 -765 -620 -731
rect -678 -799 -666 -765
rect -632 -799 -620 -765
rect -678 -833 -620 -799
rect -678 -867 -666 -833
rect -632 -867 -620 -833
rect -678 -901 -620 -867
rect -678 -935 -666 -901
rect -632 -935 -620 -901
rect -678 -969 -620 -935
rect -678 -1003 -666 -969
rect -632 -1003 -620 -969
rect -678 -1037 -620 -1003
rect -678 -1071 -666 -1037
rect -632 -1071 -620 -1037
rect -678 -1105 -620 -1071
rect -678 -1139 -666 -1105
rect -632 -1139 -620 -1105
rect -678 -1173 -620 -1139
rect -678 -1207 -666 -1173
rect -632 -1207 -620 -1173
rect -678 -1241 -620 -1207
rect -678 -1275 -666 -1241
rect -632 -1275 -620 -1241
rect -678 -1309 -620 -1275
rect -678 -1343 -666 -1309
rect -632 -1343 -620 -1309
rect -678 -1377 -620 -1343
rect -678 -1411 -666 -1377
rect -632 -1411 -620 -1377
rect -678 -1445 -620 -1411
rect -678 -1479 -666 -1445
rect -632 -1479 -620 -1445
rect -678 -1513 -620 -1479
rect -678 -1547 -666 -1513
rect -632 -1547 -620 -1513
rect -678 -1581 -620 -1547
rect -678 -1615 -666 -1581
rect -632 -1615 -620 -1581
rect -678 -1649 -620 -1615
rect -678 -1683 -666 -1649
rect -632 -1683 -620 -1649
rect -678 -1717 -620 -1683
rect -678 -1751 -666 -1717
rect -632 -1751 -620 -1717
rect -678 -1785 -620 -1751
rect -678 -1819 -666 -1785
rect -632 -1819 -620 -1785
rect -678 -1853 -620 -1819
rect -678 -1887 -666 -1853
rect -632 -1887 -620 -1853
rect -678 -1921 -620 -1887
rect -678 -1955 -666 -1921
rect -632 -1955 -620 -1921
rect -678 -1989 -620 -1955
rect -678 -2023 -666 -1989
rect -632 -2023 -620 -1989
rect -678 -2057 -620 -2023
rect -678 -2091 -666 -2057
rect -632 -2091 -620 -2057
rect -678 -2125 -620 -2091
rect -678 -2159 -666 -2125
rect -632 -2159 -620 -2125
rect -678 -2193 -620 -2159
rect -678 -2227 -666 -2193
rect -632 -2227 -620 -2193
rect -678 -2261 -620 -2227
rect -678 -2295 -666 -2261
rect -632 -2295 -620 -2261
rect -678 -2329 -620 -2295
rect -678 -2363 -666 -2329
rect -632 -2363 -620 -2329
rect -678 -2397 -620 -2363
rect -678 -2431 -666 -2397
rect -632 -2431 -620 -2397
rect -678 -2465 -620 -2431
rect -678 -2499 -666 -2465
rect -632 -2499 -620 -2465
rect -678 -2533 -620 -2499
rect -678 -2567 -666 -2533
rect -632 -2567 -620 -2533
rect -678 -2601 -620 -2567
rect -678 -2635 -666 -2601
rect -632 -2635 -620 -2601
rect -678 -2669 -620 -2635
rect -678 -2703 -666 -2669
rect -632 -2703 -620 -2669
rect -678 -2737 -620 -2703
rect -678 -2771 -666 -2737
rect -632 -2771 -620 -2737
rect -678 -2805 -620 -2771
rect -678 -2839 -666 -2805
rect -632 -2839 -620 -2805
rect -678 -2873 -620 -2839
rect -678 -2907 -666 -2873
rect -632 -2907 -620 -2873
rect -678 -2941 -620 -2907
rect -678 -2975 -666 -2941
rect -632 -2975 -620 -2941
rect -678 -3009 -620 -2975
rect -678 -3043 -666 -3009
rect -632 -3043 -620 -3009
rect -678 -3077 -620 -3043
rect -678 -3111 -666 -3077
rect -632 -3111 -620 -3077
rect -678 -3145 -620 -3111
rect -678 -3179 -666 -3145
rect -632 -3179 -620 -3145
rect -678 -3213 -620 -3179
rect -678 -3247 -666 -3213
rect -632 -3247 -620 -3213
rect -678 -3281 -620 -3247
rect -678 -3315 -666 -3281
rect -632 -3315 -620 -3281
rect -678 -3349 -620 -3315
rect -678 -3383 -666 -3349
rect -632 -3383 -620 -3349
rect -678 -3417 -620 -3383
rect -678 -3451 -666 -3417
rect -632 -3451 -620 -3417
rect -678 -3485 -620 -3451
rect -678 -3519 -666 -3485
rect -632 -3519 -620 -3485
rect -678 -3553 -620 -3519
rect -678 -3587 -666 -3553
rect -632 -3587 -620 -3553
rect -678 -3621 -620 -3587
rect -678 -3655 -666 -3621
rect -632 -3655 -620 -3621
rect -678 -3689 -620 -3655
rect -678 -3723 -666 -3689
rect -632 -3723 -620 -3689
rect -678 -3757 -620 -3723
rect -678 -3791 -666 -3757
rect -632 -3791 -620 -3757
rect -678 -3825 -620 -3791
rect -678 -3859 -666 -3825
rect -632 -3859 -620 -3825
rect -678 -3893 -620 -3859
rect -678 -3927 -666 -3893
rect -632 -3927 -620 -3893
rect -678 -3961 -620 -3927
rect -678 -3995 -666 -3961
rect -632 -3995 -620 -3961
rect -678 -4029 -620 -3995
rect -678 -4063 -666 -4029
rect -632 -4063 -620 -4029
rect -678 -4097 -620 -4063
rect -678 -4131 -666 -4097
rect -632 -4131 -620 -4097
rect -678 -4165 -620 -4131
rect -678 -4199 -666 -4165
rect -632 -4199 -620 -4165
rect -678 -4233 -620 -4199
rect -678 -4267 -666 -4233
rect -632 -4267 -620 -4233
rect -678 -4301 -620 -4267
rect -678 -4335 -666 -4301
rect -632 -4335 -620 -4301
rect -678 -4369 -620 -4335
rect -678 -4403 -666 -4369
rect -632 -4403 -620 -4369
rect -678 -4437 -620 -4403
rect -678 -4471 -666 -4437
rect -632 -4471 -620 -4437
rect -678 -4505 -620 -4471
rect -678 -4539 -666 -4505
rect -632 -4539 -620 -4505
rect -678 -4573 -620 -4539
rect -678 -4607 -666 -4573
rect -632 -4607 -620 -4573
rect -678 -4641 -620 -4607
rect -678 -4675 -666 -4641
rect -632 -4675 -620 -4641
rect -678 -4709 -620 -4675
rect -678 -4743 -666 -4709
rect -632 -4743 -620 -4709
rect -678 -4777 -620 -4743
rect -678 -4811 -666 -4777
rect -632 -4811 -620 -4777
rect -678 -4845 -620 -4811
rect -678 -4879 -666 -4845
rect -632 -4879 -620 -4845
rect -678 -4913 -620 -4879
rect -678 -4947 -666 -4913
rect -632 -4947 -620 -4913
rect -678 -4981 -620 -4947
rect -678 -5015 -666 -4981
rect -632 -5015 -620 -4981
rect -678 -5049 -620 -5015
rect -678 -5083 -666 -5049
rect -632 -5083 -620 -5049
rect -678 -5117 -620 -5083
rect -678 -5151 -666 -5117
rect -632 -5151 -620 -5117
rect -678 -5185 -620 -5151
rect -678 -5219 -666 -5185
rect -632 -5219 -620 -5185
rect -678 -5253 -620 -5219
rect -678 -5287 -666 -5253
rect -632 -5287 -620 -5253
rect -678 -5321 -620 -5287
rect -678 -5355 -666 -5321
rect -632 -5355 -620 -5321
rect -678 -5389 -620 -5355
rect -678 -5423 -666 -5389
rect -632 -5423 -620 -5389
rect -678 -5457 -620 -5423
rect -678 -5491 -666 -5457
rect -632 -5491 -620 -5457
rect -678 -5525 -620 -5491
rect -678 -5559 -666 -5525
rect -632 -5559 -620 -5525
rect -678 -5593 -620 -5559
rect -678 -5627 -666 -5593
rect -632 -5627 -620 -5593
rect -678 -5661 -620 -5627
rect -678 -5695 -666 -5661
rect -632 -5695 -620 -5661
rect -678 -5729 -620 -5695
rect -678 -5763 -666 -5729
rect -632 -5763 -620 -5729
rect -678 -5797 -620 -5763
rect -678 -5831 -666 -5797
rect -632 -5831 -620 -5797
rect -678 -5865 -620 -5831
rect -678 -5899 -666 -5865
rect -632 -5899 -620 -5865
rect -678 -5933 -620 -5899
rect -678 -5967 -666 -5933
rect -632 -5967 -620 -5933
rect -678 -6001 -620 -5967
rect -678 -6035 -666 -6001
rect -632 -6035 -620 -6001
rect -678 -6069 -620 -6035
rect -678 -6103 -666 -6069
rect -632 -6103 -620 -6069
rect -678 -6137 -620 -6103
rect -678 -6171 -666 -6137
rect -632 -6171 -620 -6137
rect -678 -6205 -620 -6171
rect -678 -6239 -666 -6205
rect -632 -6239 -620 -6205
rect -678 -6273 -620 -6239
rect -678 -6307 -666 -6273
rect -632 -6307 -620 -6273
rect -678 -6341 -620 -6307
rect -678 -6375 -666 -6341
rect -632 -6375 -620 -6341
rect -678 -6409 -620 -6375
rect -678 -6443 -666 -6409
rect -632 -6443 -620 -6409
rect -678 -6477 -620 -6443
rect -678 -6511 -666 -6477
rect -632 -6511 -620 -6477
rect -678 -6545 -620 -6511
rect -678 -6579 -666 -6545
rect -632 -6579 -620 -6545
rect -678 -6613 -620 -6579
rect -678 -6647 -666 -6613
rect -632 -6647 -620 -6613
rect -678 -6681 -620 -6647
rect -678 -6715 -666 -6681
rect -632 -6715 -620 -6681
rect -678 -6749 -620 -6715
rect -678 -6783 -666 -6749
rect -632 -6783 -620 -6749
rect -678 -6817 -620 -6783
rect -678 -6851 -666 -6817
rect -632 -6851 -620 -6817
rect -678 -6885 -620 -6851
rect -678 -6919 -666 -6885
rect -632 -6919 -620 -6885
rect -678 -6953 -620 -6919
rect -678 -6987 -666 -6953
rect -632 -6987 -620 -6953
rect -678 -7021 -620 -6987
rect -678 -7055 -666 -7021
rect -632 -7055 -620 -7021
rect -678 -7089 -620 -7055
rect -678 -7123 -666 -7089
rect -632 -7123 -620 -7089
rect -678 -7157 -620 -7123
rect -678 -7191 -666 -7157
rect -632 -7191 -620 -7157
rect -678 -7225 -620 -7191
rect -678 -7259 -666 -7225
rect -632 -7259 -620 -7225
rect -678 -7293 -620 -7259
rect -678 -7327 -666 -7293
rect -632 -7327 -620 -7293
rect -678 -7361 -620 -7327
rect -678 -7395 -666 -7361
rect -632 -7395 -620 -7361
rect -678 -7429 -620 -7395
rect -678 -7463 -666 -7429
rect -632 -7463 -620 -7429
rect -678 -7497 -620 -7463
rect -678 -7531 -666 -7497
rect -632 -7531 -620 -7497
rect -678 -7565 -620 -7531
rect -678 -7599 -666 -7565
rect -632 -7599 -620 -7565
rect -678 -7633 -620 -7599
rect -678 -7667 -666 -7633
rect -632 -7667 -620 -7633
rect -678 -7701 -620 -7667
rect -678 -7735 -666 -7701
rect -632 -7735 -620 -7701
rect -678 -7769 -620 -7735
rect -678 -7803 -666 -7769
rect -632 -7803 -620 -7769
rect -678 -7837 -620 -7803
rect -678 -7871 -666 -7837
rect -632 -7871 -620 -7837
rect -678 -7905 -620 -7871
rect -678 -7939 -666 -7905
rect -632 -7939 -620 -7905
rect -678 -7973 -620 -7939
rect -678 -8007 -666 -7973
rect -632 -8007 -620 -7973
rect -678 -8041 -620 -8007
rect -678 -8075 -666 -8041
rect -632 -8075 -620 -8041
rect -678 -8109 -620 -8075
rect -678 -8143 -666 -8109
rect -632 -8143 -620 -8109
rect -678 -8177 -620 -8143
rect -678 -8211 -666 -8177
rect -632 -8211 -620 -8177
rect -678 -8245 -620 -8211
rect -678 -8279 -666 -8245
rect -632 -8279 -620 -8245
rect -678 -8313 -620 -8279
rect -678 -8347 -666 -8313
rect -632 -8347 -620 -8313
rect -678 -8381 -620 -8347
rect -678 -8415 -666 -8381
rect -632 -8415 -620 -8381
rect -678 -8449 -620 -8415
rect -678 -8483 -666 -8449
rect -632 -8483 -620 -8449
rect -678 -8517 -620 -8483
rect -678 -8551 -666 -8517
rect -632 -8551 -620 -8517
rect -678 -8585 -620 -8551
rect -678 -8619 -666 -8585
rect -632 -8619 -620 -8585
rect -678 -8653 -620 -8619
rect -678 -8687 -666 -8653
rect -632 -8687 -620 -8653
rect -678 -8721 -620 -8687
rect -678 -8755 -666 -8721
rect -632 -8755 -620 -8721
rect -678 -8789 -620 -8755
rect -678 -8823 -666 -8789
rect -632 -8823 -620 -8789
rect -678 -8857 -620 -8823
rect -678 -8891 -666 -8857
rect -632 -8891 -620 -8857
rect -678 -8925 -620 -8891
rect -678 -8959 -666 -8925
rect -632 -8959 -620 -8925
rect -678 -8993 -620 -8959
rect -678 -9027 -666 -8993
rect -632 -9027 -620 -8993
rect -678 -9061 -620 -9027
rect -678 -9095 -666 -9061
rect -632 -9095 -620 -9061
rect -678 -9129 -620 -9095
rect -678 -9163 -666 -9129
rect -632 -9163 -620 -9129
rect -678 -9197 -620 -9163
rect -678 -9231 -666 -9197
rect -632 -9231 -620 -9197
rect -678 -9265 -620 -9231
rect -678 -9299 -666 -9265
rect -632 -9299 -620 -9265
rect -678 -9333 -620 -9299
rect -678 -9367 -666 -9333
rect -632 -9367 -620 -9333
rect -678 -9401 -620 -9367
rect -678 -9435 -666 -9401
rect -632 -9435 -620 -9401
rect -678 -9469 -620 -9435
rect -678 -9503 -666 -9469
rect -632 -9503 -620 -9469
rect -678 -9537 -620 -9503
rect -678 -9571 -666 -9537
rect -632 -9571 -620 -9537
rect -678 -9600 -620 -9571
rect -560 9571 -502 9600
rect -560 9537 -548 9571
rect -514 9537 -502 9571
rect -560 9503 -502 9537
rect -560 9469 -548 9503
rect -514 9469 -502 9503
rect -560 9435 -502 9469
rect -560 9401 -548 9435
rect -514 9401 -502 9435
rect -560 9367 -502 9401
rect -560 9333 -548 9367
rect -514 9333 -502 9367
rect -560 9299 -502 9333
rect -560 9265 -548 9299
rect -514 9265 -502 9299
rect -560 9231 -502 9265
rect -560 9197 -548 9231
rect -514 9197 -502 9231
rect -560 9163 -502 9197
rect -560 9129 -548 9163
rect -514 9129 -502 9163
rect -560 9095 -502 9129
rect -560 9061 -548 9095
rect -514 9061 -502 9095
rect -560 9027 -502 9061
rect -560 8993 -548 9027
rect -514 8993 -502 9027
rect -560 8959 -502 8993
rect -560 8925 -548 8959
rect -514 8925 -502 8959
rect -560 8891 -502 8925
rect -560 8857 -548 8891
rect -514 8857 -502 8891
rect -560 8823 -502 8857
rect -560 8789 -548 8823
rect -514 8789 -502 8823
rect -560 8755 -502 8789
rect -560 8721 -548 8755
rect -514 8721 -502 8755
rect -560 8687 -502 8721
rect -560 8653 -548 8687
rect -514 8653 -502 8687
rect -560 8619 -502 8653
rect -560 8585 -548 8619
rect -514 8585 -502 8619
rect -560 8551 -502 8585
rect -560 8517 -548 8551
rect -514 8517 -502 8551
rect -560 8483 -502 8517
rect -560 8449 -548 8483
rect -514 8449 -502 8483
rect -560 8415 -502 8449
rect -560 8381 -548 8415
rect -514 8381 -502 8415
rect -560 8347 -502 8381
rect -560 8313 -548 8347
rect -514 8313 -502 8347
rect -560 8279 -502 8313
rect -560 8245 -548 8279
rect -514 8245 -502 8279
rect -560 8211 -502 8245
rect -560 8177 -548 8211
rect -514 8177 -502 8211
rect -560 8143 -502 8177
rect -560 8109 -548 8143
rect -514 8109 -502 8143
rect -560 8075 -502 8109
rect -560 8041 -548 8075
rect -514 8041 -502 8075
rect -560 8007 -502 8041
rect -560 7973 -548 8007
rect -514 7973 -502 8007
rect -560 7939 -502 7973
rect -560 7905 -548 7939
rect -514 7905 -502 7939
rect -560 7871 -502 7905
rect -560 7837 -548 7871
rect -514 7837 -502 7871
rect -560 7803 -502 7837
rect -560 7769 -548 7803
rect -514 7769 -502 7803
rect -560 7735 -502 7769
rect -560 7701 -548 7735
rect -514 7701 -502 7735
rect -560 7667 -502 7701
rect -560 7633 -548 7667
rect -514 7633 -502 7667
rect -560 7599 -502 7633
rect -560 7565 -548 7599
rect -514 7565 -502 7599
rect -560 7531 -502 7565
rect -560 7497 -548 7531
rect -514 7497 -502 7531
rect -560 7463 -502 7497
rect -560 7429 -548 7463
rect -514 7429 -502 7463
rect -560 7395 -502 7429
rect -560 7361 -548 7395
rect -514 7361 -502 7395
rect -560 7327 -502 7361
rect -560 7293 -548 7327
rect -514 7293 -502 7327
rect -560 7259 -502 7293
rect -560 7225 -548 7259
rect -514 7225 -502 7259
rect -560 7191 -502 7225
rect -560 7157 -548 7191
rect -514 7157 -502 7191
rect -560 7123 -502 7157
rect -560 7089 -548 7123
rect -514 7089 -502 7123
rect -560 7055 -502 7089
rect -560 7021 -548 7055
rect -514 7021 -502 7055
rect -560 6987 -502 7021
rect -560 6953 -548 6987
rect -514 6953 -502 6987
rect -560 6919 -502 6953
rect -560 6885 -548 6919
rect -514 6885 -502 6919
rect -560 6851 -502 6885
rect -560 6817 -548 6851
rect -514 6817 -502 6851
rect -560 6783 -502 6817
rect -560 6749 -548 6783
rect -514 6749 -502 6783
rect -560 6715 -502 6749
rect -560 6681 -548 6715
rect -514 6681 -502 6715
rect -560 6647 -502 6681
rect -560 6613 -548 6647
rect -514 6613 -502 6647
rect -560 6579 -502 6613
rect -560 6545 -548 6579
rect -514 6545 -502 6579
rect -560 6511 -502 6545
rect -560 6477 -548 6511
rect -514 6477 -502 6511
rect -560 6443 -502 6477
rect -560 6409 -548 6443
rect -514 6409 -502 6443
rect -560 6375 -502 6409
rect -560 6341 -548 6375
rect -514 6341 -502 6375
rect -560 6307 -502 6341
rect -560 6273 -548 6307
rect -514 6273 -502 6307
rect -560 6239 -502 6273
rect -560 6205 -548 6239
rect -514 6205 -502 6239
rect -560 6171 -502 6205
rect -560 6137 -548 6171
rect -514 6137 -502 6171
rect -560 6103 -502 6137
rect -560 6069 -548 6103
rect -514 6069 -502 6103
rect -560 6035 -502 6069
rect -560 6001 -548 6035
rect -514 6001 -502 6035
rect -560 5967 -502 6001
rect -560 5933 -548 5967
rect -514 5933 -502 5967
rect -560 5899 -502 5933
rect -560 5865 -548 5899
rect -514 5865 -502 5899
rect -560 5831 -502 5865
rect -560 5797 -548 5831
rect -514 5797 -502 5831
rect -560 5763 -502 5797
rect -560 5729 -548 5763
rect -514 5729 -502 5763
rect -560 5695 -502 5729
rect -560 5661 -548 5695
rect -514 5661 -502 5695
rect -560 5627 -502 5661
rect -560 5593 -548 5627
rect -514 5593 -502 5627
rect -560 5559 -502 5593
rect -560 5525 -548 5559
rect -514 5525 -502 5559
rect -560 5491 -502 5525
rect -560 5457 -548 5491
rect -514 5457 -502 5491
rect -560 5423 -502 5457
rect -560 5389 -548 5423
rect -514 5389 -502 5423
rect -560 5355 -502 5389
rect -560 5321 -548 5355
rect -514 5321 -502 5355
rect -560 5287 -502 5321
rect -560 5253 -548 5287
rect -514 5253 -502 5287
rect -560 5219 -502 5253
rect -560 5185 -548 5219
rect -514 5185 -502 5219
rect -560 5151 -502 5185
rect -560 5117 -548 5151
rect -514 5117 -502 5151
rect -560 5083 -502 5117
rect -560 5049 -548 5083
rect -514 5049 -502 5083
rect -560 5015 -502 5049
rect -560 4981 -548 5015
rect -514 4981 -502 5015
rect -560 4947 -502 4981
rect -560 4913 -548 4947
rect -514 4913 -502 4947
rect -560 4879 -502 4913
rect -560 4845 -548 4879
rect -514 4845 -502 4879
rect -560 4811 -502 4845
rect -560 4777 -548 4811
rect -514 4777 -502 4811
rect -560 4743 -502 4777
rect -560 4709 -548 4743
rect -514 4709 -502 4743
rect -560 4675 -502 4709
rect -560 4641 -548 4675
rect -514 4641 -502 4675
rect -560 4607 -502 4641
rect -560 4573 -548 4607
rect -514 4573 -502 4607
rect -560 4539 -502 4573
rect -560 4505 -548 4539
rect -514 4505 -502 4539
rect -560 4471 -502 4505
rect -560 4437 -548 4471
rect -514 4437 -502 4471
rect -560 4403 -502 4437
rect -560 4369 -548 4403
rect -514 4369 -502 4403
rect -560 4335 -502 4369
rect -560 4301 -548 4335
rect -514 4301 -502 4335
rect -560 4267 -502 4301
rect -560 4233 -548 4267
rect -514 4233 -502 4267
rect -560 4199 -502 4233
rect -560 4165 -548 4199
rect -514 4165 -502 4199
rect -560 4131 -502 4165
rect -560 4097 -548 4131
rect -514 4097 -502 4131
rect -560 4063 -502 4097
rect -560 4029 -548 4063
rect -514 4029 -502 4063
rect -560 3995 -502 4029
rect -560 3961 -548 3995
rect -514 3961 -502 3995
rect -560 3927 -502 3961
rect -560 3893 -548 3927
rect -514 3893 -502 3927
rect -560 3859 -502 3893
rect -560 3825 -548 3859
rect -514 3825 -502 3859
rect -560 3791 -502 3825
rect -560 3757 -548 3791
rect -514 3757 -502 3791
rect -560 3723 -502 3757
rect -560 3689 -548 3723
rect -514 3689 -502 3723
rect -560 3655 -502 3689
rect -560 3621 -548 3655
rect -514 3621 -502 3655
rect -560 3587 -502 3621
rect -560 3553 -548 3587
rect -514 3553 -502 3587
rect -560 3519 -502 3553
rect -560 3485 -548 3519
rect -514 3485 -502 3519
rect -560 3451 -502 3485
rect -560 3417 -548 3451
rect -514 3417 -502 3451
rect -560 3383 -502 3417
rect -560 3349 -548 3383
rect -514 3349 -502 3383
rect -560 3315 -502 3349
rect -560 3281 -548 3315
rect -514 3281 -502 3315
rect -560 3247 -502 3281
rect -560 3213 -548 3247
rect -514 3213 -502 3247
rect -560 3179 -502 3213
rect -560 3145 -548 3179
rect -514 3145 -502 3179
rect -560 3111 -502 3145
rect -560 3077 -548 3111
rect -514 3077 -502 3111
rect -560 3043 -502 3077
rect -560 3009 -548 3043
rect -514 3009 -502 3043
rect -560 2975 -502 3009
rect -560 2941 -548 2975
rect -514 2941 -502 2975
rect -560 2907 -502 2941
rect -560 2873 -548 2907
rect -514 2873 -502 2907
rect -560 2839 -502 2873
rect -560 2805 -548 2839
rect -514 2805 -502 2839
rect -560 2771 -502 2805
rect -560 2737 -548 2771
rect -514 2737 -502 2771
rect -560 2703 -502 2737
rect -560 2669 -548 2703
rect -514 2669 -502 2703
rect -560 2635 -502 2669
rect -560 2601 -548 2635
rect -514 2601 -502 2635
rect -560 2567 -502 2601
rect -560 2533 -548 2567
rect -514 2533 -502 2567
rect -560 2499 -502 2533
rect -560 2465 -548 2499
rect -514 2465 -502 2499
rect -560 2431 -502 2465
rect -560 2397 -548 2431
rect -514 2397 -502 2431
rect -560 2363 -502 2397
rect -560 2329 -548 2363
rect -514 2329 -502 2363
rect -560 2295 -502 2329
rect -560 2261 -548 2295
rect -514 2261 -502 2295
rect -560 2227 -502 2261
rect -560 2193 -548 2227
rect -514 2193 -502 2227
rect -560 2159 -502 2193
rect -560 2125 -548 2159
rect -514 2125 -502 2159
rect -560 2091 -502 2125
rect -560 2057 -548 2091
rect -514 2057 -502 2091
rect -560 2023 -502 2057
rect -560 1989 -548 2023
rect -514 1989 -502 2023
rect -560 1955 -502 1989
rect -560 1921 -548 1955
rect -514 1921 -502 1955
rect -560 1887 -502 1921
rect -560 1853 -548 1887
rect -514 1853 -502 1887
rect -560 1819 -502 1853
rect -560 1785 -548 1819
rect -514 1785 -502 1819
rect -560 1751 -502 1785
rect -560 1717 -548 1751
rect -514 1717 -502 1751
rect -560 1683 -502 1717
rect -560 1649 -548 1683
rect -514 1649 -502 1683
rect -560 1615 -502 1649
rect -560 1581 -548 1615
rect -514 1581 -502 1615
rect -560 1547 -502 1581
rect -560 1513 -548 1547
rect -514 1513 -502 1547
rect -560 1479 -502 1513
rect -560 1445 -548 1479
rect -514 1445 -502 1479
rect -560 1411 -502 1445
rect -560 1377 -548 1411
rect -514 1377 -502 1411
rect -560 1343 -502 1377
rect -560 1309 -548 1343
rect -514 1309 -502 1343
rect -560 1275 -502 1309
rect -560 1241 -548 1275
rect -514 1241 -502 1275
rect -560 1207 -502 1241
rect -560 1173 -548 1207
rect -514 1173 -502 1207
rect -560 1139 -502 1173
rect -560 1105 -548 1139
rect -514 1105 -502 1139
rect -560 1071 -502 1105
rect -560 1037 -548 1071
rect -514 1037 -502 1071
rect -560 1003 -502 1037
rect -560 969 -548 1003
rect -514 969 -502 1003
rect -560 935 -502 969
rect -560 901 -548 935
rect -514 901 -502 935
rect -560 867 -502 901
rect -560 833 -548 867
rect -514 833 -502 867
rect -560 799 -502 833
rect -560 765 -548 799
rect -514 765 -502 799
rect -560 731 -502 765
rect -560 697 -548 731
rect -514 697 -502 731
rect -560 663 -502 697
rect -560 629 -548 663
rect -514 629 -502 663
rect -560 595 -502 629
rect -560 561 -548 595
rect -514 561 -502 595
rect -560 527 -502 561
rect -560 493 -548 527
rect -514 493 -502 527
rect -560 459 -502 493
rect -560 425 -548 459
rect -514 425 -502 459
rect -560 391 -502 425
rect -560 357 -548 391
rect -514 357 -502 391
rect -560 323 -502 357
rect -560 289 -548 323
rect -514 289 -502 323
rect -560 255 -502 289
rect -560 221 -548 255
rect -514 221 -502 255
rect -560 187 -502 221
rect -560 153 -548 187
rect -514 153 -502 187
rect -560 119 -502 153
rect -560 85 -548 119
rect -514 85 -502 119
rect -560 51 -502 85
rect -560 17 -548 51
rect -514 17 -502 51
rect -560 -17 -502 17
rect -560 -51 -548 -17
rect -514 -51 -502 -17
rect -560 -85 -502 -51
rect -560 -119 -548 -85
rect -514 -119 -502 -85
rect -560 -153 -502 -119
rect -560 -187 -548 -153
rect -514 -187 -502 -153
rect -560 -221 -502 -187
rect -560 -255 -548 -221
rect -514 -255 -502 -221
rect -560 -289 -502 -255
rect -560 -323 -548 -289
rect -514 -323 -502 -289
rect -560 -357 -502 -323
rect -560 -391 -548 -357
rect -514 -391 -502 -357
rect -560 -425 -502 -391
rect -560 -459 -548 -425
rect -514 -459 -502 -425
rect -560 -493 -502 -459
rect -560 -527 -548 -493
rect -514 -527 -502 -493
rect -560 -561 -502 -527
rect -560 -595 -548 -561
rect -514 -595 -502 -561
rect -560 -629 -502 -595
rect -560 -663 -548 -629
rect -514 -663 -502 -629
rect -560 -697 -502 -663
rect -560 -731 -548 -697
rect -514 -731 -502 -697
rect -560 -765 -502 -731
rect -560 -799 -548 -765
rect -514 -799 -502 -765
rect -560 -833 -502 -799
rect -560 -867 -548 -833
rect -514 -867 -502 -833
rect -560 -901 -502 -867
rect -560 -935 -548 -901
rect -514 -935 -502 -901
rect -560 -969 -502 -935
rect -560 -1003 -548 -969
rect -514 -1003 -502 -969
rect -560 -1037 -502 -1003
rect -560 -1071 -548 -1037
rect -514 -1071 -502 -1037
rect -560 -1105 -502 -1071
rect -560 -1139 -548 -1105
rect -514 -1139 -502 -1105
rect -560 -1173 -502 -1139
rect -560 -1207 -548 -1173
rect -514 -1207 -502 -1173
rect -560 -1241 -502 -1207
rect -560 -1275 -548 -1241
rect -514 -1275 -502 -1241
rect -560 -1309 -502 -1275
rect -560 -1343 -548 -1309
rect -514 -1343 -502 -1309
rect -560 -1377 -502 -1343
rect -560 -1411 -548 -1377
rect -514 -1411 -502 -1377
rect -560 -1445 -502 -1411
rect -560 -1479 -548 -1445
rect -514 -1479 -502 -1445
rect -560 -1513 -502 -1479
rect -560 -1547 -548 -1513
rect -514 -1547 -502 -1513
rect -560 -1581 -502 -1547
rect -560 -1615 -548 -1581
rect -514 -1615 -502 -1581
rect -560 -1649 -502 -1615
rect -560 -1683 -548 -1649
rect -514 -1683 -502 -1649
rect -560 -1717 -502 -1683
rect -560 -1751 -548 -1717
rect -514 -1751 -502 -1717
rect -560 -1785 -502 -1751
rect -560 -1819 -548 -1785
rect -514 -1819 -502 -1785
rect -560 -1853 -502 -1819
rect -560 -1887 -548 -1853
rect -514 -1887 -502 -1853
rect -560 -1921 -502 -1887
rect -560 -1955 -548 -1921
rect -514 -1955 -502 -1921
rect -560 -1989 -502 -1955
rect -560 -2023 -548 -1989
rect -514 -2023 -502 -1989
rect -560 -2057 -502 -2023
rect -560 -2091 -548 -2057
rect -514 -2091 -502 -2057
rect -560 -2125 -502 -2091
rect -560 -2159 -548 -2125
rect -514 -2159 -502 -2125
rect -560 -2193 -502 -2159
rect -560 -2227 -548 -2193
rect -514 -2227 -502 -2193
rect -560 -2261 -502 -2227
rect -560 -2295 -548 -2261
rect -514 -2295 -502 -2261
rect -560 -2329 -502 -2295
rect -560 -2363 -548 -2329
rect -514 -2363 -502 -2329
rect -560 -2397 -502 -2363
rect -560 -2431 -548 -2397
rect -514 -2431 -502 -2397
rect -560 -2465 -502 -2431
rect -560 -2499 -548 -2465
rect -514 -2499 -502 -2465
rect -560 -2533 -502 -2499
rect -560 -2567 -548 -2533
rect -514 -2567 -502 -2533
rect -560 -2601 -502 -2567
rect -560 -2635 -548 -2601
rect -514 -2635 -502 -2601
rect -560 -2669 -502 -2635
rect -560 -2703 -548 -2669
rect -514 -2703 -502 -2669
rect -560 -2737 -502 -2703
rect -560 -2771 -548 -2737
rect -514 -2771 -502 -2737
rect -560 -2805 -502 -2771
rect -560 -2839 -548 -2805
rect -514 -2839 -502 -2805
rect -560 -2873 -502 -2839
rect -560 -2907 -548 -2873
rect -514 -2907 -502 -2873
rect -560 -2941 -502 -2907
rect -560 -2975 -548 -2941
rect -514 -2975 -502 -2941
rect -560 -3009 -502 -2975
rect -560 -3043 -548 -3009
rect -514 -3043 -502 -3009
rect -560 -3077 -502 -3043
rect -560 -3111 -548 -3077
rect -514 -3111 -502 -3077
rect -560 -3145 -502 -3111
rect -560 -3179 -548 -3145
rect -514 -3179 -502 -3145
rect -560 -3213 -502 -3179
rect -560 -3247 -548 -3213
rect -514 -3247 -502 -3213
rect -560 -3281 -502 -3247
rect -560 -3315 -548 -3281
rect -514 -3315 -502 -3281
rect -560 -3349 -502 -3315
rect -560 -3383 -548 -3349
rect -514 -3383 -502 -3349
rect -560 -3417 -502 -3383
rect -560 -3451 -548 -3417
rect -514 -3451 -502 -3417
rect -560 -3485 -502 -3451
rect -560 -3519 -548 -3485
rect -514 -3519 -502 -3485
rect -560 -3553 -502 -3519
rect -560 -3587 -548 -3553
rect -514 -3587 -502 -3553
rect -560 -3621 -502 -3587
rect -560 -3655 -548 -3621
rect -514 -3655 -502 -3621
rect -560 -3689 -502 -3655
rect -560 -3723 -548 -3689
rect -514 -3723 -502 -3689
rect -560 -3757 -502 -3723
rect -560 -3791 -548 -3757
rect -514 -3791 -502 -3757
rect -560 -3825 -502 -3791
rect -560 -3859 -548 -3825
rect -514 -3859 -502 -3825
rect -560 -3893 -502 -3859
rect -560 -3927 -548 -3893
rect -514 -3927 -502 -3893
rect -560 -3961 -502 -3927
rect -560 -3995 -548 -3961
rect -514 -3995 -502 -3961
rect -560 -4029 -502 -3995
rect -560 -4063 -548 -4029
rect -514 -4063 -502 -4029
rect -560 -4097 -502 -4063
rect -560 -4131 -548 -4097
rect -514 -4131 -502 -4097
rect -560 -4165 -502 -4131
rect -560 -4199 -548 -4165
rect -514 -4199 -502 -4165
rect -560 -4233 -502 -4199
rect -560 -4267 -548 -4233
rect -514 -4267 -502 -4233
rect -560 -4301 -502 -4267
rect -560 -4335 -548 -4301
rect -514 -4335 -502 -4301
rect -560 -4369 -502 -4335
rect -560 -4403 -548 -4369
rect -514 -4403 -502 -4369
rect -560 -4437 -502 -4403
rect -560 -4471 -548 -4437
rect -514 -4471 -502 -4437
rect -560 -4505 -502 -4471
rect -560 -4539 -548 -4505
rect -514 -4539 -502 -4505
rect -560 -4573 -502 -4539
rect -560 -4607 -548 -4573
rect -514 -4607 -502 -4573
rect -560 -4641 -502 -4607
rect -560 -4675 -548 -4641
rect -514 -4675 -502 -4641
rect -560 -4709 -502 -4675
rect -560 -4743 -548 -4709
rect -514 -4743 -502 -4709
rect -560 -4777 -502 -4743
rect -560 -4811 -548 -4777
rect -514 -4811 -502 -4777
rect -560 -4845 -502 -4811
rect -560 -4879 -548 -4845
rect -514 -4879 -502 -4845
rect -560 -4913 -502 -4879
rect -560 -4947 -548 -4913
rect -514 -4947 -502 -4913
rect -560 -4981 -502 -4947
rect -560 -5015 -548 -4981
rect -514 -5015 -502 -4981
rect -560 -5049 -502 -5015
rect -560 -5083 -548 -5049
rect -514 -5083 -502 -5049
rect -560 -5117 -502 -5083
rect -560 -5151 -548 -5117
rect -514 -5151 -502 -5117
rect -560 -5185 -502 -5151
rect -560 -5219 -548 -5185
rect -514 -5219 -502 -5185
rect -560 -5253 -502 -5219
rect -560 -5287 -548 -5253
rect -514 -5287 -502 -5253
rect -560 -5321 -502 -5287
rect -560 -5355 -548 -5321
rect -514 -5355 -502 -5321
rect -560 -5389 -502 -5355
rect -560 -5423 -548 -5389
rect -514 -5423 -502 -5389
rect -560 -5457 -502 -5423
rect -560 -5491 -548 -5457
rect -514 -5491 -502 -5457
rect -560 -5525 -502 -5491
rect -560 -5559 -548 -5525
rect -514 -5559 -502 -5525
rect -560 -5593 -502 -5559
rect -560 -5627 -548 -5593
rect -514 -5627 -502 -5593
rect -560 -5661 -502 -5627
rect -560 -5695 -548 -5661
rect -514 -5695 -502 -5661
rect -560 -5729 -502 -5695
rect -560 -5763 -548 -5729
rect -514 -5763 -502 -5729
rect -560 -5797 -502 -5763
rect -560 -5831 -548 -5797
rect -514 -5831 -502 -5797
rect -560 -5865 -502 -5831
rect -560 -5899 -548 -5865
rect -514 -5899 -502 -5865
rect -560 -5933 -502 -5899
rect -560 -5967 -548 -5933
rect -514 -5967 -502 -5933
rect -560 -6001 -502 -5967
rect -560 -6035 -548 -6001
rect -514 -6035 -502 -6001
rect -560 -6069 -502 -6035
rect -560 -6103 -548 -6069
rect -514 -6103 -502 -6069
rect -560 -6137 -502 -6103
rect -560 -6171 -548 -6137
rect -514 -6171 -502 -6137
rect -560 -6205 -502 -6171
rect -560 -6239 -548 -6205
rect -514 -6239 -502 -6205
rect -560 -6273 -502 -6239
rect -560 -6307 -548 -6273
rect -514 -6307 -502 -6273
rect -560 -6341 -502 -6307
rect -560 -6375 -548 -6341
rect -514 -6375 -502 -6341
rect -560 -6409 -502 -6375
rect -560 -6443 -548 -6409
rect -514 -6443 -502 -6409
rect -560 -6477 -502 -6443
rect -560 -6511 -548 -6477
rect -514 -6511 -502 -6477
rect -560 -6545 -502 -6511
rect -560 -6579 -548 -6545
rect -514 -6579 -502 -6545
rect -560 -6613 -502 -6579
rect -560 -6647 -548 -6613
rect -514 -6647 -502 -6613
rect -560 -6681 -502 -6647
rect -560 -6715 -548 -6681
rect -514 -6715 -502 -6681
rect -560 -6749 -502 -6715
rect -560 -6783 -548 -6749
rect -514 -6783 -502 -6749
rect -560 -6817 -502 -6783
rect -560 -6851 -548 -6817
rect -514 -6851 -502 -6817
rect -560 -6885 -502 -6851
rect -560 -6919 -548 -6885
rect -514 -6919 -502 -6885
rect -560 -6953 -502 -6919
rect -560 -6987 -548 -6953
rect -514 -6987 -502 -6953
rect -560 -7021 -502 -6987
rect -560 -7055 -548 -7021
rect -514 -7055 -502 -7021
rect -560 -7089 -502 -7055
rect -560 -7123 -548 -7089
rect -514 -7123 -502 -7089
rect -560 -7157 -502 -7123
rect -560 -7191 -548 -7157
rect -514 -7191 -502 -7157
rect -560 -7225 -502 -7191
rect -560 -7259 -548 -7225
rect -514 -7259 -502 -7225
rect -560 -7293 -502 -7259
rect -560 -7327 -548 -7293
rect -514 -7327 -502 -7293
rect -560 -7361 -502 -7327
rect -560 -7395 -548 -7361
rect -514 -7395 -502 -7361
rect -560 -7429 -502 -7395
rect -560 -7463 -548 -7429
rect -514 -7463 -502 -7429
rect -560 -7497 -502 -7463
rect -560 -7531 -548 -7497
rect -514 -7531 -502 -7497
rect -560 -7565 -502 -7531
rect -560 -7599 -548 -7565
rect -514 -7599 -502 -7565
rect -560 -7633 -502 -7599
rect -560 -7667 -548 -7633
rect -514 -7667 -502 -7633
rect -560 -7701 -502 -7667
rect -560 -7735 -548 -7701
rect -514 -7735 -502 -7701
rect -560 -7769 -502 -7735
rect -560 -7803 -548 -7769
rect -514 -7803 -502 -7769
rect -560 -7837 -502 -7803
rect -560 -7871 -548 -7837
rect -514 -7871 -502 -7837
rect -560 -7905 -502 -7871
rect -560 -7939 -548 -7905
rect -514 -7939 -502 -7905
rect -560 -7973 -502 -7939
rect -560 -8007 -548 -7973
rect -514 -8007 -502 -7973
rect -560 -8041 -502 -8007
rect -560 -8075 -548 -8041
rect -514 -8075 -502 -8041
rect -560 -8109 -502 -8075
rect -560 -8143 -548 -8109
rect -514 -8143 -502 -8109
rect -560 -8177 -502 -8143
rect -560 -8211 -548 -8177
rect -514 -8211 -502 -8177
rect -560 -8245 -502 -8211
rect -560 -8279 -548 -8245
rect -514 -8279 -502 -8245
rect -560 -8313 -502 -8279
rect -560 -8347 -548 -8313
rect -514 -8347 -502 -8313
rect -560 -8381 -502 -8347
rect -560 -8415 -548 -8381
rect -514 -8415 -502 -8381
rect -560 -8449 -502 -8415
rect -560 -8483 -548 -8449
rect -514 -8483 -502 -8449
rect -560 -8517 -502 -8483
rect -560 -8551 -548 -8517
rect -514 -8551 -502 -8517
rect -560 -8585 -502 -8551
rect -560 -8619 -548 -8585
rect -514 -8619 -502 -8585
rect -560 -8653 -502 -8619
rect -560 -8687 -548 -8653
rect -514 -8687 -502 -8653
rect -560 -8721 -502 -8687
rect -560 -8755 -548 -8721
rect -514 -8755 -502 -8721
rect -560 -8789 -502 -8755
rect -560 -8823 -548 -8789
rect -514 -8823 -502 -8789
rect -560 -8857 -502 -8823
rect -560 -8891 -548 -8857
rect -514 -8891 -502 -8857
rect -560 -8925 -502 -8891
rect -560 -8959 -548 -8925
rect -514 -8959 -502 -8925
rect -560 -8993 -502 -8959
rect -560 -9027 -548 -8993
rect -514 -9027 -502 -8993
rect -560 -9061 -502 -9027
rect -560 -9095 -548 -9061
rect -514 -9095 -502 -9061
rect -560 -9129 -502 -9095
rect -560 -9163 -548 -9129
rect -514 -9163 -502 -9129
rect -560 -9197 -502 -9163
rect -560 -9231 -548 -9197
rect -514 -9231 -502 -9197
rect -560 -9265 -502 -9231
rect -560 -9299 -548 -9265
rect -514 -9299 -502 -9265
rect -560 -9333 -502 -9299
rect -560 -9367 -548 -9333
rect -514 -9367 -502 -9333
rect -560 -9401 -502 -9367
rect -560 -9435 -548 -9401
rect -514 -9435 -502 -9401
rect -560 -9469 -502 -9435
rect -560 -9503 -548 -9469
rect -514 -9503 -502 -9469
rect -560 -9537 -502 -9503
rect -560 -9571 -548 -9537
rect -514 -9571 -502 -9537
rect -560 -9600 -502 -9571
rect -442 9571 -384 9600
rect -442 9537 -430 9571
rect -396 9537 -384 9571
rect -442 9503 -384 9537
rect -442 9469 -430 9503
rect -396 9469 -384 9503
rect -442 9435 -384 9469
rect -442 9401 -430 9435
rect -396 9401 -384 9435
rect -442 9367 -384 9401
rect -442 9333 -430 9367
rect -396 9333 -384 9367
rect -442 9299 -384 9333
rect -442 9265 -430 9299
rect -396 9265 -384 9299
rect -442 9231 -384 9265
rect -442 9197 -430 9231
rect -396 9197 -384 9231
rect -442 9163 -384 9197
rect -442 9129 -430 9163
rect -396 9129 -384 9163
rect -442 9095 -384 9129
rect -442 9061 -430 9095
rect -396 9061 -384 9095
rect -442 9027 -384 9061
rect -442 8993 -430 9027
rect -396 8993 -384 9027
rect -442 8959 -384 8993
rect -442 8925 -430 8959
rect -396 8925 -384 8959
rect -442 8891 -384 8925
rect -442 8857 -430 8891
rect -396 8857 -384 8891
rect -442 8823 -384 8857
rect -442 8789 -430 8823
rect -396 8789 -384 8823
rect -442 8755 -384 8789
rect -442 8721 -430 8755
rect -396 8721 -384 8755
rect -442 8687 -384 8721
rect -442 8653 -430 8687
rect -396 8653 -384 8687
rect -442 8619 -384 8653
rect -442 8585 -430 8619
rect -396 8585 -384 8619
rect -442 8551 -384 8585
rect -442 8517 -430 8551
rect -396 8517 -384 8551
rect -442 8483 -384 8517
rect -442 8449 -430 8483
rect -396 8449 -384 8483
rect -442 8415 -384 8449
rect -442 8381 -430 8415
rect -396 8381 -384 8415
rect -442 8347 -384 8381
rect -442 8313 -430 8347
rect -396 8313 -384 8347
rect -442 8279 -384 8313
rect -442 8245 -430 8279
rect -396 8245 -384 8279
rect -442 8211 -384 8245
rect -442 8177 -430 8211
rect -396 8177 -384 8211
rect -442 8143 -384 8177
rect -442 8109 -430 8143
rect -396 8109 -384 8143
rect -442 8075 -384 8109
rect -442 8041 -430 8075
rect -396 8041 -384 8075
rect -442 8007 -384 8041
rect -442 7973 -430 8007
rect -396 7973 -384 8007
rect -442 7939 -384 7973
rect -442 7905 -430 7939
rect -396 7905 -384 7939
rect -442 7871 -384 7905
rect -442 7837 -430 7871
rect -396 7837 -384 7871
rect -442 7803 -384 7837
rect -442 7769 -430 7803
rect -396 7769 -384 7803
rect -442 7735 -384 7769
rect -442 7701 -430 7735
rect -396 7701 -384 7735
rect -442 7667 -384 7701
rect -442 7633 -430 7667
rect -396 7633 -384 7667
rect -442 7599 -384 7633
rect -442 7565 -430 7599
rect -396 7565 -384 7599
rect -442 7531 -384 7565
rect -442 7497 -430 7531
rect -396 7497 -384 7531
rect -442 7463 -384 7497
rect -442 7429 -430 7463
rect -396 7429 -384 7463
rect -442 7395 -384 7429
rect -442 7361 -430 7395
rect -396 7361 -384 7395
rect -442 7327 -384 7361
rect -442 7293 -430 7327
rect -396 7293 -384 7327
rect -442 7259 -384 7293
rect -442 7225 -430 7259
rect -396 7225 -384 7259
rect -442 7191 -384 7225
rect -442 7157 -430 7191
rect -396 7157 -384 7191
rect -442 7123 -384 7157
rect -442 7089 -430 7123
rect -396 7089 -384 7123
rect -442 7055 -384 7089
rect -442 7021 -430 7055
rect -396 7021 -384 7055
rect -442 6987 -384 7021
rect -442 6953 -430 6987
rect -396 6953 -384 6987
rect -442 6919 -384 6953
rect -442 6885 -430 6919
rect -396 6885 -384 6919
rect -442 6851 -384 6885
rect -442 6817 -430 6851
rect -396 6817 -384 6851
rect -442 6783 -384 6817
rect -442 6749 -430 6783
rect -396 6749 -384 6783
rect -442 6715 -384 6749
rect -442 6681 -430 6715
rect -396 6681 -384 6715
rect -442 6647 -384 6681
rect -442 6613 -430 6647
rect -396 6613 -384 6647
rect -442 6579 -384 6613
rect -442 6545 -430 6579
rect -396 6545 -384 6579
rect -442 6511 -384 6545
rect -442 6477 -430 6511
rect -396 6477 -384 6511
rect -442 6443 -384 6477
rect -442 6409 -430 6443
rect -396 6409 -384 6443
rect -442 6375 -384 6409
rect -442 6341 -430 6375
rect -396 6341 -384 6375
rect -442 6307 -384 6341
rect -442 6273 -430 6307
rect -396 6273 -384 6307
rect -442 6239 -384 6273
rect -442 6205 -430 6239
rect -396 6205 -384 6239
rect -442 6171 -384 6205
rect -442 6137 -430 6171
rect -396 6137 -384 6171
rect -442 6103 -384 6137
rect -442 6069 -430 6103
rect -396 6069 -384 6103
rect -442 6035 -384 6069
rect -442 6001 -430 6035
rect -396 6001 -384 6035
rect -442 5967 -384 6001
rect -442 5933 -430 5967
rect -396 5933 -384 5967
rect -442 5899 -384 5933
rect -442 5865 -430 5899
rect -396 5865 -384 5899
rect -442 5831 -384 5865
rect -442 5797 -430 5831
rect -396 5797 -384 5831
rect -442 5763 -384 5797
rect -442 5729 -430 5763
rect -396 5729 -384 5763
rect -442 5695 -384 5729
rect -442 5661 -430 5695
rect -396 5661 -384 5695
rect -442 5627 -384 5661
rect -442 5593 -430 5627
rect -396 5593 -384 5627
rect -442 5559 -384 5593
rect -442 5525 -430 5559
rect -396 5525 -384 5559
rect -442 5491 -384 5525
rect -442 5457 -430 5491
rect -396 5457 -384 5491
rect -442 5423 -384 5457
rect -442 5389 -430 5423
rect -396 5389 -384 5423
rect -442 5355 -384 5389
rect -442 5321 -430 5355
rect -396 5321 -384 5355
rect -442 5287 -384 5321
rect -442 5253 -430 5287
rect -396 5253 -384 5287
rect -442 5219 -384 5253
rect -442 5185 -430 5219
rect -396 5185 -384 5219
rect -442 5151 -384 5185
rect -442 5117 -430 5151
rect -396 5117 -384 5151
rect -442 5083 -384 5117
rect -442 5049 -430 5083
rect -396 5049 -384 5083
rect -442 5015 -384 5049
rect -442 4981 -430 5015
rect -396 4981 -384 5015
rect -442 4947 -384 4981
rect -442 4913 -430 4947
rect -396 4913 -384 4947
rect -442 4879 -384 4913
rect -442 4845 -430 4879
rect -396 4845 -384 4879
rect -442 4811 -384 4845
rect -442 4777 -430 4811
rect -396 4777 -384 4811
rect -442 4743 -384 4777
rect -442 4709 -430 4743
rect -396 4709 -384 4743
rect -442 4675 -384 4709
rect -442 4641 -430 4675
rect -396 4641 -384 4675
rect -442 4607 -384 4641
rect -442 4573 -430 4607
rect -396 4573 -384 4607
rect -442 4539 -384 4573
rect -442 4505 -430 4539
rect -396 4505 -384 4539
rect -442 4471 -384 4505
rect -442 4437 -430 4471
rect -396 4437 -384 4471
rect -442 4403 -384 4437
rect -442 4369 -430 4403
rect -396 4369 -384 4403
rect -442 4335 -384 4369
rect -442 4301 -430 4335
rect -396 4301 -384 4335
rect -442 4267 -384 4301
rect -442 4233 -430 4267
rect -396 4233 -384 4267
rect -442 4199 -384 4233
rect -442 4165 -430 4199
rect -396 4165 -384 4199
rect -442 4131 -384 4165
rect -442 4097 -430 4131
rect -396 4097 -384 4131
rect -442 4063 -384 4097
rect -442 4029 -430 4063
rect -396 4029 -384 4063
rect -442 3995 -384 4029
rect -442 3961 -430 3995
rect -396 3961 -384 3995
rect -442 3927 -384 3961
rect -442 3893 -430 3927
rect -396 3893 -384 3927
rect -442 3859 -384 3893
rect -442 3825 -430 3859
rect -396 3825 -384 3859
rect -442 3791 -384 3825
rect -442 3757 -430 3791
rect -396 3757 -384 3791
rect -442 3723 -384 3757
rect -442 3689 -430 3723
rect -396 3689 -384 3723
rect -442 3655 -384 3689
rect -442 3621 -430 3655
rect -396 3621 -384 3655
rect -442 3587 -384 3621
rect -442 3553 -430 3587
rect -396 3553 -384 3587
rect -442 3519 -384 3553
rect -442 3485 -430 3519
rect -396 3485 -384 3519
rect -442 3451 -384 3485
rect -442 3417 -430 3451
rect -396 3417 -384 3451
rect -442 3383 -384 3417
rect -442 3349 -430 3383
rect -396 3349 -384 3383
rect -442 3315 -384 3349
rect -442 3281 -430 3315
rect -396 3281 -384 3315
rect -442 3247 -384 3281
rect -442 3213 -430 3247
rect -396 3213 -384 3247
rect -442 3179 -384 3213
rect -442 3145 -430 3179
rect -396 3145 -384 3179
rect -442 3111 -384 3145
rect -442 3077 -430 3111
rect -396 3077 -384 3111
rect -442 3043 -384 3077
rect -442 3009 -430 3043
rect -396 3009 -384 3043
rect -442 2975 -384 3009
rect -442 2941 -430 2975
rect -396 2941 -384 2975
rect -442 2907 -384 2941
rect -442 2873 -430 2907
rect -396 2873 -384 2907
rect -442 2839 -384 2873
rect -442 2805 -430 2839
rect -396 2805 -384 2839
rect -442 2771 -384 2805
rect -442 2737 -430 2771
rect -396 2737 -384 2771
rect -442 2703 -384 2737
rect -442 2669 -430 2703
rect -396 2669 -384 2703
rect -442 2635 -384 2669
rect -442 2601 -430 2635
rect -396 2601 -384 2635
rect -442 2567 -384 2601
rect -442 2533 -430 2567
rect -396 2533 -384 2567
rect -442 2499 -384 2533
rect -442 2465 -430 2499
rect -396 2465 -384 2499
rect -442 2431 -384 2465
rect -442 2397 -430 2431
rect -396 2397 -384 2431
rect -442 2363 -384 2397
rect -442 2329 -430 2363
rect -396 2329 -384 2363
rect -442 2295 -384 2329
rect -442 2261 -430 2295
rect -396 2261 -384 2295
rect -442 2227 -384 2261
rect -442 2193 -430 2227
rect -396 2193 -384 2227
rect -442 2159 -384 2193
rect -442 2125 -430 2159
rect -396 2125 -384 2159
rect -442 2091 -384 2125
rect -442 2057 -430 2091
rect -396 2057 -384 2091
rect -442 2023 -384 2057
rect -442 1989 -430 2023
rect -396 1989 -384 2023
rect -442 1955 -384 1989
rect -442 1921 -430 1955
rect -396 1921 -384 1955
rect -442 1887 -384 1921
rect -442 1853 -430 1887
rect -396 1853 -384 1887
rect -442 1819 -384 1853
rect -442 1785 -430 1819
rect -396 1785 -384 1819
rect -442 1751 -384 1785
rect -442 1717 -430 1751
rect -396 1717 -384 1751
rect -442 1683 -384 1717
rect -442 1649 -430 1683
rect -396 1649 -384 1683
rect -442 1615 -384 1649
rect -442 1581 -430 1615
rect -396 1581 -384 1615
rect -442 1547 -384 1581
rect -442 1513 -430 1547
rect -396 1513 -384 1547
rect -442 1479 -384 1513
rect -442 1445 -430 1479
rect -396 1445 -384 1479
rect -442 1411 -384 1445
rect -442 1377 -430 1411
rect -396 1377 -384 1411
rect -442 1343 -384 1377
rect -442 1309 -430 1343
rect -396 1309 -384 1343
rect -442 1275 -384 1309
rect -442 1241 -430 1275
rect -396 1241 -384 1275
rect -442 1207 -384 1241
rect -442 1173 -430 1207
rect -396 1173 -384 1207
rect -442 1139 -384 1173
rect -442 1105 -430 1139
rect -396 1105 -384 1139
rect -442 1071 -384 1105
rect -442 1037 -430 1071
rect -396 1037 -384 1071
rect -442 1003 -384 1037
rect -442 969 -430 1003
rect -396 969 -384 1003
rect -442 935 -384 969
rect -442 901 -430 935
rect -396 901 -384 935
rect -442 867 -384 901
rect -442 833 -430 867
rect -396 833 -384 867
rect -442 799 -384 833
rect -442 765 -430 799
rect -396 765 -384 799
rect -442 731 -384 765
rect -442 697 -430 731
rect -396 697 -384 731
rect -442 663 -384 697
rect -442 629 -430 663
rect -396 629 -384 663
rect -442 595 -384 629
rect -442 561 -430 595
rect -396 561 -384 595
rect -442 527 -384 561
rect -442 493 -430 527
rect -396 493 -384 527
rect -442 459 -384 493
rect -442 425 -430 459
rect -396 425 -384 459
rect -442 391 -384 425
rect -442 357 -430 391
rect -396 357 -384 391
rect -442 323 -384 357
rect -442 289 -430 323
rect -396 289 -384 323
rect -442 255 -384 289
rect -442 221 -430 255
rect -396 221 -384 255
rect -442 187 -384 221
rect -442 153 -430 187
rect -396 153 -384 187
rect -442 119 -384 153
rect -442 85 -430 119
rect -396 85 -384 119
rect -442 51 -384 85
rect -442 17 -430 51
rect -396 17 -384 51
rect -442 -17 -384 17
rect -442 -51 -430 -17
rect -396 -51 -384 -17
rect -442 -85 -384 -51
rect -442 -119 -430 -85
rect -396 -119 -384 -85
rect -442 -153 -384 -119
rect -442 -187 -430 -153
rect -396 -187 -384 -153
rect -442 -221 -384 -187
rect -442 -255 -430 -221
rect -396 -255 -384 -221
rect -442 -289 -384 -255
rect -442 -323 -430 -289
rect -396 -323 -384 -289
rect -442 -357 -384 -323
rect -442 -391 -430 -357
rect -396 -391 -384 -357
rect -442 -425 -384 -391
rect -442 -459 -430 -425
rect -396 -459 -384 -425
rect -442 -493 -384 -459
rect -442 -527 -430 -493
rect -396 -527 -384 -493
rect -442 -561 -384 -527
rect -442 -595 -430 -561
rect -396 -595 -384 -561
rect -442 -629 -384 -595
rect -442 -663 -430 -629
rect -396 -663 -384 -629
rect -442 -697 -384 -663
rect -442 -731 -430 -697
rect -396 -731 -384 -697
rect -442 -765 -384 -731
rect -442 -799 -430 -765
rect -396 -799 -384 -765
rect -442 -833 -384 -799
rect -442 -867 -430 -833
rect -396 -867 -384 -833
rect -442 -901 -384 -867
rect -442 -935 -430 -901
rect -396 -935 -384 -901
rect -442 -969 -384 -935
rect -442 -1003 -430 -969
rect -396 -1003 -384 -969
rect -442 -1037 -384 -1003
rect -442 -1071 -430 -1037
rect -396 -1071 -384 -1037
rect -442 -1105 -384 -1071
rect -442 -1139 -430 -1105
rect -396 -1139 -384 -1105
rect -442 -1173 -384 -1139
rect -442 -1207 -430 -1173
rect -396 -1207 -384 -1173
rect -442 -1241 -384 -1207
rect -442 -1275 -430 -1241
rect -396 -1275 -384 -1241
rect -442 -1309 -384 -1275
rect -442 -1343 -430 -1309
rect -396 -1343 -384 -1309
rect -442 -1377 -384 -1343
rect -442 -1411 -430 -1377
rect -396 -1411 -384 -1377
rect -442 -1445 -384 -1411
rect -442 -1479 -430 -1445
rect -396 -1479 -384 -1445
rect -442 -1513 -384 -1479
rect -442 -1547 -430 -1513
rect -396 -1547 -384 -1513
rect -442 -1581 -384 -1547
rect -442 -1615 -430 -1581
rect -396 -1615 -384 -1581
rect -442 -1649 -384 -1615
rect -442 -1683 -430 -1649
rect -396 -1683 -384 -1649
rect -442 -1717 -384 -1683
rect -442 -1751 -430 -1717
rect -396 -1751 -384 -1717
rect -442 -1785 -384 -1751
rect -442 -1819 -430 -1785
rect -396 -1819 -384 -1785
rect -442 -1853 -384 -1819
rect -442 -1887 -430 -1853
rect -396 -1887 -384 -1853
rect -442 -1921 -384 -1887
rect -442 -1955 -430 -1921
rect -396 -1955 -384 -1921
rect -442 -1989 -384 -1955
rect -442 -2023 -430 -1989
rect -396 -2023 -384 -1989
rect -442 -2057 -384 -2023
rect -442 -2091 -430 -2057
rect -396 -2091 -384 -2057
rect -442 -2125 -384 -2091
rect -442 -2159 -430 -2125
rect -396 -2159 -384 -2125
rect -442 -2193 -384 -2159
rect -442 -2227 -430 -2193
rect -396 -2227 -384 -2193
rect -442 -2261 -384 -2227
rect -442 -2295 -430 -2261
rect -396 -2295 -384 -2261
rect -442 -2329 -384 -2295
rect -442 -2363 -430 -2329
rect -396 -2363 -384 -2329
rect -442 -2397 -384 -2363
rect -442 -2431 -430 -2397
rect -396 -2431 -384 -2397
rect -442 -2465 -384 -2431
rect -442 -2499 -430 -2465
rect -396 -2499 -384 -2465
rect -442 -2533 -384 -2499
rect -442 -2567 -430 -2533
rect -396 -2567 -384 -2533
rect -442 -2601 -384 -2567
rect -442 -2635 -430 -2601
rect -396 -2635 -384 -2601
rect -442 -2669 -384 -2635
rect -442 -2703 -430 -2669
rect -396 -2703 -384 -2669
rect -442 -2737 -384 -2703
rect -442 -2771 -430 -2737
rect -396 -2771 -384 -2737
rect -442 -2805 -384 -2771
rect -442 -2839 -430 -2805
rect -396 -2839 -384 -2805
rect -442 -2873 -384 -2839
rect -442 -2907 -430 -2873
rect -396 -2907 -384 -2873
rect -442 -2941 -384 -2907
rect -442 -2975 -430 -2941
rect -396 -2975 -384 -2941
rect -442 -3009 -384 -2975
rect -442 -3043 -430 -3009
rect -396 -3043 -384 -3009
rect -442 -3077 -384 -3043
rect -442 -3111 -430 -3077
rect -396 -3111 -384 -3077
rect -442 -3145 -384 -3111
rect -442 -3179 -430 -3145
rect -396 -3179 -384 -3145
rect -442 -3213 -384 -3179
rect -442 -3247 -430 -3213
rect -396 -3247 -384 -3213
rect -442 -3281 -384 -3247
rect -442 -3315 -430 -3281
rect -396 -3315 -384 -3281
rect -442 -3349 -384 -3315
rect -442 -3383 -430 -3349
rect -396 -3383 -384 -3349
rect -442 -3417 -384 -3383
rect -442 -3451 -430 -3417
rect -396 -3451 -384 -3417
rect -442 -3485 -384 -3451
rect -442 -3519 -430 -3485
rect -396 -3519 -384 -3485
rect -442 -3553 -384 -3519
rect -442 -3587 -430 -3553
rect -396 -3587 -384 -3553
rect -442 -3621 -384 -3587
rect -442 -3655 -430 -3621
rect -396 -3655 -384 -3621
rect -442 -3689 -384 -3655
rect -442 -3723 -430 -3689
rect -396 -3723 -384 -3689
rect -442 -3757 -384 -3723
rect -442 -3791 -430 -3757
rect -396 -3791 -384 -3757
rect -442 -3825 -384 -3791
rect -442 -3859 -430 -3825
rect -396 -3859 -384 -3825
rect -442 -3893 -384 -3859
rect -442 -3927 -430 -3893
rect -396 -3927 -384 -3893
rect -442 -3961 -384 -3927
rect -442 -3995 -430 -3961
rect -396 -3995 -384 -3961
rect -442 -4029 -384 -3995
rect -442 -4063 -430 -4029
rect -396 -4063 -384 -4029
rect -442 -4097 -384 -4063
rect -442 -4131 -430 -4097
rect -396 -4131 -384 -4097
rect -442 -4165 -384 -4131
rect -442 -4199 -430 -4165
rect -396 -4199 -384 -4165
rect -442 -4233 -384 -4199
rect -442 -4267 -430 -4233
rect -396 -4267 -384 -4233
rect -442 -4301 -384 -4267
rect -442 -4335 -430 -4301
rect -396 -4335 -384 -4301
rect -442 -4369 -384 -4335
rect -442 -4403 -430 -4369
rect -396 -4403 -384 -4369
rect -442 -4437 -384 -4403
rect -442 -4471 -430 -4437
rect -396 -4471 -384 -4437
rect -442 -4505 -384 -4471
rect -442 -4539 -430 -4505
rect -396 -4539 -384 -4505
rect -442 -4573 -384 -4539
rect -442 -4607 -430 -4573
rect -396 -4607 -384 -4573
rect -442 -4641 -384 -4607
rect -442 -4675 -430 -4641
rect -396 -4675 -384 -4641
rect -442 -4709 -384 -4675
rect -442 -4743 -430 -4709
rect -396 -4743 -384 -4709
rect -442 -4777 -384 -4743
rect -442 -4811 -430 -4777
rect -396 -4811 -384 -4777
rect -442 -4845 -384 -4811
rect -442 -4879 -430 -4845
rect -396 -4879 -384 -4845
rect -442 -4913 -384 -4879
rect -442 -4947 -430 -4913
rect -396 -4947 -384 -4913
rect -442 -4981 -384 -4947
rect -442 -5015 -430 -4981
rect -396 -5015 -384 -4981
rect -442 -5049 -384 -5015
rect -442 -5083 -430 -5049
rect -396 -5083 -384 -5049
rect -442 -5117 -384 -5083
rect -442 -5151 -430 -5117
rect -396 -5151 -384 -5117
rect -442 -5185 -384 -5151
rect -442 -5219 -430 -5185
rect -396 -5219 -384 -5185
rect -442 -5253 -384 -5219
rect -442 -5287 -430 -5253
rect -396 -5287 -384 -5253
rect -442 -5321 -384 -5287
rect -442 -5355 -430 -5321
rect -396 -5355 -384 -5321
rect -442 -5389 -384 -5355
rect -442 -5423 -430 -5389
rect -396 -5423 -384 -5389
rect -442 -5457 -384 -5423
rect -442 -5491 -430 -5457
rect -396 -5491 -384 -5457
rect -442 -5525 -384 -5491
rect -442 -5559 -430 -5525
rect -396 -5559 -384 -5525
rect -442 -5593 -384 -5559
rect -442 -5627 -430 -5593
rect -396 -5627 -384 -5593
rect -442 -5661 -384 -5627
rect -442 -5695 -430 -5661
rect -396 -5695 -384 -5661
rect -442 -5729 -384 -5695
rect -442 -5763 -430 -5729
rect -396 -5763 -384 -5729
rect -442 -5797 -384 -5763
rect -442 -5831 -430 -5797
rect -396 -5831 -384 -5797
rect -442 -5865 -384 -5831
rect -442 -5899 -430 -5865
rect -396 -5899 -384 -5865
rect -442 -5933 -384 -5899
rect -442 -5967 -430 -5933
rect -396 -5967 -384 -5933
rect -442 -6001 -384 -5967
rect -442 -6035 -430 -6001
rect -396 -6035 -384 -6001
rect -442 -6069 -384 -6035
rect -442 -6103 -430 -6069
rect -396 -6103 -384 -6069
rect -442 -6137 -384 -6103
rect -442 -6171 -430 -6137
rect -396 -6171 -384 -6137
rect -442 -6205 -384 -6171
rect -442 -6239 -430 -6205
rect -396 -6239 -384 -6205
rect -442 -6273 -384 -6239
rect -442 -6307 -430 -6273
rect -396 -6307 -384 -6273
rect -442 -6341 -384 -6307
rect -442 -6375 -430 -6341
rect -396 -6375 -384 -6341
rect -442 -6409 -384 -6375
rect -442 -6443 -430 -6409
rect -396 -6443 -384 -6409
rect -442 -6477 -384 -6443
rect -442 -6511 -430 -6477
rect -396 -6511 -384 -6477
rect -442 -6545 -384 -6511
rect -442 -6579 -430 -6545
rect -396 -6579 -384 -6545
rect -442 -6613 -384 -6579
rect -442 -6647 -430 -6613
rect -396 -6647 -384 -6613
rect -442 -6681 -384 -6647
rect -442 -6715 -430 -6681
rect -396 -6715 -384 -6681
rect -442 -6749 -384 -6715
rect -442 -6783 -430 -6749
rect -396 -6783 -384 -6749
rect -442 -6817 -384 -6783
rect -442 -6851 -430 -6817
rect -396 -6851 -384 -6817
rect -442 -6885 -384 -6851
rect -442 -6919 -430 -6885
rect -396 -6919 -384 -6885
rect -442 -6953 -384 -6919
rect -442 -6987 -430 -6953
rect -396 -6987 -384 -6953
rect -442 -7021 -384 -6987
rect -442 -7055 -430 -7021
rect -396 -7055 -384 -7021
rect -442 -7089 -384 -7055
rect -442 -7123 -430 -7089
rect -396 -7123 -384 -7089
rect -442 -7157 -384 -7123
rect -442 -7191 -430 -7157
rect -396 -7191 -384 -7157
rect -442 -7225 -384 -7191
rect -442 -7259 -430 -7225
rect -396 -7259 -384 -7225
rect -442 -7293 -384 -7259
rect -442 -7327 -430 -7293
rect -396 -7327 -384 -7293
rect -442 -7361 -384 -7327
rect -442 -7395 -430 -7361
rect -396 -7395 -384 -7361
rect -442 -7429 -384 -7395
rect -442 -7463 -430 -7429
rect -396 -7463 -384 -7429
rect -442 -7497 -384 -7463
rect -442 -7531 -430 -7497
rect -396 -7531 -384 -7497
rect -442 -7565 -384 -7531
rect -442 -7599 -430 -7565
rect -396 -7599 -384 -7565
rect -442 -7633 -384 -7599
rect -442 -7667 -430 -7633
rect -396 -7667 -384 -7633
rect -442 -7701 -384 -7667
rect -442 -7735 -430 -7701
rect -396 -7735 -384 -7701
rect -442 -7769 -384 -7735
rect -442 -7803 -430 -7769
rect -396 -7803 -384 -7769
rect -442 -7837 -384 -7803
rect -442 -7871 -430 -7837
rect -396 -7871 -384 -7837
rect -442 -7905 -384 -7871
rect -442 -7939 -430 -7905
rect -396 -7939 -384 -7905
rect -442 -7973 -384 -7939
rect -442 -8007 -430 -7973
rect -396 -8007 -384 -7973
rect -442 -8041 -384 -8007
rect -442 -8075 -430 -8041
rect -396 -8075 -384 -8041
rect -442 -8109 -384 -8075
rect -442 -8143 -430 -8109
rect -396 -8143 -384 -8109
rect -442 -8177 -384 -8143
rect -442 -8211 -430 -8177
rect -396 -8211 -384 -8177
rect -442 -8245 -384 -8211
rect -442 -8279 -430 -8245
rect -396 -8279 -384 -8245
rect -442 -8313 -384 -8279
rect -442 -8347 -430 -8313
rect -396 -8347 -384 -8313
rect -442 -8381 -384 -8347
rect -442 -8415 -430 -8381
rect -396 -8415 -384 -8381
rect -442 -8449 -384 -8415
rect -442 -8483 -430 -8449
rect -396 -8483 -384 -8449
rect -442 -8517 -384 -8483
rect -442 -8551 -430 -8517
rect -396 -8551 -384 -8517
rect -442 -8585 -384 -8551
rect -442 -8619 -430 -8585
rect -396 -8619 -384 -8585
rect -442 -8653 -384 -8619
rect -442 -8687 -430 -8653
rect -396 -8687 -384 -8653
rect -442 -8721 -384 -8687
rect -442 -8755 -430 -8721
rect -396 -8755 -384 -8721
rect -442 -8789 -384 -8755
rect -442 -8823 -430 -8789
rect -396 -8823 -384 -8789
rect -442 -8857 -384 -8823
rect -442 -8891 -430 -8857
rect -396 -8891 -384 -8857
rect -442 -8925 -384 -8891
rect -442 -8959 -430 -8925
rect -396 -8959 -384 -8925
rect -442 -8993 -384 -8959
rect -442 -9027 -430 -8993
rect -396 -9027 -384 -8993
rect -442 -9061 -384 -9027
rect -442 -9095 -430 -9061
rect -396 -9095 -384 -9061
rect -442 -9129 -384 -9095
rect -442 -9163 -430 -9129
rect -396 -9163 -384 -9129
rect -442 -9197 -384 -9163
rect -442 -9231 -430 -9197
rect -396 -9231 -384 -9197
rect -442 -9265 -384 -9231
rect -442 -9299 -430 -9265
rect -396 -9299 -384 -9265
rect -442 -9333 -384 -9299
rect -442 -9367 -430 -9333
rect -396 -9367 -384 -9333
rect -442 -9401 -384 -9367
rect -442 -9435 -430 -9401
rect -396 -9435 -384 -9401
rect -442 -9469 -384 -9435
rect -442 -9503 -430 -9469
rect -396 -9503 -384 -9469
rect -442 -9537 -384 -9503
rect -442 -9571 -430 -9537
rect -396 -9571 -384 -9537
rect -442 -9600 -384 -9571
rect -324 9571 -266 9600
rect -324 9537 -312 9571
rect -278 9537 -266 9571
rect -324 9503 -266 9537
rect -324 9469 -312 9503
rect -278 9469 -266 9503
rect -324 9435 -266 9469
rect -324 9401 -312 9435
rect -278 9401 -266 9435
rect -324 9367 -266 9401
rect -324 9333 -312 9367
rect -278 9333 -266 9367
rect -324 9299 -266 9333
rect -324 9265 -312 9299
rect -278 9265 -266 9299
rect -324 9231 -266 9265
rect -324 9197 -312 9231
rect -278 9197 -266 9231
rect -324 9163 -266 9197
rect -324 9129 -312 9163
rect -278 9129 -266 9163
rect -324 9095 -266 9129
rect -324 9061 -312 9095
rect -278 9061 -266 9095
rect -324 9027 -266 9061
rect -324 8993 -312 9027
rect -278 8993 -266 9027
rect -324 8959 -266 8993
rect -324 8925 -312 8959
rect -278 8925 -266 8959
rect -324 8891 -266 8925
rect -324 8857 -312 8891
rect -278 8857 -266 8891
rect -324 8823 -266 8857
rect -324 8789 -312 8823
rect -278 8789 -266 8823
rect -324 8755 -266 8789
rect -324 8721 -312 8755
rect -278 8721 -266 8755
rect -324 8687 -266 8721
rect -324 8653 -312 8687
rect -278 8653 -266 8687
rect -324 8619 -266 8653
rect -324 8585 -312 8619
rect -278 8585 -266 8619
rect -324 8551 -266 8585
rect -324 8517 -312 8551
rect -278 8517 -266 8551
rect -324 8483 -266 8517
rect -324 8449 -312 8483
rect -278 8449 -266 8483
rect -324 8415 -266 8449
rect -324 8381 -312 8415
rect -278 8381 -266 8415
rect -324 8347 -266 8381
rect -324 8313 -312 8347
rect -278 8313 -266 8347
rect -324 8279 -266 8313
rect -324 8245 -312 8279
rect -278 8245 -266 8279
rect -324 8211 -266 8245
rect -324 8177 -312 8211
rect -278 8177 -266 8211
rect -324 8143 -266 8177
rect -324 8109 -312 8143
rect -278 8109 -266 8143
rect -324 8075 -266 8109
rect -324 8041 -312 8075
rect -278 8041 -266 8075
rect -324 8007 -266 8041
rect -324 7973 -312 8007
rect -278 7973 -266 8007
rect -324 7939 -266 7973
rect -324 7905 -312 7939
rect -278 7905 -266 7939
rect -324 7871 -266 7905
rect -324 7837 -312 7871
rect -278 7837 -266 7871
rect -324 7803 -266 7837
rect -324 7769 -312 7803
rect -278 7769 -266 7803
rect -324 7735 -266 7769
rect -324 7701 -312 7735
rect -278 7701 -266 7735
rect -324 7667 -266 7701
rect -324 7633 -312 7667
rect -278 7633 -266 7667
rect -324 7599 -266 7633
rect -324 7565 -312 7599
rect -278 7565 -266 7599
rect -324 7531 -266 7565
rect -324 7497 -312 7531
rect -278 7497 -266 7531
rect -324 7463 -266 7497
rect -324 7429 -312 7463
rect -278 7429 -266 7463
rect -324 7395 -266 7429
rect -324 7361 -312 7395
rect -278 7361 -266 7395
rect -324 7327 -266 7361
rect -324 7293 -312 7327
rect -278 7293 -266 7327
rect -324 7259 -266 7293
rect -324 7225 -312 7259
rect -278 7225 -266 7259
rect -324 7191 -266 7225
rect -324 7157 -312 7191
rect -278 7157 -266 7191
rect -324 7123 -266 7157
rect -324 7089 -312 7123
rect -278 7089 -266 7123
rect -324 7055 -266 7089
rect -324 7021 -312 7055
rect -278 7021 -266 7055
rect -324 6987 -266 7021
rect -324 6953 -312 6987
rect -278 6953 -266 6987
rect -324 6919 -266 6953
rect -324 6885 -312 6919
rect -278 6885 -266 6919
rect -324 6851 -266 6885
rect -324 6817 -312 6851
rect -278 6817 -266 6851
rect -324 6783 -266 6817
rect -324 6749 -312 6783
rect -278 6749 -266 6783
rect -324 6715 -266 6749
rect -324 6681 -312 6715
rect -278 6681 -266 6715
rect -324 6647 -266 6681
rect -324 6613 -312 6647
rect -278 6613 -266 6647
rect -324 6579 -266 6613
rect -324 6545 -312 6579
rect -278 6545 -266 6579
rect -324 6511 -266 6545
rect -324 6477 -312 6511
rect -278 6477 -266 6511
rect -324 6443 -266 6477
rect -324 6409 -312 6443
rect -278 6409 -266 6443
rect -324 6375 -266 6409
rect -324 6341 -312 6375
rect -278 6341 -266 6375
rect -324 6307 -266 6341
rect -324 6273 -312 6307
rect -278 6273 -266 6307
rect -324 6239 -266 6273
rect -324 6205 -312 6239
rect -278 6205 -266 6239
rect -324 6171 -266 6205
rect -324 6137 -312 6171
rect -278 6137 -266 6171
rect -324 6103 -266 6137
rect -324 6069 -312 6103
rect -278 6069 -266 6103
rect -324 6035 -266 6069
rect -324 6001 -312 6035
rect -278 6001 -266 6035
rect -324 5967 -266 6001
rect -324 5933 -312 5967
rect -278 5933 -266 5967
rect -324 5899 -266 5933
rect -324 5865 -312 5899
rect -278 5865 -266 5899
rect -324 5831 -266 5865
rect -324 5797 -312 5831
rect -278 5797 -266 5831
rect -324 5763 -266 5797
rect -324 5729 -312 5763
rect -278 5729 -266 5763
rect -324 5695 -266 5729
rect -324 5661 -312 5695
rect -278 5661 -266 5695
rect -324 5627 -266 5661
rect -324 5593 -312 5627
rect -278 5593 -266 5627
rect -324 5559 -266 5593
rect -324 5525 -312 5559
rect -278 5525 -266 5559
rect -324 5491 -266 5525
rect -324 5457 -312 5491
rect -278 5457 -266 5491
rect -324 5423 -266 5457
rect -324 5389 -312 5423
rect -278 5389 -266 5423
rect -324 5355 -266 5389
rect -324 5321 -312 5355
rect -278 5321 -266 5355
rect -324 5287 -266 5321
rect -324 5253 -312 5287
rect -278 5253 -266 5287
rect -324 5219 -266 5253
rect -324 5185 -312 5219
rect -278 5185 -266 5219
rect -324 5151 -266 5185
rect -324 5117 -312 5151
rect -278 5117 -266 5151
rect -324 5083 -266 5117
rect -324 5049 -312 5083
rect -278 5049 -266 5083
rect -324 5015 -266 5049
rect -324 4981 -312 5015
rect -278 4981 -266 5015
rect -324 4947 -266 4981
rect -324 4913 -312 4947
rect -278 4913 -266 4947
rect -324 4879 -266 4913
rect -324 4845 -312 4879
rect -278 4845 -266 4879
rect -324 4811 -266 4845
rect -324 4777 -312 4811
rect -278 4777 -266 4811
rect -324 4743 -266 4777
rect -324 4709 -312 4743
rect -278 4709 -266 4743
rect -324 4675 -266 4709
rect -324 4641 -312 4675
rect -278 4641 -266 4675
rect -324 4607 -266 4641
rect -324 4573 -312 4607
rect -278 4573 -266 4607
rect -324 4539 -266 4573
rect -324 4505 -312 4539
rect -278 4505 -266 4539
rect -324 4471 -266 4505
rect -324 4437 -312 4471
rect -278 4437 -266 4471
rect -324 4403 -266 4437
rect -324 4369 -312 4403
rect -278 4369 -266 4403
rect -324 4335 -266 4369
rect -324 4301 -312 4335
rect -278 4301 -266 4335
rect -324 4267 -266 4301
rect -324 4233 -312 4267
rect -278 4233 -266 4267
rect -324 4199 -266 4233
rect -324 4165 -312 4199
rect -278 4165 -266 4199
rect -324 4131 -266 4165
rect -324 4097 -312 4131
rect -278 4097 -266 4131
rect -324 4063 -266 4097
rect -324 4029 -312 4063
rect -278 4029 -266 4063
rect -324 3995 -266 4029
rect -324 3961 -312 3995
rect -278 3961 -266 3995
rect -324 3927 -266 3961
rect -324 3893 -312 3927
rect -278 3893 -266 3927
rect -324 3859 -266 3893
rect -324 3825 -312 3859
rect -278 3825 -266 3859
rect -324 3791 -266 3825
rect -324 3757 -312 3791
rect -278 3757 -266 3791
rect -324 3723 -266 3757
rect -324 3689 -312 3723
rect -278 3689 -266 3723
rect -324 3655 -266 3689
rect -324 3621 -312 3655
rect -278 3621 -266 3655
rect -324 3587 -266 3621
rect -324 3553 -312 3587
rect -278 3553 -266 3587
rect -324 3519 -266 3553
rect -324 3485 -312 3519
rect -278 3485 -266 3519
rect -324 3451 -266 3485
rect -324 3417 -312 3451
rect -278 3417 -266 3451
rect -324 3383 -266 3417
rect -324 3349 -312 3383
rect -278 3349 -266 3383
rect -324 3315 -266 3349
rect -324 3281 -312 3315
rect -278 3281 -266 3315
rect -324 3247 -266 3281
rect -324 3213 -312 3247
rect -278 3213 -266 3247
rect -324 3179 -266 3213
rect -324 3145 -312 3179
rect -278 3145 -266 3179
rect -324 3111 -266 3145
rect -324 3077 -312 3111
rect -278 3077 -266 3111
rect -324 3043 -266 3077
rect -324 3009 -312 3043
rect -278 3009 -266 3043
rect -324 2975 -266 3009
rect -324 2941 -312 2975
rect -278 2941 -266 2975
rect -324 2907 -266 2941
rect -324 2873 -312 2907
rect -278 2873 -266 2907
rect -324 2839 -266 2873
rect -324 2805 -312 2839
rect -278 2805 -266 2839
rect -324 2771 -266 2805
rect -324 2737 -312 2771
rect -278 2737 -266 2771
rect -324 2703 -266 2737
rect -324 2669 -312 2703
rect -278 2669 -266 2703
rect -324 2635 -266 2669
rect -324 2601 -312 2635
rect -278 2601 -266 2635
rect -324 2567 -266 2601
rect -324 2533 -312 2567
rect -278 2533 -266 2567
rect -324 2499 -266 2533
rect -324 2465 -312 2499
rect -278 2465 -266 2499
rect -324 2431 -266 2465
rect -324 2397 -312 2431
rect -278 2397 -266 2431
rect -324 2363 -266 2397
rect -324 2329 -312 2363
rect -278 2329 -266 2363
rect -324 2295 -266 2329
rect -324 2261 -312 2295
rect -278 2261 -266 2295
rect -324 2227 -266 2261
rect -324 2193 -312 2227
rect -278 2193 -266 2227
rect -324 2159 -266 2193
rect -324 2125 -312 2159
rect -278 2125 -266 2159
rect -324 2091 -266 2125
rect -324 2057 -312 2091
rect -278 2057 -266 2091
rect -324 2023 -266 2057
rect -324 1989 -312 2023
rect -278 1989 -266 2023
rect -324 1955 -266 1989
rect -324 1921 -312 1955
rect -278 1921 -266 1955
rect -324 1887 -266 1921
rect -324 1853 -312 1887
rect -278 1853 -266 1887
rect -324 1819 -266 1853
rect -324 1785 -312 1819
rect -278 1785 -266 1819
rect -324 1751 -266 1785
rect -324 1717 -312 1751
rect -278 1717 -266 1751
rect -324 1683 -266 1717
rect -324 1649 -312 1683
rect -278 1649 -266 1683
rect -324 1615 -266 1649
rect -324 1581 -312 1615
rect -278 1581 -266 1615
rect -324 1547 -266 1581
rect -324 1513 -312 1547
rect -278 1513 -266 1547
rect -324 1479 -266 1513
rect -324 1445 -312 1479
rect -278 1445 -266 1479
rect -324 1411 -266 1445
rect -324 1377 -312 1411
rect -278 1377 -266 1411
rect -324 1343 -266 1377
rect -324 1309 -312 1343
rect -278 1309 -266 1343
rect -324 1275 -266 1309
rect -324 1241 -312 1275
rect -278 1241 -266 1275
rect -324 1207 -266 1241
rect -324 1173 -312 1207
rect -278 1173 -266 1207
rect -324 1139 -266 1173
rect -324 1105 -312 1139
rect -278 1105 -266 1139
rect -324 1071 -266 1105
rect -324 1037 -312 1071
rect -278 1037 -266 1071
rect -324 1003 -266 1037
rect -324 969 -312 1003
rect -278 969 -266 1003
rect -324 935 -266 969
rect -324 901 -312 935
rect -278 901 -266 935
rect -324 867 -266 901
rect -324 833 -312 867
rect -278 833 -266 867
rect -324 799 -266 833
rect -324 765 -312 799
rect -278 765 -266 799
rect -324 731 -266 765
rect -324 697 -312 731
rect -278 697 -266 731
rect -324 663 -266 697
rect -324 629 -312 663
rect -278 629 -266 663
rect -324 595 -266 629
rect -324 561 -312 595
rect -278 561 -266 595
rect -324 527 -266 561
rect -324 493 -312 527
rect -278 493 -266 527
rect -324 459 -266 493
rect -324 425 -312 459
rect -278 425 -266 459
rect -324 391 -266 425
rect -324 357 -312 391
rect -278 357 -266 391
rect -324 323 -266 357
rect -324 289 -312 323
rect -278 289 -266 323
rect -324 255 -266 289
rect -324 221 -312 255
rect -278 221 -266 255
rect -324 187 -266 221
rect -324 153 -312 187
rect -278 153 -266 187
rect -324 119 -266 153
rect -324 85 -312 119
rect -278 85 -266 119
rect -324 51 -266 85
rect -324 17 -312 51
rect -278 17 -266 51
rect -324 -17 -266 17
rect -324 -51 -312 -17
rect -278 -51 -266 -17
rect -324 -85 -266 -51
rect -324 -119 -312 -85
rect -278 -119 -266 -85
rect -324 -153 -266 -119
rect -324 -187 -312 -153
rect -278 -187 -266 -153
rect -324 -221 -266 -187
rect -324 -255 -312 -221
rect -278 -255 -266 -221
rect -324 -289 -266 -255
rect -324 -323 -312 -289
rect -278 -323 -266 -289
rect -324 -357 -266 -323
rect -324 -391 -312 -357
rect -278 -391 -266 -357
rect -324 -425 -266 -391
rect -324 -459 -312 -425
rect -278 -459 -266 -425
rect -324 -493 -266 -459
rect -324 -527 -312 -493
rect -278 -527 -266 -493
rect -324 -561 -266 -527
rect -324 -595 -312 -561
rect -278 -595 -266 -561
rect -324 -629 -266 -595
rect -324 -663 -312 -629
rect -278 -663 -266 -629
rect -324 -697 -266 -663
rect -324 -731 -312 -697
rect -278 -731 -266 -697
rect -324 -765 -266 -731
rect -324 -799 -312 -765
rect -278 -799 -266 -765
rect -324 -833 -266 -799
rect -324 -867 -312 -833
rect -278 -867 -266 -833
rect -324 -901 -266 -867
rect -324 -935 -312 -901
rect -278 -935 -266 -901
rect -324 -969 -266 -935
rect -324 -1003 -312 -969
rect -278 -1003 -266 -969
rect -324 -1037 -266 -1003
rect -324 -1071 -312 -1037
rect -278 -1071 -266 -1037
rect -324 -1105 -266 -1071
rect -324 -1139 -312 -1105
rect -278 -1139 -266 -1105
rect -324 -1173 -266 -1139
rect -324 -1207 -312 -1173
rect -278 -1207 -266 -1173
rect -324 -1241 -266 -1207
rect -324 -1275 -312 -1241
rect -278 -1275 -266 -1241
rect -324 -1309 -266 -1275
rect -324 -1343 -312 -1309
rect -278 -1343 -266 -1309
rect -324 -1377 -266 -1343
rect -324 -1411 -312 -1377
rect -278 -1411 -266 -1377
rect -324 -1445 -266 -1411
rect -324 -1479 -312 -1445
rect -278 -1479 -266 -1445
rect -324 -1513 -266 -1479
rect -324 -1547 -312 -1513
rect -278 -1547 -266 -1513
rect -324 -1581 -266 -1547
rect -324 -1615 -312 -1581
rect -278 -1615 -266 -1581
rect -324 -1649 -266 -1615
rect -324 -1683 -312 -1649
rect -278 -1683 -266 -1649
rect -324 -1717 -266 -1683
rect -324 -1751 -312 -1717
rect -278 -1751 -266 -1717
rect -324 -1785 -266 -1751
rect -324 -1819 -312 -1785
rect -278 -1819 -266 -1785
rect -324 -1853 -266 -1819
rect -324 -1887 -312 -1853
rect -278 -1887 -266 -1853
rect -324 -1921 -266 -1887
rect -324 -1955 -312 -1921
rect -278 -1955 -266 -1921
rect -324 -1989 -266 -1955
rect -324 -2023 -312 -1989
rect -278 -2023 -266 -1989
rect -324 -2057 -266 -2023
rect -324 -2091 -312 -2057
rect -278 -2091 -266 -2057
rect -324 -2125 -266 -2091
rect -324 -2159 -312 -2125
rect -278 -2159 -266 -2125
rect -324 -2193 -266 -2159
rect -324 -2227 -312 -2193
rect -278 -2227 -266 -2193
rect -324 -2261 -266 -2227
rect -324 -2295 -312 -2261
rect -278 -2295 -266 -2261
rect -324 -2329 -266 -2295
rect -324 -2363 -312 -2329
rect -278 -2363 -266 -2329
rect -324 -2397 -266 -2363
rect -324 -2431 -312 -2397
rect -278 -2431 -266 -2397
rect -324 -2465 -266 -2431
rect -324 -2499 -312 -2465
rect -278 -2499 -266 -2465
rect -324 -2533 -266 -2499
rect -324 -2567 -312 -2533
rect -278 -2567 -266 -2533
rect -324 -2601 -266 -2567
rect -324 -2635 -312 -2601
rect -278 -2635 -266 -2601
rect -324 -2669 -266 -2635
rect -324 -2703 -312 -2669
rect -278 -2703 -266 -2669
rect -324 -2737 -266 -2703
rect -324 -2771 -312 -2737
rect -278 -2771 -266 -2737
rect -324 -2805 -266 -2771
rect -324 -2839 -312 -2805
rect -278 -2839 -266 -2805
rect -324 -2873 -266 -2839
rect -324 -2907 -312 -2873
rect -278 -2907 -266 -2873
rect -324 -2941 -266 -2907
rect -324 -2975 -312 -2941
rect -278 -2975 -266 -2941
rect -324 -3009 -266 -2975
rect -324 -3043 -312 -3009
rect -278 -3043 -266 -3009
rect -324 -3077 -266 -3043
rect -324 -3111 -312 -3077
rect -278 -3111 -266 -3077
rect -324 -3145 -266 -3111
rect -324 -3179 -312 -3145
rect -278 -3179 -266 -3145
rect -324 -3213 -266 -3179
rect -324 -3247 -312 -3213
rect -278 -3247 -266 -3213
rect -324 -3281 -266 -3247
rect -324 -3315 -312 -3281
rect -278 -3315 -266 -3281
rect -324 -3349 -266 -3315
rect -324 -3383 -312 -3349
rect -278 -3383 -266 -3349
rect -324 -3417 -266 -3383
rect -324 -3451 -312 -3417
rect -278 -3451 -266 -3417
rect -324 -3485 -266 -3451
rect -324 -3519 -312 -3485
rect -278 -3519 -266 -3485
rect -324 -3553 -266 -3519
rect -324 -3587 -312 -3553
rect -278 -3587 -266 -3553
rect -324 -3621 -266 -3587
rect -324 -3655 -312 -3621
rect -278 -3655 -266 -3621
rect -324 -3689 -266 -3655
rect -324 -3723 -312 -3689
rect -278 -3723 -266 -3689
rect -324 -3757 -266 -3723
rect -324 -3791 -312 -3757
rect -278 -3791 -266 -3757
rect -324 -3825 -266 -3791
rect -324 -3859 -312 -3825
rect -278 -3859 -266 -3825
rect -324 -3893 -266 -3859
rect -324 -3927 -312 -3893
rect -278 -3927 -266 -3893
rect -324 -3961 -266 -3927
rect -324 -3995 -312 -3961
rect -278 -3995 -266 -3961
rect -324 -4029 -266 -3995
rect -324 -4063 -312 -4029
rect -278 -4063 -266 -4029
rect -324 -4097 -266 -4063
rect -324 -4131 -312 -4097
rect -278 -4131 -266 -4097
rect -324 -4165 -266 -4131
rect -324 -4199 -312 -4165
rect -278 -4199 -266 -4165
rect -324 -4233 -266 -4199
rect -324 -4267 -312 -4233
rect -278 -4267 -266 -4233
rect -324 -4301 -266 -4267
rect -324 -4335 -312 -4301
rect -278 -4335 -266 -4301
rect -324 -4369 -266 -4335
rect -324 -4403 -312 -4369
rect -278 -4403 -266 -4369
rect -324 -4437 -266 -4403
rect -324 -4471 -312 -4437
rect -278 -4471 -266 -4437
rect -324 -4505 -266 -4471
rect -324 -4539 -312 -4505
rect -278 -4539 -266 -4505
rect -324 -4573 -266 -4539
rect -324 -4607 -312 -4573
rect -278 -4607 -266 -4573
rect -324 -4641 -266 -4607
rect -324 -4675 -312 -4641
rect -278 -4675 -266 -4641
rect -324 -4709 -266 -4675
rect -324 -4743 -312 -4709
rect -278 -4743 -266 -4709
rect -324 -4777 -266 -4743
rect -324 -4811 -312 -4777
rect -278 -4811 -266 -4777
rect -324 -4845 -266 -4811
rect -324 -4879 -312 -4845
rect -278 -4879 -266 -4845
rect -324 -4913 -266 -4879
rect -324 -4947 -312 -4913
rect -278 -4947 -266 -4913
rect -324 -4981 -266 -4947
rect -324 -5015 -312 -4981
rect -278 -5015 -266 -4981
rect -324 -5049 -266 -5015
rect -324 -5083 -312 -5049
rect -278 -5083 -266 -5049
rect -324 -5117 -266 -5083
rect -324 -5151 -312 -5117
rect -278 -5151 -266 -5117
rect -324 -5185 -266 -5151
rect -324 -5219 -312 -5185
rect -278 -5219 -266 -5185
rect -324 -5253 -266 -5219
rect -324 -5287 -312 -5253
rect -278 -5287 -266 -5253
rect -324 -5321 -266 -5287
rect -324 -5355 -312 -5321
rect -278 -5355 -266 -5321
rect -324 -5389 -266 -5355
rect -324 -5423 -312 -5389
rect -278 -5423 -266 -5389
rect -324 -5457 -266 -5423
rect -324 -5491 -312 -5457
rect -278 -5491 -266 -5457
rect -324 -5525 -266 -5491
rect -324 -5559 -312 -5525
rect -278 -5559 -266 -5525
rect -324 -5593 -266 -5559
rect -324 -5627 -312 -5593
rect -278 -5627 -266 -5593
rect -324 -5661 -266 -5627
rect -324 -5695 -312 -5661
rect -278 -5695 -266 -5661
rect -324 -5729 -266 -5695
rect -324 -5763 -312 -5729
rect -278 -5763 -266 -5729
rect -324 -5797 -266 -5763
rect -324 -5831 -312 -5797
rect -278 -5831 -266 -5797
rect -324 -5865 -266 -5831
rect -324 -5899 -312 -5865
rect -278 -5899 -266 -5865
rect -324 -5933 -266 -5899
rect -324 -5967 -312 -5933
rect -278 -5967 -266 -5933
rect -324 -6001 -266 -5967
rect -324 -6035 -312 -6001
rect -278 -6035 -266 -6001
rect -324 -6069 -266 -6035
rect -324 -6103 -312 -6069
rect -278 -6103 -266 -6069
rect -324 -6137 -266 -6103
rect -324 -6171 -312 -6137
rect -278 -6171 -266 -6137
rect -324 -6205 -266 -6171
rect -324 -6239 -312 -6205
rect -278 -6239 -266 -6205
rect -324 -6273 -266 -6239
rect -324 -6307 -312 -6273
rect -278 -6307 -266 -6273
rect -324 -6341 -266 -6307
rect -324 -6375 -312 -6341
rect -278 -6375 -266 -6341
rect -324 -6409 -266 -6375
rect -324 -6443 -312 -6409
rect -278 -6443 -266 -6409
rect -324 -6477 -266 -6443
rect -324 -6511 -312 -6477
rect -278 -6511 -266 -6477
rect -324 -6545 -266 -6511
rect -324 -6579 -312 -6545
rect -278 -6579 -266 -6545
rect -324 -6613 -266 -6579
rect -324 -6647 -312 -6613
rect -278 -6647 -266 -6613
rect -324 -6681 -266 -6647
rect -324 -6715 -312 -6681
rect -278 -6715 -266 -6681
rect -324 -6749 -266 -6715
rect -324 -6783 -312 -6749
rect -278 -6783 -266 -6749
rect -324 -6817 -266 -6783
rect -324 -6851 -312 -6817
rect -278 -6851 -266 -6817
rect -324 -6885 -266 -6851
rect -324 -6919 -312 -6885
rect -278 -6919 -266 -6885
rect -324 -6953 -266 -6919
rect -324 -6987 -312 -6953
rect -278 -6987 -266 -6953
rect -324 -7021 -266 -6987
rect -324 -7055 -312 -7021
rect -278 -7055 -266 -7021
rect -324 -7089 -266 -7055
rect -324 -7123 -312 -7089
rect -278 -7123 -266 -7089
rect -324 -7157 -266 -7123
rect -324 -7191 -312 -7157
rect -278 -7191 -266 -7157
rect -324 -7225 -266 -7191
rect -324 -7259 -312 -7225
rect -278 -7259 -266 -7225
rect -324 -7293 -266 -7259
rect -324 -7327 -312 -7293
rect -278 -7327 -266 -7293
rect -324 -7361 -266 -7327
rect -324 -7395 -312 -7361
rect -278 -7395 -266 -7361
rect -324 -7429 -266 -7395
rect -324 -7463 -312 -7429
rect -278 -7463 -266 -7429
rect -324 -7497 -266 -7463
rect -324 -7531 -312 -7497
rect -278 -7531 -266 -7497
rect -324 -7565 -266 -7531
rect -324 -7599 -312 -7565
rect -278 -7599 -266 -7565
rect -324 -7633 -266 -7599
rect -324 -7667 -312 -7633
rect -278 -7667 -266 -7633
rect -324 -7701 -266 -7667
rect -324 -7735 -312 -7701
rect -278 -7735 -266 -7701
rect -324 -7769 -266 -7735
rect -324 -7803 -312 -7769
rect -278 -7803 -266 -7769
rect -324 -7837 -266 -7803
rect -324 -7871 -312 -7837
rect -278 -7871 -266 -7837
rect -324 -7905 -266 -7871
rect -324 -7939 -312 -7905
rect -278 -7939 -266 -7905
rect -324 -7973 -266 -7939
rect -324 -8007 -312 -7973
rect -278 -8007 -266 -7973
rect -324 -8041 -266 -8007
rect -324 -8075 -312 -8041
rect -278 -8075 -266 -8041
rect -324 -8109 -266 -8075
rect -324 -8143 -312 -8109
rect -278 -8143 -266 -8109
rect -324 -8177 -266 -8143
rect -324 -8211 -312 -8177
rect -278 -8211 -266 -8177
rect -324 -8245 -266 -8211
rect -324 -8279 -312 -8245
rect -278 -8279 -266 -8245
rect -324 -8313 -266 -8279
rect -324 -8347 -312 -8313
rect -278 -8347 -266 -8313
rect -324 -8381 -266 -8347
rect -324 -8415 -312 -8381
rect -278 -8415 -266 -8381
rect -324 -8449 -266 -8415
rect -324 -8483 -312 -8449
rect -278 -8483 -266 -8449
rect -324 -8517 -266 -8483
rect -324 -8551 -312 -8517
rect -278 -8551 -266 -8517
rect -324 -8585 -266 -8551
rect -324 -8619 -312 -8585
rect -278 -8619 -266 -8585
rect -324 -8653 -266 -8619
rect -324 -8687 -312 -8653
rect -278 -8687 -266 -8653
rect -324 -8721 -266 -8687
rect -324 -8755 -312 -8721
rect -278 -8755 -266 -8721
rect -324 -8789 -266 -8755
rect -324 -8823 -312 -8789
rect -278 -8823 -266 -8789
rect -324 -8857 -266 -8823
rect -324 -8891 -312 -8857
rect -278 -8891 -266 -8857
rect -324 -8925 -266 -8891
rect -324 -8959 -312 -8925
rect -278 -8959 -266 -8925
rect -324 -8993 -266 -8959
rect -324 -9027 -312 -8993
rect -278 -9027 -266 -8993
rect -324 -9061 -266 -9027
rect -324 -9095 -312 -9061
rect -278 -9095 -266 -9061
rect -324 -9129 -266 -9095
rect -324 -9163 -312 -9129
rect -278 -9163 -266 -9129
rect -324 -9197 -266 -9163
rect -324 -9231 -312 -9197
rect -278 -9231 -266 -9197
rect -324 -9265 -266 -9231
rect -324 -9299 -312 -9265
rect -278 -9299 -266 -9265
rect -324 -9333 -266 -9299
rect -324 -9367 -312 -9333
rect -278 -9367 -266 -9333
rect -324 -9401 -266 -9367
rect -324 -9435 -312 -9401
rect -278 -9435 -266 -9401
rect -324 -9469 -266 -9435
rect -324 -9503 -312 -9469
rect -278 -9503 -266 -9469
rect -324 -9537 -266 -9503
rect -324 -9571 -312 -9537
rect -278 -9571 -266 -9537
rect -324 -9600 -266 -9571
rect -206 9571 -148 9600
rect -206 9537 -194 9571
rect -160 9537 -148 9571
rect -206 9503 -148 9537
rect -206 9469 -194 9503
rect -160 9469 -148 9503
rect -206 9435 -148 9469
rect -206 9401 -194 9435
rect -160 9401 -148 9435
rect -206 9367 -148 9401
rect -206 9333 -194 9367
rect -160 9333 -148 9367
rect -206 9299 -148 9333
rect -206 9265 -194 9299
rect -160 9265 -148 9299
rect -206 9231 -148 9265
rect -206 9197 -194 9231
rect -160 9197 -148 9231
rect -206 9163 -148 9197
rect -206 9129 -194 9163
rect -160 9129 -148 9163
rect -206 9095 -148 9129
rect -206 9061 -194 9095
rect -160 9061 -148 9095
rect -206 9027 -148 9061
rect -206 8993 -194 9027
rect -160 8993 -148 9027
rect -206 8959 -148 8993
rect -206 8925 -194 8959
rect -160 8925 -148 8959
rect -206 8891 -148 8925
rect -206 8857 -194 8891
rect -160 8857 -148 8891
rect -206 8823 -148 8857
rect -206 8789 -194 8823
rect -160 8789 -148 8823
rect -206 8755 -148 8789
rect -206 8721 -194 8755
rect -160 8721 -148 8755
rect -206 8687 -148 8721
rect -206 8653 -194 8687
rect -160 8653 -148 8687
rect -206 8619 -148 8653
rect -206 8585 -194 8619
rect -160 8585 -148 8619
rect -206 8551 -148 8585
rect -206 8517 -194 8551
rect -160 8517 -148 8551
rect -206 8483 -148 8517
rect -206 8449 -194 8483
rect -160 8449 -148 8483
rect -206 8415 -148 8449
rect -206 8381 -194 8415
rect -160 8381 -148 8415
rect -206 8347 -148 8381
rect -206 8313 -194 8347
rect -160 8313 -148 8347
rect -206 8279 -148 8313
rect -206 8245 -194 8279
rect -160 8245 -148 8279
rect -206 8211 -148 8245
rect -206 8177 -194 8211
rect -160 8177 -148 8211
rect -206 8143 -148 8177
rect -206 8109 -194 8143
rect -160 8109 -148 8143
rect -206 8075 -148 8109
rect -206 8041 -194 8075
rect -160 8041 -148 8075
rect -206 8007 -148 8041
rect -206 7973 -194 8007
rect -160 7973 -148 8007
rect -206 7939 -148 7973
rect -206 7905 -194 7939
rect -160 7905 -148 7939
rect -206 7871 -148 7905
rect -206 7837 -194 7871
rect -160 7837 -148 7871
rect -206 7803 -148 7837
rect -206 7769 -194 7803
rect -160 7769 -148 7803
rect -206 7735 -148 7769
rect -206 7701 -194 7735
rect -160 7701 -148 7735
rect -206 7667 -148 7701
rect -206 7633 -194 7667
rect -160 7633 -148 7667
rect -206 7599 -148 7633
rect -206 7565 -194 7599
rect -160 7565 -148 7599
rect -206 7531 -148 7565
rect -206 7497 -194 7531
rect -160 7497 -148 7531
rect -206 7463 -148 7497
rect -206 7429 -194 7463
rect -160 7429 -148 7463
rect -206 7395 -148 7429
rect -206 7361 -194 7395
rect -160 7361 -148 7395
rect -206 7327 -148 7361
rect -206 7293 -194 7327
rect -160 7293 -148 7327
rect -206 7259 -148 7293
rect -206 7225 -194 7259
rect -160 7225 -148 7259
rect -206 7191 -148 7225
rect -206 7157 -194 7191
rect -160 7157 -148 7191
rect -206 7123 -148 7157
rect -206 7089 -194 7123
rect -160 7089 -148 7123
rect -206 7055 -148 7089
rect -206 7021 -194 7055
rect -160 7021 -148 7055
rect -206 6987 -148 7021
rect -206 6953 -194 6987
rect -160 6953 -148 6987
rect -206 6919 -148 6953
rect -206 6885 -194 6919
rect -160 6885 -148 6919
rect -206 6851 -148 6885
rect -206 6817 -194 6851
rect -160 6817 -148 6851
rect -206 6783 -148 6817
rect -206 6749 -194 6783
rect -160 6749 -148 6783
rect -206 6715 -148 6749
rect -206 6681 -194 6715
rect -160 6681 -148 6715
rect -206 6647 -148 6681
rect -206 6613 -194 6647
rect -160 6613 -148 6647
rect -206 6579 -148 6613
rect -206 6545 -194 6579
rect -160 6545 -148 6579
rect -206 6511 -148 6545
rect -206 6477 -194 6511
rect -160 6477 -148 6511
rect -206 6443 -148 6477
rect -206 6409 -194 6443
rect -160 6409 -148 6443
rect -206 6375 -148 6409
rect -206 6341 -194 6375
rect -160 6341 -148 6375
rect -206 6307 -148 6341
rect -206 6273 -194 6307
rect -160 6273 -148 6307
rect -206 6239 -148 6273
rect -206 6205 -194 6239
rect -160 6205 -148 6239
rect -206 6171 -148 6205
rect -206 6137 -194 6171
rect -160 6137 -148 6171
rect -206 6103 -148 6137
rect -206 6069 -194 6103
rect -160 6069 -148 6103
rect -206 6035 -148 6069
rect -206 6001 -194 6035
rect -160 6001 -148 6035
rect -206 5967 -148 6001
rect -206 5933 -194 5967
rect -160 5933 -148 5967
rect -206 5899 -148 5933
rect -206 5865 -194 5899
rect -160 5865 -148 5899
rect -206 5831 -148 5865
rect -206 5797 -194 5831
rect -160 5797 -148 5831
rect -206 5763 -148 5797
rect -206 5729 -194 5763
rect -160 5729 -148 5763
rect -206 5695 -148 5729
rect -206 5661 -194 5695
rect -160 5661 -148 5695
rect -206 5627 -148 5661
rect -206 5593 -194 5627
rect -160 5593 -148 5627
rect -206 5559 -148 5593
rect -206 5525 -194 5559
rect -160 5525 -148 5559
rect -206 5491 -148 5525
rect -206 5457 -194 5491
rect -160 5457 -148 5491
rect -206 5423 -148 5457
rect -206 5389 -194 5423
rect -160 5389 -148 5423
rect -206 5355 -148 5389
rect -206 5321 -194 5355
rect -160 5321 -148 5355
rect -206 5287 -148 5321
rect -206 5253 -194 5287
rect -160 5253 -148 5287
rect -206 5219 -148 5253
rect -206 5185 -194 5219
rect -160 5185 -148 5219
rect -206 5151 -148 5185
rect -206 5117 -194 5151
rect -160 5117 -148 5151
rect -206 5083 -148 5117
rect -206 5049 -194 5083
rect -160 5049 -148 5083
rect -206 5015 -148 5049
rect -206 4981 -194 5015
rect -160 4981 -148 5015
rect -206 4947 -148 4981
rect -206 4913 -194 4947
rect -160 4913 -148 4947
rect -206 4879 -148 4913
rect -206 4845 -194 4879
rect -160 4845 -148 4879
rect -206 4811 -148 4845
rect -206 4777 -194 4811
rect -160 4777 -148 4811
rect -206 4743 -148 4777
rect -206 4709 -194 4743
rect -160 4709 -148 4743
rect -206 4675 -148 4709
rect -206 4641 -194 4675
rect -160 4641 -148 4675
rect -206 4607 -148 4641
rect -206 4573 -194 4607
rect -160 4573 -148 4607
rect -206 4539 -148 4573
rect -206 4505 -194 4539
rect -160 4505 -148 4539
rect -206 4471 -148 4505
rect -206 4437 -194 4471
rect -160 4437 -148 4471
rect -206 4403 -148 4437
rect -206 4369 -194 4403
rect -160 4369 -148 4403
rect -206 4335 -148 4369
rect -206 4301 -194 4335
rect -160 4301 -148 4335
rect -206 4267 -148 4301
rect -206 4233 -194 4267
rect -160 4233 -148 4267
rect -206 4199 -148 4233
rect -206 4165 -194 4199
rect -160 4165 -148 4199
rect -206 4131 -148 4165
rect -206 4097 -194 4131
rect -160 4097 -148 4131
rect -206 4063 -148 4097
rect -206 4029 -194 4063
rect -160 4029 -148 4063
rect -206 3995 -148 4029
rect -206 3961 -194 3995
rect -160 3961 -148 3995
rect -206 3927 -148 3961
rect -206 3893 -194 3927
rect -160 3893 -148 3927
rect -206 3859 -148 3893
rect -206 3825 -194 3859
rect -160 3825 -148 3859
rect -206 3791 -148 3825
rect -206 3757 -194 3791
rect -160 3757 -148 3791
rect -206 3723 -148 3757
rect -206 3689 -194 3723
rect -160 3689 -148 3723
rect -206 3655 -148 3689
rect -206 3621 -194 3655
rect -160 3621 -148 3655
rect -206 3587 -148 3621
rect -206 3553 -194 3587
rect -160 3553 -148 3587
rect -206 3519 -148 3553
rect -206 3485 -194 3519
rect -160 3485 -148 3519
rect -206 3451 -148 3485
rect -206 3417 -194 3451
rect -160 3417 -148 3451
rect -206 3383 -148 3417
rect -206 3349 -194 3383
rect -160 3349 -148 3383
rect -206 3315 -148 3349
rect -206 3281 -194 3315
rect -160 3281 -148 3315
rect -206 3247 -148 3281
rect -206 3213 -194 3247
rect -160 3213 -148 3247
rect -206 3179 -148 3213
rect -206 3145 -194 3179
rect -160 3145 -148 3179
rect -206 3111 -148 3145
rect -206 3077 -194 3111
rect -160 3077 -148 3111
rect -206 3043 -148 3077
rect -206 3009 -194 3043
rect -160 3009 -148 3043
rect -206 2975 -148 3009
rect -206 2941 -194 2975
rect -160 2941 -148 2975
rect -206 2907 -148 2941
rect -206 2873 -194 2907
rect -160 2873 -148 2907
rect -206 2839 -148 2873
rect -206 2805 -194 2839
rect -160 2805 -148 2839
rect -206 2771 -148 2805
rect -206 2737 -194 2771
rect -160 2737 -148 2771
rect -206 2703 -148 2737
rect -206 2669 -194 2703
rect -160 2669 -148 2703
rect -206 2635 -148 2669
rect -206 2601 -194 2635
rect -160 2601 -148 2635
rect -206 2567 -148 2601
rect -206 2533 -194 2567
rect -160 2533 -148 2567
rect -206 2499 -148 2533
rect -206 2465 -194 2499
rect -160 2465 -148 2499
rect -206 2431 -148 2465
rect -206 2397 -194 2431
rect -160 2397 -148 2431
rect -206 2363 -148 2397
rect -206 2329 -194 2363
rect -160 2329 -148 2363
rect -206 2295 -148 2329
rect -206 2261 -194 2295
rect -160 2261 -148 2295
rect -206 2227 -148 2261
rect -206 2193 -194 2227
rect -160 2193 -148 2227
rect -206 2159 -148 2193
rect -206 2125 -194 2159
rect -160 2125 -148 2159
rect -206 2091 -148 2125
rect -206 2057 -194 2091
rect -160 2057 -148 2091
rect -206 2023 -148 2057
rect -206 1989 -194 2023
rect -160 1989 -148 2023
rect -206 1955 -148 1989
rect -206 1921 -194 1955
rect -160 1921 -148 1955
rect -206 1887 -148 1921
rect -206 1853 -194 1887
rect -160 1853 -148 1887
rect -206 1819 -148 1853
rect -206 1785 -194 1819
rect -160 1785 -148 1819
rect -206 1751 -148 1785
rect -206 1717 -194 1751
rect -160 1717 -148 1751
rect -206 1683 -148 1717
rect -206 1649 -194 1683
rect -160 1649 -148 1683
rect -206 1615 -148 1649
rect -206 1581 -194 1615
rect -160 1581 -148 1615
rect -206 1547 -148 1581
rect -206 1513 -194 1547
rect -160 1513 -148 1547
rect -206 1479 -148 1513
rect -206 1445 -194 1479
rect -160 1445 -148 1479
rect -206 1411 -148 1445
rect -206 1377 -194 1411
rect -160 1377 -148 1411
rect -206 1343 -148 1377
rect -206 1309 -194 1343
rect -160 1309 -148 1343
rect -206 1275 -148 1309
rect -206 1241 -194 1275
rect -160 1241 -148 1275
rect -206 1207 -148 1241
rect -206 1173 -194 1207
rect -160 1173 -148 1207
rect -206 1139 -148 1173
rect -206 1105 -194 1139
rect -160 1105 -148 1139
rect -206 1071 -148 1105
rect -206 1037 -194 1071
rect -160 1037 -148 1071
rect -206 1003 -148 1037
rect -206 969 -194 1003
rect -160 969 -148 1003
rect -206 935 -148 969
rect -206 901 -194 935
rect -160 901 -148 935
rect -206 867 -148 901
rect -206 833 -194 867
rect -160 833 -148 867
rect -206 799 -148 833
rect -206 765 -194 799
rect -160 765 -148 799
rect -206 731 -148 765
rect -206 697 -194 731
rect -160 697 -148 731
rect -206 663 -148 697
rect -206 629 -194 663
rect -160 629 -148 663
rect -206 595 -148 629
rect -206 561 -194 595
rect -160 561 -148 595
rect -206 527 -148 561
rect -206 493 -194 527
rect -160 493 -148 527
rect -206 459 -148 493
rect -206 425 -194 459
rect -160 425 -148 459
rect -206 391 -148 425
rect -206 357 -194 391
rect -160 357 -148 391
rect -206 323 -148 357
rect -206 289 -194 323
rect -160 289 -148 323
rect -206 255 -148 289
rect -206 221 -194 255
rect -160 221 -148 255
rect -206 187 -148 221
rect -206 153 -194 187
rect -160 153 -148 187
rect -206 119 -148 153
rect -206 85 -194 119
rect -160 85 -148 119
rect -206 51 -148 85
rect -206 17 -194 51
rect -160 17 -148 51
rect -206 -17 -148 17
rect -206 -51 -194 -17
rect -160 -51 -148 -17
rect -206 -85 -148 -51
rect -206 -119 -194 -85
rect -160 -119 -148 -85
rect -206 -153 -148 -119
rect -206 -187 -194 -153
rect -160 -187 -148 -153
rect -206 -221 -148 -187
rect -206 -255 -194 -221
rect -160 -255 -148 -221
rect -206 -289 -148 -255
rect -206 -323 -194 -289
rect -160 -323 -148 -289
rect -206 -357 -148 -323
rect -206 -391 -194 -357
rect -160 -391 -148 -357
rect -206 -425 -148 -391
rect -206 -459 -194 -425
rect -160 -459 -148 -425
rect -206 -493 -148 -459
rect -206 -527 -194 -493
rect -160 -527 -148 -493
rect -206 -561 -148 -527
rect -206 -595 -194 -561
rect -160 -595 -148 -561
rect -206 -629 -148 -595
rect -206 -663 -194 -629
rect -160 -663 -148 -629
rect -206 -697 -148 -663
rect -206 -731 -194 -697
rect -160 -731 -148 -697
rect -206 -765 -148 -731
rect -206 -799 -194 -765
rect -160 -799 -148 -765
rect -206 -833 -148 -799
rect -206 -867 -194 -833
rect -160 -867 -148 -833
rect -206 -901 -148 -867
rect -206 -935 -194 -901
rect -160 -935 -148 -901
rect -206 -969 -148 -935
rect -206 -1003 -194 -969
rect -160 -1003 -148 -969
rect -206 -1037 -148 -1003
rect -206 -1071 -194 -1037
rect -160 -1071 -148 -1037
rect -206 -1105 -148 -1071
rect -206 -1139 -194 -1105
rect -160 -1139 -148 -1105
rect -206 -1173 -148 -1139
rect -206 -1207 -194 -1173
rect -160 -1207 -148 -1173
rect -206 -1241 -148 -1207
rect -206 -1275 -194 -1241
rect -160 -1275 -148 -1241
rect -206 -1309 -148 -1275
rect -206 -1343 -194 -1309
rect -160 -1343 -148 -1309
rect -206 -1377 -148 -1343
rect -206 -1411 -194 -1377
rect -160 -1411 -148 -1377
rect -206 -1445 -148 -1411
rect -206 -1479 -194 -1445
rect -160 -1479 -148 -1445
rect -206 -1513 -148 -1479
rect -206 -1547 -194 -1513
rect -160 -1547 -148 -1513
rect -206 -1581 -148 -1547
rect -206 -1615 -194 -1581
rect -160 -1615 -148 -1581
rect -206 -1649 -148 -1615
rect -206 -1683 -194 -1649
rect -160 -1683 -148 -1649
rect -206 -1717 -148 -1683
rect -206 -1751 -194 -1717
rect -160 -1751 -148 -1717
rect -206 -1785 -148 -1751
rect -206 -1819 -194 -1785
rect -160 -1819 -148 -1785
rect -206 -1853 -148 -1819
rect -206 -1887 -194 -1853
rect -160 -1887 -148 -1853
rect -206 -1921 -148 -1887
rect -206 -1955 -194 -1921
rect -160 -1955 -148 -1921
rect -206 -1989 -148 -1955
rect -206 -2023 -194 -1989
rect -160 -2023 -148 -1989
rect -206 -2057 -148 -2023
rect -206 -2091 -194 -2057
rect -160 -2091 -148 -2057
rect -206 -2125 -148 -2091
rect -206 -2159 -194 -2125
rect -160 -2159 -148 -2125
rect -206 -2193 -148 -2159
rect -206 -2227 -194 -2193
rect -160 -2227 -148 -2193
rect -206 -2261 -148 -2227
rect -206 -2295 -194 -2261
rect -160 -2295 -148 -2261
rect -206 -2329 -148 -2295
rect -206 -2363 -194 -2329
rect -160 -2363 -148 -2329
rect -206 -2397 -148 -2363
rect -206 -2431 -194 -2397
rect -160 -2431 -148 -2397
rect -206 -2465 -148 -2431
rect -206 -2499 -194 -2465
rect -160 -2499 -148 -2465
rect -206 -2533 -148 -2499
rect -206 -2567 -194 -2533
rect -160 -2567 -148 -2533
rect -206 -2601 -148 -2567
rect -206 -2635 -194 -2601
rect -160 -2635 -148 -2601
rect -206 -2669 -148 -2635
rect -206 -2703 -194 -2669
rect -160 -2703 -148 -2669
rect -206 -2737 -148 -2703
rect -206 -2771 -194 -2737
rect -160 -2771 -148 -2737
rect -206 -2805 -148 -2771
rect -206 -2839 -194 -2805
rect -160 -2839 -148 -2805
rect -206 -2873 -148 -2839
rect -206 -2907 -194 -2873
rect -160 -2907 -148 -2873
rect -206 -2941 -148 -2907
rect -206 -2975 -194 -2941
rect -160 -2975 -148 -2941
rect -206 -3009 -148 -2975
rect -206 -3043 -194 -3009
rect -160 -3043 -148 -3009
rect -206 -3077 -148 -3043
rect -206 -3111 -194 -3077
rect -160 -3111 -148 -3077
rect -206 -3145 -148 -3111
rect -206 -3179 -194 -3145
rect -160 -3179 -148 -3145
rect -206 -3213 -148 -3179
rect -206 -3247 -194 -3213
rect -160 -3247 -148 -3213
rect -206 -3281 -148 -3247
rect -206 -3315 -194 -3281
rect -160 -3315 -148 -3281
rect -206 -3349 -148 -3315
rect -206 -3383 -194 -3349
rect -160 -3383 -148 -3349
rect -206 -3417 -148 -3383
rect -206 -3451 -194 -3417
rect -160 -3451 -148 -3417
rect -206 -3485 -148 -3451
rect -206 -3519 -194 -3485
rect -160 -3519 -148 -3485
rect -206 -3553 -148 -3519
rect -206 -3587 -194 -3553
rect -160 -3587 -148 -3553
rect -206 -3621 -148 -3587
rect -206 -3655 -194 -3621
rect -160 -3655 -148 -3621
rect -206 -3689 -148 -3655
rect -206 -3723 -194 -3689
rect -160 -3723 -148 -3689
rect -206 -3757 -148 -3723
rect -206 -3791 -194 -3757
rect -160 -3791 -148 -3757
rect -206 -3825 -148 -3791
rect -206 -3859 -194 -3825
rect -160 -3859 -148 -3825
rect -206 -3893 -148 -3859
rect -206 -3927 -194 -3893
rect -160 -3927 -148 -3893
rect -206 -3961 -148 -3927
rect -206 -3995 -194 -3961
rect -160 -3995 -148 -3961
rect -206 -4029 -148 -3995
rect -206 -4063 -194 -4029
rect -160 -4063 -148 -4029
rect -206 -4097 -148 -4063
rect -206 -4131 -194 -4097
rect -160 -4131 -148 -4097
rect -206 -4165 -148 -4131
rect -206 -4199 -194 -4165
rect -160 -4199 -148 -4165
rect -206 -4233 -148 -4199
rect -206 -4267 -194 -4233
rect -160 -4267 -148 -4233
rect -206 -4301 -148 -4267
rect -206 -4335 -194 -4301
rect -160 -4335 -148 -4301
rect -206 -4369 -148 -4335
rect -206 -4403 -194 -4369
rect -160 -4403 -148 -4369
rect -206 -4437 -148 -4403
rect -206 -4471 -194 -4437
rect -160 -4471 -148 -4437
rect -206 -4505 -148 -4471
rect -206 -4539 -194 -4505
rect -160 -4539 -148 -4505
rect -206 -4573 -148 -4539
rect -206 -4607 -194 -4573
rect -160 -4607 -148 -4573
rect -206 -4641 -148 -4607
rect -206 -4675 -194 -4641
rect -160 -4675 -148 -4641
rect -206 -4709 -148 -4675
rect -206 -4743 -194 -4709
rect -160 -4743 -148 -4709
rect -206 -4777 -148 -4743
rect -206 -4811 -194 -4777
rect -160 -4811 -148 -4777
rect -206 -4845 -148 -4811
rect -206 -4879 -194 -4845
rect -160 -4879 -148 -4845
rect -206 -4913 -148 -4879
rect -206 -4947 -194 -4913
rect -160 -4947 -148 -4913
rect -206 -4981 -148 -4947
rect -206 -5015 -194 -4981
rect -160 -5015 -148 -4981
rect -206 -5049 -148 -5015
rect -206 -5083 -194 -5049
rect -160 -5083 -148 -5049
rect -206 -5117 -148 -5083
rect -206 -5151 -194 -5117
rect -160 -5151 -148 -5117
rect -206 -5185 -148 -5151
rect -206 -5219 -194 -5185
rect -160 -5219 -148 -5185
rect -206 -5253 -148 -5219
rect -206 -5287 -194 -5253
rect -160 -5287 -148 -5253
rect -206 -5321 -148 -5287
rect -206 -5355 -194 -5321
rect -160 -5355 -148 -5321
rect -206 -5389 -148 -5355
rect -206 -5423 -194 -5389
rect -160 -5423 -148 -5389
rect -206 -5457 -148 -5423
rect -206 -5491 -194 -5457
rect -160 -5491 -148 -5457
rect -206 -5525 -148 -5491
rect -206 -5559 -194 -5525
rect -160 -5559 -148 -5525
rect -206 -5593 -148 -5559
rect -206 -5627 -194 -5593
rect -160 -5627 -148 -5593
rect -206 -5661 -148 -5627
rect -206 -5695 -194 -5661
rect -160 -5695 -148 -5661
rect -206 -5729 -148 -5695
rect -206 -5763 -194 -5729
rect -160 -5763 -148 -5729
rect -206 -5797 -148 -5763
rect -206 -5831 -194 -5797
rect -160 -5831 -148 -5797
rect -206 -5865 -148 -5831
rect -206 -5899 -194 -5865
rect -160 -5899 -148 -5865
rect -206 -5933 -148 -5899
rect -206 -5967 -194 -5933
rect -160 -5967 -148 -5933
rect -206 -6001 -148 -5967
rect -206 -6035 -194 -6001
rect -160 -6035 -148 -6001
rect -206 -6069 -148 -6035
rect -206 -6103 -194 -6069
rect -160 -6103 -148 -6069
rect -206 -6137 -148 -6103
rect -206 -6171 -194 -6137
rect -160 -6171 -148 -6137
rect -206 -6205 -148 -6171
rect -206 -6239 -194 -6205
rect -160 -6239 -148 -6205
rect -206 -6273 -148 -6239
rect -206 -6307 -194 -6273
rect -160 -6307 -148 -6273
rect -206 -6341 -148 -6307
rect -206 -6375 -194 -6341
rect -160 -6375 -148 -6341
rect -206 -6409 -148 -6375
rect -206 -6443 -194 -6409
rect -160 -6443 -148 -6409
rect -206 -6477 -148 -6443
rect -206 -6511 -194 -6477
rect -160 -6511 -148 -6477
rect -206 -6545 -148 -6511
rect -206 -6579 -194 -6545
rect -160 -6579 -148 -6545
rect -206 -6613 -148 -6579
rect -206 -6647 -194 -6613
rect -160 -6647 -148 -6613
rect -206 -6681 -148 -6647
rect -206 -6715 -194 -6681
rect -160 -6715 -148 -6681
rect -206 -6749 -148 -6715
rect -206 -6783 -194 -6749
rect -160 -6783 -148 -6749
rect -206 -6817 -148 -6783
rect -206 -6851 -194 -6817
rect -160 -6851 -148 -6817
rect -206 -6885 -148 -6851
rect -206 -6919 -194 -6885
rect -160 -6919 -148 -6885
rect -206 -6953 -148 -6919
rect -206 -6987 -194 -6953
rect -160 -6987 -148 -6953
rect -206 -7021 -148 -6987
rect -206 -7055 -194 -7021
rect -160 -7055 -148 -7021
rect -206 -7089 -148 -7055
rect -206 -7123 -194 -7089
rect -160 -7123 -148 -7089
rect -206 -7157 -148 -7123
rect -206 -7191 -194 -7157
rect -160 -7191 -148 -7157
rect -206 -7225 -148 -7191
rect -206 -7259 -194 -7225
rect -160 -7259 -148 -7225
rect -206 -7293 -148 -7259
rect -206 -7327 -194 -7293
rect -160 -7327 -148 -7293
rect -206 -7361 -148 -7327
rect -206 -7395 -194 -7361
rect -160 -7395 -148 -7361
rect -206 -7429 -148 -7395
rect -206 -7463 -194 -7429
rect -160 -7463 -148 -7429
rect -206 -7497 -148 -7463
rect -206 -7531 -194 -7497
rect -160 -7531 -148 -7497
rect -206 -7565 -148 -7531
rect -206 -7599 -194 -7565
rect -160 -7599 -148 -7565
rect -206 -7633 -148 -7599
rect -206 -7667 -194 -7633
rect -160 -7667 -148 -7633
rect -206 -7701 -148 -7667
rect -206 -7735 -194 -7701
rect -160 -7735 -148 -7701
rect -206 -7769 -148 -7735
rect -206 -7803 -194 -7769
rect -160 -7803 -148 -7769
rect -206 -7837 -148 -7803
rect -206 -7871 -194 -7837
rect -160 -7871 -148 -7837
rect -206 -7905 -148 -7871
rect -206 -7939 -194 -7905
rect -160 -7939 -148 -7905
rect -206 -7973 -148 -7939
rect -206 -8007 -194 -7973
rect -160 -8007 -148 -7973
rect -206 -8041 -148 -8007
rect -206 -8075 -194 -8041
rect -160 -8075 -148 -8041
rect -206 -8109 -148 -8075
rect -206 -8143 -194 -8109
rect -160 -8143 -148 -8109
rect -206 -8177 -148 -8143
rect -206 -8211 -194 -8177
rect -160 -8211 -148 -8177
rect -206 -8245 -148 -8211
rect -206 -8279 -194 -8245
rect -160 -8279 -148 -8245
rect -206 -8313 -148 -8279
rect -206 -8347 -194 -8313
rect -160 -8347 -148 -8313
rect -206 -8381 -148 -8347
rect -206 -8415 -194 -8381
rect -160 -8415 -148 -8381
rect -206 -8449 -148 -8415
rect -206 -8483 -194 -8449
rect -160 -8483 -148 -8449
rect -206 -8517 -148 -8483
rect -206 -8551 -194 -8517
rect -160 -8551 -148 -8517
rect -206 -8585 -148 -8551
rect -206 -8619 -194 -8585
rect -160 -8619 -148 -8585
rect -206 -8653 -148 -8619
rect -206 -8687 -194 -8653
rect -160 -8687 -148 -8653
rect -206 -8721 -148 -8687
rect -206 -8755 -194 -8721
rect -160 -8755 -148 -8721
rect -206 -8789 -148 -8755
rect -206 -8823 -194 -8789
rect -160 -8823 -148 -8789
rect -206 -8857 -148 -8823
rect -206 -8891 -194 -8857
rect -160 -8891 -148 -8857
rect -206 -8925 -148 -8891
rect -206 -8959 -194 -8925
rect -160 -8959 -148 -8925
rect -206 -8993 -148 -8959
rect -206 -9027 -194 -8993
rect -160 -9027 -148 -8993
rect -206 -9061 -148 -9027
rect -206 -9095 -194 -9061
rect -160 -9095 -148 -9061
rect -206 -9129 -148 -9095
rect -206 -9163 -194 -9129
rect -160 -9163 -148 -9129
rect -206 -9197 -148 -9163
rect -206 -9231 -194 -9197
rect -160 -9231 -148 -9197
rect -206 -9265 -148 -9231
rect -206 -9299 -194 -9265
rect -160 -9299 -148 -9265
rect -206 -9333 -148 -9299
rect -206 -9367 -194 -9333
rect -160 -9367 -148 -9333
rect -206 -9401 -148 -9367
rect -206 -9435 -194 -9401
rect -160 -9435 -148 -9401
rect -206 -9469 -148 -9435
rect -206 -9503 -194 -9469
rect -160 -9503 -148 -9469
rect -206 -9537 -148 -9503
rect -206 -9571 -194 -9537
rect -160 -9571 -148 -9537
rect -206 -9600 -148 -9571
rect -88 9571 -30 9600
rect -88 9537 -76 9571
rect -42 9537 -30 9571
rect -88 9503 -30 9537
rect -88 9469 -76 9503
rect -42 9469 -30 9503
rect -88 9435 -30 9469
rect -88 9401 -76 9435
rect -42 9401 -30 9435
rect -88 9367 -30 9401
rect -88 9333 -76 9367
rect -42 9333 -30 9367
rect -88 9299 -30 9333
rect -88 9265 -76 9299
rect -42 9265 -30 9299
rect -88 9231 -30 9265
rect -88 9197 -76 9231
rect -42 9197 -30 9231
rect -88 9163 -30 9197
rect -88 9129 -76 9163
rect -42 9129 -30 9163
rect -88 9095 -30 9129
rect -88 9061 -76 9095
rect -42 9061 -30 9095
rect -88 9027 -30 9061
rect -88 8993 -76 9027
rect -42 8993 -30 9027
rect -88 8959 -30 8993
rect -88 8925 -76 8959
rect -42 8925 -30 8959
rect -88 8891 -30 8925
rect -88 8857 -76 8891
rect -42 8857 -30 8891
rect -88 8823 -30 8857
rect -88 8789 -76 8823
rect -42 8789 -30 8823
rect -88 8755 -30 8789
rect -88 8721 -76 8755
rect -42 8721 -30 8755
rect -88 8687 -30 8721
rect -88 8653 -76 8687
rect -42 8653 -30 8687
rect -88 8619 -30 8653
rect -88 8585 -76 8619
rect -42 8585 -30 8619
rect -88 8551 -30 8585
rect -88 8517 -76 8551
rect -42 8517 -30 8551
rect -88 8483 -30 8517
rect -88 8449 -76 8483
rect -42 8449 -30 8483
rect -88 8415 -30 8449
rect -88 8381 -76 8415
rect -42 8381 -30 8415
rect -88 8347 -30 8381
rect -88 8313 -76 8347
rect -42 8313 -30 8347
rect -88 8279 -30 8313
rect -88 8245 -76 8279
rect -42 8245 -30 8279
rect -88 8211 -30 8245
rect -88 8177 -76 8211
rect -42 8177 -30 8211
rect -88 8143 -30 8177
rect -88 8109 -76 8143
rect -42 8109 -30 8143
rect -88 8075 -30 8109
rect -88 8041 -76 8075
rect -42 8041 -30 8075
rect -88 8007 -30 8041
rect -88 7973 -76 8007
rect -42 7973 -30 8007
rect -88 7939 -30 7973
rect -88 7905 -76 7939
rect -42 7905 -30 7939
rect -88 7871 -30 7905
rect -88 7837 -76 7871
rect -42 7837 -30 7871
rect -88 7803 -30 7837
rect -88 7769 -76 7803
rect -42 7769 -30 7803
rect -88 7735 -30 7769
rect -88 7701 -76 7735
rect -42 7701 -30 7735
rect -88 7667 -30 7701
rect -88 7633 -76 7667
rect -42 7633 -30 7667
rect -88 7599 -30 7633
rect -88 7565 -76 7599
rect -42 7565 -30 7599
rect -88 7531 -30 7565
rect -88 7497 -76 7531
rect -42 7497 -30 7531
rect -88 7463 -30 7497
rect -88 7429 -76 7463
rect -42 7429 -30 7463
rect -88 7395 -30 7429
rect -88 7361 -76 7395
rect -42 7361 -30 7395
rect -88 7327 -30 7361
rect -88 7293 -76 7327
rect -42 7293 -30 7327
rect -88 7259 -30 7293
rect -88 7225 -76 7259
rect -42 7225 -30 7259
rect -88 7191 -30 7225
rect -88 7157 -76 7191
rect -42 7157 -30 7191
rect -88 7123 -30 7157
rect -88 7089 -76 7123
rect -42 7089 -30 7123
rect -88 7055 -30 7089
rect -88 7021 -76 7055
rect -42 7021 -30 7055
rect -88 6987 -30 7021
rect -88 6953 -76 6987
rect -42 6953 -30 6987
rect -88 6919 -30 6953
rect -88 6885 -76 6919
rect -42 6885 -30 6919
rect -88 6851 -30 6885
rect -88 6817 -76 6851
rect -42 6817 -30 6851
rect -88 6783 -30 6817
rect -88 6749 -76 6783
rect -42 6749 -30 6783
rect -88 6715 -30 6749
rect -88 6681 -76 6715
rect -42 6681 -30 6715
rect -88 6647 -30 6681
rect -88 6613 -76 6647
rect -42 6613 -30 6647
rect -88 6579 -30 6613
rect -88 6545 -76 6579
rect -42 6545 -30 6579
rect -88 6511 -30 6545
rect -88 6477 -76 6511
rect -42 6477 -30 6511
rect -88 6443 -30 6477
rect -88 6409 -76 6443
rect -42 6409 -30 6443
rect -88 6375 -30 6409
rect -88 6341 -76 6375
rect -42 6341 -30 6375
rect -88 6307 -30 6341
rect -88 6273 -76 6307
rect -42 6273 -30 6307
rect -88 6239 -30 6273
rect -88 6205 -76 6239
rect -42 6205 -30 6239
rect -88 6171 -30 6205
rect -88 6137 -76 6171
rect -42 6137 -30 6171
rect -88 6103 -30 6137
rect -88 6069 -76 6103
rect -42 6069 -30 6103
rect -88 6035 -30 6069
rect -88 6001 -76 6035
rect -42 6001 -30 6035
rect -88 5967 -30 6001
rect -88 5933 -76 5967
rect -42 5933 -30 5967
rect -88 5899 -30 5933
rect -88 5865 -76 5899
rect -42 5865 -30 5899
rect -88 5831 -30 5865
rect -88 5797 -76 5831
rect -42 5797 -30 5831
rect -88 5763 -30 5797
rect -88 5729 -76 5763
rect -42 5729 -30 5763
rect -88 5695 -30 5729
rect -88 5661 -76 5695
rect -42 5661 -30 5695
rect -88 5627 -30 5661
rect -88 5593 -76 5627
rect -42 5593 -30 5627
rect -88 5559 -30 5593
rect -88 5525 -76 5559
rect -42 5525 -30 5559
rect -88 5491 -30 5525
rect -88 5457 -76 5491
rect -42 5457 -30 5491
rect -88 5423 -30 5457
rect -88 5389 -76 5423
rect -42 5389 -30 5423
rect -88 5355 -30 5389
rect -88 5321 -76 5355
rect -42 5321 -30 5355
rect -88 5287 -30 5321
rect -88 5253 -76 5287
rect -42 5253 -30 5287
rect -88 5219 -30 5253
rect -88 5185 -76 5219
rect -42 5185 -30 5219
rect -88 5151 -30 5185
rect -88 5117 -76 5151
rect -42 5117 -30 5151
rect -88 5083 -30 5117
rect -88 5049 -76 5083
rect -42 5049 -30 5083
rect -88 5015 -30 5049
rect -88 4981 -76 5015
rect -42 4981 -30 5015
rect -88 4947 -30 4981
rect -88 4913 -76 4947
rect -42 4913 -30 4947
rect -88 4879 -30 4913
rect -88 4845 -76 4879
rect -42 4845 -30 4879
rect -88 4811 -30 4845
rect -88 4777 -76 4811
rect -42 4777 -30 4811
rect -88 4743 -30 4777
rect -88 4709 -76 4743
rect -42 4709 -30 4743
rect -88 4675 -30 4709
rect -88 4641 -76 4675
rect -42 4641 -30 4675
rect -88 4607 -30 4641
rect -88 4573 -76 4607
rect -42 4573 -30 4607
rect -88 4539 -30 4573
rect -88 4505 -76 4539
rect -42 4505 -30 4539
rect -88 4471 -30 4505
rect -88 4437 -76 4471
rect -42 4437 -30 4471
rect -88 4403 -30 4437
rect -88 4369 -76 4403
rect -42 4369 -30 4403
rect -88 4335 -30 4369
rect -88 4301 -76 4335
rect -42 4301 -30 4335
rect -88 4267 -30 4301
rect -88 4233 -76 4267
rect -42 4233 -30 4267
rect -88 4199 -30 4233
rect -88 4165 -76 4199
rect -42 4165 -30 4199
rect -88 4131 -30 4165
rect -88 4097 -76 4131
rect -42 4097 -30 4131
rect -88 4063 -30 4097
rect -88 4029 -76 4063
rect -42 4029 -30 4063
rect -88 3995 -30 4029
rect -88 3961 -76 3995
rect -42 3961 -30 3995
rect -88 3927 -30 3961
rect -88 3893 -76 3927
rect -42 3893 -30 3927
rect -88 3859 -30 3893
rect -88 3825 -76 3859
rect -42 3825 -30 3859
rect -88 3791 -30 3825
rect -88 3757 -76 3791
rect -42 3757 -30 3791
rect -88 3723 -30 3757
rect -88 3689 -76 3723
rect -42 3689 -30 3723
rect -88 3655 -30 3689
rect -88 3621 -76 3655
rect -42 3621 -30 3655
rect -88 3587 -30 3621
rect -88 3553 -76 3587
rect -42 3553 -30 3587
rect -88 3519 -30 3553
rect -88 3485 -76 3519
rect -42 3485 -30 3519
rect -88 3451 -30 3485
rect -88 3417 -76 3451
rect -42 3417 -30 3451
rect -88 3383 -30 3417
rect -88 3349 -76 3383
rect -42 3349 -30 3383
rect -88 3315 -30 3349
rect -88 3281 -76 3315
rect -42 3281 -30 3315
rect -88 3247 -30 3281
rect -88 3213 -76 3247
rect -42 3213 -30 3247
rect -88 3179 -30 3213
rect -88 3145 -76 3179
rect -42 3145 -30 3179
rect -88 3111 -30 3145
rect -88 3077 -76 3111
rect -42 3077 -30 3111
rect -88 3043 -30 3077
rect -88 3009 -76 3043
rect -42 3009 -30 3043
rect -88 2975 -30 3009
rect -88 2941 -76 2975
rect -42 2941 -30 2975
rect -88 2907 -30 2941
rect -88 2873 -76 2907
rect -42 2873 -30 2907
rect -88 2839 -30 2873
rect -88 2805 -76 2839
rect -42 2805 -30 2839
rect -88 2771 -30 2805
rect -88 2737 -76 2771
rect -42 2737 -30 2771
rect -88 2703 -30 2737
rect -88 2669 -76 2703
rect -42 2669 -30 2703
rect -88 2635 -30 2669
rect -88 2601 -76 2635
rect -42 2601 -30 2635
rect -88 2567 -30 2601
rect -88 2533 -76 2567
rect -42 2533 -30 2567
rect -88 2499 -30 2533
rect -88 2465 -76 2499
rect -42 2465 -30 2499
rect -88 2431 -30 2465
rect -88 2397 -76 2431
rect -42 2397 -30 2431
rect -88 2363 -30 2397
rect -88 2329 -76 2363
rect -42 2329 -30 2363
rect -88 2295 -30 2329
rect -88 2261 -76 2295
rect -42 2261 -30 2295
rect -88 2227 -30 2261
rect -88 2193 -76 2227
rect -42 2193 -30 2227
rect -88 2159 -30 2193
rect -88 2125 -76 2159
rect -42 2125 -30 2159
rect -88 2091 -30 2125
rect -88 2057 -76 2091
rect -42 2057 -30 2091
rect -88 2023 -30 2057
rect -88 1989 -76 2023
rect -42 1989 -30 2023
rect -88 1955 -30 1989
rect -88 1921 -76 1955
rect -42 1921 -30 1955
rect -88 1887 -30 1921
rect -88 1853 -76 1887
rect -42 1853 -30 1887
rect -88 1819 -30 1853
rect -88 1785 -76 1819
rect -42 1785 -30 1819
rect -88 1751 -30 1785
rect -88 1717 -76 1751
rect -42 1717 -30 1751
rect -88 1683 -30 1717
rect -88 1649 -76 1683
rect -42 1649 -30 1683
rect -88 1615 -30 1649
rect -88 1581 -76 1615
rect -42 1581 -30 1615
rect -88 1547 -30 1581
rect -88 1513 -76 1547
rect -42 1513 -30 1547
rect -88 1479 -30 1513
rect -88 1445 -76 1479
rect -42 1445 -30 1479
rect -88 1411 -30 1445
rect -88 1377 -76 1411
rect -42 1377 -30 1411
rect -88 1343 -30 1377
rect -88 1309 -76 1343
rect -42 1309 -30 1343
rect -88 1275 -30 1309
rect -88 1241 -76 1275
rect -42 1241 -30 1275
rect -88 1207 -30 1241
rect -88 1173 -76 1207
rect -42 1173 -30 1207
rect -88 1139 -30 1173
rect -88 1105 -76 1139
rect -42 1105 -30 1139
rect -88 1071 -30 1105
rect -88 1037 -76 1071
rect -42 1037 -30 1071
rect -88 1003 -30 1037
rect -88 969 -76 1003
rect -42 969 -30 1003
rect -88 935 -30 969
rect -88 901 -76 935
rect -42 901 -30 935
rect -88 867 -30 901
rect -88 833 -76 867
rect -42 833 -30 867
rect -88 799 -30 833
rect -88 765 -76 799
rect -42 765 -30 799
rect -88 731 -30 765
rect -88 697 -76 731
rect -42 697 -30 731
rect -88 663 -30 697
rect -88 629 -76 663
rect -42 629 -30 663
rect -88 595 -30 629
rect -88 561 -76 595
rect -42 561 -30 595
rect -88 527 -30 561
rect -88 493 -76 527
rect -42 493 -30 527
rect -88 459 -30 493
rect -88 425 -76 459
rect -42 425 -30 459
rect -88 391 -30 425
rect -88 357 -76 391
rect -42 357 -30 391
rect -88 323 -30 357
rect -88 289 -76 323
rect -42 289 -30 323
rect -88 255 -30 289
rect -88 221 -76 255
rect -42 221 -30 255
rect -88 187 -30 221
rect -88 153 -76 187
rect -42 153 -30 187
rect -88 119 -30 153
rect -88 85 -76 119
rect -42 85 -30 119
rect -88 51 -30 85
rect -88 17 -76 51
rect -42 17 -30 51
rect -88 -17 -30 17
rect -88 -51 -76 -17
rect -42 -51 -30 -17
rect -88 -85 -30 -51
rect -88 -119 -76 -85
rect -42 -119 -30 -85
rect -88 -153 -30 -119
rect -88 -187 -76 -153
rect -42 -187 -30 -153
rect -88 -221 -30 -187
rect -88 -255 -76 -221
rect -42 -255 -30 -221
rect -88 -289 -30 -255
rect -88 -323 -76 -289
rect -42 -323 -30 -289
rect -88 -357 -30 -323
rect -88 -391 -76 -357
rect -42 -391 -30 -357
rect -88 -425 -30 -391
rect -88 -459 -76 -425
rect -42 -459 -30 -425
rect -88 -493 -30 -459
rect -88 -527 -76 -493
rect -42 -527 -30 -493
rect -88 -561 -30 -527
rect -88 -595 -76 -561
rect -42 -595 -30 -561
rect -88 -629 -30 -595
rect -88 -663 -76 -629
rect -42 -663 -30 -629
rect -88 -697 -30 -663
rect -88 -731 -76 -697
rect -42 -731 -30 -697
rect -88 -765 -30 -731
rect -88 -799 -76 -765
rect -42 -799 -30 -765
rect -88 -833 -30 -799
rect -88 -867 -76 -833
rect -42 -867 -30 -833
rect -88 -901 -30 -867
rect -88 -935 -76 -901
rect -42 -935 -30 -901
rect -88 -969 -30 -935
rect -88 -1003 -76 -969
rect -42 -1003 -30 -969
rect -88 -1037 -30 -1003
rect -88 -1071 -76 -1037
rect -42 -1071 -30 -1037
rect -88 -1105 -30 -1071
rect -88 -1139 -76 -1105
rect -42 -1139 -30 -1105
rect -88 -1173 -30 -1139
rect -88 -1207 -76 -1173
rect -42 -1207 -30 -1173
rect -88 -1241 -30 -1207
rect -88 -1275 -76 -1241
rect -42 -1275 -30 -1241
rect -88 -1309 -30 -1275
rect -88 -1343 -76 -1309
rect -42 -1343 -30 -1309
rect -88 -1377 -30 -1343
rect -88 -1411 -76 -1377
rect -42 -1411 -30 -1377
rect -88 -1445 -30 -1411
rect -88 -1479 -76 -1445
rect -42 -1479 -30 -1445
rect -88 -1513 -30 -1479
rect -88 -1547 -76 -1513
rect -42 -1547 -30 -1513
rect -88 -1581 -30 -1547
rect -88 -1615 -76 -1581
rect -42 -1615 -30 -1581
rect -88 -1649 -30 -1615
rect -88 -1683 -76 -1649
rect -42 -1683 -30 -1649
rect -88 -1717 -30 -1683
rect -88 -1751 -76 -1717
rect -42 -1751 -30 -1717
rect -88 -1785 -30 -1751
rect -88 -1819 -76 -1785
rect -42 -1819 -30 -1785
rect -88 -1853 -30 -1819
rect -88 -1887 -76 -1853
rect -42 -1887 -30 -1853
rect -88 -1921 -30 -1887
rect -88 -1955 -76 -1921
rect -42 -1955 -30 -1921
rect -88 -1989 -30 -1955
rect -88 -2023 -76 -1989
rect -42 -2023 -30 -1989
rect -88 -2057 -30 -2023
rect -88 -2091 -76 -2057
rect -42 -2091 -30 -2057
rect -88 -2125 -30 -2091
rect -88 -2159 -76 -2125
rect -42 -2159 -30 -2125
rect -88 -2193 -30 -2159
rect -88 -2227 -76 -2193
rect -42 -2227 -30 -2193
rect -88 -2261 -30 -2227
rect -88 -2295 -76 -2261
rect -42 -2295 -30 -2261
rect -88 -2329 -30 -2295
rect -88 -2363 -76 -2329
rect -42 -2363 -30 -2329
rect -88 -2397 -30 -2363
rect -88 -2431 -76 -2397
rect -42 -2431 -30 -2397
rect -88 -2465 -30 -2431
rect -88 -2499 -76 -2465
rect -42 -2499 -30 -2465
rect -88 -2533 -30 -2499
rect -88 -2567 -76 -2533
rect -42 -2567 -30 -2533
rect -88 -2601 -30 -2567
rect -88 -2635 -76 -2601
rect -42 -2635 -30 -2601
rect -88 -2669 -30 -2635
rect -88 -2703 -76 -2669
rect -42 -2703 -30 -2669
rect -88 -2737 -30 -2703
rect -88 -2771 -76 -2737
rect -42 -2771 -30 -2737
rect -88 -2805 -30 -2771
rect -88 -2839 -76 -2805
rect -42 -2839 -30 -2805
rect -88 -2873 -30 -2839
rect -88 -2907 -76 -2873
rect -42 -2907 -30 -2873
rect -88 -2941 -30 -2907
rect -88 -2975 -76 -2941
rect -42 -2975 -30 -2941
rect -88 -3009 -30 -2975
rect -88 -3043 -76 -3009
rect -42 -3043 -30 -3009
rect -88 -3077 -30 -3043
rect -88 -3111 -76 -3077
rect -42 -3111 -30 -3077
rect -88 -3145 -30 -3111
rect -88 -3179 -76 -3145
rect -42 -3179 -30 -3145
rect -88 -3213 -30 -3179
rect -88 -3247 -76 -3213
rect -42 -3247 -30 -3213
rect -88 -3281 -30 -3247
rect -88 -3315 -76 -3281
rect -42 -3315 -30 -3281
rect -88 -3349 -30 -3315
rect -88 -3383 -76 -3349
rect -42 -3383 -30 -3349
rect -88 -3417 -30 -3383
rect -88 -3451 -76 -3417
rect -42 -3451 -30 -3417
rect -88 -3485 -30 -3451
rect -88 -3519 -76 -3485
rect -42 -3519 -30 -3485
rect -88 -3553 -30 -3519
rect -88 -3587 -76 -3553
rect -42 -3587 -30 -3553
rect -88 -3621 -30 -3587
rect -88 -3655 -76 -3621
rect -42 -3655 -30 -3621
rect -88 -3689 -30 -3655
rect -88 -3723 -76 -3689
rect -42 -3723 -30 -3689
rect -88 -3757 -30 -3723
rect -88 -3791 -76 -3757
rect -42 -3791 -30 -3757
rect -88 -3825 -30 -3791
rect -88 -3859 -76 -3825
rect -42 -3859 -30 -3825
rect -88 -3893 -30 -3859
rect -88 -3927 -76 -3893
rect -42 -3927 -30 -3893
rect -88 -3961 -30 -3927
rect -88 -3995 -76 -3961
rect -42 -3995 -30 -3961
rect -88 -4029 -30 -3995
rect -88 -4063 -76 -4029
rect -42 -4063 -30 -4029
rect -88 -4097 -30 -4063
rect -88 -4131 -76 -4097
rect -42 -4131 -30 -4097
rect -88 -4165 -30 -4131
rect -88 -4199 -76 -4165
rect -42 -4199 -30 -4165
rect -88 -4233 -30 -4199
rect -88 -4267 -76 -4233
rect -42 -4267 -30 -4233
rect -88 -4301 -30 -4267
rect -88 -4335 -76 -4301
rect -42 -4335 -30 -4301
rect -88 -4369 -30 -4335
rect -88 -4403 -76 -4369
rect -42 -4403 -30 -4369
rect -88 -4437 -30 -4403
rect -88 -4471 -76 -4437
rect -42 -4471 -30 -4437
rect -88 -4505 -30 -4471
rect -88 -4539 -76 -4505
rect -42 -4539 -30 -4505
rect -88 -4573 -30 -4539
rect -88 -4607 -76 -4573
rect -42 -4607 -30 -4573
rect -88 -4641 -30 -4607
rect -88 -4675 -76 -4641
rect -42 -4675 -30 -4641
rect -88 -4709 -30 -4675
rect -88 -4743 -76 -4709
rect -42 -4743 -30 -4709
rect -88 -4777 -30 -4743
rect -88 -4811 -76 -4777
rect -42 -4811 -30 -4777
rect -88 -4845 -30 -4811
rect -88 -4879 -76 -4845
rect -42 -4879 -30 -4845
rect -88 -4913 -30 -4879
rect -88 -4947 -76 -4913
rect -42 -4947 -30 -4913
rect -88 -4981 -30 -4947
rect -88 -5015 -76 -4981
rect -42 -5015 -30 -4981
rect -88 -5049 -30 -5015
rect -88 -5083 -76 -5049
rect -42 -5083 -30 -5049
rect -88 -5117 -30 -5083
rect -88 -5151 -76 -5117
rect -42 -5151 -30 -5117
rect -88 -5185 -30 -5151
rect -88 -5219 -76 -5185
rect -42 -5219 -30 -5185
rect -88 -5253 -30 -5219
rect -88 -5287 -76 -5253
rect -42 -5287 -30 -5253
rect -88 -5321 -30 -5287
rect -88 -5355 -76 -5321
rect -42 -5355 -30 -5321
rect -88 -5389 -30 -5355
rect -88 -5423 -76 -5389
rect -42 -5423 -30 -5389
rect -88 -5457 -30 -5423
rect -88 -5491 -76 -5457
rect -42 -5491 -30 -5457
rect -88 -5525 -30 -5491
rect -88 -5559 -76 -5525
rect -42 -5559 -30 -5525
rect -88 -5593 -30 -5559
rect -88 -5627 -76 -5593
rect -42 -5627 -30 -5593
rect -88 -5661 -30 -5627
rect -88 -5695 -76 -5661
rect -42 -5695 -30 -5661
rect -88 -5729 -30 -5695
rect -88 -5763 -76 -5729
rect -42 -5763 -30 -5729
rect -88 -5797 -30 -5763
rect -88 -5831 -76 -5797
rect -42 -5831 -30 -5797
rect -88 -5865 -30 -5831
rect -88 -5899 -76 -5865
rect -42 -5899 -30 -5865
rect -88 -5933 -30 -5899
rect -88 -5967 -76 -5933
rect -42 -5967 -30 -5933
rect -88 -6001 -30 -5967
rect -88 -6035 -76 -6001
rect -42 -6035 -30 -6001
rect -88 -6069 -30 -6035
rect -88 -6103 -76 -6069
rect -42 -6103 -30 -6069
rect -88 -6137 -30 -6103
rect -88 -6171 -76 -6137
rect -42 -6171 -30 -6137
rect -88 -6205 -30 -6171
rect -88 -6239 -76 -6205
rect -42 -6239 -30 -6205
rect -88 -6273 -30 -6239
rect -88 -6307 -76 -6273
rect -42 -6307 -30 -6273
rect -88 -6341 -30 -6307
rect -88 -6375 -76 -6341
rect -42 -6375 -30 -6341
rect -88 -6409 -30 -6375
rect -88 -6443 -76 -6409
rect -42 -6443 -30 -6409
rect -88 -6477 -30 -6443
rect -88 -6511 -76 -6477
rect -42 -6511 -30 -6477
rect -88 -6545 -30 -6511
rect -88 -6579 -76 -6545
rect -42 -6579 -30 -6545
rect -88 -6613 -30 -6579
rect -88 -6647 -76 -6613
rect -42 -6647 -30 -6613
rect -88 -6681 -30 -6647
rect -88 -6715 -76 -6681
rect -42 -6715 -30 -6681
rect -88 -6749 -30 -6715
rect -88 -6783 -76 -6749
rect -42 -6783 -30 -6749
rect -88 -6817 -30 -6783
rect -88 -6851 -76 -6817
rect -42 -6851 -30 -6817
rect -88 -6885 -30 -6851
rect -88 -6919 -76 -6885
rect -42 -6919 -30 -6885
rect -88 -6953 -30 -6919
rect -88 -6987 -76 -6953
rect -42 -6987 -30 -6953
rect -88 -7021 -30 -6987
rect -88 -7055 -76 -7021
rect -42 -7055 -30 -7021
rect -88 -7089 -30 -7055
rect -88 -7123 -76 -7089
rect -42 -7123 -30 -7089
rect -88 -7157 -30 -7123
rect -88 -7191 -76 -7157
rect -42 -7191 -30 -7157
rect -88 -7225 -30 -7191
rect -88 -7259 -76 -7225
rect -42 -7259 -30 -7225
rect -88 -7293 -30 -7259
rect -88 -7327 -76 -7293
rect -42 -7327 -30 -7293
rect -88 -7361 -30 -7327
rect -88 -7395 -76 -7361
rect -42 -7395 -30 -7361
rect -88 -7429 -30 -7395
rect -88 -7463 -76 -7429
rect -42 -7463 -30 -7429
rect -88 -7497 -30 -7463
rect -88 -7531 -76 -7497
rect -42 -7531 -30 -7497
rect -88 -7565 -30 -7531
rect -88 -7599 -76 -7565
rect -42 -7599 -30 -7565
rect -88 -7633 -30 -7599
rect -88 -7667 -76 -7633
rect -42 -7667 -30 -7633
rect -88 -7701 -30 -7667
rect -88 -7735 -76 -7701
rect -42 -7735 -30 -7701
rect -88 -7769 -30 -7735
rect -88 -7803 -76 -7769
rect -42 -7803 -30 -7769
rect -88 -7837 -30 -7803
rect -88 -7871 -76 -7837
rect -42 -7871 -30 -7837
rect -88 -7905 -30 -7871
rect -88 -7939 -76 -7905
rect -42 -7939 -30 -7905
rect -88 -7973 -30 -7939
rect -88 -8007 -76 -7973
rect -42 -8007 -30 -7973
rect -88 -8041 -30 -8007
rect -88 -8075 -76 -8041
rect -42 -8075 -30 -8041
rect -88 -8109 -30 -8075
rect -88 -8143 -76 -8109
rect -42 -8143 -30 -8109
rect -88 -8177 -30 -8143
rect -88 -8211 -76 -8177
rect -42 -8211 -30 -8177
rect -88 -8245 -30 -8211
rect -88 -8279 -76 -8245
rect -42 -8279 -30 -8245
rect -88 -8313 -30 -8279
rect -88 -8347 -76 -8313
rect -42 -8347 -30 -8313
rect -88 -8381 -30 -8347
rect -88 -8415 -76 -8381
rect -42 -8415 -30 -8381
rect -88 -8449 -30 -8415
rect -88 -8483 -76 -8449
rect -42 -8483 -30 -8449
rect -88 -8517 -30 -8483
rect -88 -8551 -76 -8517
rect -42 -8551 -30 -8517
rect -88 -8585 -30 -8551
rect -88 -8619 -76 -8585
rect -42 -8619 -30 -8585
rect -88 -8653 -30 -8619
rect -88 -8687 -76 -8653
rect -42 -8687 -30 -8653
rect -88 -8721 -30 -8687
rect -88 -8755 -76 -8721
rect -42 -8755 -30 -8721
rect -88 -8789 -30 -8755
rect -88 -8823 -76 -8789
rect -42 -8823 -30 -8789
rect -88 -8857 -30 -8823
rect -88 -8891 -76 -8857
rect -42 -8891 -30 -8857
rect -88 -8925 -30 -8891
rect -88 -8959 -76 -8925
rect -42 -8959 -30 -8925
rect -88 -8993 -30 -8959
rect -88 -9027 -76 -8993
rect -42 -9027 -30 -8993
rect -88 -9061 -30 -9027
rect -88 -9095 -76 -9061
rect -42 -9095 -30 -9061
rect -88 -9129 -30 -9095
rect -88 -9163 -76 -9129
rect -42 -9163 -30 -9129
rect -88 -9197 -30 -9163
rect -88 -9231 -76 -9197
rect -42 -9231 -30 -9197
rect -88 -9265 -30 -9231
rect -88 -9299 -76 -9265
rect -42 -9299 -30 -9265
rect -88 -9333 -30 -9299
rect -88 -9367 -76 -9333
rect -42 -9367 -30 -9333
rect -88 -9401 -30 -9367
rect -88 -9435 -76 -9401
rect -42 -9435 -30 -9401
rect -88 -9469 -30 -9435
rect -88 -9503 -76 -9469
rect -42 -9503 -30 -9469
rect -88 -9537 -30 -9503
rect -88 -9571 -76 -9537
rect -42 -9571 -30 -9537
rect -88 -9600 -30 -9571
rect 30 9571 88 9600
rect 30 9537 42 9571
rect 76 9537 88 9571
rect 30 9503 88 9537
rect 30 9469 42 9503
rect 76 9469 88 9503
rect 30 9435 88 9469
rect 30 9401 42 9435
rect 76 9401 88 9435
rect 30 9367 88 9401
rect 30 9333 42 9367
rect 76 9333 88 9367
rect 30 9299 88 9333
rect 30 9265 42 9299
rect 76 9265 88 9299
rect 30 9231 88 9265
rect 30 9197 42 9231
rect 76 9197 88 9231
rect 30 9163 88 9197
rect 30 9129 42 9163
rect 76 9129 88 9163
rect 30 9095 88 9129
rect 30 9061 42 9095
rect 76 9061 88 9095
rect 30 9027 88 9061
rect 30 8993 42 9027
rect 76 8993 88 9027
rect 30 8959 88 8993
rect 30 8925 42 8959
rect 76 8925 88 8959
rect 30 8891 88 8925
rect 30 8857 42 8891
rect 76 8857 88 8891
rect 30 8823 88 8857
rect 30 8789 42 8823
rect 76 8789 88 8823
rect 30 8755 88 8789
rect 30 8721 42 8755
rect 76 8721 88 8755
rect 30 8687 88 8721
rect 30 8653 42 8687
rect 76 8653 88 8687
rect 30 8619 88 8653
rect 30 8585 42 8619
rect 76 8585 88 8619
rect 30 8551 88 8585
rect 30 8517 42 8551
rect 76 8517 88 8551
rect 30 8483 88 8517
rect 30 8449 42 8483
rect 76 8449 88 8483
rect 30 8415 88 8449
rect 30 8381 42 8415
rect 76 8381 88 8415
rect 30 8347 88 8381
rect 30 8313 42 8347
rect 76 8313 88 8347
rect 30 8279 88 8313
rect 30 8245 42 8279
rect 76 8245 88 8279
rect 30 8211 88 8245
rect 30 8177 42 8211
rect 76 8177 88 8211
rect 30 8143 88 8177
rect 30 8109 42 8143
rect 76 8109 88 8143
rect 30 8075 88 8109
rect 30 8041 42 8075
rect 76 8041 88 8075
rect 30 8007 88 8041
rect 30 7973 42 8007
rect 76 7973 88 8007
rect 30 7939 88 7973
rect 30 7905 42 7939
rect 76 7905 88 7939
rect 30 7871 88 7905
rect 30 7837 42 7871
rect 76 7837 88 7871
rect 30 7803 88 7837
rect 30 7769 42 7803
rect 76 7769 88 7803
rect 30 7735 88 7769
rect 30 7701 42 7735
rect 76 7701 88 7735
rect 30 7667 88 7701
rect 30 7633 42 7667
rect 76 7633 88 7667
rect 30 7599 88 7633
rect 30 7565 42 7599
rect 76 7565 88 7599
rect 30 7531 88 7565
rect 30 7497 42 7531
rect 76 7497 88 7531
rect 30 7463 88 7497
rect 30 7429 42 7463
rect 76 7429 88 7463
rect 30 7395 88 7429
rect 30 7361 42 7395
rect 76 7361 88 7395
rect 30 7327 88 7361
rect 30 7293 42 7327
rect 76 7293 88 7327
rect 30 7259 88 7293
rect 30 7225 42 7259
rect 76 7225 88 7259
rect 30 7191 88 7225
rect 30 7157 42 7191
rect 76 7157 88 7191
rect 30 7123 88 7157
rect 30 7089 42 7123
rect 76 7089 88 7123
rect 30 7055 88 7089
rect 30 7021 42 7055
rect 76 7021 88 7055
rect 30 6987 88 7021
rect 30 6953 42 6987
rect 76 6953 88 6987
rect 30 6919 88 6953
rect 30 6885 42 6919
rect 76 6885 88 6919
rect 30 6851 88 6885
rect 30 6817 42 6851
rect 76 6817 88 6851
rect 30 6783 88 6817
rect 30 6749 42 6783
rect 76 6749 88 6783
rect 30 6715 88 6749
rect 30 6681 42 6715
rect 76 6681 88 6715
rect 30 6647 88 6681
rect 30 6613 42 6647
rect 76 6613 88 6647
rect 30 6579 88 6613
rect 30 6545 42 6579
rect 76 6545 88 6579
rect 30 6511 88 6545
rect 30 6477 42 6511
rect 76 6477 88 6511
rect 30 6443 88 6477
rect 30 6409 42 6443
rect 76 6409 88 6443
rect 30 6375 88 6409
rect 30 6341 42 6375
rect 76 6341 88 6375
rect 30 6307 88 6341
rect 30 6273 42 6307
rect 76 6273 88 6307
rect 30 6239 88 6273
rect 30 6205 42 6239
rect 76 6205 88 6239
rect 30 6171 88 6205
rect 30 6137 42 6171
rect 76 6137 88 6171
rect 30 6103 88 6137
rect 30 6069 42 6103
rect 76 6069 88 6103
rect 30 6035 88 6069
rect 30 6001 42 6035
rect 76 6001 88 6035
rect 30 5967 88 6001
rect 30 5933 42 5967
rect 76 5933 88 5967
rect 30 5899 88 5933
rect 30 5865 42 5899
rect 76 5865 88 5899
rect 30 5831 88 5865
rect 30 5797 42 5831
rect 76 5797 88 5831
rect 30 5763 88 5797
rect 30 5729 42 5763
rect 76 5729 88 5763
rect 30 5695 88 5729
rect 30 5661 42 5695
rect 76 5661 88 5695
rect 30 5627 88 5661
rect 30 5593 42 5627
rect 76 5593 88 5627
rect 30 5559 88 5593
rect 30 5525 42 5559
rect 76 5525 88 5559
rect 30 5491 88 5525
rect 30 5457 42 5491
rect 76 5457 88 5491
rect 30 5423 88 5457
rect 30 5389 42 5423
rect 76 5389 88 5423
rect 30 5355 88 5389
rect 30 5321 42 5355
rect 76 5321 88 5355
rect 30 5287 88 5321
rect 30 5253 42 5287
rect 76 5253 88 5287
rect 30 5219 88 5253
rect 30 5185 42 5219
rect 76 5185 88 5219
rect 30 5151 88 5185
rect 30 5117 42 5151
rect 76 5117 88 5151
rect 30 5083 88 5117
rect 30 5049 42 5083
rect 76 5049 88 5083
rect 30 5015 88 5049
rect 30 4981 42 5015
rect 76 4981 88 5015
rect 30 4947 88 4981
rect 30 4913 42 4947
rect 76 4913 88 4947
rect 30 4879 88 4913
rect 30 4845 42 4879
rect 76 4845 88 4879
rect 30 4811 88 4845
rect 30 4777 42 4811
rect 76 4777 88 4811
rect 30 4743 88 4777
rect 30 4709 42 4743
rect 76 4709 88 4743
rect 30 4675 88 4709
rect 30 4641 42 4675
rect 76 4641 88 4675
rect 30 4607 88 4641
rect 30 4573 42 4607
rect 76 4573 88 4607
rect 30 4539 88 4573
rect 30 4505 42 4539
rect 76 4505 88 4539
rect 30 4471 88 4505
rect 30 4437 42 4471
rect 76 4437 88 4471
rect 30 4403 88 4437
rect 30 4369 42 4403
rect 76 4369 88 4403
rect 30 4335 88 4369
rect 30 4301 42 4335
rect 76 4301 88 4335
rect 30 4267 88 4301
rect 30 4233 42 4267
rect 76 4233 88 4267
rect 30 4199 88 4233
rect 30 4165 42 4199
rect 76 4165 88 4199
rect 30 4131 88 4165
rect 30 4097 42 4131
rect 76 4097 88 4131
rect 30 4063 88 4097
rect 30 4029 42 4063
rect 76 4029 88 4063
rect 30 3995 88 4029
rect 30 3961 42 3995
rect 76 3961 88 3995
rect 30 3927 88 3961
rect 30 3893 42 3927
rect 76 3893 88 3927
rect 30 3859 88 3893
rect 30 3825 42 3859
rect 76 3825 88 3859
rect 30 3791 88 3825
rect 30 3757 42 3791
rect 76 3757 88 3791
rect 30 3723 88 3757
rect 30 3689 42 3723
rect 76 3689 88 3723
rect 30 3655 88 3689
rect 30 3621 42 3655
rect 76 3621 88 3655
rect 30 3587 88 3621
rect 30 3553 42 3587
rect 76 3553 88 3587
rect 30 3519 88 3553
rect 30 3485 42 3519
rect 76 3485 88 3519
rect 30 3451 88 3485
rect 30 3417 42 3451
rect 76 3417 88 3451
rect 30 3383 88 3417
rect 30 3349 42 3383
rect 76 3349 88 3383
rect 30 3315 88 3349
rect 30 3281 42 3315
rect 76 3281 88 3315
rect 30 3247 88 3281
rect 30 3213 42 3247
rect 76 3213 88 3247
rect 30 3179 88 3213
rect 30 3145 42 3179
rect 76 3145 88 3179
rect 30 3111 88 3145
rect 30 3077 42 3111
rect 76 3077 88 3111
rect 30 3043 88 3077
rect 30 3009 42 3043
rect 76 3009 88 3043
rect 30 2975 88 3009
rect 30 2941 42 2975
rect 76 2941 88 2975
rect 30 2907 88 2941
rect 30 2873 42 2907
rect 76 2873 88 2907
rect 30 2839 88 2873
rect 30 2805 42 2839
rect 76 2805 88 2839
rect 30 2771 88 2805
rect 30 2737 42 2771
rect 76 2737 88 2771
rect 30 2703 88 2737
rect 30 2669 42 2703
rect 76 2669 88 2703
rect 30 2635 88 2669
rect 30 2601 42 2635
rect 76 2601 88 2635
rect 30 2567 88 2601
rect 30 2533 42 2567
rect 76 2533 88 2567
rect 30 2499 88 2533
rect 30 2465 42 2499
rect 76 2465 88 2499
rect 30 2431 88 2465
rect 30 2397 42 2431
rect 76 2397 88 2431
rect 30 2363 88 2397
rect 30 2329 42 2363
rect 76 2329 88 2363
rect 30 2295 88 2329
rect 30 2261 42 2295
rect 76 2261 88 2295
rect 30 2227 88 2261
rect 30 2193 42 2227
rect 76 2193 88 2227
rect 30 2159 88 2193
rect 30 2125 42 2159
rect 76 2125 88 2159
rect 30 2091 88 2125
rect 30 2057 42 2091
rect 76 2057 88 2091
rect 30 2023 88 2057
rect 30 1989 42 2023
rect 76 1989 88 2023
rect 30 1955 88 1989
rect 30 1921 42 1955
rect 76 1921 88 1955
rect 30 1887 88 1921
rect 30 1853 42 1887
rect 76 1853 88 1887
rect 30 1819 88 1853
rect 30 1785 42 1819
rect 76 1785 88 1819
rect 30 1751 88 1785
rect 30 1717 42 1751
rect 76 1717 88 1751
rect 30 1683 88 1717
rect 30 1649 42 1683
rect 76 1649 88 1683
rect 30 1615 88 1649
rect 30 1581 42 1615
rect 76 1581 88 1615
rect 30 1547 88 1581
rect 30 1513 42 1547
rect 76 1513 88 1547
rect 30 1479 88 1513
rect 30 1445 42 1479
rect 76 1445 88 1479
rect 30 1411 88 1445
rect 30 1377 42 1411
rect 76 1377 88 1411
rect 30 1343 88 1377
rect 30 1309 42 1343
rect 76 1309 88 1343
rect 30 1275 88 1309
rect 30 1241 42 1275
rect 76 1241 88 1275
rect 30 1207 88 1241
rect 30 1173 42 1207
rect 76 1173 88 1207
rect 30 1139 88 1173
rect 30 1105 42 1139
rect 76 1105 88 1139
rect 30 1071 88 1105
rect 30 1037 42 1071
rect 76 1037 88 1071
rect 30 1003 88 1037
rect 30 969 42 1003
rect 76 969 88 1003
rect 30 935 88 969
rect 30 901 42 935
rect 76 901 88 935
rect 30 867 88 901
rect 30 833 42 867
rect 76 833 88 867
rect 30 799 88 833
rect 30 765 42 799
rect 76 765 88 799
rect 30 731 88 765
rect 30 697 42 731
rect 76 697 88 731
rect 30 663 88 697
rect 30 629 42 663
rect 76 629 88 663
rect 30 595 88 629
rect 30 561 42 595
rect 76 561 88 595
rect 30 527 88 561
rect 30 493 42 527
rect 76 493 88 527
rect 30 459 88 493
rect 30 425 42 459
rect 76 425 88 459
rect 30 391 88 425
rect 30 357 42 391
rect 76 357 88 391
rect 30 323 88 357
rect 30 289 42 323
rect 76 289 88 323
rect 30 255 88 289
rect 30 221 42 255
rect 76 221 88 255
rect 30 187 88 221
rect 30 153 42 187
rect 76 153 88 187
rect 30 119 88 153
rect 30 85 42 119
rect 76 85 88 119
rect 30 51 88 85
rect 30 17 42 51
rect 76 17 88 51
rect 30 -17 88 17
rect 30 -51 42 -17
rect 76 -51 88 -17
rect 30 -85 88 -51
rect 30 -119 42 -85
rect 76 -119 88 -85
rect 30 -153 88 -119
rect 30 -187 42 -153
rect 76 -187 88 -153
rect 30 -221 88 -187
rect 30 -255 42 -221
rect 76 -255 88 -221
rect 30 -289 88 -255
rect 30 -323 42 -289
rect 76 -323 88 -289
rect 30 -357 88 -323
rect 30 -391 42 -357
rect 76 -391 88 -357
rect 30 -425 88 -391
rect 30 -459 42 -425
rect 76 -459 88 -425
rect 30 -493 88 -459
rect 30 -527 42 -493
rect 76 -527 88 -493
rect 30 -561 88 -527
rect 30 -595 42 -561
rect 76 -595 88 -561
rect 30 -629 88 -595
rect 30 -663 42 -629
rect 76 -663 88 -629
rect 30 -697 88 -663
rect 30 -731 42 -697
rect 76 -731 88 -697
rect 30 -765 88 -731
rect 30 -799 42 -765
rect 76 -799 88 -765
rect 30 -833 88 -799
rect 30 -867 42 -833
rect 76 -867 88 -833
rect 30 -901 88 -867
rect 30 -935 42 -901
rect 76 -935 88 -901
rect 30 -969 88 -935
rect 30 -1003 42 -969
rect 76 -1003 88 -969
rect 30 -1037 88 -1003
rect 30 -1071 42 -1037
rect 76 -1071 88 -1037
rect 30 -1105 88 -1071
rect 30 -1139 42 -1105
rect 76 -1139 88 -1105
rect 30 -1173 88 -1139
rect 30 -1207 42 -1173
rect 76 -1207 88 -1173
rect 30 -1241 88 -1207
rect 30 -1275 42 -1241
rect 76 -1275 88 -1241
rect 30 -1309 88 -1275
rect 30 -1343 42 -1309
rect 76 -1343 88 -1309
rect 30 -1377 88 -1343
rect 30 -1411 42 -1377
rect 76 -1411 88 -1377
rect 30 -1445 88 -1411
rect 30 -1479 42 -1445
rect 76 -1479 88 -1445
rect 30 -1513 88 -1479
rect 30 -1547 42 -1513
rect 76 -1547 88 -1513
rect 30 -1581 88 -1547
rect 30 -1615 42 -1581
rect 76 -1615 88 -1581
rect 30 -1649 88 -1615
rect 30 -1683 42 -1649
rect 76 -1683 88 -1649
rect 30 -1717 88 -1683
rect 30 -1751 42 -1717
rect 76 -1751 88 -1717
rect 30 -1785 88 -1751
rect 30 -1819 42 -1785
rect 76 -1819 88 -1785
rect 30 -1853 88 -1819
rect 30 -1887 42 -1853
rect 76 -1887 88 -1853
rect 30 -1921 88 -1887
rect 30 -1955 42 -1921
rect 76 -1955 88 -1921
rect 30 -1989 88 -1955
rect 30 -2023 42 -1989
rect 76 -2023 88 -1989
rect 30 -2057 88 -2023
rect 30 -2091 42 -2057
rect 76 -2091 88 -2057
rect 30 -2125 88 -2091
rect 30 -2159 42 -2125
rect 76 -2159 88 -2125
rect 30 -2193 88 -2159
rect 30 -2227 42 -2193
rect 76 -2227 88 -2193
rect 30 -2261 88 -2227
rect 30 -2295 42 -2261
rect 76 -2295 88 -2261
rect 30 -2329 88 -2295
rect 30 -2363 42 -2329
rect 76 -2363 88 -2329
rect 30 -2397 88 -2363
rect 30 -2431 42 -2397
rect 76 -2431 88 -2397
rect 30 -2465 88 -2431
rect 30 -2499 42 -2465
rect 76 -2499 88 -2465
rect 30 -2533 88 -2499
rect 30 -2567 42 -2533
rect 76 -2567 88 -2533
rect 30 -2601 88 -2567
rect 30 -2635 42 -2601
rect 76 -2635 88 -2601
rect 30 -2669 88 -2635
rect 30 -2703 42 -2669
rect 76 -2703 88 -2669
rect 30 -2737 88 -2703
rect 30 -2771 42 -2737
rect 76 -2771 88 -2737
rect 30 -2805 88 -2771
rect 30 -2839 42 -2805
rect 76 -2839 88 -2805
rect 30 -2873 88 -2839
rect 30 -2907 42 -2873
rect 76 -2907 88 -2873
rect 30 -2941 88 -2907
rect 30 -2975 42 -2941
rect 76 -2975 88 -2941
rect 30 -3009 88 -2975
rect 30 -3043 42 -3009
rect 76 -3043 88 -3009
rect 30 -3077 88 -3043
rect 30 -3111 42 -3077
rect 76 -3111 88 -3077
rect 30 -3145 88 -3111
rect 30 -3179 42 -3145
rect 76 -3179 88 -3145
rect 30 -3213 88 -3179
rect 30 -3247 42 -3213
rect 76 -3247 88 -3213
rect 30 -3281 88 -3247
rect 30 -3315 42 -3281
rect 76 -3315 88 -3281
rect 30 -3349 88 -3315
rect 30 -3383 42 -3349
rect 76 -3383 88 -3349
rect 30 -3417 88 -3383
rect 30 -3451 42 -3417
rect 76 -3451 88 -3417
rect 30 -3485 88 -3451
rect 30 -3519 42 -3485
rect 76 -3519 88 -3485
rect 30 -3553 88 -3519
rect 30 -3587 42 -3553
rect 76 -3587 88 -3553
rect 30 -3621 88 -3587
rect 30 -3655 42 -3621
rect 76 -3655 88 -3621
rect 30 -3689 88 -3655
rect 30 -3723 42 -3689
rect 76 -3723 88 -3689
rect 30 -3757 88 -3723
rect 30 -3791 42 -3757
rect 76 -3791 88 -3757
rect 30 -3825 88 -3791
rect 30 -3859 42 -3825
rect 76 -3859 88 -3825
rect 30 -3893 88 -3859
rect 30 -3927 42 -3893
rect 76 -3927 88 -3893
rect 30 -3961 88 -3927
rect 30 -3995 42 -3961
rect 76 -3995 88 -3961
rect 30 -4029 88 -3995
rect 30 -4063 42 -4029
rect 76 -4063 88 -4029
rect 30 -4097 88 -4063
rect 30 -4131 42 -4097
rect 76 -4131 88 -4097
rect 30 -4165 88 -4131
rect 30 -4199 42 -4165
rect 76 -4199 88 -4165
rect 30 -4233 88 -4199
rect 30 -4267 42 -4233
rect 76 -4267 88 -4233
rect 30 -4301 88 -4267
rect 30 -4335 42 -4301
rect 76 -4335 88 -4301
rect 30 -4369 88 -4335
rect 30 -4403 42 -4369
rect 76 -4403 88 -4369
rect 30 -4437 88 -4403
rect 30 -4471 42 -4437
rect 76 -4471 88 -4437
rect 30 -4505 88 -4471
rect 30 -4539 42 -4505
rect 76 -4539 88 -4505
rect 30 -4573 88 -4539
rect 30 -4607 42 -4573
rect 76 -4607 88 -4573
rect 30 -4641 88 -4607
rect 30 -4675 42 -4641
rect 76 -4675 88 -4641
rect 30 -4709 88 -4675
rect 30 -4743 42 -4709
rect 76 -4743 88 -4709
rect 30 -4777 88 -4743
rect 30 -4811 42 -4777
rect 76 -4811 88 -4777
rect 30 -4845 88 -4811
rect 30 -4879 42 -4845
rect 76 -4879 88 -4845
rect 30 -4913 88 -4879
rect 30 -4947 42 -4913
rect 76 -4947 88 -4913
rect 30 -4981 88 -4947
rect 30 -5015 42 -4981
rect 76 -5015 88 -4981
rect 30 -5049 88 -5015
rect 30 -5083 42 -5049
rect 76 -5083 88 -5049
rect 30 -5117 88 -5083
rect 30 -5151 42 -5117
rect 76 -5151 88 -5117
rect 30 -5185 88 -5151
rect 30 -5219 42 -5185
rect 76 -5219 88 -5185
rect 30 -5253 88 -5219
rect 30 -5287 42 -5253
rect 76 -5287 88 -5253
rect 30 -5321 88 -5287
rect 30 -5355 42 -5321
rect 76 -5355 88 -5321
rect 30 -5389 88 -5355
rect 30 -5423 42 -5389
rect 76 -5423 88 -5389
rect 30 -5457 88 -5423
rect 30 -5491 42 -5457
rect 76 -5491 88 -5457
rect 30 -5525 88 -5491
rect 30 -5559 42 -5525
rect 76 -5559 88 -5525
rect 30 -5593 88 -5559
rect 30 -5627 42 -5593
rect 76 -5627 88 -5593
rect 30 -5661 88 -5627
rect 30 -5695 42 -5661
rect 76 -5695 88 -5661
rect 30 -5729 88 -5695
rect 30 -5763 42 -5729
rect 76 -5763 88 -5729
rect 30 -5797 88 -5763
rect 30 -5831 42 -5797
rect 76 -5831 88 -5797
rect 30 -5865 88 -5831
rect 30 -5899 42 -5865
rect 76 -5899 88 -5865
rect 30 -5933 88 -5899
rect 30 -5967 42 -5933
rect 76 -5967 88 -5933
rect 30 -6001 88 -5967
rect 30 -6035 42 -6001
rect 76 -6035 88 -6001
rect 30 -6069 88 -6035
rect 30 -6103 42 -6069
rect 76 -6103 88 -6069
rect 30 -6137 88 -6103
rect 30 -6171 42 -6137
rect 76 -6171 88 -6137
rect 30 -6205 88 -6171
rect 30 -6239 42 -6205
rect 76 -6239 88 -6205
rect 30 -6273 88 -6239
rect 30 -6307 42 -6273
rect 76 -6307 88 -6273
rect 30 -6341 88 -6307
rect 30 -6375 42 -6341
rect 76 -6375 88 -6341
rect 30 -6409 88 -6375
rect 30 -6443 42 -6409
rect 76 -6443 88 -6409
rect 30 -6477 88 -6443
rect 30 -6511 42 -6477
rect 76 -6511 88 -6477
rect 30 -6545 88 -6511
rect 30 -6579 42 -6545
rect 76 -6579 88 -6545
rect 30 -6613 88 -6579
rect 30 -6647 42 -6613
rect 76 -6647 88 -6613
rect 30 -6681 88 -6647
rect 30 -6715 42 -6681
rect 76 -6715 88 -6681
rect 30 -6749 88 -6715
rect 30 -6783 42 -6749
rect 76 -6783 88 -6749
rect 30 -6817 88 -6783
rect 30 -6851 42 -6817
rect 76 -6851 88 -6817
rect 30 -6885 88 -6851
rect 30 -6919 42 -6885
rect 76 -6919 88 -6885
rect 30 -6953 88 -6919
rect 30 -6987 42 -6953
rect 76 -6987 88 -6953
rect 30 -7021 88 -6987
rect 30 -7055 42 -7021
rect 76 -7055 88 -7021
rect 30 -7089 88 -7055
rect 30 -7123 42 -7089
rect 76 -7123 88 -7089
rect 30 -7157 88 -7123
rect 30 -7191 42 -7157
rect 76 -7191 88 -7157
rect 30 -7225 88 -7191
rect 30 -7259 42 -7225
rect 76 -7259 88 -7225
rect 30 -7293 88 -7259
rect 30 -7327 42 -7293
rect 76 -7327 88 -7293
rect 30 -7361 88 -7327
rect 30 -7395 42 -7361
rect 76 -7395 88 -7361
rect 30 -7429 88 -7395
rect 30 -7463 42 -7429
rect 76 -7463 88 -7429
rect 30 -7497 88 -7463
rect 30 -7531 42 -7497
rect 76 -7531 88 -7497
rect 30 -7565 88 -7531
rect 30 -7599 42 -7565
rect 76 -7599 88 -7565
rect 30 -7633 88 -7599
rect 30 -7667 42 -7633
rect 76 -7667 88 -7633
rect 30 -7701 88 -7667
rect 30 -7735 42 -7701
rect 76 -7735 88 -7701
rect 30 -7769 88 -7735
rect 30 -7803 42 -7769
rect 76 -7803 88 -7769
rect 30 -7837 88 -7803
rect 30 -7871 42 -7837
rect 76 -7871 88 -7837
rect 30 -7905 88 -7871
rect 30 -7939 42 -7905
rect 76 -7939 88 -7905
rect 30 -7973 88 -7939
rect 30 -8007 42 -7973
rect 76 -8007 88 -7973
rect 30 -8041 88 -8007
rect 30 -8075 42 -8041
rect 76 -8075 88 -8041
rect 30 -8109 88 -8075
rect 30 -8143 42 -8109
rect 76 -8143 88 -8109
rect 30 -8177 88 -8143
rect 30 -8211 42 -8177
rect 76 -8211 88 -8177
rect 30 -8245 88 -8211
rect 30 -8279 42 -8245
rect 76 -8279 88 -8245
rect 30 -8313 88 -8279
rect 30 -8347 42 -8313
rect 76 -8347 88 -8313
rect 30 -8381 88 -8347
rect 30 -8415 42 -8381
rect 76 -8415 88 -8381
rect 30 -8449 88 -8415
rect 30 -8483 42 -8449
rect 76 -8483 88 -8449
rect 30 -8517 88 -8483
rect 30 -8551 42 -8517
rect 76 -8551 88 -8517
rect 30 -8585 88 -8551
rect 30 -8619 42 -8585
rect 76 -8619 88 -8585
rect 30 -8653 88 -8619
rect 30 -8687 42 -8653
rect 76 -8687 88 -8653
rect 30 -8721 88 -8687
rect 30 -8755 42 -8721
rect 76 -8755 88 -8721
rect 30 -8789 88 -8755
rect 30 -8823 42 -8789
rect 76 -8823 88 -8789
rect 30 -8857 88 -8823
rect 30 -8891 42 -8857
rect 76 -8891 88 -8857
rect 30 -8925 88 -8891
rect 30 -8959 42 -8925
rect 76 -8959 88 -8925
rect 30 -8993 88 -8959
rect 30 -9027 42 -8993
rect 76 -9027 88 -8993
rect 30 -9061 88 -9027
rect 30 -9095 42 -9061
rect 76 -9095 88 -9061
rect 30 -9129 88 -9095
rect 30 -9163 42 -9129
rect 76 -9163 88 -9129
rect 30 -9197 88 -9163
rect 30 -9231 42 -9197
rect 76 -9231 88 -9197
rect 30 -9265 88 -9231
rect 30 -9299 42 -9265
rect 76 -9299 88 -9265
rect 30 -9333 88 -9299
rect 30 -9367 42 -9333
rect 76 -9367 88 -9333
rect 30 -9401 88 -9367
rect 30 -9435 42 -9401
rect 76 -9435 88 -9401
rect 30 -9469 88 -9435
rect 30 -9503 42 -9469
rect 76 -9503 88 -9469
rect 30 -9537 88 -9503
rect 30 -9571 42 -9537
rect 76 -9571 88 -9537
rect 30 -9600 88 -9571
rect 148 9571 206 9600
rect 148 9537 160 9571
rect 194 9537 206 9571
rect 148 9503 206 9537
rect 148 9469 160 9503
rect 194 9469 206 9503
rect 148 9435 206 9469
rect 148 9401 160 9435
rect 194 9401 206 9435
rect 148 9367 206 9401
rect 148 9333 160 9367
rect 194 9333 206 9367
rect 148 9299 206 9333
rect 148 9265 160 9299
rect 194 9265 206 9299
rect 148 9231 206 9265
rect 148 9197 160 9231
rect 194 9197 206 9231
rect 148 9163 206 9197
rect 148 9129 160 9163
rect 194 9129 206 9163
rect 148 9095 206 9129
rect 148 9061 160 9095
rect 194 9061 206 9095
rect 148 9027 206 9061
rect 148 8993 160 9027
rect 194 8993 206 9027
rect 148 8959 206 8993
rect 148 8925 160 8959
rect 194 8925 206 8959
rect 148 8891 206 8925
rect 148 8857 160 8891
rect 194 8857 206 8891
rect 148 8823 206 8857
rect 148 8789 160 8823
rect 194 8789 206 8823
rect 148 8755 206 8789
rect 148 8721 160 8755
rect 194 8721 206 8755
rect 148 8687 206 8721
rect 148 8653 160 8687
rect 194 8653 206 8687
rect 148 8619 206 8653
rect 148 8585 160 8619
rect 194 8585 206 8619
rect 148 8551 206 8585
rect 148 8517 160 8551
rect 194 8517 206 8551
rect 148 8483 206 8517
rect 148 8449 160 8483
rect 194 8449 206 8483
rect 148 8415 206 8449
rect 148 8381 160 8415
rect 194 8381 206 8415
rect 148 8347 206 8381
rect 148 8313 160 8347
rect 194 8313 206 8347
rect 148 8279 206 8313
rect 148 8245 160 8279
rect 194 8245 206 8279
rect 148 8211 206 8245
rect 148 8177 160 8211
rect 194 8177 206 8211
rect 148 8143 206 8177
rect 148 8109 160 8143
rect 194 8109 206 8143
rect 148 8075 206 8109
rect 148 8041 160 8075
rect 194 8041 206 8075
rect 148 8007 206 8041
rect 148 7973 160 8007
rect 194 7973 206 8007
rect 148 7939 206 7973
rect 148 7905 160 7939
rect 194 7905 206 7939
rect 148 7871 206 7905
rect 148 7837 160 7871
rect 194 7837 206 7871
rect 148 7803 206 7837
rect 148 7769 160 7803
rect 194 7769 206 7803
rect 148 7735 206 7769
rect 148 7701 160 7735
rect 194 7701 206 7735
rect 148 7667 206 7701
rect 148 7633 160 7667
rect 194 7633 206 7667
rect 148 7599 206 7633
rect 148 7565 160 7599
rect 194 7565 206 7599
rect 148 7531 206 7565
rect 148 7497 160 7531
rect 194 7497 206 7531
rect 148 7463 206 7497
rect 148 7429 160 7463
rect 194 7429 206 7463
rect 148 7395 206 7429
rect 148 7361 160 7395
rect 194 7361 206 7395
rect 148 7327 206 7361
rect 148 7293 160 7327
rect 194 7293 206 7327
rect 148 7259 206 7293
rect 148 7225 160 7259
rect 194 7225 206 7259
rect 148 7191 206 7225
rect 148 7157 160 7191
rect 194 7157 206 7191
rect 148 7123 206 7157
rect 148 7089 160 7123
rect 194 7089 206 7123
rect 148 7055 206 7089
rect 148 7021 160 7055
rect 194 7021 206 7055
rect 148 6987 206 7021
rect 148 6953 160 6987
rect 194 6953 206 6987
rect 148 6919 206 6953
rect 148 6885 160 6919
rect 194 6885 206 6919
rect 148 6851 206 6885
rect 148 6817 160 6851
rect 194 6817 206 6851
rect 148 6783 206 6817
rect 148 6749 160 6783
rect 194 6749 206 6783
rect 148 6715 206 6749
rect 148 6681 160 6715
rect 194 6681 206 6715
rect 148 6647 206 6681
rect 148 6613 160 6647
rect 194 6613 206 6647
rect 148 6579 206 6613
rect 148 6545 160 6579
rect 194 6545 206 6579
rect 148 6511 206 6545
rect 148 6477 160 6511
rect 194 6477 206 6511
rect 148 6443 206 6477
rect 148 6409 160 6443
rect 194 6409 206 6443
rect 148 6375 206 6409
rect 148 6341 160 6375
rect 194 6341 206 6375
rect 148 6307 206 6341
rect 148 6273 160 6307
rect 194 6273 206 6307
rect 148 6239 206 6273
rect 148 6205 160 6239
rect 194 6205 206 6239
rect 148 6171 206 6205
rect 148 6137 160 6171
rect 194 6137 206 6171
rect 148 6103 206 6137
rect 148 6069 160 6103
rect 194 6069 206 6103
rect 148 6035 206 6069
rect 148 6001 160 6035
rect 194 6001 206 6035
rect 148 5967 206 6001
rect 148 5933 160 5967
rect 194 5933 206 5967
rect 148 5899 206 5933
rect 148 5865 160 5899
rect 194 5865 206 5899
rect 148 5831 206 5865
rect 148 5797 160 5831
rect 194 5797 206 5831
rect 148 5763 206 5797
rect 148 5729 160 5763
rect 194 5729 206 5763
rect 148 5695 206 5729
rect 148 5661 160 5695
rect 194 5661 206 5695
rect 148 5627 206 5661
rect 148 5593 160 5627
rect 194 5593 206 5627
rect 148 5559 206 5593
rect 148 5525 160 5559
rect 194 5525 206 5559
rect 148 5491 206 5525
rect 148 5457 160 5491
rect 194 5457 206 5491
rect 148 5423 206 5457
rect 148 5389 160 5423
rect 194 5389 206 5423
rect 148 5355 206 5389
rect 148 5321 160 5355
rect 194 5321 206 5355
rect 148 5287 206 5321
rect 148 5253 160 5287
rect 194 5253 206 5287
rect 148 5219 206 5253
rect 148 5185 160 5219
rect 194 5185 206 5219
rect 148 5151 206 5185
rect 148 5117 160 5151
rect 194 5117 206 5151
rect 148 5083 206 5117
rect 148 5049 160 5083
rect 194 5049 206 5083
rect 148 5015 206 5049
rect 148 4981 160 5015
rect 194 4981 206 5015
rect 148 4947 206 4981
rect 148 4913 160 4947
rect 194 4913 206 4947
rect 148 4879 206 4913
rect 148 4845 160 4879
rect 194 4845 206 4879
rect 148 4811 206 4845
rect 148 4777 160 4811
rect 194 4777 206 4811
rect 148 4743 206 4777
rect 148 4709 160 4743
rect 194 4709 206 4743
rect 148 4675 206 4709
rect 148 4641 160 4675
rect 194 4641 206 4675
rect 148 4607 206 4641
rect 148 4573 160 4607
rect 194 4573 206 4607
rect 148 4539 206 4573
rect 148 4505 160 4539
rect 194 4505 206 4539
rect 148 4471 206 4505
rect 148 4437 160 4471
rect 194 4437 206 4471
rect 148 4403 206 4437
rect 148 4369 160 4403
rect 194 4369 206 4403
rect 148 4335 206 4369
rect 148 4301 160 4335
rect 194 4301 206 4335
rect 148 4267 206 4301
rect 148 4233 160 4267
rect 194 4233 206 4267
rect 148 4199 206 4233
rect 148 4165 160 4199
rect 194 4165 206 4199
rect 148 4131 206 4165
rect 148 4097 160 4131
rect 194 4097 206 4131
rect 148 4063 206 4097
rect 148 4029 160 4063
rect 194 4029 206 4063
rect 148 3995 206 4029
rect 148 3961 160 3995
rect 194 3961 206 3995
rect 148 3927 206 3961
rect 148 3893 160 3927
rect 194 3893 206 3927
rect 148 3859 206 3893
rect 148 3825 160 3859
rect 194 3825 206 3859
rect 148 3791 206 3825
rect 148 3757 160 3791
rect 194 3757 206 3791
rect 148 3723 206 3757
rect 148 3689 160 3723
rect 194 3689 206 3723
rect 148 3655 206 3689
rect 148 3621 160 3655
rect 194 3621 206 3655
rect 148 3587 206 3621
rect 148 3553 160 3587
rect 194 3553 206 3587
rect 148 3519 206 3553
rect 148 3485 160 3519
rect 194 3485 206 3519
rect 148 3451 206 3485
rect 148 3417 160 3451
rect 194 3417 206 3451
rect 148 3383 206 3417
rect 148 3349 160 3383
rect 194 3349 206 3383
rect 148 3315 206 3349
rect 148 3281 160 3315
rect 194 3281 206 3315
rect 148 3247 206 3281
rect 148 3213 160 3247
rect 194 3213 206 3247
rect 148 3179 206 3213
rect 148 3145 160 3179
rect 194 3145 206 3179
rect 148 3111 206 3145
rect 148 3077 160 3111
rect 194 3077 206 3111
rect 148 3043 206 3077
rect 148 3009 160 3043
rect 194 3009 206 3043
rect 148 2975 206 3009
rect 148 2941 160 2975
rect 194 2941 206 2975
rect 148 2907 206 2941
rect 148 2873 160 2907
rect 194 2873 206 2907
rect 148 2839 206 2873
rect 148 2805 160 2839
rect 194 2805 206 2839
rect 148 2771 206 2805
rect 148 2737 160 2771
rect 194 2737 206 2771
rect 148 2703 206 2737
rect 148 2669 160 2703
rect 194 2669 206 2703
rect 148 2635 206 2669
rect 148 2601 160 2635
rect 194 2601 206 2635
rect 148 2567 206 2601
rect 148 2533 160 2567
rect 194 2533 206 2567
rect 148 2499 206 2533
rect 148 2465 160 2499
rect 194 2465 206 2499
rect 148 2431 206 2465
rect 148 2397 160 2431
rect 194 2397 206 2431
rect 148 2363 206 2397
rect 148 2329 160 2363
rect 194 2329 206 2363
rect 148 2295 206 2329
rect 148 2261 160 2295
rect 194 2261 206 2295
rect 148 2227 206 2261
rect 148 2193 160 2227
rect 194 2193 206 2227
rect 148 2159 206 2193
rect 148 2125 160 2159
rect 194 2125 206 2159
rect 148 2091 206 2125
rect 148 2057 160 2091
rect 194 2057 206 2091
rect 148 2023 206 2057
rect 148 1989 160 2023
rect 194 1989 206 2023
rect 148 1955 206 1989
rect 148 1921 160 1955
rect 194 1921 206 1955
rect 148 1887 206 1921
rect 148 1853 160 1887
rect 194 1853 206 1887
rect 148 1819 206 1853
rect 148 1785 160 1819
rect 194 1785 206 1819
rect 148 1751 206 1785
rect 148 1717 160 1751
rect 194 1717 206 1751
rect 148 1683 206 1717
rect 148 1649 160 1683
rect 194 1649 206 1683
rect 148 1615 206 1649
rect 148 1581 160 1615
rect 194 1581 206 1615
rect 148 1547 206 1581
rect 148 1513 160 1547
rect 194 1513 206 1547
rect 148 1479 206 1513
rect 148 1445 160 1479
rect 194 1445 206 1479
rect 148 1411 206 1445
rect 148 1377 160 1411
rect 194 1377 206 1411
rect 148 1343 206 1377
rect 148 1309 160 1343
rect 194 1309 206 1343
rect 148 1275 206 1309
rect 148 1241 160 1275
rect 194 1241 206 1275
rect 148 1207 206 1241
rect 148 1173 160 1207
rect 194 1173 206 1207
rect 148 1139 206 1173
rect 148 1105 160 1139
rect 194 1105 206 1139
rect 148 1071 206 1105
rect 148 1037 160 1071
rect 194 1037 206 1071
rect 148 1003 206 1037
rect 148 969 160 1003
rect 194 969 206 1003
rect 148 935 206 969
rect 148 901 160 935
rect 194 901 206 935
rect 148 867 206 901
rect 148 833 160 867
rect 194 833 206 867
rect 148 799 206 833
rect 148 765 160 799
rect 194 765 206 799
rect 148 731 206 765
rect 148 697 160 731
rect 194 697 206 731
rect 148 663 206 697
rect 148 629 160 663
rect 194 629 206 663
rect 148 595 206 629
rect 148 561 160 595
rect 194 561 206 595
rect 148 527 206 561
rect 148 493 160 527
rect 194 493 206 527
rect 148 459 206 493
rect 148 425 160 459
rect 194 425 206 459
rect 148 391 206 425
rect 148 357 160 391
rect 194 357 206 391
rect 148 323 206 357
rect 148 289 160 323
rect 194 289 206 323
rect 148 255 206 289
rect 148 221 160 255
rect 194 221 206 255
rect 148 187 206 221
rect 148 153 160 187
rect 194 153 206 187
rect 148 119 206 153
rect 148 85 160 119
rect 194 85 206 119
rect 148 51 206 85
rect 148 17 160 51
rect 194 17 206 51
rect 148 -17 206 17
rect 148 -51 160 -17
rect 194 -51 206 -17
rect 148 -85 206 -51
rect 148 -119 160 -85
rect 194 -119 206 -85
rect 148 -153 206 -119
rect 148 -187 160 -153
rect 194 -187 206 -153
rect 148 -221 206 -187
rect 148 -255 160 -221
rect 194 -255 206 -221
rect 148 -289 206 -255
rect 148 -323 160 -289
rect 194 -323 206 -289
rect 148 -357 206 -323
rect 148 -391 160 -357
rect 194 -391 206 -357
rect 148 -425 206 -391
rect 148 -459 160 -425
rect 194 -459 206 -425
rect 148 -493 206 -459
rect 148 -527 160 -493
rect 194 -527 206 -493
rect 148 -561 206 -527
rect 148 -595 160 -561
rect 194 -595 206 -561
rect 148 -629 206 -595
rect 148 -663 160 -629
rect 194 -663 206 -629
rect 148 -697 206 -663
rect 148 -731 160 -697
rect 194 -731 206 -697
rect 148 -765 206 -731
rect 148 -799 160 -765
rect 194 -799 206 -765
rect 148 -833 206 -799
rect 148 -867 160 -833
rect 194 -867 206 -833
rect 148 -901 206 -867
rect 148 -935 160 -901
rect 194 -935 206 -901
rect 148 -969 206 -935
rect 148 -1003 160 -969
rect 194 -1003 206 -969
rect 148 -1037 206 -1003
rect 148 -1071 160 -1037
rect 194 -1071 206 -1037
rect 148 -1105 206 -1071
rect 148 -1139 160 -1105
rect 194 -1139 206 -1105
rect 148 -1173 206 -1139
rect 148 -1207 160 -1173
rect 194 -1207 206 -1173
rect 148 -1241 206 -1207
rect 148 -1275 160 -1241
rect 194 -1275 206 -1241
rect 148 -1309 206 -1275
rect 148 -1343 160 -1309
rect 194 -1343 206 -1309
rect 148 -1377 206 -1343
rect 148 -1411 160 -1377
rect 194 -1411 206 -1377
rect 148 -1445 206 -1411
rect 148 -1479 160 -1445
rect 194 -1479 206 -1445
rect 148 -1513 206 -1479
rect 148 -1547 160 -1513
rect 194 -1547 206 -1513
rect 148 -1581 206 -1547
rect 148 -1615 160 -1581
rect 194 -1615 206 -1581
rect 148 -1649 206 -1615
rect 148 -1683 160 -1649
rect 194 -1683 206 -1649
rect 148 -1717 206 -1683
rect 148 -1751 160 -1717
rect 194 -1751 206 -1717
rect 148 -1785 206 -1751
rect 148 -1819 160 -1785
rect 194 -1819 206 -1785
rect 148 -1853 206 -1819
rect 148 -1887 160 -1853
rect 194 -1887 206 -1853
rect 148 -1921 206 -1887
rect 148 -1955 160 -1921
rect 194 -1955 206 -1921
rect 148 -1989 206 -1955
rect 148 -2023 160 -1989
rect 194 -2023 206 -1989
rect 148 -2057 206 -2023
rect 148 -2091 160 -2057
rect 194 -2091 206 -2057
rect 148 -2125 206 -2091
rect 148 -2159 160 -2125
rect 194 -2159 206 -2125
rect 148 -2193 206 -2159
rect 148 -2227 160 -2193
rect 194 -2227 206 -2193
rect 148 -2261 206 -2227
rect 148 -2295 160 -2261
rect 194 -2295 206 -2261
rect 148 -2329 206 -2295
rect 148 -2363 160 -2329
rect 194 -2363 206 -2329
rect 148 -2397 206 -2363
rect 148 -2431 160 -2397
rect 194 -2431 206 -2397
rect 148 -2465 206 -2431
rect 148 -2499 160 -2465
rect 194 -2499 206 -2465
rect 148 -2533 206 -2499
rect 148 -2567 160 -2533
rect 194 -2567 206 -2533
rect 148 -2601 206 -2567
rect 148 -2635 160 -2601
rect 194 -2635 206 -2601
rect 148 -2669 206 -2635
rect 148 -2703 160 -2669
rect 194 -2703 206 -2669
rect 148 -2737 206 -2703
rect 148 -2771 160 -2737
rect 194 -2771 206 -2737
rect 148 -2805 206 -2771
rect 148 -2839 160 -2805
rect 194 -2839 206 -2805
rect 148 -2873 206 -2839
rect 148 -2907 160 -2873
rect 194 -2907 206 -2873
rect 148 -2941 206 -2907
rect 148 -2975 160 -2941
rect 194 -2975 206 -2941
rect 148 -3009 206 -2975
rect 148 -3043 160 -3009
rect 194 -3043 206 -3009
rect 148 -3077 206 -3043
rect 148 -3111 160 -3077
rect 194 -3111 206 -3077
rect 148 -3145 206 -3111
rect 148 -3179 160 -3145
rect 194 -3179 206 -3145
rect 148 -3213 206 -3179
rect 148 -3247 160 -3213
rect 194 -3247 206 -3213
rect 148 -3281 206 -3247
rect 148 -3315 160 -3281
rect 194 -3315 206 -3281
rect 148 -3349 206 -3315
rect 148 -3383 160 -3349
rect 194 -3383 206 -3349
rect 148 -3417 206 -3383
rect 148 -3451 160 -3417
rect 194 -3451 206 -3417
rect 148 -3485 206 -3451
rect 148 -3519 160 -3485
rect 194 -3519 206 -3485
rect 148 -3553 206 -3519
rect 148 -3587 160 -3553
rect 194 -3587 206 -3553
rect 148 -3621 206 -3587
rect 148 -3655 160 -3621
rect 194 -3655 206 -3621
rect 148 -3689 206 -3655
rect 148 -3723 160 -3689
rect 194 -3723 206 -3689
rect 148 -3757 206 -3723
rect 148 -3791 160 -3757
rect 194 -3791 206 -3757
rect 148 -3825 206 -3791
rect 148 -3859 160 -3825
rect 194 -3859 206 -3825
rect 148 -3893 206 -3859
rect 148 -3927 160 -3893
rect 194 -3927 206 -3893
rect 148 -3961 206 -3927
rect 148 -3995 160 -3961
rect 194 -3995 206 -3961
rect 148 -4029 206 -3995
rect 148 -4063 160 -4029
rect 194 -4063 206 -4029
rect 148 -4097 206 -4063
rect 148 -4131 160 -4097
rect 194 -4131 206 -4097
rect 148 -4165 206 -4131
rect 148 -4199 160 -4165
rect 194 -4199 206 -4165
rect 148 -4233 206 -4199
rect 148 -4267 160 -4233
rect 194 -4267 206 -4233
rect 148 -4301 206 -4267
rect 148 -4335 160 -4301
rect 194 -4335 206 -4301
rect 148 -4369 206 -4335
rect 148 -4403 160 -4369
rect 194 -4403 206 -4369
rect 148 -4437 206 -4403
rect 148 -4471 160 -4437
rect 194 -4471 206 -4437
rect 148 -4505 206 -4471
rect 148 -4539 160 -4505
rect 194 -4539 206 -4505
rect 148 -4573 206 -4539
rect 148 -4607 160 -4573
rect 194 -4607 206 -4573
rect 148 -4641 206 -4607
rect 148 -4675 160 -4641
rect 194 -4675 206 -4641
rect 148 -4709 206 -4675
rect 148 -4743 160 -4709
rect 194 -4743 206 -4709
rect 148 -4777 206 -4743
rect 148 -4811 160 -4777
rect 194 -4811 206 -4777
rect 148 -4845 206 -4811
rect 148 -4879 160 -4845
rect 194 -4879 206 -4845
rect 148 -4913 206 -4879
rect 148 -4947 160 -4913
rect 194 -4947 206 -4913
rect 148 -4981 206 -4947
rect 148 -5015 160 -4981
rect 194 -5015 206 -4981
rect 148 -5049 206 -5015
rect 148 -5083 160 -5049
rect 194 -5083 206 -5049
rect 148 -5117 206 -5083
rect 148 -5151 160 -5117
rect 194 -5151 206 -5117
rect 148 -5185 206 -5151
rect 148 -5219 160 -5185
rect 194 -5219 206 -5185
rect 148 -5253 206 -5219
rect 148 -5287 160 -5253
rect 194 -5287 206 -5253
rect 148 -5321 206 -5287
rect 148 -5355 160 -5321
rect 194 -5355 206 -5321
rect 148 -5389 206 -5355
rect 148 -5423 160 -5389
rect 194 -5423 206 -5389
rect 148 -5457 206 -5423
rect 148 -5491 160 -5457
rect 194 -5491 206 -5457
rect 148 -5525 206 -5491
rect 148 -5559 160 -5525
rect 194 -5559 206 -5525
rect 148 -5593 206 -5559
rect 148 -5627 160 -5593
rect 194 -5627 206 -5593
rect 148 -5661 206 -5627
rect 148 -5695 160 -5661
rect 194 -5695 206 -5661
rect 148 -5729 206 -5695
rect 148 -5763 160 -5729
rect 194 -5763 206 -5729
rect 148 -5797 206 -5763
rect 148 -5831 160 -5797
rect 194 -5831 206 -5797
rect 148 -5865 206 -5831
rect 148 -5899 160 -5865
rect 194 -5899 206 -5865
rect 148 -5933 206 -5899
rect 148 -5967 160 -5933
rect 194 -5967 206 -5933
rect 148 -6001 206 -5967
rect 148 -6035 160 -6001
rect 194 -6035 206 -6001
rect 148 -6069 206 -6035
rect 148 -6103 160 -6069
rect 194 -6103 206 -6069
rect 148 -6137 206 -6103
rect 148 -6171 160 -6137
rect 194 -6171 206 -6137
rect 148 -6205 206 -6171
rect 148 -6239 160 -6205
rect 194 -6239 206 -6205
rect 148 -6273 206 -6239
rect 148 -6307 160 -6273
rect 194 -6307 206 -6273
rect 148 -6341 206 -6307
rect 148 -6375 160 -6341
rect 194 -6375 206 -6341
rect 148 -6409 206 -6375
rect 148 -6443 160 -6409
rect 194 -6443 206 -6409
rect 148 -6477 206 -6443
rect 148 -6511 160 -6477
rect 194 -6511 206 -6477
rect 148 -6545 206 -6511
rect 148 -6579 160 -6545
rect 194 -6579 206 -6545
rect 148 -6613 206 -6579
rect 148 -6647 160 -6613
rect 194 -6647 206 -6613
rect 148 -6681 206 -6647
rect 148 -6715 160 -6681
rect 194 -6715 206 -6681
rect 148 -6749 206 -6715
rect 148 -6783 160 -6749
rect 194 -6783 206 -6749
rect 148 -6817 206 -6783
rect 148 -6851 160 -6817
rect 194 -6851 206 -6817
rect 148 -6885 206 -6851
rect 148 -6919 160 -6885
rect 194 -6919 206 -6885
rect 148 -6953 206 -6919
rect 148 -6987 160 -6953
rect 194 -6987 206 -6953
rect 148 -7021 206 -6987
rect 148 -7055 160 -7021
rect 194 -7055 206 -7021
rect 148 -7089 206 -7055
rect 148 -7123 160 -7089
rect 194 -7123 206 -7089
rect 148 -7157 206 -7123
rect 148 -7191 160 -7157
rect 194 -7191 206 -7157
rect 148 -7225 206 -7191
rect 148 -7259 160 -7225
rect 194 -7259 206 -7225
rect 148 -7293 206 -7259
rect 148 -7327 160 -7293
rect 194 -7327 206 -7293
rect 148 -7361 206 -7327
rect 148 -7395 160 -7361
rect 194 -7395 206 -7361
rect 148 -7429 206 -7395
rect 148 -7463 160 -7429
rect 194 -7463 206 -7429
rect 148 -7497 206 -7463
rect 148 -7531 160 -7497
rect 194 -7531 206 -7497
rect 148 -7565 206 -7531
rect 148 -7599 160 -7565
rect 194 -7599 206 -7565
rect 148 -7633 206 -7599
rect 148 -7667 160 -7633
rect 194 -7667 206 -7633
rect 148 -7701 206 -7667
rect 148 -7735 160 -7701
rect 194 -7735 206 -7701
rect 148 -7769 206 -7735
rect 148 -7803 160 -7769
rect 194 -7803 206 -7769
rect 148 -7837 206 -7803
rect 148 -7871 160 -7837
rect 194 -7871 206 -7837
rect 148 -7905 206 -7871
rect 148 -7939 160 -7905
rect 194 -7939 206 -7905
rect 148 -7973 206 -7939
rect 148 -8007 160 -7973
rect 194 -8007 206 -7973
rect 148 -8041 206 -8007
rect 148 -8075 160 -8041
rect 194 -8075 206 -8041
rect 148 -8109 206 -8075
rect 148 -8143 160 -8109
rect 194 -8143 206 -8109
rect 148 -8177 206 -8143
rect 148 -8211 160 -8177
rect 194 -8211 206 -8177
rect 148 -8245 206 -8211
rect 148 -8279 160 -8245
rect 194 -8279 206 -8245
rect 148 -8313 206 -8279
rect 148 -8347 160 -8313
rect 194 -8347 206 -8313
rect 148 -8381 206 -8347
rect 148 -8415 160 -8381
rect 194 -8415 206 -8381
rect 148 -8449 206 -8415
rect 148 -8483 160 -8449
rect 194 -8483 206 -8449
rect 148 -8517 206 -8483
rect 148 -8551 160 -8517
rect 194 -8551 206 -8517
rect 148 -8585 206 -8551
rect 148 -8619 160 -8585
rect 194 -8619 206 -8585
rect 148 -8653 206 -8619
rect 148 -8687 160 -8653
rect 194 -8687 206 -8653
rect 148 -8721 206 -8687
rect 148 -8755 160 -8721
rect 194 -8755 206 -8721
rect 148 -8789 206 -8755
rect 148 -8823 160 -8789
rect 194 -8823 206 -8789
rect 148 -8857 206 -8823
rect 148 -8891 160 -8857
rect 194 -8891 206 -8857
rect 148 -8925 206 -8891
rect 148 -8959 160 -8925
rect 194 -8959 206 -8925
rect 148 -8993 206 -8959
rect 148 -9027 160 -8993
rect 194 -9027 206 -8993
rect 148 -9061 206 -9027
rect 148 -9095 160 -9061
rect 194 -9095 206 -9061
rect 148 -9129 206 -9095
rect 148 -9163 160 -9129
rect 194 -9163 206 -9129
rect 148 -9197 206 -9163
rect 148 -9231 160 -9197
rect 194 -9231 206 -9197
rect 148 -9265 206 -9231
rect 148 -9299 160 -9265
rect 194 -9299 206 -9265
rect 148 -9333 206 -9299
rect 148 -9367 160 -9333
rect 194 -9367 206 -9333
rect 148 -9401 206 -9367
rect 148 -9435 160 -9401
rect 194 -9435 206 -9401
rect 148 -9469 206 -9435
rect 148 -9503 160 -9469
rect 194 -9503 206 -9469
rect 148 -9537 206 -9503
rect 148 -9571 160 -9537
rect 194 -9571 206 -9537
rect 148 -9600 206 -9571
rect 266 9571 324 9600
rect 266 9537 278 9571
rect 312 9537 324 9571
rect 266 9503 324 9537
rect 266 9469 278 9503
rect 312 9469 324 9503
rect 266 9435 324 9469
rect 266 9401 278 9435
rect 312 9401 324 9435
rect 266 9367 324 9401
rect 266 9333 278 9367
rect 312 9333 324 9367
rect 266 9299 324 9333
rect 266 9265 278 9299
rect 312 9265 324 9299
rect 266 9231 324 9265
rect 266 9197 278 9231
rect 312 9197 324 9231
rect 266 9163 324 9197
rect 266 9129 278 9163
rect 312 9129 324 9163
rect 266 9095 324 9129
rect 266 9061 278 9095
rect 312 9061 324 9095
rect 266 9027 324 9061
rect 266 8993 278 9027
rect 312 8993 324 9027
rect 266 8959 324 8993
rect 266 8925 278 8959
rect 312 8925 324 8959
rect 266 8891 324 8925
rect 266 8857 278 8891
rect 312 8857 324 8891
rect 266 8823 324 8857
rect 266 8789 278 8823
rect 312 8789 324 8823
rect 266 8755 324 8789
rect 266 8721 278 8755
rect 312 8721 324 8755
rect 266 8687 324 8721
rect 266 8653 278 8687
rect 312 8653 324 8687
rect 266 8619 324 8653
rect 266 8585 278 8619
rect 312 8585 324 8619
rect 266 8551 324 8585
rect 266 8517 278 8551
rect 312 8517 324 8551
rect 266 8483 324 8517
rect 266 8449 278 8483
rect 312 8449 324 8483
rect 266 8415 324 8449
rect 266 8381 278 8415
rect 312 8381 324 8415
rect 266 8347 324 8381
rect 266 8313 278 8347
rect 312 8313 324 8347
rect 266 8279 324 8313
rect 266 8245 278 8279
rect 312 8245 324 8279
rect 266 8211 324 8245
rect 266 8177 278 8211
rect 312 8177 324 8211
rect 266 8143 324 8177
rect 266 8109 278 8143
rect 312 8109 324 8143
rect 266 8075 324 8109
rect 266 8041 278 8075
rect 312 8041 324 8075
rect 266 8007 324 8041
rect 266 7973 278 8007
rect 312 7973 324 8007
rect 266 7939 324 7973
rect 266 7905 278 7939
rect 312 7905 324 7939
rect 266 7871 324 7905
rect 266 7837 278 7871
rect 312 7837 324 7871
rect 266 7803 324 7837
rect 266 7769 278 7803
rect 312 7769 324 7803
rect 266 7735 324 7769
rect 266 7701 278 7735
rect 312 7701 324 7735
rect 266 7667 324 7701
rect 266 7633 278 7667
rect 312 7633 324 7667
rect 266 7599 324 7633
rect 266 7565 278 7599
rect 312 7565 324 7599
rect 266 7531 324 7565
rect 266 7497 278 7531
rect 312 7497 324 7531
rect 266 7463 324 7497
rect 266 7429 278 7463
rect 312 7429 324 7463
rect 266 7395 324 7429
rect 266 7361 278 7395
rect 312 7361 324 7395
rect 266 7327 324 7361
rect 266 7293 278 7327
rect 312 7293 324 7327
rect 266 7259 324 7293
rect 266 7225 278 7259
rect 312 7225 324 7259
rect 266 7191 324 7225
rect 266 7157 278 7191
rect 312 7157 324 7191
rect 266 7123 324 7157
rect 266 7089 278 7123
rect 312 7089 324 7123
rect 266 7055 324 7089
rect 266 7021 278 7055
rect 312 7021 324 7055
rect 266 6987 324 7021
rect 266 6953 278 6987
rect 312 6953 324 6987
rect 266 6919 324 6953
rect 266 6885 278 6919
rect 312 6885 324 6919
rect 266 6851 324 6885
rect 266 6817 278 6851
rect 312 6817 324 6851
rect 266 6783 324 6817
rect 266 6749 278 6783
rect 312 6749 324 6783
rect 266 6715 324 6749
rect 266 6681 278 6715
rect 312 6681 324 6715
rect 266 6647 324 6681
rect 266 6613 278 6647
rect 312 6613 324 6647
rect 266 6579 324 6613
rect 266 6545 278 6579
rect 312 6545 324 6579
rect 266 6511 324 6545
rect 266 6477 278 6511
rect 312 6477 324 6511
rect 266 6443 324 6477
rect 266 6409 278 6443
rect 312 6409 324 6443
rect 266 6375 324 6409
rect 266 6341 278 6375
rect 312 6341 324 6375
rect 266 6307 324 6341
rect 266 6273 278 6307
rect 312 6273 324 6307
rect 266 6239 324 6273
rect 266 6205 278 6239
rect 312 6205 324 6239
rect 266 6171 324 6205
rect 266 6137 278 6171
rect 312 6137 324 6171
rect 266 6103 324 6137
rect 266 6069 278 6103
rect 312 6069 324 6103
rect 266 6035 324 6069
rect 266 6001 278 6035
rect 312 6001 324 6035
rect 266 5967 324 6001
rect 266 5933 278 5967
rect 312 5933 324 5967
rect 266 5899 324 5933
rect 266 5865 278 5899
rect 312 5865 324 5899
rect 266 5831 324 5865
rect 266 5797 278 5831
rect 312 5797 324 5831
rect 266 5763 324 5797
rect 266 5729 278 5763
rect 312 5729 324 5763
rect 266 5695 324 5729
rect 266 5661 278 5695
rect 312 5661 324 5695
rect 266 5627 324 5661
rect 266 5593 278 5627
rect 312 5593 324 5627
rect 266 5559 324 5593
rect 266 5525 278 5559
rect 312 5525 324 5559
rect 266 5491 324 5525
rect 266 5457 278 5491
rect 312 5457 324 5491
rect 266 5423 324 5457
rect 266 5389 278 5423
rect 312 5389 324 5423
rect 266 5355 324 5389
rect 266 5321 278 5355
rect 312 5321 324 5355
rect 266 5287 324 5321
rect 266 5253 278 5287
rect 312 5253 324 5287
rect 266 5219 324 5253
rect 266 5185 278 5219
rect 312 5185 324 5219
rect 266 5151 324 5185
rect 266 5117 278 5151
rect 312 5117 324 5151
rect 266 5083 324 5117
rect 266 5049 278 5083
rect 312 5049 324 5083
rect 266 5015 324 5049
rect 266 4981 278 5015
rect 312 4981 324 5015
rect 266 4947 324 4981
rect 266 4913 278 4947
rect 312 4913 324 4947
rect 266 4879 324 4913
rect 266 4845 278 4879
rect 312 4845 324 4879
rect 266 4811 324 4845
rect 266 4777 278 4811
rect 312 4777 324 4811
rect 266 4743 324 4777
rect 266 4709 278 4743
rect 312 4709 324 4743
rect 266 4675 324 4709
rect 266 4641 278 4675
rect 312 4641 324 4675
rect 266 4607 324 4641
rect 266 4573 278 4607
rect 312 4573 324 4607
rect 266 4539 324 4573
rect 266 4505 278 4539
rect 312 4505 324 4539
rect 266 4471 324 4505
rect 266 4437 278 4471
rect 312 4437 324 4471
rect 266 4403 324 4437
rect 266 4369 278 4403
rect 312 4369 324 4403
rect 266 4335 324 4369
rect 266 4301 278 4335
rect 312 4301 324 4335
rect 266 4267 324 4301
rect 266 4233 278 4267
rect 312 4233 324 4267
rect 266 4199 324 4233
rect 266 4165 278 4199
rect 312 4165 324 4199
rect 266 4131 324 4165
rect 266 4097 278 4131
rect 312 4097 324 4131
rect 266 4063 324 4097
rect 266 4029 278 4063
rect 312 4029 324 4063
rect 266 3995 324 4029
rect 266 3961 278 3995
rect 312 3961 324 3995
rect 266 3927 324 3961
rect 266 3893 278 3927
rect 312 3893 324 3927
rect 266 3859 324 3893
rect 266 3825 278 3859
rect 312 3825 324 3859
rect 266 3791 324 3825
rect 266 3757 278 3791
rect 312 3757 324 3791
rect 266 3723 324 3757
rect 266 3689 278 3723
rect 312 3689 324 3723
rect 266 3655 324 3689
rect 266 3621 278 3655
rect 312 3621 324 3655
rect 266 3587 324 3621
rect 266 3553 278 3587
rect 312 3553 324 3587
rect 266 3519 324 3553
rect 266 3485 278 3519
rect 312 3485 324 3519
rect 266 3451 324 3485
rect 266 3417 278 3451
rect 312 3417 324 3451
rect 266 3383 324 3417
rect 266 3349 278 3383
rect 312 3349 324 3383
rect 266 3315 324 3349
rect 266 3281 278 3315
rect 312 3281 324 3315
rect 266 3247 324 3281
rect 266 3213 278 3247
rect 312 3213 324 3247
rect 266 3179 324 3213
rect 266 3145 278 3179
rect 312 3145 324 3179
rect 266 3111 324 3145
rect 266 3077 278 3111
rect 312 3077 324 3111
rect 266 3043 324 3077
rect 266 3009 278 3043
rect 312 3009 324 3043
rect 266 2975 324 3009
rect 266 2941 278 2975
rect 312 2941 324 2975
rect 266 2907 324 2941
rect 266 2873 278 2907
rect 312 2873 324 2907
rect 266 2839 324 2873
rect 266 2805 278 2839
rect 312 2805 324 2839
rect 266 2771 324 2805
rect 266 2737 278 2771
rect 312 2737 324 2771
rect 266 2703 324 2737
rect 266 2669 278 2703
rect 312 2669 324 2703
rect 266 2635 324 2669
rect 266 2601 278 2635
rect 312 2601 324 2635
rect 266 2567 324 2601
rect 266 2533 278 2567
rect 312 2533 324 2567
rect 266 2499 324 2533
rect 266 2465 278 2499
rect 312 2465 324 2499
rect 266 2431 324 2465
rect 266 2397 278 2431
rect 312 2397 324 2431
rect 266 2363 324 2397
rect 266 2329 278 2363
rect 312 2329 324 2363
rect 266 2295 324 2329
rect 266 2261 278 2295
rect 312 2261 324 2295
rect 266 2227 324 2261
rect 266 2193 278 2227
rect 312 2193 324 2227
rect 266 2159 324 2193
rect 266 2125 278 2159
rect 312 2125 324 2159
rect 266 2091 324 2125
rect 266 2057 278 2091
rect 312 2057 324 2091
rect 266 2023 324 2057
rect 266 1989 278 2023
rect 312 1989 324 2023
rect 266 1955 324 1989
rect 266 1921 278 1955
rect 312 1921 324 1955
rect 266 1887 324 1921
rect 266 1853 278 1887
rect 312 1853 324 1887
rect 266 1819 324 1853
rect 266 1785 278 1819
rect 312 1785 324 1819
rect 266 1751 324 1785
rect 266 1717 278 1751
rect 312 1717 324 1751
rect 266 1683 324 1717
rect 266 1649 278 1683
rect 312 1649 324 1683
rect 266 1615 324 1649
rect 266 1581 278 1615
rect 312 1581 324 1615
rect 266 1547 324 1581
rect 266 1513 278 1547
rect 312 1513 324 1547
rect 266 1479 324 1513
rect 266 1445 278 1479
rect 312 1445 324 1479
rect 266 1411 324 1445
rect 266 1377 278 1411
rect 312 1377 324 1411
rect 266 1343 324 1377
rect 266 1309 278 1343
rect 312 1309 324 1343
rect 266 1275 324 1309
rect 266 1241 278 1275
rect 312 1241 324 1275
rect 266 1207 324 1241
rect 266 1173 278 1207
rect 312 1173 324 1207
rect 266 1139 324 1173
rect 266 1105 278 1139
rect 312 1105 324 1139
rect 266 1071 324 1105
rect 266 1037 278 1071
rect 312 1037 324 1071
rect 266 1003 324 1037
rect 266 969 278 1003
rect 312 969 324 1003
rect 266 935 324 969
rect 266 901 278 935
rect 312 901 324 935
rect 266 867 324 901
rect 266 833 278 867
rect 312 833 324 867
rect 266 799 324 833
rect 266 765 278 799
rect 312 765 324 799
rect 266 731 324 765
rect 266 697 278 731
rect 312 697 324 731
rect 266 663 324 697
rect 266 629 278 663
rect 312 629 324 663
rect 266 595 324 629
rect 266 561 278 595
rect 312 561 324 595
rect 266 527 324 561
rect 266 493 278 527
rect 312 493 324 527
rect 266 459 324 493
rect 266 425 278 459
rect 312 425 324 459
rect 266 391 324 425
rect 266 357 278 391
rect 312 357 324 391
rect 266 323 324 357
rect 266 289 278 323
rect 312 289 324 323
rect 266 255 324 289
rect 266 221 278 255
rect 312 221 324 255
rect 266 187 324 221
rect 266 153 278 187
rect 312 153 324 187
rect 266 119 324 153
rect 266 85 278 119
rect 312 85 324 119
rect 266 51 324 85
rect 266 17 278 51
rect 312 17 324 51
rect 266 -17 324 17
rect 266 -51 278 -17
rect 312 -51 324 -17
rect 266 -85 324 -51
rect 266 -119 278 -85
rect 312 -119 324 -85
rect 266 -153 324 -119
rect 266 -187 278 -153
rect 312 -187 324 -153
rect 266 -221 324 -187
rect 266 -255 278 -221
rect 312 -255 324 -221
rect 266 -289 324 -255
rect 266 -323 278 -289
rect 312 -323 324 -289
rect 266 -357 324 -323
rect 266 -391 278 -357
rect 312 -391 324 -357
rect 266 -425 324 -391
rect 266 -459 278 -425
rect 312 -459 324 -425
rect 266 -493 324 -459
rect 266 -527 278 -493
rect 312 -527 324 -493
rect 266 -561 324 -527
rect 266 -595 278 -561
rect 312 -595 324 -561
rect 266 -629 324 -595
rect 266 -663 278 -629
rect 312 -663 324 -629
rect 266 -697 324 -663
rect 266 -731 278 -697
rect 312 -731 324 -697
rect 266 -765 324 -731
rect 266 -799 278 -765
rect 312 -799 324 -765
rect 266 -833 324 -799
rect 266 -867 278 -833
rect 312 -867 324 -833
rect 266 -901 324 -867
rect 266 -935 278 -901
rect 312 -935 324 -901
rect 266 -969 324 -935
rect 266 -1003 278 -969
rect 312 -1003 324 -969
rect 266 -1037 324 -1003
rect 266 -1071 278 -1037
rect 312 -1071 324 -1037
rect 266 -1105 324 -1071
rect 266 -1139 278 -1105
rect 312 -1139 324 -1105
rect 266 -1173 324 -1139
rect 266 -1207 278 -1173
rect 312 -1207 324 -1173
rect 266 -1241 324 -1207
rect 266 -1275 278 -1241
rect 312 -1275 324 -1241
rect 266 -1309 324 -1275
rect 266 -1343 278 -1309
rect 312 -1343 324 -1309
rect 266 -1377 324 -1343
rect 266 -1411 278 -1377
rect 312 -1411 324 -1377
rect 266 -1445 324 -1411
rect 266 -1479 278 -1445
rect 312 -1479 324 -1445
rect 266 -1513 324 -1479
rect 266 -1547 278 -1513
rect 312 -1547 324 -1513
rect 266 -1581 324 -1547
rect 266 -1615 278 -1581
rect 312 -1615 324 -1581
rect 266 -1649 324 -1615
rect 266 -1683 278 -1649
rect 312 -1683 324 -1649
rect 266 -1717 324 -1683
rect 266 -1751 278 -1717
rect 312 -1751 324 -1717
rect 266 -1785 324 -1751
rect 266 -1819 278 -1785
rect 312 -1819 324 -1785
rect 266 -1853 324 -1819
rect 266 -1887 278 -1853
rect 312 -1887 324 -1853
rect 266 -1921 324 -1887
rect 266 -1955 278 -1921
rect 312 -1955 324 -1921
rect 266 -1989 324 -1955
rect 266 -2023 278 -1989
rect 312 -2023 324 -1989
rect 266 -2057 324 -2023
rect 266 -2091 278 -2057
rect 312 -2091 324 -2057
rect 266 -2125 324 -2091
rect 266 -2159 278 -2125
rect 312 -2159 324 -2125
rect 266 -2193 324 -2159
rect 266 -2227 278 -2193
rect 312 -2227 324 -2193
rect 266 -2261 324 -2227
rect 266 -2295 278 -2261
rect 312 -2295 324 -2261
rect 266 -2329 324 -2295
rect 266 -2363 278 -2329
rect 312 -2363 324 -2329
rect 266 -2397 324 -2363
rect 266 -2431 278 -2397
rect 312 -2431 324 -2397
rect 266 -2465 324 -2431
rect 266 -2499 278 -2465
rect 312 -2499 324 -2465
rect 266 -2533 324 -2499
rect 266 -2567 278 -2533
rect 312 -2567 324 -2533
rect 266 -2601 324 -2567
rect 266 -2635 278 -2601
rect 312 -2635 324 -2601
rect 266 -2669 324 -2635
rect 266 -2703 278 -2669
rect 312 -2703 324 -2669
rect 266 -2737 324 -2703
rect 266 -2771 278 -2737
rect 312 -2771 324 -2737
rect 266 -2805 324 -2771
rect 266 -2839 278 -2805
rect 312 -2839 324 -2805
rect 266 -2873 324 -2839
rect 266 -2907 278 -2873
rect 312 -2907 324 -2873
rect 266 -2941 324 -2907
rect 266 -2975 278 -2941
rect 312 -2975 324 -2941
rect 266 -3009 324 -2975
rect 266 -3043 278 -3009
rect 312 -3043 324 -3009
rect 266 -3077 324 -3043
rect 266 -3111 278 -3077
rect 312 -3111 324 -3077
rect 266 -3145 324 -3111
rect 266 -3179 278 -3145
rect 312 -3179 324 -3145
rect 266 -3213 324 -3179
rect 266 -3247 278 -3213
rect 312 -3247 324 -3213
rect 266 -3281 324 -3247
rect 266 -3315 278 -3281
rect 312 -3315 324 -3281
rect 266 -3349 324 -3315
rect 266 -3383 278 -3349
rect 312 -3383 324 -3349
rect 266 -3417 324 -3383
rect 266 -3451 278 -3417
rect 312 -3451 324 -3417
rect 266 -3485 324 -3451
rect 266 -3519 278 -3485
rect 312 -3519 324 -3485
rect 266 -3553 324 -3519
rect 266 -3587 278 -3553
rect 312 -3587 324 -3553
rect 266 -3621 324 -3587
rect 266 -3655 278 -3621
rect 312 -3655 324 -3621
rect 266 -3689 324 -3655
rect 266 -3723 278 -3689
rect 312 -3723 324 -3689
rect 266 -3757 324 -3723
rect 266 -3791 278 -3757
rect 312 -3791 324 -3757
rect 266 -3825 324 -3791
rect 266 -3859 278 -3825
rect 312 -3859 324 -3825
rect 266 -3893 324 -3859
rect 266 -3927 278 -3893
rect 312 -3927 324 -3893
rect 266 -3961 324 -3927
rect 266 -3995 278 -3961
rect 312 -3995 324 -3961
rect 266 -4029 324 -3995
rect 266 -4063 278 -4029
rect 312 -4063 324 -4029
rect 266 -4097 324 -4063
rect 266 -4131 278 -4097
rect 312 -4131 324 -4097
rect 266 -4165 324 -4131
rect 266 -4199 278 -4165
rect 312 -4199 324 -4165
rect 266 -4233 324 -4199
rect 266 -4267 278 -4233
rect 312 -4267 324 -4233
rect 266 -4301 324 -4267
rect 266 -4335 278 -4301
rect 312 -4335 324 -4301
rect 266 -4369 324 -4335
rect 266 -4403 278 -4369
rect 312 -4403 324 -4369
rect 266 -4437 324 -4403
rect 266 -4471 278 -4437
rect 312 -4471 324 -4437
rect 266 -4505 324 -4471
rect 266 -4539 278 -4505
rect 312 -4539 324 -4505
rect 266 -4573 324 -4539
rect 266 -4607 278 -4573
rect 312 -4607 324 -4573
rect 266 -4641 324 -4607
rect 266 -4675 278 -4641
rect 312 -4675 324 -4641
rect 266 -4709 324 -4675
rect 266 -4743 278 -4709
rect 312 -4743 324 -4709
rect 266 -4777 324 -4743
rect 266 -4811 278 -4777
rect 312 -4811 324 -4777
rect 266 -4845 324 -4811
rect 266 -4879 278 -4845
rect 312 -4879 324 -4845
rect 266 -4913 324 -4879
rect 266 -4947 278 -4913
rect 312 -4947 324 -4913
rect 266 -4981 324 -4947
rect 266 -5015 278 -4981
rect 312 -5015 324 -4981
rect 266 -5049 324 -5015
rect 266 -5083 278 -5049
rect 312 -5083 324 -5049
rect 266 -5117 324 -5083
rect 266 -5151 278 -5117
rect 312 -5151 324 -5117
rect 266 -5185 324 -5151
rect 266 -5219 278 -5185
rect 312 -5219 324 -5185
rect 266 -5253 324 -5219
rect 266 -5287 278 -5253
rect 312 -5287 324 -5253
rect 266 -5321 324 -5287
rect 266 -5355 278 -5321
rect 312 -5355 324 -5321
rect 266 -5389 324 -5355
rect 266 -5423 278 -5389
rect 312 -5423 324 -5389
rect 266 -5457 324 -5423
rect 266 -5491 278 -5457
rect 312 -5491 324 -5457
rect 266 -5525 324 -5491
rect 266 -5559 278 -5525
rect 312 -5559 324 -5525
rect 266 -5593 324 -5559
rect 266 -5627 278 -5593
rect 312 -5627 324 -5593
rect 266 -5661 324 -5627
rect 266 -5695 278 -5661
rect 312 -5695 324 -5661
rect 266 -5729 324 -5695
rect 266 -5763 278 -5729
rect 312 -5763 324 -5729
rect 266 -5797 324 -5763
rect 266 -5831 278 -5797
rect 312 -5831 324 -5797
rect 266 -5865 324 -5831
rect 266 -5899 278 -5865
rect 312 -5899 324 -5865
rect 266 -5933 324 -5899
rect 266 -5967 278 -5933
rect 312 -5967 324 -5933
rect 266 -6001 324 -5967
rect 266 -6035 278 -6001
rect 312 -6035 324 -6001
rect 266 -6069 324 -6035
rect 266 -6103 278 -6069
rect 312 -6103 324 -6069
rect 266 -6137 324 -6103
rect 266 -6171 278 -6137
rect 312 -6171 324 -6137
rect 266 -6205 324 -6171
rect 266 -6239 278 -6205
rect 312 -6239 324 -6205
rect 266 -6273 324 -6239
rect 266 -6307 278 -6273
rect 312 -6307 324 -6273
rect 266 -6341 324 -6307
rect 266 -6375 278 -6341
rect 312 -6375 324 -6341
rect 266 -6409 324 -6375
rect 266 -6443 278 -6409
rect 312 -6443 324 -6409
rect 266 -6477 324 -6443
rect 266 -6511 278 -6477
rect 312 -6511 324 -6477
rect 266 -6545 324 -6511
rect 266 -6579 278 -6545
rect 312 -6579 324 -6545
rect 266 -6613 324 -6579
rect 266 -6647 278 -6613
rect 312 -6647 324 -6613
rect 266 -6681 324 -6647
rect 266 -6715 278 -6681
rect 312 -6715 324 -6681
rect 266 -6749 324 -6715
rect 266 -6783 278 -6749
rect 312 -6783 324 -6749
rect 266 -6817 324 -6783
rect 266 -6851 278 -6817
rect 312 -6851 324 -6817
rect 266 -6885 324 -6851
rect 266 -6919 278 -6885
rect 312 -6919 324 -6885
rect 266 -6953 324 -6919
rect 266 -6987 278 -6953
rect 312 -6987 324 -6953
rect 266 -7021 324 -6987
rect 266 -7055 278 -7021
rect 312 -7055 324 -7021
rect 266 -7089 324 -7055
rect 266 -7123 278 -7089
rect 312 -7123 324 -7089
rect 266 -7157 324 -7123
rect 266 -7191 278 -7157
rect 312 -7191 324 -7157
rect 266 -7225 324 -7191
rect 266 -7259 278 -7225
rect 312 -7259 324 -7225
rect 266 -7293 324 -7259
rect 266 -7327 278 -7293
rect 312 -7327 324 -7293
rect 266 -7361 324 -7327
rect 266 -7395 278 -7361
rect 312 -7395 324 -7361
rect 266 -7429 324 -7395
rect 266 -7463 278 -7429
rect 312 -7463 324 -7429
rect 266 -7497 324 -7463
rect 266 -7531 278 -7497
rect 312 -7531 324 -7497
rect 266 -7565 324 -7531
rect 266 -7599 278 -7565
rect 312 -7599 324 -7565
rect 266 -7633 324 -7599
rect 266 -7667 278 -7633
rect 312 -7667 324 -7633
rect 266 -7701 324 -7667
rect 266 -7735 278 -7701
rect 312 -7735 324 -7701
rect 266 -7769 324 -7735
rect 266 -7803 278 -7769
rect 312 -7803 324 -7769
rect 266 -7837 324 -7803
rect 266 -7871 278 -7837
rect 312 -7871 324 -7837
rect 266 -7905 324 -7871
rect 266 -7939 278 -7905
rect 312 -7939 324 -7905
rect 266 -7973 324 -7939
rect 266 -8007 278 -7973
rect 312 -8007 324 -7973
rect 266 -8041 324 -8007
rect 266 -8075 278 -8041
rect 312 -8075 324 -8041
rect 266 -8109 324 -8075
rect 266 -8143 278 -8109
rect 312 -8143 324 -8109
rect 266 -8177 324 -8143
rect 266 -8211 278 -8177
rect 312 -8211 324 -8177
rect 266 -8245 324 -8211
rect 266 -8279 278 -8245
rect 312 -8279 324 -8245
rect 266 -8313 324 -8279
rect 266 -8347 278 -8313
rect 312 -8347 324 -8313
rect 266 -8381 324 -8347
rect 266 -8415 278 -8381
rect 312 -8415 324 -8381
rect 266 -8449 324 -8415
rect 266 -8483 278 -8449
rect 312 -8483 324 -8449
rect 266 -8517 324 -8483
rect 266 -8551 278 -8517
rect 312 -8551 324 -8517
rect 266 -8585 324 -8551
rect 266 -8619 278 -8585
rect 312 -8619 324 -8585
rect 266 -8653 324 -8619
rect 266 -8687 278 -8653
rect 312 -8687 324 -8653
rect 266 -8721 324 -8687
rect 266 -8755 278 -8721
rect 312 -8755 324 -8721
rect 266 -8789 324 -8755
rect 266 -8823 278 -8789
rect 312 -8823 324 -8789
rect 266 -8857 324 -8823
rect 266 -8891 278 -8857
rect 312 -8891 324 -8857
rect 266 -8925 324 -8891
rect 266 -8959 278 -8925
rect 312 -8959 324 -8925
rect 266 -8993 324 -8959
rect 266 -9027 278 -8993
rect 312 -9027 324 -8993
rect 266 -9061 324 -9027
rect 266 -9095 278 -9061
rect 312 -9095 324 -9061
rect 266 -9129 324 -9095
rect 266 -9163 278 -9129
rect 312 -9163 324 -9129
rect 266 -9197 324 -9163
rect 266 -9231 278 -9197
rect 312 -9231 324 -9197
rect 266 -9265 324 -9231
rect 266 -9299 278 -9265
rect 312 -9299 324 -9265
rect 266 -9333 324 -9299
rect 266 -9367 278 -9333
rect 312 -9367 324 -9333
rect 266 -9401 324 -9367
rect 266 -9435 278 -9401
rect 312 -9435 324 -9401
rect 266 -9469 324 -9435
rect 266 -9503 278 -9469
rect 312 -9503 324 -9469
rect 266 -9537 324 -9503
rect 266 -9571 278 -9537
rect 312 -9571 324 -9537
rect 266 -9600 324 -9571
rect 384 9571 442 9600
rect 384 9537 396 9571
rect 430 9537 442 9571
rect 384 9503 442 9537
rect 384 9469 396 9503
rect 430 9469 442 9503
rect 384 9435 442 9469
rect 384 9401 396 9435
rect 430 9401 442 9435
rect 384 9367 442 9401
rect 384 9333 396 9367
rect 430 9333 442 9367
rect 384 9299 442 9333
rect 384 9265 396 9299
rect 430 9265 442 9299
rect 384 9231 442 9265
rect 384 9197 396 9231
rect 430 9197 442 9231
rect 384 9163 442 9197
rect 384 9129 396 9163
rect 430 9129 442 9163
rect 384 9095 442 9129
rect 384 9061 396 9095
rect 430 9061 442 9095
rect 384 9027 442 9061
rect 384 8993 396 9027
rect 430 8993 442 9027
rect 384 8959 442 8993
rect 384 8925 396 8959
rect 430 8925 442 8959
rect 384 8891 442 8925
rect 384 8857 396 8891
rect 430 8857 442 8891
rect 384 8823 442 8857
rect 384 8789 396 8823
rect 430 8789 442 8823
rect 384 8755 442 8789
rect 384 8721 396 8755
rect 430 8721 442 8755
rect 384 8687 442 8721
rect 384 8653 396 8687
rect 430 8653 442 8687
rect 384 8619 442 8653
rect 384 8585 396 8619
rect 430 8585 442 8619
rect 384 8551 442 8585
rect 384 8517 396 8551
rect 430 8517 442 8551
rect 384 8483 442 8517
rect 384 8449 396 8483
rect 430 8449 442 8483
rect 384 8415 442 8449
rect 384 8381 396 8415
rect 430 8381 442 8415
rect 384 8347 442 8381
rect 384 8313 396 8347
rect 430 8313 442 8347
rect 384 8279 442 8313
rect 384 8245 396 8279
rect 430 8245 442 8279
rect 384 8211 442 8245
rect 384 8177 396 8211
rect 430 8177 442 8211
rect 384 8143 442 8177
rect 384 8109 396 8143
rect 430 8109 442 8143
rect 384 8075 442 8109
rect 384 8041 396 8075
rect 430 8041 442 8075
rect 384 8007 442 8041
rect 384 7973 396 8007
rect 430 7973 442 8007
rect 384 7939 442 7973
rect 384 7905 396 7939
rect 430 7905 442 7939
rect 384 7871 442 7905
rect 384 7837 396 7871
rect 430 7837 442 7871
rect 384 7803 442 7837
rect 384 7769 396 7803
rect 430 7769 442 7803
rect 384 7735 442 7769
rect 384 7701 396 7735
rect 430 7701 442 7735
rect 384 7667 442 7701
rect 384 7633 396 7667
rect 430 7633 442 7667
rect 384 7599 442 7633
rect 384 7565 396 7599
rect 430 7565 442 7599
rect 384 7531 442 7565
rect 384 7497 396 7531
rect 430 7497 442 7531
rect 384 7463 442 7497
rect 384 7429 396 7463
rect 430 7429 442 7463
rect 384 7395 442 7429
rect 384 7361 396 7395
rect 430 7361 442 7395
rect 384 7327 442 7361
rect 384 7293 396 7327
rect 430 7293 442 7327
rect 384 7259 442 7293
rect 384 7225 396 7259
rect 430 7225 442 7259
rect 384 7191 442 7225
rect 384 7157 396 7191
rect 430 7157 442 7191
rect 384 7123 442 7157
rect 384 7089 396 7123
rect 430 7089 442 7123
rect 384 7055 442 7089
rect 384 7021 396 7055
rect 430 7021 442 7055
rect 384 6987 442 7021
rect 384 6953 396 6987
rect 430 6953 442 6987
rect 384 6919 442 6953
rect 384 6885 396 6919
rect 430 6885 442 6919
rect 384 6851 442 6885
rect 384 6817 396 6851
rect 430 6817 442 6851
rect 384 6783 442 6817
rect 384 6749 396 6783
rect 430 6749 442 6783
rect 384 6715 442 6749
rect 384 6681 396 6715
rect 430 6681 442 6715
rect 384 6647 442 6681
rect 384 6613 396 6647
rect 430 6613 442 6647
rect 384 6579 442 6613
rect 384 6545 396 6579
rect 430 6545 442 6579
rect 384 6511 442 6545
rect 384 6477 396 6511
rect 430 6477 442 6511
rect 384 6443 442 6477
rect 384 6409 396 6443
rect 430 6409 442 6443
rect 384 6375 442 6409
rect 384 6341 396 6375
rect 430 6341 442 6375
rect 384 6307 442 6341
rect 384 6273 396 6307
rect 430 6273 442 6307
rect 384 6239 442 6273
rect 384 6205 396 6239
rect 430 6205 442 6239
rect 384 6171 442 6205
rect 384 6137 396 6171
rect 430 6137 442 6171
rect 384 6103 442 6137
rect 384 6069 396 6103
rect 430 6069 442 6103
rect 384 6035 442 6069
rect 384 6001 396 6035
rect 430 6001 442 6035
rect 384 5967 442 6001
rect 384 5933 396 5967
rect 430 5933 442 5967
rect 384 5899 442 5933
rect 384 5865 396 5899
rect 430 5865 442 5899
rect 384 5831 442 5865
rect 384 5797 396 5831
rect 430 5797 442 5831
rect 384 5763 442 5797
rect 384 5729 396 5763
rect 430 5729 442 5763
rect 384 5695 442 5729
rect 384 5661 396 5695
rect 430 5661 442 5695
rect 384 5627 442 5661
rect 384 5593 396 5627
rect 430 5593 442 5627
rect 384 5559 442 5593
rect 384 5525 396 5559
rect 430 5525 442 5559
rect 384 5491 442 5525
rect 384 5457 396 5491
rect 430 5457 442 5491
rect 384 5423 442 5457
rect 384 5389 396 5423
rect 430 5389 442 5423
rect 384 5355 442 5389
rect 384 5321 396 5355
rect 430 5321 442 5355
rect 384 5287 442 5321
rect 384 5253 396 5287
rect 430 5253 442 5287
rect 384 5219 442 5253
rect 384 5185 396 5219
rect 430 5185 442 5219
rect 384 5151 442 5185
rect 384 5117 396 5151
rect 430 5117 442 5151
rect 384 5083 442 5117
rect 384 5049 396 5083
rect 430 5049 442 5083
rect 384 5015 442 5049
rect 384 4981 396 5015
rect 430 4981 442 5015
rect 384 4947 442 4981
rect 384 4913 396 4947
rect 430 4913 442 4947
rect 384 4879 442 4913
rect 384 4845 396 4879
rect 430 4845 442 4879
rect 384 4811 442 4845
rect 384 4777 396 4811
rect 430 4777 442 4811
rect 384 4743 442 4777
rect 384 4709 396 4743
rect 430 4709 442 4743
rect 384 4675 442 4709
rect 384 4641 396 4675
rect 430 4641 442 4675
rect 384 4607 442 4641
rect 384 4573 396 4607
rect 430 4573 442 4607
rect 384 4539 442 4573
rect 384 4505 396 4539
rect 430 4505 442 4539
rect 384 4471 442 4505
rect 384 4437 396 4471
rect 430 4437 442 4471
rect 384 4403 442 4437
rect 384 4369 396 4403
rect 430 4369 442 4403
rect 384 4335 442 4369
rect 384 4301 396 4335
rect 430 4301 442 4335
rect 384 4267 442 4301
rect 384 4233 396 4267
rect 430 4233 442 4267
rect 384 4199 442 4233
rect 384 4165 396 4199
rect 430 4165 442 4199
rect 384 4131 442 4165
rect 384 4097 396 4131
rect 430 4097 442 4131
rect 384 4063 442 4097
rect 384 4029 396 4063
rect 430 4029 442 4063
rect 384 3995 442 4029
rect 384 3961 396 3995
rect 430 3961 442 3995
rect 384 3927 442 3961
rect 384 3893 396 3927
rect 430 3893 442 3927
rect 384 3859 442 3893
rect 384 3825 396 3859
rect 430 3825 442 3859
rect 384 3791 442 3825
rect 384 3757 396 3791
rect 430 3757 442 3791
rect 384 3723 442 3757
rect 384 3689 396 3723
rect 430 3689 442 3723
rect 384 3655 442 3689
rect 384 3621 396 3655
rect 430 3621 442 3655
rect 384 3587 442 3621
rect 384 3553 396 3587
rect 430 3553 442 3587
rect 384 3519 442 3553
rect 384 3485 396 3519
rect 430 3485 442 3519
rect 384 3451 442 3485
rect 384 3417 396 3451
rect 430 3417 442 3451
rect 384 3383 442 3417
rect 384 3349 396 3383
rect 430 3349 442 3383
rect 384 3315 442 3349
rect 384 3281 396 3315
rect 430 3281 442 3315
rect 384 3247 442 3281
rect 384 3213 396 3247
rect 430 3213 442 3247
rect 384 3179 442 3213
rect 384 3145 396 3179
rect 430 3145 442 3179
rect 384 3111 442 3145
rect 384 3077 396 3111
rect 430 3077 442 3111
rect 384 3043 442 3077
rect 384 3009 396 3043
rect 430 3009 442 3043
rect 384 2975 442 3009
rect 384 2941 396 2975
rect 430 2941 442 2975
rect 384 2907 442 2941
rect 384 2873 396 2907
rect 430 2873 442 2907
rect 384 2839 442 2873
rect 384 2805 396 2839
rect 430 2805 442 2839
rect 384 2771 442 2805
rect 384 2737 396 2771
rect 430 2737 442 2771
rect 384 2703 442 2737
rect 384 2669 396 2703
rect 430 2669 442 2703
rect 384 2635 442 2669
rect 384 2601 396 2635
rect 430 2601 442 2635
rect 384 2567 442 2601
rect 384 2533 396 2567
rect 430 2533 442 2567
rect 384 2499 442 2533
rect 384 2465 396 2499
rect 430 2465 442 2499
rect 384 2431 442 2465
rect 384 2397 396 2431
rect 430 2397 442 2431
rect 384 2363 442 2397
rect 384 2329 396 2363
rect 430 2329 442 2363
rect 384 2295 442 2329
rect 384 2261 396 2295
rect 430 2261 442 2295
rect 384 2227 442 2261
rect 384 2193 396 2227
rect 430 2193 442 2227
rect 384 2159 442 2193
rect 384 2125 396 2159
rect 430 2125 442 2159
rect 384 2091 442 2125
rect 384 2057 396 2091
rect 430 2057 442 2091
rect 384 2023 442 2057
rect 384 1989 396 2023
rect 430 1989 442 2023
rect 384 1955 442 1989
rect 384 1921 396 1955
rect 430 1921 442 1955
rect 384 1887 442 1921
rect 384 1853 396 1887
rect 430 1853 442 1887
rect 384 1819 442 1853
rect 384 1785 396 1819
rect 430 1785 442 1819
rect 384 1751 442 1785
rect 384 1717 396 1751
rect 430 1717 442 1751
rect 384 1683 442 1717
rect 384 1649 396 1683
rect 430 1649 442 1683
rect 384 1615 442 1649
rect 384 1581 396 1615
rect 430 1581 442 1615
rect 384 1547 442 1581
rect 384 1513 396 1547
rect 430 1513 442 1547
rect 384 1479 442 1513
rect 384 1445 396 1479
rect 430 1445 442 1479
rect 384 1411 442 1445
rect 384 1377 396 1411
rect 430 1377 442 1411
rect 384 1343 442 1377
rect 384 1309 396 1343
rect 430 1309 442 1343
rect 384 1275 442 1309
rect 384 1241 396 1275
rect 430 1241 442 1275
rect 384 1207 442 1241
rect 384 1173 396 1207
rect 430 1173 442 1207
rect 384 1139 442 1173
rect 384 1105 396 1139
rect 430 1105 442 1139
rect 384 1071 442 1105
rect 384 1037 396 1071
rect 430 1037 442 1071
rect 384 1003 442 1037
rect 384 969 396 1003
rect 430 969 442 1003
rect 384 935 442 969
rect 384 901 396 935
rect 430 901 442 935
rect 384 867 442 901
rect 384 833 396 867
rect 430 833 442 867
rect 384 799 442 833
rect 384 765 396 799
rect 430 765 442 799
rect 384 731 442 765
rect 384 697 396 731
rect 430 697 442 731
rect 384 663 442 697
rect 384 629 396 663
rect 430 629 442 663
rect 384 595 442 629
rect 384 561 396 595
rect 430 561 442 595
rect 384 527 442 561
rect 384 493 396 527
rect 430 493 442 527
rect 384 459 442 493
rect 384 425 396 459
rect 430 425 442 459
rect 384 391 442 425
rect 384 357 396 391
rect 430 357 442 391
rect 384 323 442 357
rect 384 289 396 323
rect 430 289 442 323
rect 384 255 442 289
rect 384 221 396 255
rect 430 221 442 255
rect 384 187 442 221
rect 384 153 396 187
rect 430 153 442 187
rect 384 119 442 153
rect 384 85 396 119
rect 430 85 442 119
rect 384 51 442 85
rect 384 17 396 51
rect 430 17 442 51
rect 384 -17 442 17
rect 384 -51 396 -17
rect 430 -51 442 -17
rect 384 -85 442 -51
rect 384 -119 396 -85
rect 430 -119 442 -85
rect 384 -153 442 -119
rect 384 -187 396 -153
rect 430 -187 442 -153
rect 384 -221 442 -187
rect 384 -255 396 -221
rect 430 -255 442 -221
rect 384 -289 442 -255
rect 384 -323 396 -289
rect 430 -323 442 -289
rect 384 -357 442 -323
rect 384 -391 396 -357
rect 430 -391 442 -357
rect 384 -425 442 -391
rect 384 -459 396 -425
rect 430 -459 442 -425
rect 384 -493 442 -459
rect 384 -527 396 -493
rect 430 -527 442 -493
rect 384 -561 442 -527
rect 384 -595 396 -561
rect 430 -595 442 -561
rect 384 -629 442 -595
rect 384 -663 396 -629
rect 430 -663 442 -629
rect 384 -697 442 -663
rect 384 -731 396 -697
rect 430 -731 442 -697
rect 384 -765 442 -731
rect 384 -799 396 -765
rect 430 -799 442 -765
rect 384 -833 442 -799
rect 384 -867 396 -833
rect 430 -867 442 -833
rect 384 -901 442 -867
rect 384 -935 396 -901
rect 430 -935 442 -901
rect 384 -969 442 -935
rect 384 -1003 396 -969
rect 430 -1003 442 -969
rect 384 -1037 442 -1003
rect 384 -1071 396 -1037
rect 430 -1071 442 -1037
rect 384 -1105 442 -1071
rect 384 -1139 396 -1105
rect 430 -1139 442 -1105
rect 384 -1173 442 -1139
rect 384 -1207 396 -1173
rect 430 -1207 442 -1173
rect 384 -1241 442 -1207
rect 384 -1275 396 -1241
rect 430 -1275 442 -1241
rect 384 -1309 442 -1275
rect 384 -1343 396 -1309
rect 430 -1343 442 -1309
rect 384 -1377 442 -1343
rect 384 -1411 396 -1377
rect 430 -1411 442 -1377
rect 384 -1445 442 -1411
rect 384 -1479 396 -1445
rect 430 -1479 442 -1445
rect 384 -1513 442 -1479
rect 384 -1547 396 -1513
rect 430 -1547 442 -1513
rect 384 -1581 442 -1547
rect 384 -1615 396 -1581
rect 430 -1615 442 -1581
rect 384 -1649 442 -1615
rect 384 -1683 396 -1649
rect 430 -1683 442 -1649
rect 384 -1717 442 -1683
rect 384 -1751 396 -1717
rect 430 -1751 442 -1717
rect 384 -1785 442 -1751
rect 384 -1819 396 -1785
rect 430 -1819 442 -1785
rect 384 -1853 442 -1819
rect 384 -1887 396 -1853
rect 430 -1887 442 -1853
rect 384 -1921 442 -1887
rect 384 -1955 396 -1921
rect 430 -1955 442 -1921
rect 384 -1989 442 -1955
rect 384 -2023 396 -1989
rect 430 -2023 442 -1989
rect 384 -2057 442 -2023
rect 384 -2091 396 -2057
rect 430 -2091 442 -2057
rect 384 -2125 442 -2091
rect 384 -2159 396 -2125
rect 430 -2159 442 -2125
rect 384 -2193 442 -2159
rect 384 -2227 396 -2193
rect 430 -2227 442 -2193
rect 384 -2261 442 -2227
rect 384 -2295 396 -2261
rect 430 -2295 442 -2261
rect 384 -2329 442 -2295
rect 384 -2363 396 -2329
rect 430 -2363 442 -2329
rect 384 -2397 442 -2363
rect 384 -2431 396 -2397
rect 430 -2431 442 -2397
rect 384 -2465 442 -2431
rect 384 -2499 396 -2465
rect 430 -2499 442 -2465
rect 384 -2533 442 -2499
rect 384 -2567 396 -2533
rect 430 -2567 442 -2533
rect 384 -2601 442 -2567
rect 384 -2635 396 -2601
rect 430 -2635 442 -2601
rect 384 -2669 442 -2635
rect 384 -2703 396 -2669
rect 430 -2703 442 -2669
rect 384 -2737 442 -2703
rect 384 -2771 396 -2737
rect 430 -2771 442 -2737
rect 384 -2805 442 -2771
rect 384 -2839 396 -2805
rect 430 -2839 442 -2805
rect 384 -2873 442 -2839
rect 384 -2907 396 -2873
rect 430 -2907 442 -2873
rect 384 -2941 442 -2907
rect 384 -2975 396 -2941
rect 430 -2975 442 -2941
rect 384 -3009 442 -2975
rect 384 -3043 396 -3009
rect 430 -3043 442 -3009
rect 384 -3077 442 -3043
rect 384 -3111 396 -3077
rect 430 -3111 442 -3077
rect 384 -3145 442 -3111
rect 384 -3179 396 -3145
rect 430 -3179 442 -3145
rect 384 -3213 442 -3179
rect 384 -3247 396 -3213
rect 430 -3247 442 -3213
rect 384 -3281 442 -3247
rect 384 -3315 396 -3281
rect 430 -3315 442 -3281
rect 384 -3349 442 -3315
rect 384 -3383 396 -3349
rect 430 -3383 442 -3349
rect 384 -3417 442 -3383
rect 384 -3451 396 -3417
rect 430 -3451 442 -3417
rect 384 -3485 442 -3451
rect 384 -3519 396 -3485
rect 430 -3519 442 -3485
rect 384 -3553 442 -3519
rect 384 -3587 396 -3553
rect 430 -3587 442 -3553
rect 384 -3621 442 -3587
rect 384 -3655 396 -3621
rect 430 -3655 442 -3621
rect 384 -3689 442 -3655
rect 384 -3723 396 -3689
rect 430 -3723 442 -3689
rect 384 -3757 442 -3723
rect 384 -3791 396 -3757
rect 430 -3791 442 -3757
rect 384 -3825 442 -3791
rect 384 -3859 396 -3825
rect 430 -3859 442 -3825
rect 384 -3893 442 -3859
rect 384 -3927 396 -3893
rect 430 -3927 442 -3893
rect 384 -3961 442 -3927
rect 384 -3995 396 -3961
rect 430 -3995 442 -3961
rect 384 -4029 442 -3995
rect 384 -4063 396 -4029
rect 430 -4063 442 -4029
rect 384 -4097 442 -4063
rect 384 -4131 396 -4097
rect 430 -4131 442 -4097
rect 384 -4165 442 -4131
rect 384 -4199 396 -4165
rect 430 -4199 442 -4165
rect 384 -4233 442 -4199
rect 384 -4267 396 -4233
rect 430 -4267 442 -4233
rect 384 -4301 442 -4267
rect 384 -4335 396 -4301
rect 430 -4335 442 -4301
rect 384 -4369 442 -4335
rect 384 -4403 396 -4369
rect 430 -4403 442 -4369
rect 384 -4437 442 -4403
rect 384 -4471 396 -4437
rect 430 -4471 442 -4437
rect 384 -4505 442 -4471
rect 384 -4539 396 -4505
rect 430 -4539 442 -4505
rect 384 -4573 442 -4539
rect 384 -4607 396 -4573
rect 430 -4607 442 -4573
rect 384 -4641 442 -4607
rect 384 -4675 396 -4641
rect 430 -4675 442 -4641
rect 384 -4709 442 -4675
rect 384 -4743 396 -4709
rect 430 -4743 442 -4709
rect 384 -4777 442 -4743
rect 384 -4811 396 -4777
rect 430 -4811 442 -4777
rect 384 -4845 442 -4811
rect 384 -4879 396 -4845
rect 430 -4879 442 -4845
rect 384 -4913 442 -4879
rect 384 -4947 396 -4913
rect 430 -4947 442 -4913
rect 384 -4981 442 -4947
rect 384 -5015 396 -4981
rect 430 -5015 442 -4981
rect 384 -5049 442 -5015
rect 384 -5083 396 -5049
rect 430 -5083 442 -5049
rect 384 -5117 442 -5083
rect 384 -5151 396 -5117
rect 430 -5151 442 -5117
rect 384 -5185 442 -5151
rect 384 -5219 396 -5185
rect 430 -5219 442 -5185
rect 384 -5253 442 -5219
rect 384 -5287 396 -5253
rect 430 -5287 442 -5253
rect 384 -5321 442 -5287
rect 384 -5355 396 -5321
rect 430 -5355 442 -5321
rect 384 -5389 442 -5355
rect 384 -5423 396 -5389
rect 430 -5423 442 -5389
rect 384 -5457 442 -5423
rect 384 -5491 396 -5457
rect 430 -5491 442 -5457
rect 384 -5525 442 -5491
rect 384 -5559 396 -5525
rect 430 -5559 442 -5525
rect 384 -5593 442 -5559
rect 384 -5627 396 -5593
rect 430 -5627 442 -5593
rect 384 -5661 442 -5627
rect 384 -5695 396 -5661
rect 430 -5695 442 -5661
rect 384 -5729 442 -5695
rect 384 -5763 396 -5729
rect 430 -5763 442 -5729
rect 384 -5797 442 -5763
rect 384 -5831 396 -5797
rect 430 -5831 442 -5797
rect 384 -5865 442 -5831
rect 384 -5899 396 -5865
rect 430 -5899 442 -5865
rect 384 -5933 442 -5899
rect 384 -5967 396 -5933
rect 430 -5967 442 -5933
rect 384 -6001 442 -5967
rect 384 -6035 396 -6001
rect 430 -6035 442 -6001
rect 384 -6069 442 -6035
rect 384 -6103 396 -6069
rect 430 -6103 442 -6069
rect 384 -6137 442 -6103
rect 384 -6171 396 -6137
rect 430 -6171 442 -6137
rect 384 -6205 442 -6171
rect 384 -6239 396 -6205
rect 430 -6239 442 -6205
rect 384 -6273 442 -6239
rect 384 -6307 396 -6273
rect 430 -6307 442 -6273
rect 384 -6341 442 -6307
rect 384 -6375 396 -6341
rect 430 -6375 442 -6341
rect 384 -6409 442 -6375
rect 384 -6443 396 -6409
rect 430 -6443 442 -6409
rect 384 -6477 442 -6443
rect 384 -6511 396 -6477
rect 430 -6511 442 -6477
rect 384 -6545 442 -6511
rect 384 -6579 396 -6545
rect 430 -6579 442 -6545
rect 384 -6613 442 -6579
rect 384 -6647 396 -6613
rect 430 -6647 442 -6613
rect 384 -6681 442 -6647
rect 384 -6715 396 -6681
rect 430 -6715 442 -6681
rect 384 -6749 442 -6715
rect 384 -6783 396 -6749
rect 430 -6783 442 -6749
rect 384 -6817 442 -6783
rect 384 -6851 396 -6817
rect 430 -6851 442 -6817
rect 384 -6885 442 -6851
rect 384 -6919 396 -6885
rect 430 -6919 442 -6885
rect 384 -6953 442 -6919
rect 384 -6987 396 -6953
rect 430 -6987 442 -6953
rect 384 -7021 442 -6987
rect 384 -7055 396 -7021
rect 430 -7055 442 -7021
rect 384 -7089 442 -7055
rect 384 -7123 396 -7089
rect 430 -7123 442 -7089
rect 384 -7157 442 -7123
rect 384 -7191 396 -7157
rect 430 -7191 442 -7157
rect 384 -7225 442 -7191
rect 384 -7259 396 -7225
rect 430 -7259 442 -7225
rect 384 -7293 442 -7259
rect 384 -7327 396 -7293
rect 430 -7327 442 -7293
rect 384 -7361 442 -7327
rect 384 -7395 396 -7361
rect 430 -7395 442 -7361
rect 384 -7429 442 -7395
rect 384 -7463 396 -7429
rect 430 -7463 442 -7429
rect 384 -7497 442 -7463
rect 384 -7531 396 -7497
rect 430 -7531 442 -7497
rect 384 -7565 442 -7531
rect 384 -7599 396 -7565
rect 430 -7599 442 -7565
rect 384 -7633 442 -7599
rect 384 -7667 396 -7633
rect 430 -7667 442 -7633
rect 384 -7701 442 -7667
rect 384 -7735 396 -7701
rect 430 -7735 442 -7701
rect 384 -7769 442 -7735
rect 384 -7803 396 -7769
rect 430 -7803 442 -7769
rect 384 -7837 442 -7803
rect 384 -7871 396 -7837
rect 430 -7871 442 -7837
rect 384 -7905 442 -7871
rect 384 -7939 396 -7905
rect 430 -7939 442 -7905
rect 384 -7973 442 -7939
rect 384 -8007 396 -7973
rect 430 -8007 442 -7973
rect 384 -8041 442 -8007
rect 384 -8075 396 -8041
rect 430 -8075 442 -8041
rect 384 -8109 442 -8075
rect 384 -8143 396 -8109
rect 430 -8143 442 -8109
rect 384 -8177 442 -8143
rect 384 -8211 396 -8177
rect 430 -8211 442 -8177
rect 384 -8245 442 -8211
rect 384 -8279 396 -8245
rect 430 -8279 442 -8245
rect 384 -8313 442 -8279
rect 384 -8347 396 -8313
rect 430 -8347 442 -8313
rect 384 -8381 442 -8347
rect 384 -8415 396 -8381
rect 430 -8415 442 -8381
rect 384 -8449 442 -8415
rect 384 -8483 396 -8449
rect 430 -8483 442 -8449
rect 384 -8517 442 -8483
rect 384 -8551 396 -8517
rect 430 -8551 442 -8517
rect 384 -8585 442 -8551
rect 384 -8619 396 -8585
rect 430 -8619 442 -8585
rect 384 -8653 442 -8619
rect 384 -8687 396 -8653
rect 430 -8687 442 -8653
rect 384 -8721 442 -8687
rect 384 -8755 396 -8721
rect 430 -8755 442 -8721
rect 384 -8789 442 -8755
rect 384 -8823 396 -8789
rect 430 -8823 442 -8789
rect 384 -8857 442 -8823
rect 384 -8891 396 -8857
rect 430 -8891 442 -8857
rect 384 -8925 442 -8891
rect 384 -8959 396 -8925
rect 430 -8959 442 -8925
rect 384 -8993 442 -8959
rect 384 -9027 396 -8993
rect 430 -9027 442 -8993
rect 384 -9061 442 -9027
rect 384 -9095 396 -9061
rect 430 -9095 442 -9061
rect 384 -9129 442 -9095
rect 384 -9163 396 -9129
rect 430 -9163 442 -9129
rect 384 -9197 442 -9163
rect 384 -9231 396 -9197
rect 430 -9231 442 -9197
rect 384 -9265 442 -9231
rect 384 -9299 396 -9265
rect 430 -9299 442 -9265
rect 384 -9333 442 -9299
rect 384 -9367 396 -9333
rect 430 -9367 442 -9333
rect 384 -9401 442 -9367
rect 384 -9435 396 -9401
rect 430 -9435 442 -9401
rect 384 -9469 442 -9435
rect 384 -9503 396 -9469
rect 430 -9503 442 -9469
rect 384 -9537 442 -9503
rect 384 -9571 396 -9537
rect 430 -9571 442 -9537
rect 384 -9600 442 -9571
rect 502 9571 560 9600
rect 502 9537 514 9571
rect 548 9537 560 9571
rect 502 9503 560 9537
rect 502 9469 514 9503
rect 548 9469 560 9503
rect 502 9435 560 9469
rect 502 9401 514 9435
rect 548 9401 560 9435
rect 502 9367 560 9401
rect 502 9333 514 9367
rect 548 9333 560 9367
rect 502 9299 560 9333
rect 502 9265 514 9299
rect 548 9265 560 9299
rect 502 9231 560 9265
rect 502 9197 514 9231
rect 548 9197 560 9231
rect 502 9163 560 9197
rect 502 9129 514 9163
rect 548 9129 560 9163
rect 502 9095 560 9129
rect 502 9061 514 9095
rect 548 9061 560 9095
rect 502 9027 560 9061
rect 502 8993 514 9027
rect 548 8993 560 9027
rect 502 8959 560 8993
rect 502 8925 514 8959
rect 548 8925 560 8959
rect 502 8891 560 8925
rect 502 8857 514 8891
rect 548 8857 560 8891
rect 502 8823 560 8857
rect 502 8789 514 8823
rect 548 8789 560 8823
rect 502 8755 560 8789
rect 502 8721 514 8755
rect 548 8721 560 8755
rect 502 8687 560 8721
rect 502 8653 514 8687
rect 548 8653 560 8687
rect 502 8619 560 8653
rect 502 8585 514 8619
rect 548 8585 560 8619
rect 502 8551 560 8585
rect 502 8517 514 8551
rect 548 8517 560 8551
rect 502 8483 560 8517
rect 502 8449 514 8483
rect 548 8449 560 8483
rect 502 8415 560 8449
rect 502 8381 514 8415
rect 548 8381 560 8415
rect 502 8347 560 8381
rect 502 8313 514 8347
rect 548 8313 560 8347
rect 502 8279 560 8313
rect 502 8245 514 8279
rect 548 8245 560 8279
rect 502 8211 560 8245
rect 502 8177 514 8211
rect 548 8177 560 8211
rect 502 8143 560 8177
rect 502 8109 514 8143
rect 548 8109 560 8143
rect 502 8075 560 8109
rect 502 8041 514 8075
rect 548 8041 560 8075
rect 502 8007 560 8041
rect 502 7973 514 8007
rect 548 7973 560 8007
rect 502 7939 560 7973
rect 502 7905 514 7939
rect 548 7905 560 7939
rect 502 7871 560 7905
rect 502 7837 514 7871
rect 548 7837 560 7871
rect 502 7803 560 7837
rect 502 7769 514 7803
rect 548 7769 560 7803
rect 502 7735 560 7769
rect 502 7701 514 7735
rect 548 7701 560 7735
rect 502 7667 560 7701
rect 502 7633 514 7667
rect 548 7633 560 7667
rect 502 7599 560 7633
rect 502 7565 514 7599
rect 548 7565 560 7599
rect 502 7531 560 7565
rect 502 7497 514 7531
rect 548 7497 560 7531
rect 502 7463 560 7497
rect 502 7429 514 7463
rect 548 7429 560 7463
rect 502 7395 560 7429
rect 502 7361 514 7395
rect 548 7361 560 7395
rect 502 7327 560 7361
rect 502 7293 514 7327
rect 548 7293 560 7327
rect 502 7259 560 7293
rect 502 7225 514 7259
rect 548 7225 560 7259
rect 502 7191 560 7225
rect 502 7157 514 7191
rect 548 7157 560 7191
rect 502 7123 560 7157
rect 502 7089 514 7123
rect 548 7089 560 7123
rect 502 7055 560 7089
rect 502 7021 514 7055
rect 548 7021 560 7055
rect 502 6987 560 7021
rect 502 6953 514 6987
rect 548 6953 560 6987
rect 502 6919 560 6953
rect 502 6885 514 6919
rect 548 6885 560 6919
rect 502 6851 560 6885
rect 502 6817 514 6851
rect 548 6817 560 6851
rect 502 6783 560 6817
rect 502 6749 514 6783
rect 548 6749 560 6783
rect 502 6715 560 6749
rect 502 6681 514 6715
rect 548 6681 560 6715
rect 502 6647 560 6681
rect 502 6613 514 6647
rect 548 6613 560 6647
rect 502 6579 560 6613
rect 502 6545 514 6579
rect 548 6545 560 6579
rect 502 6511 560 6545
rect 502 6477 514 6511
rect 548 6477 560 6511
rect 502 6443 560 6477
rect 502 6409 514 6443
rect 548 6409 560 6443
rect 502 6375 560 6409
rect 502 6341 514 6375
rect 548 6341 560 6375
rect 502 6307 560 6341
rect 502 6273 514 6307
rect 548 6273 560 6307
rect 502 6239 560 6273
rect 502 6205 514 6239
rect 548 6205 560 6239
rect 502 6171 560 6205
rect 502 6137 514 6171
rect 548 6137 560 6171
rect 502 6103 560 6137
rect 502 6069 514 6103
rect 548 6069 560 6103
rect 502 6035 560 6069
rect 502 6001 514 6035
rect 548 6001 560 6035
rect 502 5967 560 6001
rect 502 5933 514 5967
rect 548 5933 560 5967
rect 502 5899 560 5933
rect 502 5865 514 5899
rect 548 5865 560 5899
rect 502 5831 560 5865
rect 502 5797 514 5831
rect 548 5797 560 5831
rect 502 5763 560 5797
rect 502 5729 514 5763
rect 548 5729 560 5763
rect 502 5695 560 5729
rect 502 5661 514 5695
rect 548 5661 560 5695
rect 502 5627 560 5661
rect 502 5593 514 5627
rect 548 5593 560 5627
rect 502 5559 560 5593
rect 502 5525 514 5559
rect 548 5525 560 5559
rect 502 5491 560 5525
rect 502 5457 514 5491
rect 548 5457 560 5491
rect 502 5423 560 5457
rect 502 5389 514 5423
rect 548 5389 560 5423
rect 502 5355 560 5389
rect 502 5321 514 5355
rect 548 5321 560 5355
rect 502 5287 560 5321
rect 502 5253 514 5287
rect 548 5253 560 5287
rect 502 5219 560 5253
rect 502 5185 514 5219
rect 548 5185 560 5219
rect 502 5151 560 5185
rect 502 5117 514 5151
rect 548 5117 560 5151
rect 502 5083 560 5117
rect 502 5049 514 5083
rect 548 5049 560 5083
rect 502 5015 560 5049
rect 502 4981 514 5015
rect 548 4981 560 5015
rect 502 4947 560 4981
rect 502 4913 514 4947
rect 548 4913 560 4947
rect 502 4879 560 4913
rect 502 4845 514 4879
rect 548 4845 560 4879
rect 502 4811 560 4845
rect 502 4777 514 4811
rect 548 4777 560 4811
rect 502 4743 560 4777
rect 502 4709 514 4743
rect 548 4709 560 4743
rect 502 4675 560 4709
rect 502 4641 514 4675
rect 548 4641 560 4675
rect 502 4607 560 4641
rect 502 4573 514 4607
rect 548 4573 560 4607
rect 502 4539 560 4573
rect 502 4505 514 4539
rect 548 4505 560 4539
rect 502 4471 560 4505
rect 502 4437 514 4471
rect 548 4437 560 4471
rect 502 4403 560 4437
rect 502 4369 514 4403
rect 548 4369 560 4403
rect 502 4335 560 4369
rect 502 4301 514 4335
rect 548 4301 560 4335
rect 502 4267 560 4301
rect 502 4233 514 4267
rect 548 4233 560 4267
rect 502 4199 560 4233
rect 502 4165 514 4199
rect 548 4165 560 4199
rect 502 4131 560 4165
rect 502 4097 514 4131
rect 548 4097 560 4131
rect 502 4063 560 4097
rect 502 4029 514 4063
rect 548 4029 560 4063
rect 502 3995 560 4029
rect 502 3961 514 3995
rect 548 3961 560 3995
rect 502 3927 560 3961
rect 502 3893 514 3927
rect 548 3893 560 3927
rect 502 3859 560 3893
rect 502 3825 514 3859
rect 548 3825 560 3859
rect 502 3791 560 3825
rect 502 3757 514 3791
rect 548 3757 560 3791
rect 502 3723 560 3757
rect 502 3689 514 3723
rect 548 3689 560 3723
rect 502 3655 560 3689
rect 502 3621 514 3655
rect 548 3621 560 3655
rect 502 3587 560 3621
rect 502 3553 514 3587
rect 548 3553 560 3587
rect 502 3519 560 3553
rect 502 3485 514 3519
rect 548 3485 560 3519
rect 502 3451 560 3485
rect 502 3417 514 3451
rect 548 3417 560 3451
rect 502 3383 560 3417
rect 502 3349 514 3383
rect 548 3349 560 3383
rect 502 3315 560 3349
rect 502 3281 514 3315
rect 548 3281 560 3315
rect 502 3247 560 3281
rect 502 3213 514 3247
rect 548 3213 560 3247
rect 502 3179 560 3213
rect 502 3145 514 3179
rect 548 3145 560 3179
rect 502 3111 560 3145
rect 502 3077 514 3111
rect 548 3077 560 3111
rect 502 3043 560 3077
rect 502 3009 514 3043
rect 548 3009 560 3043
rect 502 2975 560 3009
rect 502 2941 514 2975
rect 548 2941 560 2975
rect 502 2907 560 2941
rect 502 2873 514 2907
rect 548 2873 560 2907
rect 502 2839 560 2873
rect 502 2805 514 2839
rect 548 2805 560 2839
rect 502 2771 560 2805
rect 502 2737 514 2771
rect 548 2737 560 2771
rect 502 2703 560 2737
rect 502 2669 514 2703
rect 548 2669 560 2703
rect 502 2635 560 2669
rect 502 2601 514 2635
rect 548 2601 560 2635
rect 502 2567 560 2601
rect 502 2533 514 2567
rect 548 2533 560 2567
rect 502 2499 560 2533
rect 502 2465 514 2499
rect 548 2465 560 2499
rect 502 2431 560 2465
rect 502 2397 514 2431
rect 548 2397 560 2431
rect 502 2363 560 2397
rect 502 2329 514 2363
rect 548 2329 560 2363
rect 502 2295 560 2329
rect 502 2261 514 2295
rect 548 2261 560 2295
rect 502 2227 560 2261
rect 502 2193 514 2227
rect 548 2193 560 2227
rect 502 2159 560 2193
rect 502 2125 514 2159
rect 548 2125 560 2159
rect 502 2091 560 2125
rect 502 2057 514 2091
rect 548 2057 560 2091
rect 502 2023 560 2057
rect 502 1989 514 2023
rect 548 1989 560 2023
rect 502 1955 560 1989
rect 502 1921 514 1955
rect 548 1921 560 1955
rect 502 1887 560 1921
rect 502 1853 514 1887
rect 548 1853 560 1887
rect 502 1819 560 1853
rect 502 1785 514 1819
rect 548 1785 560 1819
rect 502 1751 560 1785
rect 502 1717 514 1751
rect 548 1717 560 1751
rect 502 1683 560 1717
rect 502 1649 514 1683
rect 548 1649 560 1683
rect 502 1615 560 1649
rect 502 1581 514 1615
rect 548 1581 560 1615
rect 502 1547 560 1581
rect 502 1513 514 1547
rect 548 1513 560 1547
rect 502 1479 560 1513
rect 502 1445 514 1479
rect 548 1445 560 1479
rect 502 1411 560 1445
rect 502 1377 514 1411
rect 548 1377 560 1411
rect 502 1343 560 1377
rect 502 1309 514 1343
rect 548 1309 560 1343
rect 502 1275 560 1309
rect 502 1241 514 1275
rect 548 1241 560 1275
rect 502 1207 560 1241
rect 502 1173 514 1207
rect 548 1173 560 1207
rect 502 1139 560 1173
rect 502 1105 514 1139
rect 548 1105 560 1139
rect 502 1071 560 1105
rect 502 1037 514 1071
rect 548 1037 560 1071
rect 502 1003 560 1037
rect 502 969 514 1003
rect 548 969 560 1003
rect 502 935 560 969
rect 502 901 514 935
rect 548 901 560 935
rect 502 867 560 901
rect 502 833 514 867
rect 548 833 560 867
rect 502 799 560 833
rect 502 765 514 799
rect 548 765 560 799
rect 502 731 560 765
rect 502 697 514 731
rect 548 697 560 731
rect 502 663 560 697
rect 502 629 514 663
rect 548 629 560 663
rect 502 595 560 629
rect 502 561 514 595
rect 548 561 560 595
rect 502 527 560 561
rect 502 493 514 527
rect 548 493 560 527
rect 502 459 560 493
rect 502 425 514 459
rect 548 425 560 459
rect 502 391 560 425
rect 502 357 514 391
rect 548 357 560 391
rect 502 323 560 357
rect 502 289 514 323
rect 548 289 560 323
rect 502 255 560 289
rect 502 221 514 255
rect 548 221 560 255
rect 502 187 560 221
rect 502 153 514 187
rect 548 153 560 187
rect 502 119 560 153
rect 502 85 514 119
rect 548 85 560 119
rect 502 51 560 85
rect 502 17 514 51
rect 548 17 560 51
rect 502 -17 560 17
rect 502 -51 514 -17
rect 548 -51 560 -17
rect 502 -85 560 -51
rect 502 -119 514 -85
rect 548 -119 560 -85
rect 502 -153 560 -119
rect 502 -187 514 -153
rect 548 -187 560 -153
rect 502 -221 560 -187
rect 502 -255 514 -221
rect 548 -255 560 -221
rect 502 -289 560 -255
rect 502 -323 514 -289
rect 548 -323 560 -289
rect 502 -357 560 -323
rect 502 -391 514 -357
rect 548 -391 560 -357
rect 502 -425 560 -391
rect 502 -459 514 -425
rect 548 -459 560 -425
rect 502 -493 560 -459
rect 502 -527 514 -493
rect 548 -527 560 -493
rect 502 -561 560 -527
rect 502 -595 514 -561
rect 548 -595 560 -561
rect 502 -629 560 -595
rect 502 -663 514 -629
rect 548 -663 560 -629
rect 502 -697 560 -663
rect 502 -731 514 -697
rect 548 -731 560 -697
rect 502 -765 560 -731
rect 502 -799 514 -765
rect 548 -799 560 -765
rect 502 -833 560 -799
rect 502 -867 514 -833
rect 548 -867 560 -833
rect 502 -901 560 -867
rect 502 -935 514 -901
rect 548 -935 560 -901
rect 502 -969 560 -935
rect 502 -1003 514 -969
rect 548 -1003 560 -969
rect 502 -1037 560 -1003
rect 502 -1071 514 -1037
rect 548 -1071 560 -1037
rect 502 -1105 560 -1071
rect 502 -1139 514 -1105
rect 548 -1139 560 -1105
rect 502 -1173 560 -1139
rect 502 -1207 514 -1173
rect 548 -1207 560 -1173
rect 502 -1241 560 -1207
rect 502 -1275 514 -1241
rect 548 -1275 560 -1241
rect 502 -1309 560 -1275
rect 502 -1343 514 -1309
rect 548 -1343 560 -1309
rect 502 -1377 560 -1343
rect 502 -1411 514 -1377
rect 548 -1411 560 -1377
rect 502 -1445 560 -1411
rect 502 -1479 514 -1445
rect 548 -1479 560 -1445
rect 502 -1513 560 -1479
rect 502 -1547 514 -1513
rect 548 -1547 560 -1513
rect 502 -1581 560 -1547
rect 502 -1615 514 -1581
rect 548 -1615 560 -1581
rect 502 -1649 560 -1615
rect 502 -1683 514 -1649
rect 548 -1683 560 -1649
rect 502 -1717 560 -1683
rect 502 -1751 514 -1717
rect 548 -1751 560 -1717
rect 502 -1785 560 -1751
rect 502 -1819 514 -1785
rect 548 -1819 560 -1785
rect 502 -1853 560 -1819
rect 502 -1887 514 -1853
rect 548 -1887 560 -1853
rect 502 -1921 560 -1887
rect 502 -1955 514 -1921
rect 548 -1955 560 -1921
rect 502 -1989 560 -1955
rect 502 -2023 514 -1989
rect 548 -2023 560 -1989
rect 502 -2057 560 -2023
rect 502 -2091 514 -2057
rect 548 -2091 560 -2057
rect 502 -2125 560 -2091
rect 502 -2159 514 -2125
rect 548 -2159 560 -2125
rect 502 -2193 560 -2159
rect 502 -2227 514 -2193
rect 548 -2227 560 -2193
rect 502 -2261 560 -2227
rect 502 -2295 514 -2261
rect 548 -2295 560 -2261
rect 502 -2329 560 -2295
rect 502 -2363 514 -2329
rect 548 -2363 560 -2329
rect 502 -2397 560 -2363
rect 502 -2431 514 -2397
rect 548 -2431 560 -2397
rect 502 -2465 560 -2431
rect 502 -2499 514 -2465
rect 548 -2499 560 -2465
rect 502 -2533 560 -2499
rect 502 -2567 514 -2533
rect 548 -2567 560 -2533
rect 502 -2601 560 -2567
rect 502 -2635 514 -2601
rect 548 -2635 560 -2601
rect 502 -2669 560 -2635
rect 502 -2703 514 -2669
rect 548 -2703 560 -2669
rect 502 -2737 560 -2703
rect 502 -2771 514 -2737
rect 548 -2771 560 -2737
rect 502 -2805 560 -2771
rect 502 -2839 514 -2805
rect 548 -2839 560 -2805
rect 502 -2873 560 -2839
rect 502 -2907 514 -2873
rect 548 -2907 560 -2873
rect 502 -2941 560 -2907
rect 502 -2975 514 -2941
rect 548 -2975 560 -2941
rect 502 -3009 560 -2975
rect 502 -3043 514 -3009
rect 548 -3043 560 -3009
rect 502 -3077 560 -3043
rect 502 -3111 514 -3077
rect 548 -3111 560 -3077
rect 502 -3145 560 -3111
rect 502 -3179 514 -3145
rect 548 -3179 560 -3145
rect 502 -3213 560 -3179
rect 502 -3247 514 -3213
rect 548 -3247 560 -3213
rect 502 -3281 560 -3247
rect 502 -3315 514 -3281
rect 548 -3315 560 -3281
rect 502 -3349 560 -3315
rect 502 -3383 514 -3349
rect 548 -3383 560 -3349
rect 502 -3417 560 -3383
rect 502 -3451 514 -3417
rect 548 -3451 560 -3417
rect 502 -3485 560 -3451
rect 502 -3519 514 -3485
rect 548 -3519 560 -3485
rect 502 -3553 560 -3519
rect 502 -3587 514 -3553
rect 548 -3587 560 -3553
rect 502 -3621 560 -3587
rect 502 -3655 514 -3621
rect 548 -3655 560 -3621
rect 502 -3689 560 -3655
rect 502 -3723 514 -3689
rect 548 -3723 560 -3689
rect 502 -3757 560 -3723
rect 502 -3791 514 -3757
rect 548 -3791 560 -3757
rect 502 -3825 560 -3791
rect 502 -3859 514 -3825
rect 548 -3859 560 -3825
rect 502 -3893 560 -3859
rect 502 -3927 514 -3893
rect 548 -3927 560 -3893
rect 502 -3961 560 -3927
rect 502 -3995 514 -3961
rect 548 -3995 560 -3961
rect 502 -4029 560 -3995
rect 502 -4063 514 -4029
rect 548 -4063 560 -4029
rect 502 -4097 560 -4063
rect 502 -4131 514 -4097
rect 548 -4131 560 -4097
rect 502 -4165 560 -4131
rect 502 -4199 514 -4165
rect 548 -4199 560 -4165
rect 502 -4233 560 -4199
rect 502 -4267 514 -4233
rect 548 -4267 560 -4233
rect 502 -4301 560 -4267
rect 502 -4335 514 -4301
rect 548 -4335 560 -4301
rect 502 -4369 560 -4335
rect 502 -4403 514 -4369
rect 548 -4403 560 -4369
rect 502 -4437 560 -4403
rect 502 -4471 514 -4437
rect 548 -4471 560 -4437
rect 502 -4505 560 -4471
rect 502 -4539 514 -4505
rect 548 -4539 560 -4505
rect 502 -4573 560 -4539
rect 502 -4607 514 -4573
rect 548 -4607 560 -4573
rect 502 -4641 560 -4607
rect 502 -4675 514 -4641
rect 548 -4675 560 -4641
rect 502 -4709 560 -4675
rect 502 -4743 514 -4709
rect 548 -4743 560 -4709
rect 502 -4777 560 -4743
rect 502 -4811 514 -4777
rect 548 -4811 560 -4777
rect 502 -4845 560 -4811
rect 502 -4879 514 -4845
rect 548 -4879 560 -4845
rect 502 -4913 560 -4879
rect 502 -4947 514 -4913
rect 548 -4947 560 -4913
rect 502 -4981 560 -4947
rect 502 -5015 514 -4981
rect 548 -5015 560 -4981
rect 502 -5049 560 -5015
rect 502 -5083 514 -5049
rect 548 -5083 560 -5049
rect 502 -5117 560 -5083
rect 502 -5151 514 -5117
rect 548 -5151 560 -5117
rect 502 -5185 560 -5151
rect 502 -5219 514 -5185
rect 548 -5219 560 -5185
rect 502 -5253 560 -5219
rect 502 -5287 514 -5253
rect 548 -5287 560 -5253
rect 502 -5321 560 -5287
rect 502 -5355 514 -5321
rect 548 -5355 560 -5321
rect 502 -5389 560 -5355
rect 502 -5423 514 -5389
rect 548 -5423 560 -5389
rect 502 -5457 560 -5423
rect 502 -5491 514 -5457
rect 548 -5491 560 -5457
rect 502 -5525 560 -5491
rect 502 -5559 514 -5525
rect 548 -5559 560 -5525
rect 502 -5593 560 -5559
rect 502 -5627 514 -5593
rect 548 -5627 560 -5593
rect 502 -5661 560 -5627
rect 502 -5695 514 -5661
rect 548 -5695 560 -5661
rect 502 -5729 560 -5695
rect 502 -5763 514 -5729
rect 548 -5763 560 -5729
rect 502 -5797 560 -5763
rect 502 -5831 514 -5797
rect 548 -5831 560 -5797
rect 502 -5865 560 -5831
rect 502 -5899 514 -5865
rect 548 -5899 560 -5865
rect 502 -5933 560 -5899
rect 502 -5967 514 -5933
rect 548 -5967 560 -5933
rect 502 -6001 560 -5967
rect 502 -6035 514 -6001
rect 548 -6035 560 -6001
rect 502 -6069 560 -6035
rect 502 -6103 514 -6069
rect 548 -6103 560 -6069
rect 502 -6137 560 -6103
rect 502 -6171 514 -6137
rect 548 -6171 560 -6137
rect 502 -6205 560 -6171
rect 502 -6239 514 -6205
rect 548 -6239 560 -6205
rect 502 -6273 560 -6239
rect 502 -6307 514 -6273
rect 548 -6307 560 -6273
rect 502 -6341 560 -6307
rect 502 -6375 514 -6341
rect 548 -6375 560 -6341
rect 502 -6409 560 -6375
rect 502 -6443 514 -6409
rect 548 -6443 560 -6409
rect 502 -6477 560 -6443
rect 502 -6511 514 -6477
rect 548 -6511 560 -6477
rect 502 -6545 560 -6511
rect 502 -6579 514 -6545
rect 548 -6579 560 -6545
rect 502 -6613 560 -6579
rect 502 -6647 514 -6613
rect 548 -6647 560 -6613
rect 502 -6681 560 -6647
rect 502 -6715 514 -6681
rect 548 -6715 560 -6681
rect 502 -6749 560 -6715
rect 502 -6783 514 -6749
rect 548 -6783 560 -6749
rect 502 -6817 560 -6783
rect 502 -6851 514 -6817
rect 548 -6851 560 -6817
rect 502 -6885 560 -6851
rect 502 -6919 514 -6885
rect 548 -6919 560 -6885
rect 502 -6953 560 -6919
rect 502 -6987 514 -6953
rect 548 -6987 560 -6953
rect 502 -7021 560 -6987
rect 502 -7055 514 -7021
rect 548 -7055 560 -7021
rect 502 -7089 560 -7055
rect 502 -7123 514 -7089
rect 548 -7123 560 -7089
rect 502 -7157 560 -7123
rect 502 -7191 514 -7157
rect 548 -7191 560 -7157
rect 502 -7225 560 -7191
rect 502 -7259 514 -7225
rect 548 -7259 560 -7225
rect 502 -7293 560 -7259
rect 502 -7327 514 -7293
rect 548 -7327 560 -7293
rect 502 -7361 560 -7327
rect 502 -7395 514 -7361
rect 548 -7395 560 -7361
rect 502 -7429 560 -7395
rect 502 -7463 514 -7429
rect 548 -7463 560 -7429
rect 502 -7497 560 -7463
rect 502 -7531 514 -7497
rect 548 -7531 560 -7497
rect 502 -7565 560 -7531
rect 502 -7599 514 -7565
rect 548 -7599 560 -7565
rect 502 -7633 560 -7599
rect 502 -7667 514 -7633
rect 548 -7667 560 -7633
rect 502 -7701 560 -7667
rect 502 -7735 514 -7701
rect 548 -7735 560 -7701
rect 502 -7769 560 -7735
rect 502 -7803 514 -7769
rect 548 -7803 560 -7769
rect 502 -7837 560 -7803
rect 502 -7871 514 -7837
rect 548 -7871 560 -7837
rect 502 -7905 560 -7871
rect 502 -7939 514 -7905
rect 548 -7939 560 -7905
rect 502 -7973 560 -7939
rect 502 -8007 514 -7973
rect 548 -8007 560 -7973
rect 502 -8041 560 -8007
rect 502 -8075 514 -8041
rect 548 -8075 560 -8041
rect 502 -8109 560 -8075
rect 502 -8143 514 -8109
rect 548 -8143 560 -8109
rect 502 -8177 560 -8143
rect 502 -8211 514 -8177
rect 548 -8211 560 -8177
rect 502 -8245 560 -8211
rect 502 -8279 514 -8245
rect 548 -8279 560 -8245
rect 502 -8313 560 -8279
rect 502 -8347 514 -8313
rect 548 -8347 560 -8313
rect 502 -8381 560 -8347
rect 502 -8415 514 -8381
rect 548 -8415 560 -8381
rect 502 -8449 560 -8415
rect 502 -8483 514 -8449
rect 548 -8483 560 -8449
rect 502 -8517 560 -8483
rect 502 -8551 514 -8517
rect 548 -8551 560 -8517
rect 502 -8585 560 -8551
rect 502 -8619 514 -8585
rect 548 -8619 560 -8585
rect 502 -8653 560 -8619
rect 502 -8687 514 -8653
rect 548 -8687 560 -8653
rect 502 -8721 560 -8687
rect 502 -8755 514 -8721
rect 548 -8755 560 -8721
rect 502 -8789 560 -8755
rect 502 -8823 514 -8789
rect 548 -8823 560 -8789
rect 502 -8857 560 -8823
rect 502 -8891 514 -8857
rect 548 -8891 560 -8857
rect 502 -8925 560 -8891
rect 502 -8959 514 -8925
rect 548 -8959 560 -8925
rect 502 -8993 560 -8959
rect 502 -9027 514 -8993
rect 548 -9027 560 -8993
rect 502 -9061 560 -9027
rect 502 -9095 514 -9061
rect 548 -9095 560 -9061
rect 502 -9129 560 -9095
rect 502 -9163 514 -9129
rect 548 -9163 560 -9129
rect 502 -9197 560 -9163
rect 502 -9231 514 -9197
rect 548 -9231 560 -9197
rect 502 -9265 560 -9231
rect 502 -9299 514 -9265
rect 548 -9299 560 -9265
rect 502 -9333 560 -9299
rect 502 -9367 514 -9333
rect 548 -9367 560 -9333
rect 502 -9401 560 -9367
rect 502 -9435 514 -9401
rect 548 -9435 560 -9401
rect 502 -9469 560 -9435
rect 502 -9503 514 -9469
rect 548 -9503 560 -9469
rect 502 -9537 560 -9503
rect 502 -9571 514 -9537
rect 548 -9571 560 -9537
rect 502 -9600 560 -9571
rect 620 9571 678 9600
rect 620 9537 632 9571
rect 666 9537 678 9571
rect 620 9503 678 9537
rect 620 9469 632 9503
rect 666 9469 678 9503
rect 620 9435 678 9469
rect 620 9401 632 9435
rect 666 9401 678 9435
rect 620 9367 678 9401
rect 620 9333 632 9367
rect 666 9333 678 9367
rect 620 9299 678 9333
rect 620 9265 632 9299
rect 666 9265 678 9299
rect 620 9231 678 9265
rect 620 9197 632 9231
rect 666 9197 678 9231
rect 620 9163 678 9197
rect 620 9129 632 9163
rect 666 9129 678 9163
rect 620 9095 678 9129
rect 620 9061 632 9095
rect 666 9061 678 9095
rect 620 9027 678 9061
rect 620 8993 632 9027
rect 666 8993 678 9027
rect 620 8959 678 8993
rect 620 8925 632 8959
rect 666 8925 678 8959
rect 620 8891 678 8925
rect 620 8857 632 8891
rect 666 8857 678 8891
rect 620 8823 678 8857
rect 620 8789 632 8823
rect 666 8789 678 8823
rect 620 8755 678 8789
rect 620 8721 632 8755
rect 666 8721 678 8755
rect 620 8687 678 8721
rect 620 8653 632 8687
rect 666 8653 678 8687
rect 620 8619 678 8653
rect 620 8585 632 8619
rect 666 8585 678 8619
rect 620 8551 678 8585
rect 620 8517 632 8551
rect 666 8517 678 8551
rect 620 8483 678 8517
rect 620 8449 632 8483
rect 666 8449 678 8483
rect 620 8415 678 8449
rect 620 8381 632 8415
rect 666 8381 678 8415
rect 620 8347 678 8381
rect 620 8313 632 8347
rect 666 8313 678 8347
rect 620 8279 678 8313
rect 620 8245 632 8279
rect 666 8245 678 8279
rect 620 8211 678 8245
rect 620 8177 632 8211
rect 666 8177 678 8211
rect 620 8143 678 8177
rect 620 8109 632 8143
rect 666 8109 678 8143
rect 620 8075 678 8109
rect 620 8041 632 8075
rect 666 8041 678 8075
rect 620 8007 678 8041
rect 620 7973 632 8007
rect 666 7973 678 8007
rect 620 7939 678 7973
rect 620 7905 632 7939
rect 666 7905 678 7939
rect 620 7871 678 7905
rect 620 7837 632 7871
rect 666 7837 678 7871
rect 620 7803 678 7837
rect 620 7769 632 7803
rect 666 7769 678 7803
rect 620 7735 678 7769
rect 620 7701 632 7735
rect 666 7701 678 7735
rect 620 7667 678 7701
rect 620 7633 632 7667
rect 666 7633 678 7667
rect 620 7599 678 7633
rect 620 7565 632 7599
rect 666 7565 678 7599
rect 620 7531 678 7565
rect 620 7497 632 7531
rect 666 7497 678 7531
rect 620 7463 678 7497
rect 620 7429 632 7463
rect 666 7429 678 7463
rect 620 7395 678 7429
rect 620 7361 632 7395
rect 666 7361 678 7395
rect 620 7327 678 7361
rect 620 7293 632 7327
rect 666 7293 678 7327
rect 620 7259 678 7293
rect 620 7225 632 7259
rect 666 7225 678 7259
rect 620 7191 678 7225
rect 620 7157 632 7191
rect 666 7157 678 7191
rect 620 7123 678 7157
rect 620 7089 632 7123
rect 666 7089 678 7123
rect 620 7055 678 7089
rect 620 7021 632 7055
rect 666 7021 678 7055
rect 620 6987 678 7021
rect 620 6953 632 6987
rect 666 6953 678 6987
rect 620 6919 678 6953
rect 620 6885 632 6919
rect 666 6885 678 6919
rect 620 6851 678 6885
rect 620 6817 632 6851
rect 666 6817 678 6851
rect 620 6783 678 6817
rect 620 6749 632 6783
rect 666 6749 678 6783
rect 620 6715 678 6749
rect 620 6681 632 6715
rect 666 6681 678 6715
rect 620 6647 678 6681
rect 620 6613 632 6647
rect 666 6613 678 6647
rect 620 6579 678 6613
rect 620 6545 632 6579
rect 666 6545 678 6579
rect 620 6511 678 6545
rect 620 6477 632 6511
rect 666 6477 678 6511
rect 620 6443 678 6477
rect 620 6409 632 6443
rect 666 6409 678 6443
rect 620 6375 678 6409
rect 620 6341 632 6375
rect 666 6341 678 6375
rect 620 6307 678 6341
rect 620 6273 632 6307
rect 666 6273 678 6307
rect 620 6239 678 6273
rect 620 6205 632 6239
rect 666 6205 678 6239
rect 620 6171 678 6205
rect 620 6137 632 6171
rect 666 6137 678 6171
rect 620 6103 678 6137
rect 620 6069 632 6103
rect 666 6069 678 6103
rect 620 6035 678 6069
rect 620 6001 632 6035
rect 666 6001 678 6035
rect 620 5967 678 6001
rect 620 5933 632 5967
rect 666 5933 678 5967
rect 620 5899 678 5933
rect 620 5865 632 5899
rect 666 5865 678 5899
rect 620 5831 678 5865
rect 620 5797 632 5831
rect 666 5797 678 5831
rect 620 5763 678 5797
rect 620 5729 632 5763
rect 666 5729 678 5763
rect 620 5695 678 5729
rect 620 5661 632 5695
rect 666 5661 678 5695
rect 620 5627 678 5661
rect 620 5593 632 5627
rect 666 5593 678 5627
rect 620 5559 678 5593
rect 620 5525 632 5559
rect 666 5525 678 5559
rect 620 5491 678 5525
rect 620 5457 632 5491
rect 666 5457 678 5491
rect 620 5423 678 5457
rect 620 5389 632 5423
rect 666 5389 678 5423
rect 620 5355 678 5389
rect 620 5321 632 5355
rect 666 5321 678 5355
rect 620 5287 678 5321
rect 620 5253 632 5287
rect 666 5253 678 5287
rect 620 5219 678 5253
rect 620 5185 632 5219
rect 666 5185 678 5219
rect 620 5151 678 5185
rect 620 5117 632 5151
rect 666 5117 678 5151
rect 620 5083 678 5117
rect 620 5049 632 5083
rect 666 5049 678 5083
rect 620 5015 678 5049
rect 620 4981 632 5015
rect 666 4981 678 5015
rect 620 4947 678 4981
rect 620 4913 632 4947
rect 666 4913 678 4947
rect 620 4879 678 4913
rect 620 4845 632 4879
rect 666 4845 678 4879
rect 620 4811 678 4845
rect 620 4777 632 4811
rect 666 4777 678 4811
rect 620 4743 678 4777
rect 620 4709 632 4743
rect 666 4709 678 4743
rect 620 4675 678 4709
rect 620 4641 632 4675
rect 666 4641 678 4675
rect 620 4607 678 4641
rect 620 4573 632 4607
rect 666 4573 678 4607
rect 620 4539 678 4573
rect 620 4505 632 4539
rect 666 4505 678 4539
rect 620 4471 678 4505
rect 620 4437 632 4471
rect 666 4437 678 4471
rect 620 4403 678 4437
rect 620 4369 632 4403
rect 666 4369 678 4403
rect 620 4335 678 4369
rect 620 4301 632 4335
rect 666 4301 678 4335
rect 620 4267 678 4301
rect 620 4233 632 4267
rect 666 4233 678 4267
rect 620 4199 678 4233
rect 620 4165 632 4199
rect 666 4165 678 4199
rect 620 4131 678 4165
rect 620 4097 632 4131
rect 666 4097 678 4131
rect 620 4063 678 4097
rect 620 4029 632 4063
rect 666 4029 678 4063
rect 620 3995 678 4029
rect 620 3961 632 3995
rect 666 3961 678 3995
rect 620 3927 678 3961
rect 620 3893 632 3927
rect 666 3893 678 3927
rect 620 3859 678 3893
rect 620 3825 632 3859
rect 666 3825 678 3859
rect 620 3791 678 3825
rect 620 3757 632 3791
rect 666 3757 678 3791
rect 620 3723 678 3757
rect 620 3689 632 3723
rect 666 3689 678 3723
rect 620 3655 678 3689
rect 620 3621 632 3655
rect 666 3621 678 3655
rect 620 3587 678 3621
rect 620 3553 632 3587
rect 666 3553 678 3587
rect 620 3519 678 3553
rect 620 3485 632 3519
rect 666 3485 678 3519
rect 620 3451 678 3485
rect 620 3417 632 3451
rect 666 3417 678 3451
rect 620 3383 678 3417
rect 620 3349 632 3383
rect 666 3349 678 3383
rect 620 3315 678 3349
rect 620 3281 632 3315
rect 666 3281 678 3315
rect 620 3247 678 3281
rect 620 3213 632 3247
rect 666 3213 678 3247
rect 620 3179 678 3213
rect 620 3145 632 3179
rect 666 3145 678 3179
rect 620 3111 678 3145
rect 620 3077 632 3111
rect 666 3077 678 3111
rect 620 3043 678 3077
rect 620 3009 632 3043
rect 666 3009 678 3043
rect 620 2975 678 3009
rect 620 2941 632 2975
rect 666 2941 678 2975
rect 620 2907 678 2941
rect 620 2873 632 2907
rect 666 2873 678 2907
rect 620 2839 678 2873
rect 620 2805 632 2839
rect 666 2805 678 2839
rect 620 2771 678 2805
rect 620 2737 632 2771
rect 666 2737 678 2771
rect 620 2703 678 2737
rect 620 2669 632 2703
rect 666 2669 678 2703
rect 620 2635 678 2669
rect 620 2601 632 2635
rect 666 2601 678 2635
rect 620 2567 678 2601
rect 620 2533 632 2567
rect 666 2533 678 2567
rect 620 2499 678 2533
rect 620 2465 632 2499
rect 666 2465 678 2499
rect 620 2431 678 2465
rect 620 2397 632 2431
rect 666 2397 678 2431
rect 620 2363 678 2397
rect 620 2329 632 2363
rect 666 2329 678 2363
rect 620 2295 678 2329
rect 620 2261 632 2295
rect 666 2261 678 2295
rect 620 2227 678 2261
rect 620 2193 632 2227
rect 666 2193 678 2227
rect 620 2159 678 2193
rect 620 2125 632 2159
rect 666 2125 678 2159
rect 620 2091 678 2125
rect 620 2057 632 2091
rect 666 2057 678 2091
rect 620 2023 678 2057
rect 620 1989 632 2023
rect 666 1989 678 2023
rect 620 1955 678 1989
rect 620 1921 632 1955
rect 666 1921 678 1955
rect 620 1887 678 1921
rect 620 1853 632 1887
rect 666 1853 678 1887
rect 620 1819 678 1853
rect 620 1785 632 1819
rect 666 1785 678 1819
rect 620 1751 678 1785
rect 620 1717 632 1751
rect 666 1717 678 1751
rect 620 1683 678 1717
rect 620 1649 632 1683
rect 666 1649 678 1683
rect 620 1615 678 1649
rect 620 1581 632 1615
rect 666 1581 678 1615
rect 620 1547 678 1581
rect 620 1513 632 1547
rect 666 1513 678 1547
rect 620 1479 678 1513
rect 620 1445 632 1479
rect 666 1445 678 1479
rect 620 1411 678 1445
rect 620 1377 632 1411
rect 666 1377 678 1411
rect 620 1343 678 1377
rect 620 1309 632 1343
rect 666 1309 678 1343
rect 620 1275 678 1309
rect 620 1241 632 1275
rect 666 1241 678 1275
rect 620 1207 678 1241
rect 620 1173 632 1207
rect 666 1173 678 1207
rect 620 1139 678 1173
rect 620 1105 632 1139
rect 666 1105 678 1139
rect 620 1071 678 1105
rect 620 1037 632 1071
rect 666 1037 678 1071
rect 620 1003 678 1037
rect 620 969 632 1003
rect 666 969 678 1003
rect 620 935 678 969
rect 620 901 632 935
rect 666 901 678 935
rect 620 867 678 901
rect 620 833 632 867
rect 666 833 678 867
rect 620 799 678 833
rect 620 765 632 799
rect 666 765 678 799
rect 620 731 678 765
rect 620 697 632 731
rect 666 697 678 731
rect 620 663 678 697
rect 620 629 632 663
rect 666 629 678 663
rect 620 595 678 629
rect 620 561 632 595
rect 666 561 678 595
rect 620 527 678 561
rect 620 493 632 527
rect 666 493 678 527
rect 620 459 678 493
rect 620 425 632 459
rect 666 425 678 459
rect 620 391 678 425
rect 620 357 632 391
rect 666 357 678 391
rect 620 323 678 357
rect 620 289 632 323
rect 666 289 678 323
rect 620 255 678 289
rect 620 221 632 255
rect 666 221 678 255
rect 620 187 678 221
rect 620 153 632 187
rect 666 153 678 187
rect 620 119 678 153
rect 620 85 632 119
rect 666 85 678 119
rect 620 51 678 85
rect 620 17 632 51
rect 666 17 678 51
rect 620 -17 678 17
rect 620 -51 632 -17
rect 666 -51 678 -17
rect 620 -85 678 -51
rect 620 -119 632 -85
rect 666 -119 678 -85
rect 620 -153 678 -119
rect 620 -187 632 -153
rect 666 -187 678 -153
rect 620 -221 678 -187
rect 620 -255 632 -221
rect 666 -255 678 -221
rect 620 -289 678 -255
rect 620 -323 632 -289
rect 666 -323 678 -289
rect 620 -357 678 -323
rect 620 -391 632 -357
rect 666 -391 678 -357
rect 620 -425 678 -391
rect 620 -459 632 -425
rect 666 -459 678 -425
rect 620 -493 678 -459
rect 620 -527 632 -493
rect 666 -527 678 -493
rect 620 -561 678 -527
rect 620 -595 632 -561
rect 666 -595 678 -561
rect 620 -629 678 -595
rect 620 -663 632 -629
rect 666 -663 678 -629
rect 620 -697 678 -663
rect 620 -731 632 -697
rect 666 -731 678 -697
rect 620 -765 678 -731
rect 620 -799 632 -765
rect 666 -799 678 -765
rect 620 -833 678 -799
rect 620 -867 632 -833
rect 666 -867 678 -833
rect 620 -901 678 -867
rect 620 -935 632 -901
rect 666 -935 678 -901
rect 620 -969 678 -935
rect 620 -1003 632 -969
rect 666 -1003 678 -969
rect 620 -1037 678 -1003
rect 620 -1071 632 -1037
rect 666 -1071 678 -1037
rect 620 -1105 678 -1071
rect 620 -1139 632 -1105
rect 666 -1139 678 -1105
rect 620 -1173 678 -1139
rect 620 -1207 632 -1173
rect 666 -1207 678 -1173
rect 620 -1241 678 -1207
rect 620 -1275 632 -1241
rect 666 -1275 678 -1241
rect 620 -1309 678 -1275
rect 620 -1343 632 -1309
rect 666 -1343 678 -1309
rect 620 -1377 678 -1343
rect 620 -1411 632 -1377
rect 666 -1411 678 -1377
rect 620 -1445 678 -1411
rect 620 -1479 632 -1445
rect 666 -1479 678 -1445
rect 620 -1513 678 -1479
rect 620 -1547 632 -1513
rect 666 -1547 678 -1513
rect 620 -1581 678 -1547
rect 620 -1615 632 -1581
rect 666 -1615 678 -1581
rect 620 -1649 678 -1615
rect 620 -1683 632 -1649
rect 666 -1683 678 -1649
rect 620 -1717 678 -1683
rect 620 -1751 632 -1717
rect 666 -1751 678 -1717
rect 620 -1785 678 -1751
rect 620 -1819 632 -1785
rect 666 -1819 678 -1785
rect 620 -1853 678 -1819
rect 620 -1887 632 -1853
rect 666 -1887 678 -1853
rect 620 -1921 678 -1887
rect 620 -1955 632 -1921
rect 666 -1955 678 -1921
rect 620 -1989 678 -1955
rect 620 -2023 632 -1989
rect 666 -2023 678 -1989
rect 620 -2057 678 -2023
rect 620 -2091 632 -2057
rect 666 -2091 678 -2057
rect 620 -2125 678 -2091
rect 620 -2159 632 -2125
rect 666 -2159 678 -2125
rect 620 -2193 678 -2159
rect 620 -2227 632 -2193
rect 666 -2227 678 -2193
rect 620 -2261 678 -2227
rect 620 -2295 632 -2261
rect 666 -2295 678 -2261
rect 620 -2329 678 -2295
rect 620 -2363 632 -2329
rect 666 -2363 678 -2329
rect 620 -2397 678 -2363
rect 620 -2431 632 -2397
rect 666 -2431 678 -2397
rect 620 -2465 678 -2431
rect 620 -2499 632 -2465
rect 666 -2499 678 -2465
rect 620 -2533 678 -2499
rect 620 -2567 632 -2533
rect 666 -2567 678 -2533
rect 620 -2601 678 -2567
rect 620 -2635 632 -2601
rect 666 -2635 678 -2601
rect 620 -2669 678 -2635
rect 620 -2703 632 -2669
rect 666 -2703 678 -2669
rect 620 -2737 678 -2703
rect 620 -2771 632 -2737
rect 666 -2771 678 -2737
rect 620 -2805 678 -2771
rect 620 -2839 632 -2805
rect 666 -2839 678 -2805
rect 620 -2873 678 -2839
rect 620 -2907 632 -2873
rect 666 -2907 678 -2873
rect 620 -2941 678 -2907
rect 620 -2975 632 -2941
rect 666 -2975 678 -2941
rect 620 -3009 678 -2975
rect 620 -3043 632 -3009
rect 666 -3043 678 -3009
rect 620 -3077 678 -3043
rect 620 -3111 632 -3077
rect 666 -3111 678 -3077
rect 620 -3145 678 -3111
rect 620 -3179 632 -3145
rect 666 -3179 678 -3145
rect 620 -3213 678 -3179
rect 620 -3247 632 -3213
rect 666 -3247 678 -3213
rect 620 -3281 678 -3247
rect 620 -3315 632 -3281
rect 666 -3315 678 -3281
rect 620 -3349 678 -3315
rect 620 -3383 632 -3349
rect 666 -3383 678 -3349
rect 620 -3417 678 -3383
rect 620 -3451 632 -3417
rect 666 -3451 678 -3417
rect 620 -3485 678 -3451
rect 620 -3519 632 -3485
rect 666 -3519 678 -3485
rect 620 -3553 678 -3519
rect 620 -3587 632 -3553
rect 666 -3587 678 -3553
rect 620 -3621 678 -3587
rect 620 -3655 632 -3621
rect 666 -3655 678 -3621
rect 620 -3689 678 -3655
rect 620 -3723 632 -3689
rect 666 -3723 678 -3689
rect 620 -3757 678 -3723
rect 620 -3791 632 -3757
rect 666 -3791 678 -3757
rect 620 -3825 678 -3791
rect 620 -3859 632 -3825
rect 666 -3859 678 -3825
rect 620 -3893 678 -3859
rect 620 -3927 632 -3893
rect 666 -3927 678 -3893
rect 620 -3961 678 -3927
rect 620 -3995 632 -3961
rect 666 -3995 678 -3961
rect 620 -4029 678 -3995
rect 620 -4063 632 -4029
rect 666 -4063 678 -4029
rect 620 -4097 678 -4063
rect 620 -4131 632 -4097
rect 666 -4131 678 -4097
rect 620 -4165 678 -4131
rect 620 -4199 632 -4165
rect 666 -4199 678 -4165
rect 620 -4233 678 -4199
rect 620 -4267 632 -4233
rect 666 -4267 678 -4233
rect 620 -4301 678 -4267
rect 620 -4335 632 -4301
rect 666 -4335 678 -4301
rect 620 -4369 678 -4335
rect 620 -4403 632 -4369
rect 666 -4403 678 -4369
rect 620 -4437 678 -4403
rect 620 -4471 632 -4437
rect 666 -4471 678 -4437
rect 620 -4505 678 -4471
rect 620 -4539 632 -4505
rect 666 -4539 678 -4505
rect 620 -4573 678 -4539
rect 620 -4607 632 -4573
rect 666 -4607 678 -4573
rect 620 -4641 678 -4607
rect 620 -4675 632 -4641
rect 666 -4675 678 -4641
rect 620 -4709 678 -4675
rect 620 -4743 632 -4709
rect 666 -4743 678 -4709
rect 620 -4777 678 -4743
rect 620 -4811 632 -4777
rect 666 -4811 678 -4777
rect 620 -4845 678 -4811
rect 620 -4879 632 -4845
rect 666 -4879 678 -4845
rect 620 -4913 678 -4879
rect 620 -4947 632 -4913
rect 666 -4947 678 -4913
rect 620 -4981 678 -4947
rect 620 -5015 632 -4981
rect 666 -5015 678 -4981
rect 620 -5049 678 -5015
rect 620 -5083 632 -5049
rect 666 -5083 678 -5049
rect 620 -5117 678 -5083
rect 620 -5151 632 -5117
rect 666 -5151 678 -5117
rect 620 -5185 678 -5151
rect 620 -5219 632 -5185
rect 666 -5219 678 -5185
rect 620 -5253 678 -5219
rect 620 -5287 632 -5253
rect 666 -5287 678 -5253
rect 620 -5321 678 -5287
rect 620 -5355 632 -5321
rect 666 -5355 678 -5321
rect 620 -5389 678 -5355
rect 620 -5423 632 -5389
rect 666 -5423 678 -5389
rect 620 -5457 678 -5423
rect 620 -5491 632 -5457
rect 666 -5491 678 -5457
rect 620 -5525 678 -5491
rect 620 -5559 632 -5525
rect 666 -5559 678 -5525
rect 620 -5593 678 -5559
rect 620 -5627 632 -5593
rect 666 -5627 678 -5593
rect 620 -5661 678 -5627
rect 620 -5695 632 -5661
rect 666 -5695 678 -5661
rect 620 -5729 678 -5695
rect 620 -5763 632 -5729
rect 666 -5763 678 -5729
rect 620 -5797 678 -5763
rect 620 -5831 632 -5797
rect 666 -5831 678 -5797
rect 620 -5865 678 -5831
rect 620 -5899 632 -5865
rect 666 -5899 678 -5865
rect 620 -5933 678 -5899
rect 620 -5967 632 -5933
rect 666 -5967 678 -5933
rect 620 -6001 678 -5967
rect 620 -6035 632 -6001
rect 666 -6035 678 -6001
rect 620 -6069 678 -6035
rect 620 -6103 632 -6069
rect 666 -6103 678 -6069
rect 620 -6137 678 -6103
rect 620 -6171 632 -6137
rect 666 -6171 678 -6137
rect 620 -6205 678 -6171
rect 620 -6239 632 -6205
rect 666 -6239 678 -6205
rect 620 -6273 678 -6239
rect 620 -6307 632 -6273
rect 666 -6307 678 -6273
rect 620 -6341 678 -6307
rect 620 -6375 632 -6341
rect 666 -6375 678 -6341
rect 620 -6409 678 -6375
rect 620 -6443 632 -6409
rect 666 -6443 678 -6409
rect 620 -6477 678 -6443
rect 620 -6511 632 -6477
rect 666 -6511 678 -6477
rect 620 -6545 678 -6511
rect 620 -6579 632 -6545
rect 666 -6579 678 -6545
rect 620 -6613 678 -6579
rect 620 -6647 632 -6613
rect 666 -6647 678 -6613
rect 620 -6681 678 -6647
rect 620 -6715 632 -6681
rect 666 -6715 678 -6681
rect 620 -6749 678 -6715
rect 620 -6783 632 -6749
rect 666 -6783 678 -6749
rect 620 -6817 678 -6783
rect 620 -6851 632 -6817
rect 666 -6851 678 -6817
rect 620 -6885 678 -6851
rect 620 -6919 632 -6885
rect 666 -6919 678 -6885
rect 620 -6953 678 -6919
rect 620 -6987 632 -6953
rect 666 -6987 678 -6953
rect 620 -7021 678 -6987
rect 620 -7055 632 -7021
rect 666 -7055 678 -7021
rect 620 -7089 678 -7055
rect 620 -7123 632 -7089
rect 666 -7123 678 -7089
rect 620 -7157 678 -7123
rect 620 -7191 632 -7157
rect 666 -7191 678 -7157
rect 620 -7225 678 -7191
rect 620 -7259 632 -7225
rect 666 -7259 678 -7225
rect 620 -7293 678 -7259
rect 620 -7327 632 -7293
rect 666 -7327 678 -7293
rect 620 -7361 678 -7327
rect 620 -7395 632 -7361
rect 666 -7395 678 -7361
rect 620 -7429 678 -7395
rect 620 -7463 632 -7429
rect 666 -7463 678 -7429
rect 620 -7497 678 -7463
rect 620 -7531 632 -7497
rect 666 -7531 678 -7497
rect 620 -7565 678 -7531
rect 620 -7599 632 -7565
rect 666 -7599 678 -7565
rect 620 -7633 678 -7599
rect 620 -7667 632 -7633
rect 666 -7667 678 -7633
rect 620 -7701 678 -7667
rect 620 -7735 632 -7701
rect 666 -7735 678 -7701
rect 620 -7769 678 -7735
rect 620 -7803 632 -7769
rect 666 -7803 678 -7769
rect 620 -7837 678 -7803
rect 620 -7871 632 -7837
rect 666 -7871 678 -7837
rect 620 -7905 678 -7871
rect 620 -7939 632 -7905
rect 666 -7939 678 -7905
rect 620 -7973 678 -7939
rect 620 -8007 632 -7973
rect 666 -8007 678 -7973
rect 620 -8041 678 -8007
rect 620 -8075 632 -8041
rect 666 -8075 678 -8041
rect 620 -8109 678 -8075
rect 620 -8143 632 -8109
rect 666 -8143 678 -8109
rect 620 -8177 678 -8143
rect 620 -8211 632 -8177
rect 666 -8211 678 -8177
rect 620 -8245 678 -8211
rect 620 -8279 632 -8245
rect 666 -8279 678 -8245
rect 620 -8313 678 -8279
rect 620 -8347 632 -8313
rect 666 -8347 678 -8313
rect 620 -8381 678 -8347
rect 620 -8415 632 -8381
rect 666 -8415 678 -8381
rect 620 -8449 678 -8415
rect 620 -8483 632 -8449
rect 666 -8483 678 -8449
rect 620 -8517 678 -8483
rect 620 -8551 632 -8517
rect 666 -8551 678 -8517
rect 620 -8585 678 -8551
rect 620 -8619 632 -8585
rect 666 -8619 678 -8585
rect 620 -8653 678 -8619
rect 620 -8687 632 -8653
rect 666 -8687 678 -8653
rect 620 -8721 678 -8687
rect 620 -8755 632 -8721
rect 666 -8755 678 -8721
rect 620 -8789 678 -8755
rect 620 -8823 632 -8789
rect 666 -8823 678 -8789
rect 620 -8857 678 -8823
rect 620 -8891 632 -8857
rect 666 -8891 678 -8857
rect 620 -8925 678 -8891
rect 620 -8959 632 -8925
rect 666 -8959 678 -8925
rect 620 -8993 678 -8959
rect 620 -9027 632 -8993
rect 666 -9027 678 -8993
rect 620 -9061 678 -9027
rect 620 -9095 632 -9061
rect 666 -9095 678 -9061
rect 620 -9129 678 -9095
rect 620 -9163 632 -9129
rect 666 -9163 678 -9129
rect 620 -9197 678 -9163
rect 620 -9231 632 -9197
rect 666 -9231 678 -9197
rect 620 -9265 678 -9231
rect 620 -9299 632 -9265
rect 666 -9299 678 -9265
rect 620 -9333 678 -9299
rect 620 -9367 632 -9333
rect 666 -9367 678 -9333
rect 620 -9401 678 -9367
rect 620 -9435 632 -9401
rect 666 -9435 678 -9401
rect 620 -9469 678 -9435
rect 620 -9503 632 -9469
rect 666 -9503 678 -9469
rect 620 -9537 678 -9503
rect 620 -9571 632 -9537
rect 666 -9571 678 -9537
rect 620 -9600 678 -9571
rect 738 9571 796 9600
rect 738 9537 750 9571
rect 784 9537 796 9571
rect 738 9503 796 9537
rect 738 9469 750 9503
rect 784 9469 796 9503
rect 738 9435 796 9469
rect 738 9401 750 9435
rect 784 9401 796 9435
rect 738 9367 796 9401
rect 738 9333 750 9367
rect 784 9333 796 9367
rect 738 9299 796 9333
rect 738 9265 750 9299
rect 784 9265 796 9299
rect 738 9231 796 9265
rect 738 9197 750 9231
rect 784 9197 796 9231
rect 738 9163 796 9197
rect 738 9129 750 9163
rect 784 9129 796 9163
rect 738 9095 796 9129
rect 738 9061 750 9095
rect 784 9061 796 9095
rect 738 9027 796 9061
rect 738 8993 750 9027
rect 784 8993 796 9027
rect 738 8959 796 8993
rect 738 8925 750 8959
rect 784 8925 796 8959
rect 738 8891 796 8925
rect 738 8857 750 8891
rect 784 8857 796 8891
rect 738 8823 796 8857
rect 738 8789 750 8823
rect 784 8789 796 8823
rect 738 8755 796 8789
rect 738 8721 750 8755
rect 784 8721 796 8755
rect 738 8687 796 8721
rect 738 8653 750 8687
rect 784 8653 796 8687
rect 738 8619 796 8653
rect 738 8585 750 8619
rect 784 8585 796 8619
rect 738 8551 796 8585
rect 738 8517 750 8551
rect 784 8517 796 8551
rect 738 8483 796 8517
rect 738 8449 750 8483
rect 784 8449 796 8483
rect 738 8415 796 8449
rect 738 8381 750 8415
rect 784 8381 796 8415
rect 738 8347 796 8381
rect 738 8313 750 8347
rect 784 8313 796 8347
rect 738 8279 796 8313
rect 738 8245 750 8279
rect 784 8245 796 8279
rect 738 8211 796 8245
rect 738 8177 750 8211
rect 784 8177 796 8211
rect 738 8143 796 8177
rect 738 8109 750 8143
rect 784 8109 796 8143
rect 738 8075 796 8109
rect 738 8041 750 8075
rect 784 8041 796 8075
rect 738 8007 796 8041
rect 738 7973 750 8007
rect 784 7973 796 8007
rect 738 7939 796 7973
rect 738 7905 750 7939
rect 784 7905 796 7939
rect 738 7871 796 7905
rect 738 7837 750 7871
rect 784 7837 796 7871
rect 738 7803 796 7837
rect 738 7769 750 7803
rect 784 7769 796 7803
rect 738 7735 796 7769
rect 738 7701 750 7735
rect 784 7701 796 7735
rect 738 7667 796 7701
rect 738 7633 750 7667
rect 784 7633 796 7667
rect 738 7599 796 7633
rect 738 7565 750 7599
rect 784 7565 796 7599
rect 738 7531 796 7565
rect 738 7497 750 7531
rect 784 7497 796 7531
rect 738 7463 796 7497
rect 738 7429 750 7463
rect 784 7429 796 7463
rect 738 7395 796 7429
rect 738 7361 750 7395
rect 784 7361 796 7395
rect 738 7327 796 7361
rect 738 7293 750 7327
rect 784 7293 796 7327
rect 738 7259 796 7293
rect 738 7225 750 7259
rect 784 7225 796 7259
rect 738 7191 796 7225
rect 738 7157 750 7191
rect 784 7157 796 7191
rect 738 7123 796 7157
rect 738 7089 750 7123
rect 784 7089 796 7123
rect 738 7055 796 7089
rect 738 7021 750 7055
rect 784 7021 796 7055
rect 738 6987 796 7021
rect 738 6953 750 6987
rect 784 6953 796 6987
rect 738 6919 796 6953
rect 738 6885 750 6919
rect 784 6885 796 6919
rect 738 6851 796 6885
rect 738 6817 750 6851
rect 784 6817 796 6851
rect 738 6783 796 6817
rect 738 6749 750 6783
rect 784 6749 796 6783
rect 738 6715 796 6749
rect 738 6681 750 6715
rect 784 6681 796 6715
rect 738 6647 796 6681
rect 738 6613 750 6647
rect 784 6613 796 6647
rect 738 6579 796 6613
rect 738 6545 750 6579
rect 784 6545 796 6579
rect 738 6511 796 6545
rect 738 6477 750 6511
rect 784 6477 796 6511
rect 738 6443 796 6477
rect 738 6409 750 6443
rect 784 6409 796 6443
rect 738 6375 796 6409
rect 738 6341 750 6375
rect 784 6341 796 6375
rect 738 6307 796 6341
rect 738 6273 750 6307
rect 784 6273 796 6307
rect 738 6239 796 6273
rect 738 6205 750 6239
rect 784 6205 796 6239
rect 738 6171 796 6205
rect 738 6137 750 6171
rect 784 6137 796 6171
rect 738 6103 796 6137
rect 738 6069 750 6103
rect 784 6069 796 6103
rect 738 6035 796 6069
rect 738 6001 750 6035
rect 784 6001 796 6035
rect 738 5967 796 6001
rect 738 5933 750 5967
rect 784 5933 796 5967
rect 738 5899 796 5933
rect 738 5865 750 5899
rect 784 5865 796 5899
rect 738 5831 796 5865
rect 738 5797 750 5831
rect 784 5797 796 5831
rect 738 5763 796 5797
rect 738 5729 750 5763
rect 784 5729 796 5763
rect 738 5695 796 5729
rect 738 5661 750 5695
rect 784 5661 796 5695
rect 738 5627 796 5661
rect 738 5593 750 5627
rect 784 5593 796 5627
rect 738 5559 796 5593
rect 738 5525 750 5559
rect 784 5525 796 5559
rect 738 5491 796 5525
rect 738 5457 750 5491
rect 784 5457 796 5491
rect 738 5423 796 5457
rect 738 5389 750 5423
rect 784 5389 796 5423
rect 738 5355 796 5389
rect 738 5321 750 5355
rect 784 5321 796 5355
rect 738 5287 796 5321
rect 738 5253 750 5287
rect 784 5253 796 5287
rect 738 5219 796 5253
rect 738 5185 750 5219
rect 784 5185 796 5219
rect 738 5151 796 5185
rect 738 5117 750 5151
rect 784 5117 796 5151
rect 738 5083 796 5117
rect 738 5049 750 5083
rect 784 5049 796 5083
rect 738 5015 796 5049
rect 738 4981 750 5015
rect 784 4981 796 5015
rect 738 4947 796 4981
rect 738 4913 750 4947
rect 784 4913 796 4947
rect 738 4879 796 4913
rect 738 4845 750 4879
rect 784 4845 796 4879
rect 738 4811 796 4845
rect 738 4777 750 4811
rect 784 4777 796 4811
rect 738 4743 796 4777
rect 738 4709 750 4743
rect 784 4709 796 4743
rect 738 4675 796 4709
rect 738 4641 750 4675
rect 784 4641 796 4675
rect 738 4607 796 4641
rect 738 4573 750 4607
rect 784 4573 796 4607
rect 738 4539 796 4573
rect 738 4505 750 4539
rect 784 4505 796 4539
rect 738 4471 796 4505
rect 738 4437 750 4471
rect 784 4437 796 4471
rect 738 4403 796 4437
rect 738 4369 750 4403
rect 784 4369 796 4403
rect 738 4335 796 4369
rect 738 4301 750 4335
rect 784 4301 796 4335
rect 738 4267 796 4301
rect 738 4233 750 4267
rect 784 4233 796 4267
rect 738 4199 796 4233
rect 738 4165 750 4199
rect 784 4165 796 4199
rect 738 4131 796 4165
rect 738 4097 750 4131
rect 784 4097 796 4131
rect 738 4063 796 4097
rect 738 4029 750 4063
rect 784 4029 796 4063
rect 738 3995 796 4029
rect 738 3961 750 3995
rect 784 3961 796 3995
rect 738 3927 796 3961
rect 738 3893 750 3927
rect 784 3893 796 3927
rect 738 3859 796 3893
rect 738 3825 750 3859
rect 784 3825 796 3859
rect 738 3791 796 3825
rect 738 3757 750 3791
rect 784 3757 796 3791
rect 738 3723 796 3757
rect 738 3689 750 3723
rect 784 3689 796 3723
rect 738 3655 796 3689
rect 738 3621 750 3655
rect 784 3621 796 3655
rect 738 3587 796 3621
rect 738 3553 750 3587
rect 784 3553 796 3587
rect 738 3519 796 3553
rect 738 3485 750 3519
rect 784 3485 796 3519
rect 738 3451 796 3485
rect 738 3417 750 3451
rect 784 3417 796 3451
rect 738 3383 796 3417
rect 738 3349 750 3383
rect 784 3349 796 3383
rect 738 3315 796 3349
rect 738 3281 750 3315
rect 784 3281 796 3315
rect 738 3247 796 3281
rect 738 3213 750 3247
rect 784 3213 796 3247
rect 738 3179 796 3213
rect 738 3145 750 3179
rect 784 3145 796 3179
rect 738 3111 796 3145
rect 738 3077 750 3111
rect 784 3077 796 3111
rect 738 3043 796 3077
rect 738 3009 750 3043
rect 784 3009 796 3043
rect 738 2975 796 3009
rect 738 2941 750 2975
rect 784 2941 796 2975
rect 738 2907 796 2941
rect 738 2873 750 2907
rect 784 2873 796 2907
rect 738 2839 796 2873
rect 738 2805 750 2839
rect 784 2805 796 2839
rect 738 2771 796 2805
rect 738 2737 750 2771
rect 784 2737 796 2771
rect 738 2703 796 2737
rect 738 2669 750 2703
rect 784 2669 796 2703
rect 738 2635 796 2669
rect 738 2601 750 2635
rect 784 2601 796 2635
rect 738 2567 796 2601
rect 738 2533 750 2567
rect 784 2533 796 2567
rect 738 2499 796 2533
rect 738 2465 750 2499
rect 784 2465 796 2499
rect 738 2431 796 2465
rect 738 2397 750 2431
rect 784 2397 796 2431
rect 738 2363 796 2397
rect 738 2329 750 2363
rect 784 2329 796 2363
rect 738 2295 796 2329
rect 738 2261 750 2295
rect 784 2261 796 2295
rect 738 2227 796 2261
rect 738 2193 750 2227
rect 784 2193 796 2227
rect 738 2159 796 2193
rect 738 2125 750 2159
rect 784 2125 796 2159
rect 738 2091 796 2125
rect 738 2057 750 2091
rect 784 2057 796 2091
rect 738 2023 796 2057
rect 738 1989 750 2023
rect 784 1989 796 2023
rect 738 1955 796 1989
rect 738 1921 750 1955
rect 784 1921 796 1955
rect 738 1887 796 1921
rect 738 1853 750 1887
rect 784 1853 796 1887
rect 738 1819 796 1853
rect 738 1785 750 1819
rect 784 1785 796 1819
rect 738 1751 796 1785
rect 738 1717 750 1751
rect 784 1717 796 1751
rect 738 1683 796 1717
rect 738 1649 750 1683
rect 784 1649 796 1683
rect 738 1615 796 1649
rect 738 1581 750 1615
rect 784 1581 796 1615
rect 738 1547 796 1581
rect 738 1513 750 1547
rect 784 1513 796 1547
rect 738 1479 796 1513
rect 738 1445 750 1479
rect 784 1445 796 1479
rect 738 1411 796 1445
rect 738 1377 750 1411
rect 784 1377 796 1411
rect 738 1343 796 1377
rect 738 1309 750 1343
rect 784 1309 796 1343
rect 738 1275 796 1309
rect 738 1241 750 1275
rect 784 1241 796 1275
rect 738 1207 796 1241
rect 738 1173 750 1207
rect 784 1173 796 1207
rect 738 1139 796 1173
rect 738 1105 750 1139
rect 784 1105 796 1139
rect 738 1071 796 1105
rect 738 1037 750 1071
rect 784 1037 796 1071
rect 738 1003 796 1037
rect 738 969 750 1003
rect 784 969 796 1003
rect 738 935 796 969
rect 738 901 750 935
rect 784 901 796 935
rect 738 867 796 901
rect 738 833 750 867
rect 784 833 796 867
rect 738 799 796 833
rect 738 765 750 799
rect 784 765 796 799
rect 738 731 796 765
rect 738 697 750 731
rect 784 697 796 731
rect 738 663 796 697
rect 738 629 750 663
rect 784 629 796 663
rect 738 595 796 629
rect 738 561 750 595
rect 784 561 796 595
rect 738 527 796 561
rect 738 493 750 527
rect 784 493 796 527
rect 738 459 796 493
rect 738 425 750 459
rect 784 425 796 459
rect 738 391 796 425
rect 738 357 750 391
rect 784 357 796 391
rect 738 323 796 357
rect 738 289 750 323
rect 784 289 796 323
rect 738 255 796 289
rect 738 221 750 255
rect 784 221 796 255
rect 738 187 796 221
rect 738 153 750 187
rect 784 153 796 187
rect 738 119 796 153
rect 738 85 750 119
rect 784 85 796 119
rect 738 51 796 85
rect 738 17 750 51
rect 784 17 796 51
rect 738 -17 796 17
rect 738 -51 750 -17
rect 784 -51 796 -17
rect 738 -85 796 -51
rect 738 -119 750 -85
rect 784 -119 796 -85
rect 738 -153 796 -119
rect 738 -187 750 -153
rect 784 -187 796 -153
rect 738 -221 796 -187
rect 738 -255 750 -221
rect 784 -255 796 -221
rect 738 -289 796 -255
rect 738 -323 750 -289
rect 784 -323 796 -289
rect 738 -357 796 -323
rect 738 -391 750 -357
rect 784 -391 796 -357
rect 738 -425 796 -391
rect 738 -459 750 -425
rect 784 -459 796 -425
rect 738 -493 796 -459
rect 738 -527 750 -493
rect 784 -527 796 -493
rect 738 -561 796 -527
rect 738 -595 750 -561
rect 784 -595 796 -561
rect 738 -629 796 -595
rect 738 -663 750 -629
rect 784 -663 796 -629
rect 738 -697 796 -663
rect 738 -731 750 -697
rect 784 -731 796 -697
rect 738 -765 796 -731
rect 738 -799 750 -765
rect 784 -799 796 -765
rect 738 -833 796 -799
rect 738 -867 750 -833
rect 784 -867 796 -833
rect 738 -901 796 -867
rect 738 -935 750 -901
rect 784 -935 796 -901
rect 738 -969 796 -935
rect 738 -1003 750 -969
rect 784 -1003 796 -969
rect 738 -1037 796 -1003
rect 738 -1071 750 -1037
rect 784 -1071 796 -1037
rect 738 -1105 796 -1071
rect 738 -1139 750 -1105
rect 784 -1139 796 -1105
rect 738 -1173 796 -1139
rect 738 -1207 750 -1173
rect 784 -1207 796 -1173
rect 738 -1241 796 -1207
rect 738 -1275 750 -1241
rect 784 -1275 796 -1241
rect 738 -1309 796 -1275
rect 738 -1343 750 -1309
rect 784 -1343 796 -1309
rect 738 -1377 796 -1343
rect 738 -1411 750 -1377
rect 784 -1411 796 -1377
rect 738 -1445 796 -1411
rect 738 -1479 750 -1445
rect 784 -1479 796 -1445
rect 738 -1513 796 -1479
rect 738 -1547 750 -1513
rect 784 -1547 796 -1513
rect 738 -1581 796 -1547
rect 738 -1615 750 -1581
rect 784 -1615 796 -1581
rect 738 -1649 796 -1615
rect 738 -1683 750 -1649
rect 784 -1683 796 -1649
rect 738 -1717 796 -1683
rect 738 -1751 750 -1717
rect 784 -1751 796 -1717
rect 738 -1785 796 -1751
rect 738 -1819 750 -1785
rect 784 -1819 796 -1785
rect 738 -1853 796 -1819
rect 738 -1887 750 -1853
rect 784 -1887 796 -1853
rect 738 -1921 796 -1887
rect 738 -1955 750 -1921
rect 784 -1955 796 -1921
rect 738 -1989 796 -1955
rect 738 -2023 750 -1989
rect 784 -2023 796 -1989
rect 738 -2057 796 -2023
rect 738 -2091 750 -2057
rect 784 -2091 796 -2057
rect 738 -2125 796 -2091
rect 738 -2159 750 -2125
rect 784 -2159 796 -2125
rect 738 -2193 796 -2159
rect 738 -2227 750 -2193
rect 784 -2227 796 -2193
rect 738 -2261 796 -2227
rect 738 -2295 750 -2261
rect 784 -2295 796 -2261
rect 738 -2329 796 -2295
rect 738 -2363 750 -2329
rect 784 -2363 796 -2329
rect 738 -2397 796 -2363
rect 738 -2431 750 -2397
rect 784 -2431 796 -2397
rect 738 -2465 796 -2431
rect 738 -2499 750 -2465
rect 784 -2499 796 -2465
rect 738 -2533 796 -2499
rect 738 -2567 750 -2533
rect 784 -2567 796 -2533
rect 738 -2601 796 -2567
rect 738 -2635 750 -2601
rect 784 -2635 796 -2601
rect 738 -2669 796 -2635
rect 738 -2703 750 -2669
rect 784 -2703 796 -2669
rect 738 -2737 796 -2703
rect 738 -2771 750 -2737
rect 784 -2771 796 -2737
rect 738 -2805 796 -2771
rect 738 -2839 750 -2805
rect 784 -2839 796 -2805
rect 738 -2873 796 -2839
rect 738 -2907 750 -2873
rect 784 -2907 796 -2873
rect 738 -2941 796 -2907
rect 738 -2975 750 -2941
rect 784 -2975 796 -2941
rect 738 -3009 796 -2975
rect 738 -3043 750 -3009
rect 784 -3043 796 -3009
rect 738 -3077 796 -3043
rect 738 -3111 750 -3077
rect 784 -3111 796 -3077
rect 738 -3145 796 -3111
rect 738 -3179 750 -3145
rect 784 -3179 796 -3145
rect 738 -3213 796 -3179
rect 738 -3247 750 -3213
rect 784 -3247 796 -3213
rect 738 -3281 796 -3247
rect 738 -3315 750 -3281
rect 784 -3315 796 -3281
rect 738 -3349 796 -3315
rect 738 -3383 750 -3349
rect 784 -3383 796 -3349
rect 738 -3417 796 -3383
rect 738 -3451 750 -3417
rect 784 -3451 796 -3417
rect 738 -3485 796 -3451
rect 738 -3519 750 -3485
rect 784 -3519 796 -3485
rect 738 -3553 796 -3519
rect 738 -3587 750 -3553
rect 784 -3587 796 -3553
rect 738 -3621 796 -3587
rect 738 -3655 750 -3621
rect 784 -3655 796 -3621
rect 738 -3689 796 -3655
rect 738 -3723 750 -3689
rect 784 -3723 796 -3689
rect 738 -3757 796 -3723
rect 738 -3791 750 -3757
rect 784 -3791 796 -3757
rect 738 -3825 796 -3791
rect 738 -3859 750 -3825
rect 784 -3859 796 -3825
rect 738 -3893 796 -3859
rect 738 -3927 750 -3893
rect 784 -3927 796 -3893
rect 738 -3961 796 -3927
rect 738 -3995 750 -3961
rect 784 -3995 796 -3961
rect 738 -4029 796 -3995
rect 738 -4063 750 -4029
rect 784 -4063 796 -4029
rect 738 -4097 796 -4063
rect 738 -4131 750 -4097
rect 784 -4131 796 -4097
rect 738 -4165 796 -4131
rect 738 -4199 750 -4165
rect 784 -4199 796 -4165
rect 738 -4233 796 -4199
rect 738 -4267 750 -4233
rect 784 -4267 796 -4233
rect 738 -4301 796 -4267
rect 738 -4335 750 -4301
rect 784 -4335 796 -4301
rect 738 -4369 796 -4335
rect 738 -4403 750 -4369
rect 784 -4403 796 -4369
rect 738 -4437 796 -4403
rect 738 -4471 750 -4437
rect 784 -4471 796 -4437
rect 738 -4505 796 -4471
rect 738 -4539 750 -4505
rect 784 -4539 796 -4505
rect 738 -4573 796 -4539
rect 738 -4607 750 -4573
rect 784 -4607 796 -4573
rect 738 -4641 796 -4607
rect 738 -4675 750 -4641
rect 784 -4675 796 -4641
rect 738 -4709 796 -4675
rect 738 -4743 750 -4709
rect 784 -4743 796 -4709
rect 738 -4777 796 -4743
rect 738 -4811 750 -4777
rect 784 -4811 796 -4777
rect 738 -4845 796 -4811
rect 738 -4879 750 -4845
rect 784 -4879 796 -4845
rect 738 -4913 796 -4879
rect 738 -4947 750 -4913
rect 784 -4947 796 -4913
rect 738 -4981 796 -4947
rect 738 -5015 750 -4981
rect 784 -5015 796 -4981
rect 738 -5049 796 -5015
rect 738 -5083 750 -5049
rect 784 -5083 796 -5049
rect 738 -5117 796 -5083
rect 738 -5151 750 -5117
rect 784 -5151 796 -5117
rect 738 -5185 796 -5151
rect 738 -5219 750 -5185
rect 784 -5219 796 -5185
rect 738 -5253 796 -5219
rect 738 -5287 750 -5253
rect 784 -5287 796 -5253
rect 738 -5321 796 -5287
rect 738 -5355 750 -5321
rect 784 -5355 796 -5321
rect 738 -5389 796 -5355
rect 738 -5423 750 -5389
rect 784 -5423 796 -5389
rect 738 -5457 796 -5423
rect 738 -5491 750 -5457
rect 784 -5491 796 -5457
rect 738 -5525 796 -5491
rect 738 -5559 750 -5525
rect 784 -5559 796 -5525
rect 738 -5593 796 -5559
rect 738 -5627 750 -5593
rect 784 -5627 796 -5593
rect 738 -5661 796 -5627
rect 738 -5695 750 -5661
rect 784 -5695 796 -5661
rect 738 -5729 796 -5695
rect 738 -5763 750 -5729
rect 784 -5763 796 -5729
rect 738 -5797 796 -5763
rect 738 -5831 750 -5797
rect 784 -5831 796 -5797
rect 738 -5865 796 -5831
rect 738 -5899 750 -5865
rect 784 -5899 796 -5865
rect 738 -5933 796 -5899
rect 738 -5967 750 -5933
rect 784 -5967 796 -5933
rect 738 -6001 796 -5967
rect 738 -6035 750 -6001
rect 784 -6035 796 -6001
rect 738 -6069 796 -6035
rect 738 -6103 750 -6069
rect 784 -6103 796 -6069
rect 738 -6137 796 -6103
rect 738 -6171 750 -6137
rect 784 -6171 796 -6137
rect 738 -6205 796 -6171
rect 738 -6239 750 -6205
rect 784 -6239 796 -6205
rect 738 -6273 796 -6239
rect 738 -6307 750 -6273
rect 784 -6307 796 -6273
rect 738 -6341 796 -6307
rect 738 -6375 750 -6341
rect 784 -6375 796 -6341
rect 738 -6409 796 -6375
rect 738 -6443 750 -6409
rect 784 -6443 796 -6409
rect 738 -6477 796 -6443
rect 738 -6511 750 -6477
rect 784 -6511 796 -6477
rect 738 -6545 796 -6511
rect 738 -6579 750 -6545
rect 784 -6579 796 -6545
rect 738 -6613 796 -6579
rect 738 -6647 750 -6613
rect 784 -6647 796 -6613
rect 738 -6681 796 -6647
rect 738 -6715 750 -6681
rect 784 -6715 796 -6681
rect 738 -6749 796 -6715
rect 738 -6783 750 -6749
rect 784 -6783 796 -6749
rect 738 -6817 796 -6783
rect 738 -6851 750 -6817
rect 784 -6851 796 -6817
rect 738 -6885 796 -6851
rect 738 -6919 750 -6885
rect 784 -6919 796 -6885
rect 738 -6953 796 -6919
rect 738 -6987 750 -6953
rect 784 -6987 796 -6953
rect 738 -7021 796 -6987
rect 738 -7055 750 -7021
rect 784 -7055 796 -7021
rect 738 -7089 796 -7055
rect 738 -7123 750 -7089
rect 784 -7123 796 -7089
rect 738 -7157 796 -7123
rect 738 -7191 750 -7157
rect 784 -7191 796 -7157
rect 738 -7225 796 -7191
rect 738 -7259 750 -7225
rect 784 -7259 796 -7225
rect 738 -7293 796 -7259
rect 738 -7327 750 -7293
rect 784 -7327 796 -7293
rect 738 -7361 796 -7327
rect 738 -7395 750 -7361
rect 784 -7395 796 -7361
rect 738 -7429 796 -7395
rect 738 -7463 750 -7429
rect 784 -7463 796 -7429
rect 738 -7497 796 -7463
rect 738 -7531 750 -7497
rect 784 -7531 796 -7497
rect 738 -7565 796 -7531
rect 738 -7599 750 -7565
rect 784 -7599 796 -7565
rect 738 -7633 796 -7599
rect 738 -7667 750 -7633
rect 784 -7667 796 -7633
rect 738 -7701 796 -7667
rect 738 -7735 750 -7701
rect 784 -7735 796 -7701
rect 738 -7769 796 -7735
rect 738 -7803 750 -7769
rect 784 -7803 796 -7769
rect 738 -7837 796 -7803
rect 738 -7871 750 -7837
rect 784 -7871 796 -7837
rect 738 -7905 796 -7871
rect 738 -7939 750 -7905
rect 784 -7939 796 -7905
rect 738 -7973 796 -7939
rect 738 -8007 750 -7973
rect 784 -8007 796 -7973
rect 738 -8041 796 -8007
rect 738 -8075 750 -8041
rect 784 -8075 796 -8041
rect 738 -8109 796 -8075
rect 738 -8143 750 -8109
rect 784 -8143 796 -8109
rect 738 -8177 796 -8143
rect 738 -8211 750 -8177
rect 784 -8211 796 -8177
rect 738 -8245 796 -8211
rect 738 -8279 750 -8245
rect 784 -8279 796 -8245
rect 738 -8313 796 -8279
rect 738 -8347 750 -8313
rect 784 -8347 796 -8313
rect 738 -8381 796 -8347
rect 738 -8415 750 -8381
rect 784 -8415 796 -8381
rect 738 -8449 796 -8415
rect 738 -8483 750 -8449
rect 784 -8483 796 -8449
rect 738 -8517 796 -8483
rect 738 -8551 750 -8517
rect 784 -8551 796 -8517
rect 738 -8585 796 -8551
rect 738 -8619 750 -8585
rect 784 -8619 796 -8585
rect 738 -8653 796 -8619
rect 738 -8687 750 -8653
rect 784 -8687 796 -8653
rect 738 -8721 796 -8687
rect 738 -8755 750 -8721
rect 784 -8755 796 -8721
rect 738 -8789 796 -8755
rect 738 -8823 750 -8789
rect 784 -8823 796 -8789
rect 738 -8857 796 -8823
rect 738 -8891 750 -8857
rect 784 -8891 796 -8857
rect 738 -8925 796 -8891
rect 738 -8959 750 -8925
rect 784 -8959 796 -8925
rect 738 -8993 796 -8959
rect 738 -9027 750 -8993
rect 784 -9027 796 -8993
rect 738 -9061 796 -9027
rect 738 -9095 750 -9061
rect 784 -9095 796 -9061
rect 738 -9129 796 -9095
rect 738 -9163 750 -9129
rect 784 -9163 796 -9129
rect 738 -9197 796 -9163
rect 738 -9231 750 -9197
rect 784 -9231 796 -9197
rect 738 -9265 796 -9231
rect 738 -9299 750 -9265
rect 784 -9299 796 -9265
rect 738 -9333 796 -9299
rect 738 -9367 750 -9333
rect 784 -9367 796 -9333
rect 738 -9401 796 -9367
rect 738 -9435 750 -9401
rect 784 -9435 796 -9401
rect 738 -9469 796 -9435
rect 738 -9503 750 -9469
rect 784 -9503 796 -9469
rect 738 -9537 796 -9503
rect 738 -9571 750 -9537
rect 784 -9571 796 -9537
rect 738 -9600 796 -9571
rect 856 9571 914 9600
rect 856 9537 868 9571
rect 902 9537 914 9571
rect 856 9503 914 9537
rect 856 9469 868 9503
rect 902 9469 914 9503
rect 856 9435 914 9469
rect 856 9401 868 9435
rect 902 9401 914 9435
rect 856 9367 914 9401
rect 856 9333 868 9367
rect 902 9333 914 9367
rect 856 9299 914 9333
rect 856 9265 868 9299
rect 902 9265 914 9299
rect 856 9231 914 9265
rect 856 9197 868 9231
rect 902 9197 914 9231
rect 856 9163 914 9197
rect 856 9129 868 9163
rect 902 9129 914 9163
rect 856 9095 914 9129
rect 856 9061 868 9095
rect 902 9061 914 9095
rect 856 9027 914 9061
rect 856 8993 868 9027
rect 902 8993 914 9027
rect 856 8959 914 8993
rect 856 8925 868 8959
rect 902 8925 914 8959
rect 856 8891 914 8925
rect 856 8857 868 8891
rect 902 8857 914 8891
rect 856 8823 914 8857
rect 856 8789 868 8823
rect 902 8789 914 8823
rect 856 8755 914 8789
rect 856 8721 868 8755
rect 902 8721 914 8755
rect 856 8687 914 8721
rect 856 8653 868 8687
rect 902 8653 914 8687
rect 856 8619 914 8653
rect 856 8585 868 8619
rect 902 8585 914 8619
rect 856 8551 914 8585
rect 856 8517 868 8551
rect 902 8517 914 8551
rect 856 8483 914 8517
rect 856 8449 868 8483
rect 902 8449 914 8483
rect 856 8415 914 8449
rect 856 8381 868 8415
rect 902 8381 914 8415
rect 856 8347 914 8381
rect 856 8313 868 8347
rect 902 8313 914 8347
rect 856 8279 914 8313
rect 856 8245 868 8279
rect 902 8245 914 8279
rect 856 8211 914 8245
rect 856 8177 868 8211
rect 902 8177 914 8211
rect 856 8143 914 8177
rect 856 8109 868 8143
rect 902 8109 914 8143
rect 856 8075 914 8109
rect 856 8041 868 8075
rect 902 8041 914 8075
rect 856 8007 914 8041
rect 856 7973 868 8007
rect 902 7973 914 8007
rect 856 7939 914 7973
rect 856 7905 868 7939
rect 902 7905 914 7939
rect 856 7871 914 7905
rect 856 7837 868 7871
rect 902 7837 914 7871
rect 856 7803 914 7837
rect 856 7769 868 7803
rect 902 7769 914 7803
rect 856 7735 914 7769
rect 856 7701 868 7735
rect 902 7701 914 7735
rect 856 7667 914 7701
rect 856 7633 868 7667
rect 902 7633 914 7667
rect 856 7599 914 7633
rect 856 7565 868 7599
rect 902 7565 914 7599
rect 856 7531 914 7565
rect 856 7497 868 7531
rect 902 7497 914 7531
rect 856 7463 914 7497
rect 856 7429 868 7463
rect 902 7429 914 7463
rect 856 7395 914 7429
rect 856 7361 868 7395
rect 902 7361 914 7395
rect 856 7327 914 7361
rect 856 7293 868 7327
rect 902 7293 914 7327
rect 856 7259 914 7293
rect 856 7225 868 7259
rect 902 7225 914 7259
rect 856 7191 914 7225
rect 856 7157 868 7191
rect 902 7157 914 7191
rect 856 7123 914 7157
rect 856 7089 868 7123
rect 902 7089 914 7123
rect 856 7055 914 7089
rect 856 7021 868 7055
rect 902 7021 914 7055
rect 856 6987 914 7021
rect 856 6953 868 6987
rect 902 6953 914 6987
rect 856 6919 914 6953
rect 856 6885 868 6919
rect 902 6885 914 6919
rect 856 6851 914 6885
rect 856 6817 868 6851
rect 902 6817 914 6851
rect 856 6783 914 6817
rect 856 6749 868 6783
rect 902 6749 914 6783
rect 856 6715 914 6749
rect 856 6681 868 6715
rect 902 6681 914 6715
rect 856 6647 914 6681
rect 856 6613 868 6647
rect 902 6613 914 6647
rect 856 6579 914 6613
rect 856 6545 868 6579
rect 902 6545 914 6579
rect 856 6511 914 6545
rect 856 6477 868 6511
rect 902 6477 914 6511
rect 856 6443 914 6477
rect 856 6409 868 6443
rect 902 6409 914 6443
rect 856 6375 914 6409
rect 856 6341 868 6375
rect 902 6341 914 6375
rect 856 6307 914 6341
rect 856 6273 868 6307
rect 902 6273 914 6307
rect 856 6239 914 6273
rect 856 6205 868 6239
rect 902 6205 914 6239
rect 856 6171 914 6205
rect 856 6137 868 6171
rect 902 6137 914 6171
rect 856 6103 914 6137
rect 856 6069 868 6103
rect 902 6069 914 6103
rect 856 6035 914 6069
rect 856 6001 868 6035
rect 902 6001 914 6035
rect 856 5967 914 6001
rect 856 5933 868 5967
rect 902 5933 914 5967
rect 856 5899 914 5933
rect 856 5865 868 5899
rect 902 5865 914 5899
rect 856 5831 914 5865
rect 856 5797 868 5831
rect 902 5797 914 5831
rect 856 5763 914 5797
rect 856 5729 868 5763
rect 902 5729 914 5763
rect 856 5695 914 5729
rect 856 5661 868 5695
rect 902 5661 914 5695
rect 856 5627 914 5661
rect 856 5593 868 5627
rect 902 5593 914 5627
rect 856 5559 914 5593
rect 856 5525 868 5559
rect 902 5525 914 5559
rect 856 5491 914 5525
rect 856 5457 868 5491
rect 902 5457 914 5491
rect 856 5423 914 5457
rect 856 5389 868 5423
rect 902 5389 914 5423
rect 856 5355 914 5389
rect 856 5321 868 5355
rect 902 5321 914 5355
rect 856 5287 914 5321
rect 856 5253 868 5287
rect 902 5253 914 5287
rect 856 5219 914 5253
rect 856 5185 868 5219
rect 902 5185 914 5219
rect 856 5151 914 5185
rect 856 5117 868 5151
rect 902 5117 914 5151
rect 856 5083 914 5117
rect 856 5049 868 5083
rect 902 5049 914 5083
rect 856 5015 914 5049
rect 856 4981 868 5015
rect 902 4981 914 5015
rect 856 4947 914 4981
rect 856 4913 868 4947
rect 902 4913 914 4947
rect 856 4879 914 4913
rect 856 4845 868 4879
rect 902 4845 914 4879
rect 856 4811 914 4845
rect 856 4777 868 4811
rect 902 4777 914 4811
rect 856 4743 914 4777
rect 856 4709 868 4743
rect 902 4709 914 4743
rect 856 4675 914 4709
rect 856 4641 868 4675
rect 902 4641 914 4675
rect 856 4607 914 4641
rect 856 4573 868 4607
rect 902 4573 914 4607
rect 856 4539 914 4573
rect 856 4505 868 4539
rect 902 4505 914 4539
rect 856 4471 914 4505
rect 856 4437 868 4471
rect 902 4437 914 4471
rect 856 4403 914 4437
rect 856 4369 868 4403
rect 902 4369 914 4403
rect 856 4335 914 4369
rect 856 4301 868 4335
rect 902 4301 914 4335
rect 856 4267 914 4301
rect 856 4233 868 4267
rect 902 4233 914 4267
rect 856 4199 914 4233
rect 856 4165 868 4199
rect 902 4165 914 4199
rect 856 4131 914 4165
rect 856 4097 868 4131
rect 902 4097 914 4131
rect 856 4063 914 4097
rect 856 4029 868 4063
rect 902 4029 914 4063
rect 856 3995 914 4029
rect 856 3961 868 3995
rect 902 3961 914 3995
rect 856 3927 914 3961
rect 856 3893 868 3927
rect 902 3893 914 3927
rect 856 3859 914 3893
rect 856 3825 868 3859
rect 902 3825 914 3859
rect 856 3791 914 3825
rect 856 3757 868 3791
rect 902 3757 914 3791
rect 856 3723 914 3757
rect 856 3689 868 3723
rect 902 3689 914 3723
rect 856 3655 914 3689
rect 856 3621 868 3655
rect 902 3621 914 3655
rect 856 3587 914 3621
rect 856 3553 868 3587
rect 902 3553 914 3587
rect 856 3519 914 3553
rect 856 3485 868 3519
rect 902 3485 914 3519
rect 856 3451 914 3485
rect 856 3417 868 3451
rect 902 3417 914 3451
rect 856 3383 914 3417
rect 856 3349 868 3383
rect 902 3349 914 3383
rect 856 3315 914 3349
rect 856 3281 868 3315
rect 902 3281 914 3315
rect 856 3247 914 3281
rect 856 3213 868 3247
rect 902 3213 914 3247
rect 856 3179 914 3213
rect 856 3145 868 3179
rect 902 3145 914 3179
rect 856 3111 914 3145
rect 856 3077 868 3111
rect 902 3077 914 3111
rect 856 3043 914 3077
rect 856 3009 868 3043
rect 902 3009 914 3043
rect 856 2975 914 3009
rect 856 2941 868 2975
rect 902 2941 914 2975
rect 856 2907 914 2941
rect 856 2873 868 2907
rect 902 2873 914 2907
rect 856 2839 914 2873
rect 856 2805 868 2839
rect 902 2805 914 2839
rect 856 2771 914 2805
rect 856 2737 868 2771
rect 902 2737 914 2771
rect 856 2703 914 2737
rect 856 2669 868 2703
rect 902 2669 914 2703
rect 856 2635 914 2669
rect 856 2601 868 2635
rect 902 2601 914 2635
rect 856 2567 914 2601
rect 856 2533 868 2567
rect 902 2533 914 2567
rect 856 2499 914 2533
rect 856 2465 868 2499
rect 902 2465 914 2499
rect 856 2431 914 2465
rect 856 2397 868 2431
rect 902 2397 914 2431
rect 856 2363 914 2397
rect 856 2329 868 2363
rect 902 2329 914 2363
rect 856 2295 914 2329
rect 856 2261 868 2295
rect 902 2261 914 2295
rect 856 2227 914 2261
rect 856 2193 868 2227
rect 902 2193 914 2227
rect 856 2159 914 2193
rect 856 2125 868 2159
rect 902 2125 914 2159
rect 856 2091 914 2125
rect 856 2057 868 2091
rect 902 2057 914 2091
rect 856 2023 914 2057
rect 856 1989 868 2023
rect 902 1989 914 2023
rect 856 1955 914 1989
rect 856 1921 868 1955
rect 902 1921 914 1955
rect 856 1887 914 1921
rect 856 1853 868 1887
rect 902 1853 914 1887
rect 856 1819 914 1853
rect 856 1785 868 1819
rect 902 1785 914 1819
rect 856 1751 914 1785
rect 856 1717 868 1751
rect 902 1717 914 1751
rect 856 1683 914 1717
rect 856 1649 868 1683
rect 902 1649 914 1683
rect 856 1615 914 1649
rect 856 1581 868 1615
rect 902 1581 914 1615
rect 856 1547 914 1581
rect 856 1513 868 1547
rect 902 1513 914 1547
rect 856 1479 914 1513
rect 856 1445 868 1479
rect 902 1445 914 1479
rect 856 1411 914 1445
rect 856 1377 868 1411
rect 902 1377 914 1411
rect 856 1343 914 1377
rect 856 1309 868 1343
rect 902 1309 914 1343
rect 856 1275 914 1309
rect 856 1241 868 1275
rect 902 1241 914 1275
rect 856 1207 914 1241
rect 856 1173 868 1207
rect 902 1173 914 1207
rect 856 1139 914 1173
rect 856 1105 868 1139
rect 902 1105 914 1139
rect 856 1071 914 1105
rect 856 1037 868 1071
rect 902 1037 914 1071
rect 856 1003 914 1037
rect 856 969 868 1003
rect 902 969 914 1003
rect 856 935 914 969
rect 856 901 868 935
rect 902 901 914 935
rect 856 867 914 901
rect 856 833 868 867
rect 902 833 914 867
rect 856 799 914 833
rect 856 765 868 799
rect 902 765 914 799
rect 856 731 914 765
rect 856 697 868 731
rect 902 697 914 731
rect 856 663 914 697
rect 856 629 868 663
rect 902 629 914 663
rect 856 595 914 629
rect 856 561 868 595
rect 902 561 914 595
rect 856 527 914 561
rect 856 493 868 527
rect 902 493 914 527
rect 856 459 914 493
rect 856 425 868 459
rect 902 425 914 459
rect 856 391 914 425
rect 856 357 868 391
rect 902 357 914 391
rect 856 323 914 357
rect 856 289 868 323
rect 902 289 914 323
rect 856 255 914 289
rect 856 221 868 255
rect 902 221 914 255
rect 856 187 914 221
rect 856 153 868 187
rect 902 153 914 187
rect 856 119 914 153
rect 856 85 868 119
rect 902 85 914 119
rect 856 51 914 85
rect 856 17 868 51
rect 902 17 914 51
rect 856 -17 914 17
rect 856 -51 868 -17
rect 902 -51 914 -17
rect 856 -85 914 -51
rect 856 -119 868 -85
rect 902 -119 914 -85
rect 856 -153 914 -119
rect 856 -187 868 -153
rect 902 -187 914 -153
rect 856 -221 914 -187
rect 856 -255 868 -221
rect 902 -255 914 -221
rect 856 -289 914 -255
rect 856 -323 868 -289
rect 902 -323 914 -289
rect 856 -357 914 -323
rect 856 -391 868 -357
rect 902 -391 914 -357
rect 856 -425 914 -391
rect 856 -459 868 -425
rect 902 -459 914 -425
rect 856 -493 914 -459
rect 856 -527 868 -493
rect 902 -527 914 -493
rect 856 -561 914 -527
rect 856 -595 868 -561
rect 902 -595 914 -561
rect 856 -629 914 -595
rect 856 -663 868 -629
rect 902 -663 914 -629
rect 856 -697 914 -663
rect 856 -731 868 -697
rect 902 -731 914 -697
rect 856 -765 914 -731
rect 856 -799 868 -765
rect 902 -799 914 -765
rect 856 -833 914 -799
rect 856 -867 868 -833
rect 902 -867 914 -833
rect 856 -901 914 -867
rect 856 -935 868 -901
rect 902 -935 914 -901
rect 856 -969 914 -935
rect 856 -1003 868 -969
rect 902 -1003 914 -969
rect 856 -1037 914 -1003
rect 856 -1071 868 -1037
rect 902 -1071 914 -1037
rect 856 -1105 914 -1071
rect 856 -1139 868 -1105
rect 902 -1139 914 -1105
rect 856 -1173 914 -1139
rect 856 -1207 868 -1173
rect 902 -1207 914 -1173
rect 856 -1241 914 -1207
rect 856 -1275 868 -1241
rect 902 -1275 914 -1241
rect 856 -1309 914 -1275
rect 856 -1343 868 -1309
rect 902 -1343 914 -1309
rect 856 -1377 914 -1343
rect 856 -1411 868 -1377
rect 902 -1411 914 -1377
rect 856 -1445 914 -1411
rect 856 -1479 868 -1445
rect 902 -1479 914 -1445
rect 856 -1513 914 -1479
rect 856 -1547 868 -1513
rect 902 -1547 914 -1513
rect 856 -1581 914 -1547
rect 856 -1615 868 -1581
rect 902 -1615 914 -1581
rect 856 -1649 914 -1615
rect 856 -1683 868 -1649
rect 902 -1683 914 -1649
rect 856 -1717 914 -1683
rect 856 -1751 868 -1717
rect 902 -1751 914 -1717
rect 856 -1785 914 -1751
rect 856 -1819 868 -1785
rect 902 -1819 914 -1785
rect 856 -1853 914 -1819
rect 856 -1887 868 -1853
rect 902 -1887 914 -1853
rect 856 -1921 914 -1887
rect 856 -1955 868 -1921
rect 902 -1955 914 -1921
rect 856 -1989 914 -1955
rect 856 -2023 868 -1989
rect 902 -2023 914 -1989
rect 856 -2057 914 -2023
rect 856 -2091 868 -2057
rect 902 -2091 914 -2057
rect 856 -2125 914 -2091
rect 856 -2159 868 -2125
rect 902 -2159 914 -2125
rect 856 -2193 914 -2159
rect 856 -2227 868 -2193
rect 902 -2227 914 -2193
rect 856 -2261 914 -2227
rect 856 -2295 868 -2261
rect 902 -2295 914 -2261
rect 856 -2329 914 -2295
rect 856 -2363 868 -2329
rect 902 -2363 914 -2329
rect 856 -2397 914 -2363
rect 856 -2431 868 -2397
rect 902 -2431 914 -2397
rect 856 -2465 914 -2431
rect 856 -2499 868 -2465
rect 902 -2499 914 -2465
rect 856 -2533 914 -2499
rect 856 -2567 868 -2533
rect 902 -2567 914 -2533
rect 856 -2601 914 -2567
rect 856 -2635 868 -2601
rect 902 -2635 914 -2601
rect 856 -2669 914 -2635
rect 856 -2703 868 -2669
rect 902 -2703 914 -2669
rect 856 -2737 914 -2703
rect 856 -2771 868 -2737
rect 902 -2771 914 -2737
rect 856 -2805 914 -2771
rect 856 -2839 868 -2805
rect 902 -2839 914 -2805
rect 856 -2873 914 -2839
rect 856 -2907 868 -2873
rect 902 -2907 914 -2873
rect 856 -2941 914 -2907
rect 856 -2975 868 -2941
rect 902 -2975 914 -2941
rect 856 -3009 914 -2975
rect 856 -3043 868 -3009
rect 902 -3043 914 -3009
rect 856 -3077 914 -3043
rect 856 -3111 868 -3077
rect 902 -3111 914 -3077
rect 856 -3145 914 -3111
rect 856 -3179 868 -3145
rect 902 -3179 914 -3145
rect 856 -3213 914 -3179
rect 856 -3247 868 -3213
rect 902 -3247 914 -3213
rect 856 -3281 914 -3247
rect 856 -3315 868 -3281
rect 902 -3315 914 -3281
rect 856 -3349 914 -3315
rect 856 -3383 868 -3349
rect 902 -3383 914 -3349
rect 856 -3417 914 -3383
rect 856 -3451 868 -3417
rect 902 -3451 914 -3417
rect 856 -3485 914 -3451
rect 856 -3519 868 -3485
rect 902 -3519 914 -3485
rect 856 -3553 914 -3519
rect 856 -3587 868 -3553
rect 902 -3587 914 -3553
rect 856 -3621 914 -3587
rect 856 -3655 868 -3621
rect 902 -3655 914 -3621
rect 856 -3689 914 -3655
rect 856 -3723 868 -3689
rect 902 -3723 914 -3689
rect 856 -3757 914 -3723
rect 856 -3791 868 -3757
rect 902 -3791 914 -3757
rect 856 -3825 914 -3791
rect 856 -3859 868 -3825
rect 902 -3859 914 -3825
rect 856 -3893 914 -3859
rect 856 -3927 868 -3893
rect 902 -3927 914 -3893
rect 856 -3961 914 -3927
rect 856 -3995 868 -3961
rect 902 -3995 914 -3961
rect 856 -4029 914 -3995
rect 856 -4063 868 -4029
rect 902 -4063 914 -4029
rect 856 -4097 914 -4063
rect 856 -4131 868 -4097
rect 902 -4131 914 -4097
rect 856 -4165 914 -4131
rect 856 -4199 868 -4165
rect 902 -4199 914 -4165
rect 856 -4233 914 -4199
rect 856 -4267 868 -4233
rect 902 -4267 914 -4233
rect 856 -4301 914 -4267
rect 856 -4335 868 -4301
rect 902 -4335 914 -4301
rect 856 -4369 914 -4335
rect 856 -4403 868 -4369
rect 902 -4403 914 -4369
rect 856 -4437 914 -4403
rect 856 -4471 868 -4437
rect 902 -4471 914 -4437
rect 856 -4505 914 -4471
rect 856 -4539 868 -4505
rect 902 -4539 914 -4505
rect 856 -4573 914 -4539
rect 856 -4607 868 -4573
rect 902 -4607 914 -4573
rect 856 -4641 914 -4607
rect 856 -4675 868 -4641
rect 902 -4675 914 -4641
rect 856 -4709 914 -4675
rect 856 -4743 868 -4709
rect 902 -4743 914 -4709
rect 856 -4777 914 -4743
rect 856 -4811 868 -4777
rect 902 -4811 914 -4777
rect 856 -4845 914 -4811
rect 856 -4879 868 -4845
rect 902 -4879 914 -4845
rect 856 -4913 914 -4879
rect 856 -4947 868 -4913
rect 902 -4947 914 -4913
rect 856 -4981 914 -4947
rect 856 -5015 868 -4981
rect 902 -5015 914 -4981
rect 856 -5049 914 -5015
rect 856 -5083 868 -5049
rect 902 -5083 914 -5049
rect 856 -5117 914 -5083
rect 856 -5151 868 -5117
rect 902 -5151 914 -5117
rect 856 -5185 914 -5151
rect 856 -5219 868 -5185
rect 902 -5219 914 -5185
rect 856 -5253 914 -5219
rect 856 -5287 868 -5253
rect 902 -5287 914 -5253
rect 856 -5321 914 -5287
rect 856 -5355 868 -5321
rect 902 -5355 914 -5321
rect 856 -5389 914 -5355
rect 856 -5423 868 -5389
rect 902 -5423 914 -5389
rect 856 -5457 914 -5423
rect 856 -5491 868 -5457
rect 902 -5491 914 -5457
rect 856 -5525 914 -5491
rect 856 -5559 868 -5525
rect 902 -5559 914 -5525
rect 856 -5593 914 -5559
rect 856 -5627 868 -5593
rect 902 -5627 914 -5593
rect 856 -5661 914 -5627
rect 856 -5695 868 -5661
rect 902 -5695 914 -5661
rect 856 -5729 914 -5695
rect 856 -5763 868 -5729
rect 902 -5763 914 -5729
rect 856 -5797 914 -5763
rect 856 -5831 868 -5797
rect 902 -5831 914 -5797
rect 856 -5865 914 -5831
rect 856 -5899 868 -5865
rect 902 -5899 914 -5865
rect 856 -5933 914 -5899
rect 856 -5967 868 -5933
rect 902 -5967 914 -5933
rect 856 -6001 914 -5967
rect 856 -6035 868 -6001
rect 902 -6035 914 -6001
rect 856 -6069 914 -6035
rect 856 -6103 868 -6069
rect 902 -6103 914 -6069
rect 856 -6137 914 -6103
rect 856 -6171 868 -6137
rect 902 -6171 914 -6137
rect 856 -6205 914 -6171
rect 856 -6239 868 -6205
rect 902 -6239 914 -6205
rect 856 -6273 914 -6239
rect 856 -6307 868 -6273
rect 902 -6307 914 -6273
rect 856 -6341 914 -6307
rect 856 -6375 868 -6341
rect 902 -6375 914 -6341
rect 856 -6409 914 -6375
rect 856 -6443 868 -6409
rect 902 -6443 914 -6409
rect 856 -6477 914 -6443
rect 856 -6511 868 -6477
rect 902 -6511 914 -6477
rect 856 -6545 914 -6511
rect 856 -6579 868 -6545
rect 902 -6579 914 -6545
rect 856 -6613 914 -6579
rect 856 -6647 868 -6613
rect 902 -6647 914 -6613
rect 856 -6681 914 -6647
rect 856 -6715 868 -6681
rect 902 -6715 914 -6681
rect 856 -6749 914 -6715
rect 856 -6783 868 -6749
rect 902 -6783 914 -6749
rect 856 -6817 914 -6783
rect 856 -6851 868 -6817
rect 902 -6851 914 -6817
rect 856 -6885 914 -6851
rect 856 -6919 868 -6885
rect 902 -6919 914 -6885
rect 856 -6953 914 -6919
rect 856 -6987 868 -6953
rect 902 -6987 914 -6953
rect 856 -7021 914 -6987
rect 856 -7055 868 -7021
rect 902 -7055 914 -7021
rect 856 -7089 914 -7055
rect 856 -7123 868 -7089
rect 902 -7123 914 -7089
rect 856 -7157 914 -7123
rect 856 -7191 868 -7157
rect 902 -7191 914 -7157
rect 856 -7225 914 -7191
rect 856 -7259 868 -7225
rect 902 -7259 914 -7225
rect 856 -7293 914 -7259
rect 856 -7327 868 -7293
rect 902 -7327 914 -7293
rect 856 -7361 914 -7327
rect 856 -7395 868 -7361
rect 902 -7395 914 -7361
rect 856 -7429 914 -7395
rect 856 -7463 868 -7429
rect 902 -7463 914 -7429
rect 856 -7497 914 -7463
rect 856 -7531 868 -7497
rect 902 -7531 914 -7497
rect 856 -7565 914 -7531
rect 856 -7599 868 -7565
rect 902 -7599 914 -7565
rect 856 -7633 914 -7599
rect 856 -7667 868 -7633
rect 902 -7667 914 -7633
rect 856 -7701 914 -7667
rect 856 -7735 868 -7701
rect 902 -7735 914 -7701
rect 856 -7769 914 -7735
rect 856 -7803 868 -7769
rect 902 -7803 914 -7769
rect 856 -7837 914 -7803
rect 856 -7871 868 -7837
rect 902 -7871 914 -7837
rect 856 -7905 914 -7871
rect 856 -7939 868 -7905
rect 902 -7939 914 -7905
rect 856 -7973 914 -7939
rect 856 -8007 868 -7973
rect 902 -8007 914 -7973
rect 856 -8041 914 -8007
rect 856 -8075 868 -8041
rect 902 -8075 914 -8041
rect 856 -8109 914 -8075
rect 856 -8143 868 -8109
rect 902 -8143 914 -8109
rect 856 -8177 914 -8143
rect 856 -8211 868 -8177
rect 902 -8211 914 -8177
rect 856 -8245 914 -8211
rect 856 -8279 868 -8245
rect 902 -8279 914 -8245
rect 856 -8313 914 -8279
rect 856 -8347 868 -8313
rect 902 -8347 914 -8313
rect 856 -8381 914 -8347
rect 856 -8415 868 -8381
rect 902 -8415 914 -8381
rect 856 -8449 914 -8415
rect 856 -8483 868 -8449
rect 902 -8483 914 -8449
rect 856 -8517 914 -8483
rect 856 -8551 868 -8517
rect 902 -8551 914 -8517
rect 856 -8585 914 -8551
rect 856 -8619 868 -8585
rect 902 -8619 914 -8585
rect 856 -8653 914 -8619
rect 856 -8687 868 -8653
rect 902 -8687 914 -8653
rect 856 -8721 914 -8687
rect 856 -8755 868 -8721
rect 902 -8755 914 -8721
rect 856 -8789 914 -8755
rect 856 -8823 868 -8789
rect 902 -8823 914 -8789
rect 856 -8857 914 -8823
rect 856 -8891 868 -8857
rect 902 -8891 914 -8857
rect 856 -8925 914 -8891
rect 856 -8959 868 -8925
rect 902 -8959 914 -8925
rect 856 -8993 914 -8959
rect 856 -9027 868 -8993
rect 902 -9027 914 -8993
rect 856 -9061 914 -9027
rect 856 -9095 868 -9061
rect 902 -9095 914 -9061
rect 856 -9129 914 -9095
rect 856 -9163 868 -9129
rect 902 -9163 914 -9129
rect 856 -9197 914 -9163
rect 856 -9231 868 -9197
rect 902 -9231 914 -9197
rect 856 -9265 914 -9231
rect 856 -9299 868 -9265
rect 902 -9299 914 -9265
rect 856 -9333 914 -9299
rect 856 -9367 868 -9333
rect 902 -9367 914 -9333
rect 856 -9401 914 -9367
rect 856 -9435 868 -9401
rect 902 -9435 914 -9401
rect 856 -9469 914 -9435
rect 856 -9503 868 -9469
rect 902 -9503 914 -9469
rect 856 -9537 914 -9503
rect 856 -9571 868 -9537
rect 902 -9571 914 -9537
rect 856 -9600 914 -9571
rect 974 9571 1032 9600
rect 974 9537 986 9571
rect 1020 9537 1032 9571
rect 974 9503 1032 9537
rect 974 9469 986 9503
rect 1020 9469 1032 9503
rect 974 9435 1032 9469
rect 974 9401 986 9435
rect 1020 9401 1032 9435
rect 974 9367 1032 9401
rect 974 9333 986 9367
rect 1020 9333 1032 9367
rect 974 9299 1032 9333
rect 974 9265 986 9299
rect 1020 9265 1032 9299
rect 974 9231 1032 9265
rect 974 9197 986 9231
rect 1020 9197 1032 9231
rect 974 9163 1032 9197
rect 974 9129 986 9163
rect 1020 9129 1032 9163
rect 974 9095 1032 9129
rect 974 9061 986 9095
rect 1020 9061 1032 9095
rect 974 9027 1032 9061
rect 974 8993 986 9027
rect 1020 8993 1032 9027
rect 974 8959 1032 8993
rect 974 8925 986 8959
rect 1020 8925 1032 8959
rect 974 8891 1032 8925
rect 974 8857 986 8891
rect 1020 8857 1032 8891
rect 974 8823 1032 8857
rect 974 8789 986 8823
rect 1020 8789 1032 8823
rect 974 8755 1032 8789
rect 974 8721 986 8755
rect 1020 8721 1032 8755
rect 974 8687 1032 8721
rect 974 8653 986 8687
rect 1020 8653 1032 8687
rect 974 8619 1032 8653
rect 974 8585 986 8619
rect 1020 8585 1032 8619
rect 974 8551 1032 8585
rect 974 8517 986 8551
rect 1020 8517 1032 8551
rect 974 8483 1032 8517
rect 974 8449 986 8483
rect 1020 8449 1032 8483
rect 974 8415 1032 8449
rect 974 8381 986 8415
rect 1020 8381 1032 8415
rect 974 8347 1032 8381
rect 974 8313 986 8347
rect 1020 8313 1032 8347
rect 974 8279 1032 8313
rect 974 8245 986 8279
rect 1020 8245 1032 8279
rect 974 8211 1032 8245
rect 974 8177 986 8211
rect 1020 8177 1032 8211
rect 974 8143 1032 8177
rect 974 8109 986 8143
rect 1020 8109 1032 8143
rect 974 8075 1032 8109
rect 974 8041 986 8075
rect 1020 8041 1032 8075
rect 974 8007 1032 8041
rect 974 7973 986 8007
rect 1020 7973 1032 8007
rect 974 7939 1032 7973
rect 974 7905 986 7939
rect 1020 7905 1032 7939
rect 974 7871 1032 7905
rect 974 7837 986 7871
rect 1020 7837 1032 7871
rect 974 7803 1032 7837
rect 974 7769 986 7803
rect 1020 7769 1032 7803
rect 974 7735 1032 7769
rect 974 7701 986 7735
rect 1020 7701 1032 7735
rect 974 7667 1032 7701
rect 974 7633 986 7667
rect 1020 7633 1032 7667
rect 974 7599 1032 7633
rect 974 7565 986 7599
rect 1020 7565 1032 7599
rect 974 7531 1032 7565
rect 974 7497 986 7531
rect 1020 7497 1032 7531
rect 974 7463 1032 7497
rect 974 7429 986 7463
rect 1020 7429 1032 7463
rect 974 7395 1032 7429
rect 974 7361 986 7395
rect 1020 7361 1032 7395
rect 974 7327 1032 7361
rect 974 7293 986 7327
rect 1020 7293 1032 7327
rect 974 7259 1032 7293
rect 974 7225 986 7259
rect 1020 7225 1032 7259
rect 974 7191 1032 7225
rect 974 7157 986 7191
rect 1020 7157 1032 7191
rect 974 7123 1032 7157
rect 974 7089 986 7123
rect 1020 7089 1032 7123
rect 974 7055 1032 7089
rect 974 7021 986 7055
rect 1020 7021 1032 7055
rect 974 6987 1032 7021
rect 974 6953 986 6987
rect 1020 6953 1032 6987
rect 974 6919 1032 6953
rect 974 6885 986 6919
rect 1020 6885 1032 6919
rect 974 6851 1032 6885
rect 974 6817 986 6851
rect 1020 6817 1032 6851
rect 974 6783 1032 6817
rect 974 6749 986 6783
rect 1020 6749 1032 6783
rect 974 6715 1032 6749
rect 974 6681 986 6715
rect 1020 6681 1032 6715
rect 974 6647 1032 6681
rect 974 6613 986 6647
rect 1020 6613 1032 6647
rect 974 6579 1032 6613
rect 974 6545 986 6579
rect 1020 6545 1032 6579
rect 974 6511 1032 6545
rect 974 6477 986 6511
rect 1020 6477 1032 6511
rect 974 6443 1032 6477
rect 974 6409 986 6443
rect 1020 6409 1032 6443
rect 974 6375 1032 6409
rect 974 6341 986 6375
rect 1020 6341 1032 6375
rect 974 6307 1032 6341
rect 974 6273 986 6307
rect 1020 6273 1032 6307
rect 974 6239 1032 6273
rect 974 6205 986 6239
rect 1020 6205 1032 6239
rect 974 6171 1032 6205
rect 974 6137 986 6171
rect 1020 6137 1032 6171
rect 974 6103 1032 6137
rect 974 6069 986 6103
rect 1020 6069 1032 6103
rect 974 6035 1032 6069
rect 974 6001 986 6035
rect 1020 6001 1032 6035
rect 974 5967 1032 6001
rect 974 5933 986 5967
rect 1020 5933 1032 5967
rect 974 5899 1032 5933
rect 974 5865 986 5899
rect 1020 5865 1032 5899
rect 974 5831 1032 5865
rect 974 5797 986 5831
rect 1020 5797 1032 5831
rect 974 5763 1032 5797
rect 974 5729 986 5763
rect 1020 5729 1032 5763
rect 974 5695 1032 5729
rect 974 5661 986 5695
rect 1020 5661 1032 5695
rect 974 5627 1032 5661
rect 974 5593 986 5627
rect 1020 5593 1032 5627
rect 974 5559 1032 5593
rect 974 5525 986 5559
rect 1020 5525 1032 5559
rect 974 5491 1032 5525
rect 974 5457 986 5491
rect 1020 5457 1032 5491
rect 974 5423 1032 5457
rect 974 5389 986 5423
rect 1020 5389 1032 5423
rect 974 5355 1032 5389
rect 974 5321 986 5355
rect 1020 5321 1032 5355
rect 974 5287 1032 5321
rect 974 5253 986 5287
rect 1020 5253 1032 5287
rect 974 5219 1032 5253
rect 974 5185 986 5219
rect 1020 5185 1032 5219
rect 974 5151 1032 5185
rect 974 5117 986 5151
rect 1020 5117 1032 5151
rect 974 5083 1032 5117
rect 974 5049 986 5083
rect 1020 5049 1032 5083
rect 974 5015 1032 5049
rect 974 4981 986 5015
rect 1020 4981 1032 5015
rect 974 4947 1032 4981
rect 974 4913 986 4947
rect 1020 4913 1032 4947
rect 974 4879 1032 4913
rect 974 4845 986 4879
rect 1020 4845 1032 4879
rect 974 4811 1032 4845
rect 974 4777 986 4811
rect 1020 4777 1032 4811
rect 974 4743 1032 4777
rect 974 4709 986 4743
rect 1020 4709 1032 4743
rect 974 4675 1032 4709
rect 974 4641 986 4675
rect 1020 4641 1032 4675
rect 974 4607 1032 4641
rect 974 4573 986 4607
rect 1020 4573 1032 4607
rect 974 4539 1032 4573
rect 974 4505 986 4539
rect 1020 4505 1032 4539
rect 974 4471 1032 4505
rect 974 4437 986 4471
rect 1020 4437 1032 4471
rect 974 4403 1032 4437
rect 974 4369 986 4403
rect 1020 4369 1032 4403
rect 974 4335 1032 4369
rect 974 4301 986 4335
rect 1020 4301 1032 4335
rect 974 4267 1032 4301
rect 974 4233 986 4267
rect 1020 4233 1032 4267
rect 974 4199 1032 4233
rect 974 4165 986 4199
rect 1020 4165 1032 4199
rect 974 4131 1032 4165
rect 974 4097 986 4131
rect 1020 4097 1032 4131
rect 974 4063 1032 4097
rect 974 4029 986 4063
rect 1020 4029 1032 4063
rect 974 3995 1032 4029
rect 974 3961 986 3995
rect 1020 3961 1032 3995
rect 974 3927 1032 3961
rect 974 3893 986 3927
rect 1020 3893 1032 3927
rect 974 3859 1032 3893
rect 974 3825 986 3859
rect 1020 3825 1032 3859
rect 974 3791 1032 3825
rect 974 3757 986 3791
rect 1020 3757 1032 3791
rect 974 3723 1032 3757
rect 974 3689 986 3723
rect 1020 3689 1032 3723
rect 974 3655 1032 3689
rect 974 3621 986 3655
rect 1020 3621 1032 3655
rect 974 3587 1032 3621
rect 974 3553 986 3587
rect 1020 3553 1032 3587
rect 974 3519 1032 3553
rect 974 3485 986 3519
rect 1020 3485 1032 3519
rect 974 3451 1032 3485
rect 974 3417 986 3451
rect 1020 3417 1032 3451
rect 974 3383 1032 3417
rect 974 3349 986 3383
rect 1020 3349 1032 3383
rect 974 3315 1032 3349
rect 974 3281 986 3315
rect 1020 3281 1032 3315
rect 974 3247 1032 3281
rect 974 3213 986 3247
rect 1020 3213 1032 3247
rect 974 3179 1032 3213
rect 974 3145 986 3179
rect 1020 3145 1032 3179
rect 974 3111 1032 3145
rect 974 3077 986 3111
rect 1020 3077 1032 3111
rect 974 3043 1032 3077
rect 974 3009 986 3043
rect 1020 3009 1032 3043
rect 974 2975 1032 3009
rect 974 2941 986 2975
rect 1020 2941 1032 2975
rect 974 2907 1032 2941
rect 974 2873 986 2907
rect 1020 2873 1032 2907
rect 974 2839 1032 2873
rect 974 2805 986 2839
rect 1020 2805 1032 2839
rect 974 2771 1032 2805
rect 974 2737 986 2771
rect 1020 2737 1032 2771
rect 974 2703 1032 2737
rect 974 2669 986 2703
rect 1020 2669 1032 2703
rect 974 2635 1032 2669
rect 974 2601 986 2635
rect 1020 2601 1032 2635
rect 974 2567 1032 2601
rect 974 2533 986 2567
rect 1020 2533 1032 2567
rect 974 2499 1032 2533
rect 974 2465 986 2499
rect 1020 2465 1032 2499
rect 974 2431 1032 2465
rect 974 2397 986 2431
rect 1020 2397 1032 2431
rect 974 2363 1032 2397
rect 974 2329 986 2363
rect 1020 2329 1032 2363
rect 974 2295 1032 2329
rect 974 2261 986 2295
rect 1020 2261 1032 2295
rect 974 2227 1032 2261
rect 974 2193 986 2227
rect 1020 2193 1032 2227
rect 974 2159 1032 2193
rect 974 2125 986 2159
rect 1020 2125 1032 2159
rect 974 2091 1032 2125
rect 974 2057 986 2091
rect 1020 2057 1032 2091
rect 974 2023 1032 2057
rect 974 1989 986 2023
rect 1020 1989 1032 2023
rect 974 1955 1032 1989
rect 974 1921 986 1955
rect 1020 1921 1032 1955
rect 974 1887 1032 1921
rect 974 1853 986 1887
rect 1020 1853 1032 1887
rect 974 1819 1032 1853
rect 974 1785 986 1819
rect 1020 1785 1032 1819
rect 974 1751 1032 1785
rect 974 1717 986 1751
rect 1020 1717 1032 1751
rect 974 1683 1032 1717
rect 974 1649 986 1683
rect 1020 1649 1032 1683
rect 974 1615 1032 1649
rect 974 1581 986 1615
rect 1020 1581 1032 1615
rect 974 1547 1032 1581
rect 974 1513 986 1547
rect 1020 1513 1032 1547
rect 974 1479 1032 1513
rect 974 1445 986 1479
rect 1020 1445 1032 1479
rect 974 1411 1032 1445
rect 974 1377 986 1411
rect 1020 1377 1032 1411
rect 974 1343 1032 1377
rect 974 1309 986 1343
rect 1020 1309 1032 1343
rect 974 1275 1032 1309
rect 974 1241 986 1275
rect 1020 1241 1032 1275
rect 974 1207 1032 1241
rect 974 1173 986 1207
rect 1020 1173 1032 1207
rect 974 1139 1032 1173
rect 974 1105 986 1139
rect 1020 1105 1032 1139
rect 974 1071 1032 1105
rect 974 1037 986 1071
rect 1020 1037 1032 1071
rect 974 1003 1032 1037
rect 974 969 986 1003
rect 1020 969 1032 1003
rect 974 935 1032 969
rect 974 901 986 935
rect 1020 901 1032 935
rect 974 867 1032 901
rect 974 833 986 867
rect 1020 833 1032 867
rect 974 799 1032 833
rect 974 765 986 799
rect 1020 765 1032 799
rect 974 731 1032 765
rect 974 697 986 731
rect 1020 697 1032 731
rect 974 663 1032 697
rect 974 629 986 663
rect 1020 629 1032 663
rect 974 595 1032 629
rect 974 561 986 595
rect 1020 561 1032 595
rect 974 527 1032 561
rect 974 493 986 527
rect 1020 493 1032 527
rect 974 459 1032 493
rect 974 425 986 459
rect 1020 425 1032 459
rect 974 391 1032 425
rect 974 357 986 391
rect 1020 357 1032 391
rect 974 323 1032 357
rect 974 289 986 323
rect 1020 289 1032 323
rect 974 255 1032 289
rect 974 221 986 255
rect 1020 221 1032 255
rect 974 187 1032 221
rect 974 153 986 187
rect 1020 153 1032 187
rect 974 119 1032 153
rect 974 85 986 119
rect 1020 85 1032 119
rect 974 51 1032 85
rect 974 17 986 51
rect 1020 17 1032 51
rect 974 -17 1032 17
rect 974 -51 986 -17
rect 1020 -51 1032 -17
rect 974 -85 1032 -51
rect 974 -119 986 -85
rect 1020 -119 1032 -85
rect 974 -153 1032 -119
rect 974 -187 986 -153
rect 1020 -187 1032 -153
rect 974 -221 1032 -187
rect 974 -255 986 -221
rect 1020 -255 1032 -221
rect 974 -289 1032 -255
rect 974 -323 986 -289
rect 1020 -323 1032 -289
rect 974 -357 1032 -323
rect 974 -391 986 -357
rect 1020 -391 1032 -357
rect 974 -425 1032 -391
rect 974 -459 986 -425
rect 1020 -459 1032 -425
rect 974 -493 1032 -459
rect 974 -527 986 -493
rect 1020 -527 1032 -493
rect 974 -561 1032 -527
rect 974 -595 986 -561
rect 1020 -595 1032 -561
rect 974 -629 1032 -595
rect 974 -663 986 -629
rect 1020 -663 1032 -629
rect 974 -697 1032 -663
rect 974 -731 986 -697
rect 1020 -731 1032 -697
rect 974 -765 1032 -731
rect 974 -799 986 -765
rect 1020 -799 1032 -765
rect 974 -833 1032 -799
rect 974 -867 986 -833
rect 1020 -867 1032 -833
rect 974 -901 1032 -867
rect 974 -935 986 -901
rect 1020 -935 1032 -901
rect 974 -969 1032 -935
rect 974 -1003 986 -969
rect 1020 -1003 1032 -969
rect 974 -1037 1032 -1003
rect 974 -1071 986 -1037
rect 1020 -1071 1032 -1037
rect 974 -1105 1032 -1071
rect 974 -1139 986 -1105
rect 1020 -1139 1032 -1105
rect 974 -1173 1032 -1139
rect 974 -1207 986 -1173
rect 1020 -1207 1032 -1173
rect 974 -1241 1032 -1207
rect 974 -1275 986 -1241
rect 1020 -1275 1032 -1241
rect 974 -1309 1032 -1275
rect 974 -1343 986 -1309
rect 1020 -1343 1032 -1309
rect 974 -1377 1032 -1343
rect 974 -1411 986 -1377
rect 1020 -1411 1032 -1377
rect 974 -1445 1032 -1411
rect 974 -1479 986 -1445
rect 1020 -1479 1032 -1445
rect 974 -1513 1032 -1479
rect 974 -1547 986 -1513
rect 1020 -1547 1032 -1513
rect 974 -1581 1032 -1547
rect 974 -1615 986 -1581
rect 1020 -1615 1032 -1581
rect 974 -1649 1032 -1615
rect 974 -1683 986 -1649
rect 1020 -1683 1032 -1649
rect 974 -1717 1032 -1683
rect 974 -1751 986 -1717
rect 1020 -1751 1032 -1717
rect 974 -1785 1032 -1751
rect 974 -1819 986 -1785
rect 1020 -1819 1032 -1785
rect 974 -1853 1032 -1819
rect 974 -1887 986 -1853
rect 1020 -1887 1032 -1853
rect 974 -1921 1032 -1887
rect 974 -1955 986 -1921
rect 1020 -1955 1032 -1921
rect 974 -1989 1032 -1955
rect 974 -2023 986 -1989
rect 1020 -2023 1032 -1989
rect 974 -2057 1032 -2023
rect 974 -2091 986 -2057
rect 1020 -2091 1032 -2057
rect 974 -2125 1032 -2091
rect 974 -2159 986 -2125
rect 1020 -2159 1032 -2125
rect 974 -2193 1032 -2159
rect 974 -2227 986 -2193
rect 1020 -2227 1032 -2193
rect 974 -2261 1032 -2227
rect 974 -2295 986 -2261
rect 1020 -2295 1032 -2261
rect 974 -2329 1032 -2295
rect 974 -2363 986 -2329
rect 1020 -2363 1032 -2329
rect 974 -2397 1032 -2363
rect 974 -2431 986 -2397
rect 1020 -2431 1032 -2397
rect 974 -2465 1032 -2431
rect 974 -2499 986 -2465
rect 1020 -2499 1032 -2465
rect 974 -2533 1032 -2499
rect 974 -2567 986 -2533
rect 1020 -2567 1032 -2533
rect 974 -2601 1032 -2567
rect 974 -2635 986 -2601
rect 1020 -2635 1032 -2601
rect 974 -2669 1032 -2635
rect 974 -2703 986 -2669
rect 1020 -2703 1032 -2669
rect 974 -2737 1032 -2703
rect 974 -2771 986 -2737
rect 1020 -2771 1032 -2737
rect 974 -2805 1032 -2771
rect 974 -2839 986 -2805
rect 1020 -2839 1032 -2805
rect 974 -2873 1032 -2839
rect 974 -2907 986 -2873
rect 1020 -2907 1032 -2873
rect 974 -2941 1032 -2907
rect 974 -2975 986 -2941
rect 1020 -2975 1032 -2941
rect 974 -3009 1032 -2975
rect 974 -3043 986 -3009
rect 1020 -3043 1032 -3009
rect 974 -3077 1032 -3043
rect 974 -3111 986 -3077
rect 1020 -3111 1032 -3077
rect 974 -3145 1032 -3111
rect 974 -3179 986 -3145
rect 1020 -3179 1032 -3145
rect 974 -3213 1032 -3179
rect 974 -3247 986 -3213
rect 1020 -3247 1032 -3213
rect 974 -3281 1032 -3247
rect 974 -3315 986 -3281
rect 1020 -3315 1032 -3281
rect 974 -3349 1032 -3315
rect 974 -3383 986 -3349
rect 1020 -3383 1032 -3349
rect 974 -3417 1032 -3383
rect 974 -3451 986 -3417
rect 1020 -3451 1032 -3417
rect 974 -3485 1032 -3451
rect 974 -3519 986 -3485
rect 1020 -3519 1032 -3485
rect 974 -3553 1032 -3519
rect 974 -3587 986 -3553
rect 1020 -3587 1032 -3553
rect 974 -3621 1032 -3587
rect 974 -3655 986 -3621
rect 1020 -3655 1032 -3621
rect 974 -3689 1032 -3655
rect 974 -3723 986 -3689
rect 1020 -3723 1032 -3689
rect 974 -3757 1032 -3723
rect 974 -3791 986 -3757
rect 1020 -3791 1032 -3757
rect 974 -3825 1032 -3791
rect 974 -3859 986 -3825
rect 1020 -3859 1032 -3825
rect 974 -3893 1032 -3859
rect 974 -3927 986 -3893
rect 1020 -3927 1032 -3893
rect 974 -3961 1032 -3927
rect 974 -3995 986 -3961
rect 1020 -3995 1032 -3961
rect 974 -4029 1032 -3995
rect 974 -4063 986 -4029
rect 1020 -4063 1032 -4029
rect 974 -4097 1032 -4063
rect 974 -4131 986 -4097
rect 1020 -4131 1032 -4097
rect 974 -4165 1032 -4131
rect 974 -4199 986 -4165
rect 1020 -4199 1032 -4165
rect 974 -4233 1032 -4199
rect 974 -4267 986 -4233
rect 1020 -4267 1032 -4233
rect 974 -4301 1032 -4267
rect 974 -4335 986 -4301
rect 1020 -4335 1032 -4301
rect 974 -4369 1032 -4335
rect 974 -4403 986 -4369
rect 1020 -4403 1032 -4369
rect 974 -4437 1032 -4403
rect 974 -4471 986 -4437
rect 1020 -4471 1032 -4437
rect 974 -4505 1032 -4471
rect 974 -4539 986 -4505
rect 1020 -4539 1032 -4505
rect 974 -4573 1032 -4539
rect 974 -4607 986 -4573
rect 1020 -4607 1032 -4573
rect 974 -4641 1032 -4607
rect 974 -4675 986 -4641
rect 1020 -4675 1032 -4641
rect 974 -4709 1032 -4675
rect 974 -4743 986 -4709
rect 1020 -4743 1032 -4709
rect 974 -4777 1032 -4743
rect 974 -4811 986 -4777
rect 1020 -4811 1032 -4777
rect 974 -4845 1032 -4811
rect 974 -4879 986 -4845
rect 1020 -4879 1032 -4845
rect 974 -4913 1032 -4879
rect 974 -4947 986 -4913
rect 1020 -4947 1032 -4913
rect 974 -4981 1032 -4947
rect 974 -5015 986 -4981
rect 1020 -5015 1032 -4981
rect 974 -5049 1032 -5015
rect 974 -5083 986 -5049
rect 1020 -5083 1032 -5049
rect 974 -5117 1032 -5083
rect 974 -5151 986 -5117
rect 1020 -5151 1032 -5117
rect 974 -5185 1032 -5151
rect 974 -5219 986 -5185
rect 1020 -5219 1032 -5185
rect 974 -5253 1032 -5219
rect 974 -5287 986 -5253
rect 1020 -5287 1032 -5253
rect 974 -5321 1032 -5287
rect 974 -5355 986 -5321
rect 1020 -5355 1032 -5321
rect 974 -5389 1032 -5355
rect 974 -5423 986 -5389
rect 1020 -5423 1032 -5389
rect 974 -5457 1032 -5423
rect 974 -5491 986 -5457
rect 1020 -5491 1032 -5457
rect 974 -5525 1032 -5491
rect 974 -5559 986 -5525
rect 1020 -5559 1032 -5525
rect 974 -5593 1032 -5559
rect 974 -5627 986 -5593
rect 1020 -5627 1032 -5593
rect 974 -5661 1032 -5627
rect 974 -5695 986 -5661
rect 1020 -5695 1032 -5661
rect 974 -5729 1032 -5695
rect 974 -5763 986 -5729
rect 1020 -5763 1032 -5729
rect 974 -5797 1032 -5763
rect 974 -5831 986 -5797
rect 1020 -5831 1032 -5797
rect 974 -5865 1032 -5831
rect 974 -5899 986 -5865
rect 1020 -5899 1032 -5865
rect 974 -5933 1032 -5899
rect 974 -5967 986 -5933
rect 1020 -5967 1032 -5933
rect 974 -6001 1032 -5967
rect 974 -6035 986 -6001
rect 1020 -6035 1032 -6001
rect 974 -6069 1032 -6035
rect 974 -6103 986 -6069
rect 1020 -6103 1032 -6069
rect 974 -6137 1032 -6103
rect 974 -6171 986 -6137
rect 1020 -6171 1032 -6137
rect 974 -6205 1032 -6171
rect 974 -6239 986 -6205
rect 1020 -6239 1032 -6205
rect 974 -6273 1032 -6239
rect 974 -6307 986 -6273
rect 1020 -6307 1032 -6273
rect 974 -6341 1032 -6307
rect 974 -6375 986 -6341
rect 1020 -6375 1032 -6341
rect 974 -6409 1032 -6375
rect 974 -6443 986 -6409
rect 1020 -6443 1032 -6409
rect 974 -6477 1032 -6443
rect 974 -6511 986 -6477
rect 1020 -6511 1032 -6477
rect 974 -6545 1032 -6511
rect 974 -6579 986 -6545
rect 1020 -6579 1032 -6545
rect 974 -6613 1032 -6579
rect 974 -6647 986 -6613
rect 1020 -6647 1032 -6613
rect 974 -6681 1032 -6647
rect 974 -6715 986 -6681
rect 1020 -6715 1032 -6681
rect 974 -6749 1032 -6715
rect 974 -6783 986 -6749
rect 1020 -6783 1032 -6749
rect 974 -6817 1032 -6783
rect 974 -6851 986 -6817
rect 1020 -6851 1032 -6817
rect 974 -6885 1032 -6851
rect 974 -6919 986 -6885
rect 1020 -6919 1032 -6885
rect 974 -6953 1032 -6919
rect 974 -6987 986 -6953
rect 1020 -6987 1032 -6953
rect 974 -7021 1032 -6987
rect 974 -7055 986 -7021
rect 1020 -7055 1032 -7021
rect 974 -7089 1032 -7055
rect 974 -7123 986 -7089
rect 1020 -7123 1032 -7089
rect 974 -7157 1032 -7123
rect 974 -7191 986 -7157
rect 1020 -7191 1032 -7157
rect 974 -7225 1032 -7191
rect 974 -7259 986 -7225
rect 1020 -7259 1032 -7225
rect 974 -7293 1032 -7259
rect 974 -7327 986 -7293
rect 1020 -7327 1032 -7293
rect 974 -7361 1032 -7327
rect 974 -7395 986 -7361
rect 1020 -7395 1032 -7361
rect 974 -7429 1032 -7395
rect 974 -7463 986 -7429
rect 1020 -7463 1032 -7429
rect 974 -7497 1032 -7463
rect 974 -7531 986 -7497
rect 1020 -7531 1032 -7497
rect 974 -7565 1032 -7531
rect 974 -7599 986 -7565
rect 1020 -7599 1032 -7565
rect 974 -7633 1032 -7599
rect 974 -7667 986 -7633
rect 1020 -7667 1032 -7633
rect 974 -7701 1032 -7667
rect 974 -7735 986 -7701
rect 1020 -7735 1032 -7701
rect 974 -7769 1032 -7735
rect 974 -7803 986 -7769
rect 1020 -7803 1032 -7769
rect 974 -7837 1032 -7803
rect 974 -7871 986 -7837
rect 1020 -7871 1032 -7837
rect 974 -7905 1032 -7871
rect 974 -7939 986 -7905
rect 1020 -7939 1032 -7905
rect 974 -7973 1032 -7939
rect 974 -8007 986 -7973
rect 1020 -8007 1032 -7973
rect 974 -8041 1032 -8007
rect 974 -8075 986 -8041
rect 1020 -8075 1032 -8041
rect 974 -8109 1032 -8075
rect 974 -8143 986 -8109
rect 1020 -8143 1032 -8109
rect 974 -8177 1032 -8143
rect 974 -8211 986 -8177
rect 1020 -8211 1032 -8177
rect 974 -8245 1032 -8211
rect 974 -8279 986 -8245
rect 1020 -8279 1032 -8245
rect 974 -8313 1032 -8279
rect 974 -8347 986 -8313
rect 1020 -8347 1032 -8313
rect 974 -8381 1032 -8347
rect 974 -8415 986 -8381
rect 1020 -8415 1032 -8381
rect 974 -8449 1032 -8415
rect 974 -8483 986 -8449
rect 1020 -8483 1032 -8449
rect 974 -8517 1032 -8483
rect 974 -8551 986 -8517
rect 1020 -8551 1032 -8517
rect 974 -8585 1032 -8551
rect 974 -8619 986 -8585
rect 1020 -8619 1032 -8585
rect 974 -8653 1032 -8619
rect 974 -8687 986 -8653
rect 1020 -8687 1032 -8653
rect 974 -8721 1032 -8687
rect 974 -8755 986 -8721
rect 1020 -8755 1032 -8721
rect 974 -8789 1032 -8755
rect 974 -8823 986 -8789
rect 1020 -8823 1032 -8789
rect 974 -8857 1032 -8823
rect 974 -8891 986 -8857
rect 1020 -8891 1032 -8857
rect 974 -8925 1032 -8891
rect 974 -8959 986 -8925
rect 1020 -8959 1032 -8925
rect 974 -8993 1032 -8959
rect 974 -9027 986 -8993
rect 1020 -9027 1032 -8993
rect 974 -9061 1032 -9027
rect 974 -9095 986 -9061
rect 1020 -9095 1032 -9061
rect 974 -9129 1032 -9095
rect 974 -9163 986 -9129
rect 1020 -9163 1032 -9129
rect 974 -9197 1032 -9163
rect 974 -9231 986 -9197
rect 1020 -9231 1032 -9197
rect 974 -9265 1032 -9231
rect 974 -9299 986 -9265
rect 1020 -9299 1032 -9265
rect 974 -9333 1032 -9299
rect 974 -9367 986 -9333
rect 1020 -9367 1032 -9333
rect 974 -9401 1032 -9367
rect 974 -9435 986 -9401
rect 1020 -9435 1032 -9401
rect 974 -9469 1032 -9435
rect 974 -9503 986 -9469
rect 1020 -9503 1032 -9469
rect 974 -9537 1032 -9503
rect 974 -9571 986 -9537
rect 1020 -9571 1032 -9537
rect 974 -9600 1032 -9571
rect 1092 9571 1150 9600
rect 1092 9537 1104 9571
rect 1138 9537 1150 9571
rect 1092 9503 1150 9537
rect 1092 9469 1104 9503
rect 1138 9469 1150 9503
rect 1092 9435 1150 9469
rect 1092 9401 1104 9435
rect 1138 9401 1150 9435
rect 1092 9367 1150 9401
rect 1092 9333 1104 9367
rect 1138 9333 1150 9367
rect 1092 9299 1150 9333
rect 1092 9265 1104 9299
rect 1138 9265 1150 9299
rect 1092 9231 1150 9265
rect 1092 9197 1104 9231
rect 1138 9197 1150 9231
rect 1092 9163 1150 9197
rect 1092 9129 1104 9163
rect 1138 9129 1150 9163
rect 1092 9095 1150 9129
rect 1092 9061 1104 9095
rect 1138 9061 1150 9095
rect 1092 9027 1150 9061
rect 1092 8993 1104 9027
rect 1138 8993 1150 9027
rect 1092 8959 1150 8993
rect 1092 8925 1104 8959
rect 1138 8925 1150 8959
rect 1092 8891 1150 8925
rect 1092 8857 1104 8891
rect 1138 8857 1150 8891
rect 1092 8823 1150 8857
rect 1092 8789 1104 8823
rect 1138 8789 1150 8823
rect 1092 8755 1150 8789
rect 1092 8721 1104 8755
rect 1138 8721 1150 8755
rect 1092 8687 1150 8721
rect 1092 8653 1104 8687
rect 1138 8653 1150 8687
rect 1092 8619 1150 8653
rect 1092 8585 1104 8619
rect 1138 8585 1150 8619
rect 1092 8551 1150 8585
rect 1092 8517 1104 8551
rect 1138 8517 1150 8551
rect 1092 8483 1150 8517
rect 1092 8449 1104 8483
rect 1138 8449 1150 8483
rect 1092 8415 1150 8449
rect 1092 8381 1104 8415
rect 1138 8381 1150 8415
rect 1092 8347 1150 8381
rect 1092 8313 1104 8347
rect 1138 8313 1150 8347
rect 1092 8279 1150 8313
rect 1092 8245 1104 8279
rect 1138 8245 1150 8279
rect 1092 8211 1150 8245
rect 1092 8177 1104 8211
rect 1138 8177 1150 8211
rect 1092 8143 1150 8177
rect 1092 8109 1104 8143
rect 1138 8109 1150 8143
rect 1092 8075 1150 8109
rect 1092 8041 1104 8075
rect 1138 8041 1150 8075
rect 1092 8007 1150 8041
rect 1092 7973 1104 8007
rect 1138 7973 1150 8007
rect 1092 7939 1150 7973
rect 1092 7905 1104 7939
rect 1138 7905 1150 7939
rect 1092 7871 1150 7905
rect 1092 7837 1104 7871
rect 1138 7837 1150 7871
rect 1092 7803 1150 7837
rect 1092 7769 1104 7803
rect 1138 7769 1150 7803
rect 1092 7735 1150 7769
rect 1092 7701 1104 7735
rect 1138 7701 1150 7735
rect 1092 7667 1150 7701
rect 1092 7633 1104 7667
rect 1138 7633 1150 7667
rect 1092 7599 1150 7633
rect 1092 7565 1104 7599
rect 1138 7565 1150 7599
rect 1092 7531 1150 7565
rect 1092 7497 1104 7531
rect 1138 7497 1150 7531
rect 1092 7463 1150 7497
rect 1092 7429 1104 7463
rect 1138 7429 1150 7463
rect 1092 7395 1150 7429
rect 1092 7361 1104 7395
rect 1138 7361 1150 7395
rect 1092 7327 1150 7361
rect 1092 7293 1104 7327
rect 1138 7293 1150 7327
rect 1092 7259 1150 7293
rect 1092 7225 1104 7259
rect 1138 7225 1150 7259
rect 1092 7191 1150 7225
rect 1092 7157 1104 7191
rect 1138 7157 1150 7191
rect 1092 7123 1150 7157
rect 1092 7089 1104 7123
rect 1138 7089 1150 7123
rect 1092 7055 1150 7089
rect 1092 7021 1104 7055
rect 1138 7021 1150 7055
rect 1092 6987 1150 7021
rect 1092 6953 1104 6987
rect 1138 6953 1150 6987
rect 1092 6919 1150 6953
rect 1092 6885 1104 6919
rect 1138 6885 1150 6919
rect 1092 6851 1150 6885
rect 1092 6817 1104 6851
rect 1138 6817 1150 6851
rect 1092 6783 1150 6817
rect 1092 6749 1104 6783
rect 1138 6749 1150 6783
rect 1092 6715 1150 6749
rect 1092 6681 1104 6715
rect 1138 6681 1150 6715
rect 1092 6647 1150 6681
rect 1092 6613 1104 6647
rect 1138 6613 1150 6647
rect 1092 6579 1150 6613
rect 1092 6545 1104 6579
rect 1138 6545 1150 6579
rect 1092 6511 1150 6545
rect 1092 6477 1104 6511
rect 1138 6477 1150 6511
rect 1092 6443 1150 6477
rect 1092 6409 1104 6443
rect 1138 6409 1150 6443
rect 1092 6375 1150 6409
rect 1092 6341 1104 6375
rect 1138 6341 1150 6375
rect 1092 6307 1150 6341
rect 1092 6273 1104 6307
rect 1138 6273 1150 6307
rect 1092 6239 1150 6273
rect 1092 6205 1104 6239
rect 1138 6205 1150 6239
rect 1092 6171 1150 6205
rect 1092 6137 1104 6171
rect 1138 6137 1150 6171
rect 1092 6103 1150 6137
rect 1092 6069 1104 6103
rect 1138 6069 1150 6103
rect 1092 6035 1150 6069
rect 1092 6001 1104 6035
rect 1138 6001 1150 6035
rect 1092 5967 1150 6001
rect 1092 5933 1104 5967
rect 1138 5933 1150 5967
rect 1092 5899 1150 5933
rect 1092 5865 1104 5899
rect 1138 5865 1150 5899
rect 1092 5831 1150 5865
rect 1092 5797 1104 5831
rect 1138 5797 1150 5831
rect 1092 5763 1150 5797
rect 1092 5729 1104 5763
rect 1138 5729 1150 5763
rect 1092 5695 1150 5729
rect 1092 5661 1104 5695
rect 1138 5661 1150 5695
rect 1092 5627 1150 5661
rect 1092 5593 1104 5627
rect 1138 5593 1150 5627
rect 1092 5559 1150 5593
rect 1092 5525 1104 5559
rect 1138 5525 1150 5559
rect 1092 5491 1150 5525
rect 1092 5457 1104 5491
rect 1138 5457 1150 5491
rect 1092 5423 1150 5457
rect 1092 5389 1104 5423
rect 1138 5389 1150 5423
rect 1092 5355 1150 5389
rect 1092 5321 1104 5355
rect 1138 5321 1150 5355
rect 1092 5287 1150 5321
rect 1092 5253 1104 5287
rect 1138 5253 1150 5287
rect 1092 5219 1150 5253
rect 1092 5185 1104 5219
rect 1138 5185 1150 5219
rect 1092 5151 1150 5185
rect 1092 5117 1104 5151
rect 1138 5117 1150 5151
rect 1092 5083 1150 5117
rect 1092 5049 1104 5083
rect 1138 5049 1150 5083
rect 1092 5015 1150 5049
rect 1092 4981 1104 5015
rect 1138 4981 1150 5015
rect 1092 4947 1150 4981
rect 1092 4913 1104 4947
rect 1138 4913 1150 4947
rect 1092 4879 1150 4913
rect 1092 4845 1104 4879
rect 1138 4845 1150 4879
rect 1092 4811 1150 4845
rect 1092 4777 1104 4811
rect 1138 4777 1150 4811
rect 1092 4743 1150 4777
rect 1092 4709 1104 4743
rect 1138 4709 1150 4743
rect 1092 4675 1150 4709
rect 1092 4641 1104 4675
rect 1138 4641 1150 4675
rect 1092 4607 1150 4641
rect 1092 4573 1104 4607
rect 1138 4573 1150 4607
rect 1092 4539 1150 4573
rect 1092 4505 1104 4539
rect 1138 4505 1150 4539
rect 1092 4471 1150 4505
rect 1092 4437 1104 4471
rect 1138 4437 1150 4471
rect 1092 4403 1150 4437
rect 1092 4369 1104 4403
rect 1138 4369 1150 4403
rect 1092 4335 1150 4369
rect 1092 4301 1104 4335
rect 1138 4301 1150 4335
rect 1092 4267 1150 4301
rect 1092 4233 1104 4267
rect 1138 4233 1150 4267
rect 1092 4199 1150 4233
rect 1092 4165 1104 4199
rect 1138 4165 1150 4199
rect 1092 4131 1150 4165
rect 1092 4097 1104 4131
rect 1138 4097 1150 4131
rect 1092 4063 1150 4097
rect 1092 4029 1104 4063
rect 1138 4029 1150 4063
rect 1092 3995 1150 4029
rect 1092 3961 1104 3995
rect 1138 3961 1150 3995
rect 1092 3927 1150 3961
rect 1092 3893 1104 3927
rect 1138 3893 1150 3927
rect 1092 3859 1150 3893
rect 1092 3825 1104 3859
rect 1138 3825 1150 3859
rect 1092 3791 1150 3825
rect 1092 3757 1104 3791
rect 1138 3757 1150 3791
rect 1092 3723 1150 3757
rect 1092 3689 1104 3723
rect 1138 3689 1150 3723
rect 1092 3655 1150 3689
rect 1092 3621 1104 3655
rect 1138 3621 1150 3655
rect 1092 3587 1150 3621
rect 1092 3553 1104 3587
rect 1138 3553 1150 3587
rect 1092 3519 1150 3553
rect 1092 3485 1104 3519
rect 1138 3485 1150 3519
rect 1092 3451 1150 3485
rect 1092 3417 1104 3451
rect 1138 3417 1150 3451
rect 1092 3383 1150 3417
rect 1092 3349 1104 3383
rect 1138 3349 1150 3383
rect 1092 3315 1150 3349
rect 1092 3281 1104 3315
rect 1138 3281 1150 3315
rect 1092 3247 1150 3281
rect 1092 3213 1104 3247
rect 1138 3213 1150 3247
rect 1092 3179 1150 3213
rect 1092 3145 1104 3179
rect 1138 3145 1150 3179
rect 1092 3111 1150 3145
rect 1092 3077 1104 3111
rect 1138 3077 1150 3111
rect 1092 3043 1150 3077
rect 1092 3009 1104 3043
rect 1138 3009 1150 3043
rect 1092 2975 1150 3009
rect 1092 2941 1104 2975
rect 1138 2941 1150 2975
rect 1092 2907 1150 2941
rect 1092 2873 1104 2907
rect 1138 2873 1150 2907
rect 1092 2839 1150 2873
rect 1092 2805 1104 2839
rect 1138 2805 1150 2839
rect 1092 2771 1150 2805
rect 1092 2737 1104 2771
rect 1138 2737 1150 2771
rect 1092 2703 1150 2737
rect 1092 2669 1104 2703
rect 1138 2669 1150 2703
rect 1092 2635 1150 2669
rect 1092 2601 1104 2635
rect 1138 2601 1150 2635
rect 1092 2567 1150 2601
rect 1092 2533 1104 2567
rect 1138 2533 1150 2567
rect 1092 2499 1150 2533
rect 1092 2465 1104 2499
rect 1138 2465 1150 2499
rect 1092 2431 1150 2465
rect 1092 2397 1104 2431
rect 1138 2397 1150 2431
rect 1092 2363 1150 2397
rect 1092 2329 1104 2363
rect 1138 2329 1150 2363
rect 1092 2295 1150 2329
rect 1092 2261 1104 2295
rect 1138 2261 1150 2295
rect 1092 2227 1150 2261
rect 1092 2193 1104 2227
rect 1138 2193 1150 2227
rect 1092 2159 1150 2193
rect 1092 2125 1104 2159
rect 1138 2125 1150 2159
rect 1092 2091 1150 2125
rect 1092 2057 1104 2091
rect 1138 2057 1150 2091
rect 1092 2023 1150 2057
rect 1092 1989 1104 2023
rect 1138 1989 1150 2023
rect 1092 1955 1150 1989
rect 1092 1921 1104 1955
rect 1138 1921 1150 1955
rect 1092 1887 1150 1921
rect 1092 1853 1104 1887
rect 1138 1853 1150 1887
rect 1092 1819 1150 1853
rect 1092 1785 1104 1819
rect 1138 1785 1150 1819
rect 1092 1751 1150 1785
rect 1092 1717 1104 1751
rect 1138 1717 1150 1751
rect 1092 1683 1150 1717
rect 1092 1649 1104 1683
rect 1138 1649 1150 1683
rect 1092 1615 1150 1649
rect 1092 1581 1104 1615
rect 1138 1581 1150 1615
rect 1092 1547 1150 1581
rect 1092 1513 1104 1547
rect 1138 1513 1150 1547
rect 1092 1479 1150 1513
rect 1092 1445 1104 1479
rect 1138 1445 1150 1479
rect 1092 1411 1150 1445
rect 1092 1377 1104 1411
rect 1138 1377 1150 1411
rect 1092 1343 1150 1377
rect 1092 1309 1104 1343
rect 1138 1309 1150 1343
rect 1092 1275 1150 1309
rect 1092 1241 1104 1275
rect 1138 1241 1150 1275
rect 1092 1207 1150 1241
rect 1092 1173 1104 1207
rect 1138 1173 1150 1207
rect 1092 1139 1150 1173
rect 1092 1105 1104 1139
rect 1138 1105 1150 1139
rect 1092 1071 1150 1105
rect 1092 1037 1104 1071
rect 1138 1037 1150 1071
rect 1092 1003 1150 1037
rect 1092 969 1104 1003
rect 1138 969 1150 1003
rect 1092 935 1150 969
rect 1092 901 1104 935
rect 1138 901 1150 935
rect 1092 867 1150 901
rect 1092 833 1104 867
rect 1138 833 1150 867
rect 1092 799 1150 833
rect 1092 765 1104 799
rect 1138 765 1150 799
rect 1092 731 1150 765
rect 1092 697 1104 731
rect 1138 697 1150 731
rect 1092 663 1150 697
rect 1092 629 1104 663
rect 1138 629 1150 663
rect 1092 595 1150 629
rect 1092 561 1104 595
rect 1138 561 1150 595
rect 1092 527 1150 561
rect 1092 493 1104 527
rect 1138 493 1150 527
rect 1092 459 1150 493
rect 1092 425 1104 459
rect 1138 425 1150 459
rect 1092 391 1150 425
rect 1092 357 1104 391
rect 1138 357 1150 391
rect 1092 323 1150 357
rect 1092 289 1104 323
rect 1138 289 1150 323
rect 1092 255 1150 289
rect 1092 221 1104 255
rect 1138 221 1150 255
rect 1092 187 1150 221
rect 1092 153 1104 187
rect 1138 153 1150 187
rect 1092 119 1150 153
rect 1092 85 1104 119
rect 1138 85 1150 119
rect 1092 51 1150 85
rect 1092 17 1104 51
rect 1138 17 1150 51
rect 1092 -17 1150 17
rect 1092 -51 1104 -17
rect 1138 -51 1150 -17
rect 1092 -85 1150 -51
rect 1092 -119 1104 -85
rect 1138 -119 1150 -85
rect 1092 -153 1150 -119
rect 1092 -187 1104 -153
rect 1138 -187 1150 -153
rect 1092 -221 1150 -187
rect 1092 -255 1104 -221
rect 1138 -255 1150 -221
rect 1092 -289 1150 -255
rect 1092 -323 1104 -289
rect 1138 -323 1150 -289
rect 1092 -357 1150 -323
rect 1092 -391 1104 -357
rect 1138 -391 1150 -357
rect 1092 -425 1150 -391
rect 1092 -459 1104 -425
rect 1138 -459 1150 -425
rect 1092 -493 1150 -459
rect 1092 -527 1104 -493
rect 1138 -527 1150 -493
rect 1092 -561 1150 -527
rect 1092 -595 1104 -561
rect 1138 -595 1150 -561
rect 1092 -629 1150 -595
rect 1092 -663 1104 -629
rect 1138 -663 1150 -629
rect 1092 -697 1150 -663
rect 1092 -731 1104 -697
rect 1138 -731 1150 -697
rect 1092 -765 1150 -731
rect 1092 -799 1104 -765
rect 1138 -799 1150 -765
rect 1092 -833 1150 -799
rect 1092 -867 1104 -833
rect 1138 -867 1150 -833
rect 1092 -901 1150 -867
rect 1092 -935 1104 -901
rect 1138 -935 1150 -901
rect 1092 -969 1150 -935
rect 1092 -1003 1104 -969
rect 1138 -1003 1150 -969
rect 1092 -1037 1150 -1003
rect 1092 -1071 1104 -1037
rect 1138 -1071 1150 -1037
rect 1092 -1105 1150 -1071
rect 1092 -1139 1104 -1105
rect 1138 -1139 1150 -1105
rect 1092 -1173 1150 -1139
rect 1092 -1207 1104 -1173
rect 1138 -1207 1150 -1173
rect 1092 -1241 1150 -1207
rect 1092 -1275 1104 -1241
rect 1138 -1275 1150 -1241
rect 1092 -1309 1150 -1275
rect 1092 -1343 1104 -1309
rect 1138 -1343 1150 -1309
rect 1092 -1377 1150 -1343
rect 1092 -1411 1104 -1377
rect 1138 -1411 1150 -1377
rect 1092 -1445 1150 -1411
rect 1092 -1479 1104 -1445
rect 1138 -1479 1150 -1445
rect 1092 -1513 1150 -1479
rect 1092 -1547 1104 -1513
rect 1138 -1547 1150 -1513
rect 1092 -1581 1150 -1547
rect 1092 -1615 1104 -1581
rect 1138 -1615 1150 -1581
rect 1092 -1649 1150 -1615
rect 1092 -1683 1104 -1649
rect 1138 -1683 1150 -1649
rect 1092 -1717 1150 -1683
rect 1092 -1751 1104 -1717
rect 1138 -1751 1150 -1717
rect 1092 -1785 1150 -1751
rect 1092 -1819 1104 -1785
rect 1138 -1819 1150 -1785
rect 1092 -1853 1150 -1819
rect 1092 -1887 1104 -1853
rect 1138 -1887 1150 -1853
rect 1092 -1921 1150 -1887
rect 1092 -1955 1104 -1921
rect 1138 -1955 1150 -1921
rect 1092 -1989 1150 -1955
rect 1092 -2023 1104 -1989
rect 1138 -2023 1150 -1989
rect 1092 -2057 1150 -2023
rect 1092 -2091 1104 -2057
rect 1138 -2091 1150 -2057
rect 1092 -2125 1150 -2091
rect 1092 -2159 1104 -2125
rect 1138 -2159 1150 -2125
rect 1092 -2193 1150 -2159
rect 1092 -2227 1104 -2193
rect 1138 -2227 1150 -2193
rect 1092 -2261 1150 -2227
rect 1092 -2295 1104 -2261
rect 1138 -2295 1150 -2261
rect 1092 -2329 1150 -2295
rect 1092 -2363 1104 -2329
rect 1138 -2363 1150 -2329
rect 1092 -2397 1150 -2363
rect 1092 -2431 1104 -2397
rect 1138 -2431 1150 -2397
rect 1092 -2465 1150 -2431
rect 1092 -2499 1104 -2465
rect 1138 -2499 1150 -2465
rect 1092 -2533 1150 -2499
rect 1092 -2567 1104 -2533
rect 1138 -2567 1150 -2533
rect 1092 -2601 1150 -2567
rect 1092 -2635 1104 -2601
rect 1138 -2635 1150 -2601
rect 1092 -2669 1150 -2635
rect 1092 -2703 1104 -2669
rect 1138 -2703 1150 -2669
rect 1092 -2737 1150 -2703
rect 1092 -2771 1104 -2737
rect 1138 -2771 1150 -2737
rect 1092 -2805 1150 -2771
rect 1092 -2839 1104 -2805
rect 1138 -2839 1150 -2805
rect 1092 -2873 1150 -2839
rect 1092 -2907 1104 -2873
rect 1138 -2907 1150 -2873
rect 1092 -2941 1150 -2907
rect 1092 -2975 1104 -2941
rect 1138 -2975 1150 -2941
rect 1092 -3009 1150 -2975
rect 1092 -3043 1104 -3009
rect 1138 -3043 1150 -3009
rect 1092 -3077 1150 -3043
rect 1092 -3111 1104 -3077
rect 1138 -3111 1150 -3077
rect 1092 -3145 1150 -3111
rect 1092 -3179 1104 -3145
rect 1138 -3179 1150 -3145
rect 1092 -3213 1150 -3179
rect 1092 -3247 1104 -3213
rect 1138 -3247 1150 -3213
rect 1092 -3281 1150 -3247
rect 1092 -3315 1104 -3281
rect 1138 -3315 1150 -3281
rect 1092 -3349 1150 -3315
rect 1092 -3383 1104 -3349
rect 1138 -3383 1150 -3349
rect 1092 -3417 1150 -3383
rect 1092 -3451 1104 -3417
rect 1138 -3451 1150 -3417
rect 1092 -3485 1150 -3451
rect 1092 -3519 1104 -3485
rect 1138 -3519 1150 -3485
rect 1092 -3553 1150 -3519
rect 1092 -3587 1104 -3553
rect 1138 -3587 1150 -3553
rect 1092 -3621 1150 -3587
rect 1092 -3655 1104 -3621
rect 1138 -3655 1150 -3621
rect 1092 -3689 1150 -3655
rect 1092 -3723 1104 -3689
rect 1138 -3723 1150 -3689
rect 1092 -3757 1150 -3723
rect 1092 -3791 1104 -3757
rect 1138 -3791 1150 -3757
rect 1092 -3825 1150 -3791
rect 1092 -3859 1104 -3825
rect 1138 -3859 1150 -3825
rect 1092 -3893 1150 -3859
rect 1092 -3927 1104 -3893
rect 1138 -3927 1150 -3893
rect 1092 -3961 1150 -3927
rect 1092 -3995 1104 -3961
rect 1138 -3995 1150 -3961
rect 1092 -4029 1150 -3995
rect 1092 -4063 1104 -4029
rect 1138 -4063 1150 -4029
rect 1092 -4097 1150 -4063
rect 1092 -4131 1104 -4097
rect 1138 -4131 1150 -4097
rect 1092 -4165 1150 -4131
rect 1092 -4199 1104 -4165
rect 1138 -4199 1150 -4165
rect 1092 -4233 1150 -4199
rect 1092 -4267 1104 -4233
rect 1138 -4267 1150 -4233
rect 1092 -4301 1150 -4267
rect 1092 -4335 1104 -4301
rect 1138 -4335 1150 -4301
rect 1092 -4369 1150 -4335
rect 1092 -4403 1104 -4369
rect 1138 -4403 1150 -4369
rect 1092 -4437 1150 -4403
rect 1092 -4471 1104 -4437
rect 1138 -4471 1150 -4437
rect 1092 -4505 1150 -4471
rect 1092 -4539 1104 -4505
rect 1138 -4539 1150 -4505
rect 1092 -4573 1150 -4539
rect 1092 -4607 1104 -4573
rect 1138 -4607 1150 -4573
rect 1092 -4641 1150 -4607
rect 1092 -4675 1104 -4641
rect 1138 -4675 1150 -4641
rect 1092 -4709 1150 -4675
rect 1092 -4743 1104 -4709
rect 1138 -4743 1150 -4709
rect 1092 -4777 1150 -4743
rect 1092 -4811 1104 -4777
rect 1138 -4811 1150 -4777
rect 1092 -4845 1150 -4811
rect 1092 -4879 1104 -4845
rect 1138 -4879 1150 -4845
rect 1092 -4913 1150 -4879
rect 1092 -4947 1104 -4913
rect 1138 -4947 1150 -4913
rect 1092 -4981 1150 -4947
rect 1092 -5015 1104 -4981
rect 1138 -5015 1150 -4981
rect 1092 -5049 1150 -5015
rect 1092 -5083 1104 -5049
rect 1138 -5083 1150 -5049
rect 1092 -5117 1150 -5083
rect 1092 -5151 1104 -5117
rect 1138 -5151 1150 -5117
rect 1092 -5185 1150 -5151
rect 1092 -5219 1104 -5185
rect 1138 -5219 1150 -5185
rect 1092 -5253 1150 -5219
rect 1092 -5287 1104 -5253
rect 1138 -5287 1150 -5253
rect 1092 -5321 1150 -5287
rect 1092 -5355 1104 -5321
rect 1138 -5355 1150 -5321
rect 1092 -5389 1150 -5355
rect 1092 -5423 1104 -5389
rect 1138 -5423 1150 -5389
rect 1092 -5457 1150 -5423
rect 1092 -5491 1104 -5457
rect 1138 -5491 1150 -5457
rect 1092 -5525 1150 -5491
rect 1092 -5559 1104 -5525
rect 1138 -5559 1150 -5525
rect 1092 -5593 1150 -5559
rect 1092 -5627 1104 -5593
rect 1138 -5627 1150 -5593
rect 1092 -5661 1150 -5627
rect 1092 -5695 1104 -5661
rect 1138 -5695 1150 -5661
rect 1092 -5729 1150 -5695
rect 1092 -5763 1104 -5729
rect 1138 -5763 1150 -5729
rect 1092 -5797 1150 -5763
rect 1092 -5831 1104 -5797
rect 1138 -5831 1150 -5797
rect 1092 -5865 1150 -5831
rect 1092 -5899 1104 -5865
rect 1138 -5899 1150 -5865
rect 1092 -5933 1150 -5899
rect 1092 -5967 1104 -5933
rect 1138 -5967 1150 -5933
rect 1092 -6001 1150 -5967
rect 1092 -6035 1104 -6001
rect 1138 -6035 1150 -6001
rect 1092 -6069 1150 -6035
rect 1092 -6103 1104 -6069
rect 1138 -6103 1150 -6069
rect 1092 -6137 1150 -6103
rect 1092 -6171 1104 -6137
rect 1138 -6171 1150 -6137
rect 1092 -6205 1150 -6171
rect 1092 -6239 1104 -6205
rect 1138 -6239 1150 -6205
rect 1092 -6273 1150 -6239
rect 1092 -6307 1104 -6273
rect 1138 -6307 1150 -6273
rect 1092 -6341 1150 -6307
rect 1092 -6375 1104 -6341
rect 1138 -6375 1150 -6341
rect 1092 -6409 1150 -6375
rect 1092 -6443 1104 -6409
rect 1138 -6443 1150 -6409
rect 1092 -6477 1150 -6443
rect 1092 -6511 1104 -6477
rect 1138 -6511 1150 -6477
rect 1092 -6545 1150 -6511
rect 1092 -6579 1104 -6545
rect 1138 -6579 1150 -6545
rect 1092 -6613 1150 -6579
rect 1092 -6647 1104 -6613
rect 1138 -6647 1150 -6613
rect 1092 -6681 1150 -6647
rect 1092 -6715 1104 -6681
rect 1138 -6715 1150 -6681
rect 1092 -6749 1150 -6715
rect 1092 -6783 1104 -6749
rect 1138 -6783 1150 -6749
rect 1092 -6817 1150 -6783
rect 1092 -6851 1104 -6817
rect 1138 -6851 1150 -6817
rect 1092 -6885 1150 -6851
rect 1092 -6919 1104 -6885
rect 1138 -6919 1150 -6885
rect 1092 -6953 1150 -6919
rect 1092 -6987 1104 -6953
rect 1138 -6987 1150 -6953
rect 1092 -7021 1150 -6987
rect 1092 -7055 1104 -7021
rect 1138 -7055 1150 -7021
rect 1092 -7089 1150 -7055
rect 1092 -7123 1104 -7089
rect 1138 -7123 1150 -7089
rect 1092 -7157 1150 -7123
rect 1092 -7191 1104 -7157
rect 1138 -7191 1150 -7157
rect 1092 -7225 1150 -7191
rect 1092 -7259 1104 -7225
rect 1138 -7259 1150 -7225
rect 1092 -7293 1150 -7259
rect 1092 -7327 1104 -7293
rect 1138 -7327 1150 -7293
rect 1092 -7361 1150 -7327
rect 1092 -7395 1104 -7361
rect 1138 -7395 1150 -7361
rect 1092 -7429 1150 -7395
rect 1092 -7463 1104 -7429
rect 1138 -7463 1150 -7429
rect 1092 -7497 1150 -7463
rect 1092 -7531 1104 -7497
rect 1138 -7531 1150 -7497
rect 1092 -7565 1150 -7531
rect 1092 -7599 1104 -7565
rect 1138 -7599 1150 -7565
rect 1092 -7633 1150 -7599
rect 1092 -7667 1104 -7633
rect 1138 -7667 1150 -7633
rect 1092 -7701 1150 -7667
rect 1092 -7735 1104 -7701
rect 1138 -7735 1150 -7701
rect 1092 -7769 1150 -7735
rect 1092 -7803 1104 -7769
rect 1138 -7803 1150 -7769
rect 1092 -7837 1150 -7803
rect 1092 -7871 1104 -7837
rect 1138 -7871 1150 -7837
rect 1092 -7905 1150 -7871
rect 1092 -7939 1104 -7905
rect 1138 -7939 1150 -7905
rect 1092 -7973 1150 -7939
rect 1092 -8007 1104 -7973
rect 1138 -8007 1150 -7973
rect 1092 -8041 1150 -8007
rect 1092 -8075 1104 -8041
rect 1138 -8075 1150 -8041
rect 1092 -8109 1150 -8075
rect 1092 -8143 1104 -8109
rect 1138 -8143 1150 -8109
rect 1092 -8177 1150 -8143
rect 1092 -8211 1104 -8177
rect 1138 -8211 1150 -8177
rect 1092 -8245 1150 -8211
rect 1092 -8279 1104 -8245
rect 1138 -8279 1150 -8245
rect 1092 -8313 1150 -8279
rect 1092 -8347 1104 -8313
rect 1138 -8347 1150 -8313
rect 1092 -8381 1150 -8347
rect 1092 -8415 1104 -8381
rect 1138 -8415 1150 -8381
rect 1092 -8449 1150 -8415
rect 1092 -8483 1104 -8449
rect 1138 -8483 1150 -8449
rect 1092 -8517 1150 -8483
rect 1092 -8551 1104 -8517
rect 1138 -8551 1150 -8517
rect 1092 -8585 1150 -8551
rect 1092 -8619 1104 -8585
rect 1138 -8619 1150 -8585
rect 1092 -8653 1150 -8619
rect 1092 -8687 1104 -8653
rect 1138 -8687 1150 -8653
rect 1092 -8721 1150 -8687
rect 1092 -8755 1104 -8721
rect 1138 -8755 1150 -8721
rect 1092 -8789 1150 -8755
rect 1092 -8823 1104 -8789
rect 1138 -8823 1150 -8789
rect 1092 -8857 1150 -8823
rect 1092 -8891 1104 -8857
rect 1138 -8891 1150 -8857
rect 1092 -8925 1150 -8891
rect 1092 -8959 1104 -8925
rect 1138 -8959 1150 -8925
rect 1092 -8993 1150 -8959
rect 1092 -9027 1104 -8993
rect 1138 -9027 1150 -8993
rect 1092 -9061 1150 -9027
rect 1092 -9095 1104 -9061
rect 1138 -9095 1150 -9061
rect 1092 -9129 1150 -9095
rect 1092 -9163 1104 -9129
rect 1138 -9163 1150 -9129
rect 1092 -9197 1150 -9163
rect 1092 -9231 1104 -9197
rect 1138 -9231 1150 -9197
rect 1092 -9265 1150 -9231
rect 1092 -9299 1104 -9265
rect 1138 -9299 1150 -9265
rect 1092 -9333 1150 -9299
rect 1092 -9367 1104 -9333
rect 1138 -9367 1150 -9333
rect 1092 -9401 1150 -9367
rect 1092 -9435 1104 -9401
rect 1138 -9435 1150 -9401
rect 1092 -9469 1150 -9435
rect 1092 -9503 1104 -9469
rect 1138 -9503 1150 -9469
rect 1092 -9537 1150 -9503
rect 1092 -9571 1104 -9537
rect 1138 -9571 1150 -9537
rect 1092 -9600 1150 -9571
rect 1210 9571 1268 9600
rect 1210 9537 1222 9571
rect 1256 9537 1268 9571
rect 1210 9503 1268 9537
rect 1210 9469 1222 9503
rect 1256 9469 1268 9503
rect 1210 9435 1268 9469
rect 1210 9401 1222 9435
rect 1256 9401 1268 9435
rect 1210 9367 1268 9401
rect 1210 9333 1222 9367
rect 1256 9333 1268 9367
rect 1210 9299 1268 9333
rect 1210 9265 1222 9299
rect 1256 9265 1268 9299
rect 1210 9231 1268 9265
rect 1210 9197 1222 9231
rect 1256 9197 1268 9231
rect 1210 9163 1268 9197
rect 1210 9129 1222 9163
rect 1256 9129 1268 9163
rect 1210 9095 1268 9129
rect 1210 9061 1222 9095
rect 1256 9061 1268 9095
rect 1210 9027 1268 9061
rect 1210 8993 1222 9027
rect 1256 8993 1268 9027
rect 1210 8959 1268 8993
rect 1210 8925 1222 8959
rect 1256 8925 1268 8959
rect 1210 8891 1268 8925
rect 1210 8857 1222 8891
rect 1256 8857 1268 8891
rect 1210 8823 1268 8857
rect 1210 8789 1222 8823
rect 1256 8789 1268 8823
rect 1210 8755 1268 8789
rect 1210 8721 1222 8755
rect 1256 8721 1268 8755
rect 1210 8687 1268 8721
rect 1210 8653 1222 8687
rect 1256 8653 1268 8687
rect 1210 8619 1268 8653
rect 1210 8585 1222 8619
rect 1256 8585 1268 8619
rect 1210 8551 1268 8585
rect 1210 8517 1222 8551
rect 1256 8517 1268 8551
rect 1210 8483 1268 8517
rect 1210 8449 1222 8483
rect 1256 8449 1268 8483
rect 1210 8415 1268 8449
rect 1210 8381 1222 8415
rect 1256 8381 1268 8415
rect 1210 8347 1268 8381
rect 1210 8313 1222 8347
rect 1256 8313 1268 8347
rect 1210 8279 1268 8313
rect 1210 8245 1222 8279
rect 1256 8245 1268 8279
rect 1210 8211 1268 8245
rect 1210 8177 1222 8211
rect 1256 8177 1268 8211
rect 1210 8143 1268 8177
rect 1210 8109 1222 8143
rect 1256 8109 1268 8143
rect 1210 8075 1268 8109
rect 1210 8041 1222 8075
rect 1256 8041 1268 8075
rect 1210 8007 1268 8041
rect 1210 7973 1222 8007
rect 1256 7973 1268 8007
rect 1210 7939 1268 7973
rect 1210 7905 1222 7939
rect 1256 7905 1268 7939
rect 1210 7871 1268 7905
rect 1210 7837 1222 7871
rect 1256 7837 1268 7871
rect 1210 7803 1268 7837
rect 1210 7769 1222 7803
rect 1256 7769 1268 7803
rect 1210 7735 1268 7769
rect 1210 7701 1222 7735
rect 1256 7701 1268 7735
rect 1210 7667 1268 7701
rect 1210 7633 1222 7667
rect 1256 7633 1268 7667
rect 1210 7599 1268 7633
rect 1210 7565 1222 7599
rect 1256 7565 1268 7599
rect 1210 7531 1268 7565
rect 1210 7497 1222 7531
rect 1256 7497 1268 7531
rect 1210 7463 1268 7497
rect 1210 7429 1222 7463
rect 1256 7429 1268 7463
rect 1210 7395 1268 7429
rect 1210 7361 1222 7395
rect 1256 7361 1268 7395
rect 1210 7327 1268 7361
rect 1210 7293 1222 7327
rect 1256 7293 1268 7327
rect 1210 7259 1268 7293
rect 1210 7225 1222 7259
rect 1256 7225 1268 7259
rect 1210 7191 1268 7225
rect 1210 7157 1222 7191
rect 1256 7157 1268 7191
rect 1210 7123 1268 7157
rect 1210 7089 1222 7123
rect 1256 7089 1268 7123
rect 1210 7055 1268 7089
rect 1210 7021 1222 7055
rect 1256 7021 1268 7055
rect 1210 6987 1268 7021
rect 1210 6953 1222 6987
rect 1256 6953 1268 6987
rect 1210 6919 1268 6953
rect 1210 6885 1222 6919
rect 1256 6885 1268 6919
rect 1210 6851 1268 6885
rect 1210 6817 1222 6851
rect 1256 6817 1268 6851
rect 1210 6783 1268 6817
rect 1210 6749 1222 6783
rect 1256 6749 1268 6783
rect 1210 6715 1268 6749
rect 1210 6681 1222 6715
rect 1256 6681 1268 6715
rect 1210 6647 1268 6681
rect 1210 6613 1222 6647
rect 1256 6613 1268 6647
rect 1210 6579 1268 6613
rect 1210 6545 1222 6579
rect 1256 6545 1268 6579
rect 1210 6511 1268 6545
rect 1210 6477 1222 6511
rect 1256 6477 1268 6511
rect 1210 6443 1268 6477
rect 1210 6409 1222 6443
rect 1256 6409 1268 6443
rect 1210 6375 1268 6409
rect 1210 6341 1222 6375
rect 1256 6341 1268 6375
rect 1210 6307 1268 6341
rect 1210 6273 1222 6307
rect 1256 6273 1268 6307
rect 1210 6239 1268 6273
rect 1210 6205 1222 6239
rect 1256 6205 1268 6239
rect 1210 6171 1268 6205
rect 1210 6137 1222 6171
rect 1256 6137 1268 6171
rect 1210 6103 1268 6137
rect 1210 6069 1222 6103
rect 1256 6069 1268 6103
rect 1210 6035 1268 6069
rect 1210 6001 1222 6035
rect 1256 6001 1268 6035
rect 1210 5967 1268 6001
rect 1210 5933 1222 5967
rect 1256 5933 1268 5967
rect 1210 5899 1268 5933
rect 1210 5865 1222 5899
rect 1256 5865 1268 5899
rect 1210 5831 1268 5865
rect 1210 5797 1222 5831
rect 1256 5797 1268 5831
rect 1210 5763 1268 5797
rect 1210 5729 1222 5763
rect 1256 5729 1268 5763
rect 1210 5695 1268 5729
rect 1210 5661 1222 5695
rect 1256 5661 1268 5695
rect 1210 5627 1268 5661
rect 1210 5593 1222 5627
rect 1256 5593 1268 5627
rect 1210 5559 1268 5593
rect 1210 5525 1222 5559
rect 1256 5525 1268 5559
rect 1210 5491 1268 5525
rect 1210 5457 1222 5491
rect 1256 5457 1268 5491
rect 1210 5423 1268 5457
rect 1210 5389 1222 5423
rect 1256 5389 1268 5423
rect 1210 5355 1268 5389
rect 1210 5321 1222 5355
rect 1256 5321 1268 5355
rect 1210 5287 1268 5321
rect 1210 5253 1222 5287
rect 1256 5253 1268 5287
rect 1210 5219 1268 5253
rect 1210 5185 1222 5219
rect 1256 5185 1268 5219
rect 1210 5151 1268 5185
rect 1210 5117 1222 5151
rect 1256 5117 1268 5151
rect 1210 5083 1268 5117
rect 1210 5049 1222 5083
rect 1256 5049 1268 5083
rect 1210 5015 1268 5049
rect 1210 4981 1222 5015
rect 1256 4981 1268 5015
rect 1210 4947 1268 4981
rect 1210 4913 1222 4947
rect 1256 4913 1268 4947
rect 1210 4879 1268 4913
rect 1210 4845 1222 4879
rect 1256 4845 1268 4879
rect 1210 4811 1268 4845
rect 1210 4777 1222 4811
rect 1256 4777 1268 4811
rect 1210 4743 1268 4777
rect 1210 4709 1222 4743
rect 1256 4709 1268 4743
rect 1210 4675 1268 4709
rect 1210 4641 1222 4675
rect 1256 4641 1268 4675
rect 1210 4607 1268 4641
rect 1210 4573 1222 4607
rect 1256 4573 1268 4607
rect 1210 4539 1268 4573
rect 1210 4505 1222 4539
rect 1256 4505 1268 4539
rect 1210 4471 1268 4505
rect 1210 4437 1222 4471
rect 1256 4437 1268 4471
rect 1210 4403 1268 4437
rect 1210 4369 1222 4403
rect 1256 4369 1268 4403
rect 1210 4335 1268 4369
rect 1210 4301 1222 4335
rect 1256 4301 1268 4335
rect 1210 4267 1268 4301
rect 1210 4233 1222 4267
rect 1256 4233 1268 4267
rect 1210 4199 1268 4233
rect 1210 4165 1222 4199
rect 1256 4165 1268 4199
rect 1210 4131 1268 4165
rect 1210 4097 1222 4131
rect 1256 4097 1268 4131
rect 1210 4063 1268 4097
rect 1210 4029 1222 4063
rect 1256 4029 1268 4063
rect 1210 3995 1268 4029
rect 1210 3961 1222 3995
rect 1256 3961 1268 3995
rect 1210 3927 1268 3961
rect 1210 3893 1222 3927
rect 1256 3893 1268 3927
rect 1210 3859 1268 3893
rect 1210 3825 1222 3859
rect 1256 3825 1268 3859
rect 1210 3791 1268 3825
rect 1210 3757 1222 3791
rect 1256 3757 1268 3791
rect 1210 3723 1268 3757
rect 1210 3689 1222 3723
rect 1256 3689 1268 3723
rect 1210 3655 1268 3689
rect 1210 3621 1222 3655
rect 1256 3621 1268 3655
rect 1210 3587 1268 3621
rect 1210 3553 1222 3587
rect 1256 3553 1268 3587
rect 1210 3519 1268 3553
rect 1210 3485 1222 3519
rect 1256 3485 1268 3519
rect 1210 3451 1268 3485
rect 1210 3417 1222 3451
rect 1256 3417 1268 3451
rect 1210 3383 1268 3417
rect 1210 3349 1222 3383
rect 1256 3349 1268 3383
rect 1210 3315 1268 3349
rect 1210 3281 1222 3315
rect 1256 3281 1268 3315
rect 1210 3247 1268 3281
rect 1210 3213 1222 3247
rect 1256 3213 1268 3247
rect 1210 3179 1268 3213
rect 1210 3145 1222 3179
rect 1256 3145 1268 3179
rect 1210 3111 1268 3145
rect 1210 3077 1222 3111
rect 1256 3077 1268 3111
rect 1210 3043 1268 3077
rect 1210 3009 1222 3043
rect 1256 3009 1268 3043
rect 1210 2975 1268 3009
rect 1210 2941 1222 2975
rect 1256 2941 1268 2975
rect 1210 2907 1268 2941
rect 1210 2873 1222 2907
rect 1256 2873 1268 2907
rect 1210 2839 1268 2873
rect 1210 2805 1222 2839
rect 1256 2805 1268 2839
rect 1210 2771 1268 2805
rect 1210 2737 1222 2771
rect 1256 2737 1268 2771
rect 1210 2703 1268 2737
rect 1210 2669 1222 2703
rect 1256 2669 1268 2703
rect 1210 2635 1268 2669
rect 1210 2601 1222 2635
rect 1256 2601 1268 2635
rect 1210 2567 1268 2601
rect 1210 2533 1222 2567
rect 1256 2533 1268 2567
rect 1210 2499 1268 2533
rect 1210 2465 1222 2499
rect 1256 2465 1268 2499
rect 1210 2431 1268 2465
rect 1210 2397 1222 2431
rect 1256 2397 1268 2431
rect 1210 2363 1268 2397
rect 1210 2329 1222 2363
rect 1256 2329 1268 2363
rect 1210 2295 1268 2329
rect 1210 2261 1222 2295
rect 1256 2261 1268 2295
rect 1210 2227 1268 2261
rect 1210 2193 1222 2227
rect 1256 2193 1268 2227
rect 1210 2159 1268 2193
rect 1210 2125 1222 2159
rect 1256 2125 1268 2159
rect 1210 2091 1268 2125
rect 1210 2057 1222 2091
rect 1256 2057 1268 2091
rect 1210 2023 1268 2057
rect 1210 1989 1222 2023
rect 1256 1989 1268 2023
rect 1210 1955 1268 1989
rect 1210 1921 1222 1955
rect 1256 1921 1268 1955
rect 1210 1887 1268 1921
rect 1210 1853 1222 1887
rect 1256 1853 1268 1887
rect 1210 1819 1268 1853
rect 1210 1785 1222 1819
rect 1256 1785 1268 1819
rect 1210 1751 1268 1785
rect 1210 1717 1222 1751
rect 1256 1717 1268 1751
rect 1210 1683 1268 1717
rect 1210 1649 1222 1683
rect 1256 1649 1268 1683
rect 1210 1615 1268 1649
rect 1210 1581 1222 1615
rect 1256 1581 1268 1615
rect 1210 1547 1268 1581
rect 1210 1513 1222 1547
rect 1256 1513 1268 1547
rect 1210 1479 1268 1513
rect 1210 1445 1222 1479
rect 1256 1445 1268 1479
rect 1210 1411 1268 1445
rect 1210 1377 1222 1411
rect 1256 1377 1268 1411
rect 1210 1343 1268 1377
rect 1210 1309 1222 1343
rect 1256 1309 1268 1343
rect 1210 1275 1268 1309
rect 1210 1241 1222 1275
rect 1256 1241 1268 1275
rect 1210 1207 1268 1241
rect 1210 1173 1222 1207
rect 1256 1173 1268 1207
rect 1210 1139 1268 1173
rect 1210 1105 1222 1139
rect 1256 1105 1268 1139
rect 1210 1071 1268 1105
rect 1210 1037 1222 1071
rect 1256 1037 1268 1071
rect 1210 1003 1268 1037
rect 1210 969 1222 1003
rect 1256 969 1268 1003
rect 1210 935 1268 969
rect 1210 901 1222 935
rect 1256 901 1268 935
rect 1210 867 1268 901
rect 1210 833 1222 867
rect 1256 833 1268 867
rect 1210 799 1268 833
rect 1210 765 1222 799
rect 1256 765 1268 799
rect 1210 731 1268 765
rect 1210 697 1222 731
rect 1256 697 1268 731
rect 1210 663 1268 697
rect 1210 629 1222 663
rect 1256 629 1268 663
rect 1210 595 1268 629
rect 1210 561 1222 595
rect 1256 561 1268 595
rect 1210 527 1268 561
rect 1210 493 1222 527
rect 1256 493 1268 527
rect 1210 459 1268 493
rect 1210 425 1222 459
rect 1256 425 1268 459
rect 1210 391 1268 425
rect 1210 357 1222 391
rect 1256 357 1268 391
rect 1210 323 1268 357
rect 1210 289 1222 323
rect 1256 289 1268 323
rect 1210 255 1268 289
rect 1210 221 1222 255
rect 1256 221 1268 255
rect 1210 187 1268 221
rect 1210 153 1222 187
rect 1256 153 1268 187
rect 1210 119 1268 153
rect 1210 85 1222 119
rect 1256 85 1268 119
rect 1210 51 1268 85
rect 1210 17 1222 51
rect 1256 17 1268 51
rect 1210 -17 1268 17
rect 1210 -51 1222 -17
rect 1256 -51 1268 -17
rect 1210 -85 1268 -51
rect 1210 -119 1222 -85
rect 1256 -119 1268 -85
rect 1210 -153 1268 -119
rect 1210 -187 1222 -153
rect 1256 -187 1268 -153
rect 1210 -221 1268 -187
rect 1210 -255 1222 -221
rect 1256 -255 1268 -221
rect 1210 -289 1268 -255
rect 1210 -323 1222 -289
rect 1256 -323 1268 -289
rect 1210 -357 1268 -323
rect 1210 -391 1222 -357
rect 1256 -391 1268 -357
rect 1210 -425 1268 -391
rect 1210 -459 1222 -425
rect 1256 -459 1268 -425
rect 1210 -493 1268 -459
rect 1210 -527 1222 -493
rect 1256 -527 1268 -493
rect 1210 -561 1268 -527
rect 1210 -595 1222 -561
rect 1256 -595 1268 -561
rect 1210 -629 1268 -595
rect 1210 -663 1222 -629
rect 1256 -663 1268 -629
rect 1210 -697 1268 -663
rect 1210 -731 1222 -697
rect 1256 -731 1268 -697
rect 1210 -765 1268 -731
rect 1210 -799 1222 -765
rect 1256 -799 1268 -765
rect 1210 -833 1268 -799
rect 1210 -867 1222 -833
rect 1256 -867 1268 -833
rect 1210 -901 1268 -867
rect 1210 -935 1222 -901
rect 1256 -935 1268 -901
rect 1210 -969 1268 -935
rect 1210 -1003 1222 -969
rect 1256 -1003 1268 -969
rect 1210 -1037 1268 -1003
rect 1210 -1071 1222 -1037
rect 1256 -1071 1268 -1037
rect 1210 -1105 1268 -1071
rect 1210 -1139 1222 -1105
rect 1256 -1139 1268 -1105
rect 1210 -1173 1268 -1139
rect 1210 -1207 1222 -1173
rect 1256 -1207 1268 -1173
rect 1210 -1241 1268 -1207
rect 1210 -1275 1222 -1241
rect 1256 -1275 1268 -1241
rect 1210 -1309 1268 -1275
rect 1210 -1343 1222 -1309
rect 1256 -1343 1268 -1309
rect 1210 -1377 1268 -1343
rect 1210 -1411 1222 -1377
rect 1256 -1411 1268 -1377
rect 1210 -1445 1268 -1411
rect 1210 -1479 1222 -1445
rect 1256 -1479 1268 -1445
rect 1210 -1513 1268 -1479
rect 1210 -1547 1222 -1513
rect 1256 -1547 1268 -1513
rect 1210 -1581 1268 -1547
rect 1210 -1615 1222 -1581
rect 1256 -1615 1268 -1581
rect 1210 -1649 1268 -1615
rect 1210 -1683 1222 -1649
rect 1256 -1683 1268 -1649
rect 1210 -1717 1268 -1683
rect 1210 -1751 1222 -1717
rect 1256 -1751 1268 -1717
rect 1210 -1785 1268 -1751
rect 1210 -1819 1222 -1785
rect 1256 -1819 1268 -1785
rect 1210 -1853 1268 -1819
rect 1210 -1887 1222 -1853
rect 1256 -1887 1268 -1853
rect 1210 -1921 1268 -1887
rect 1210 -1955 1222 -1921
rect 1256 -1955 1268 -1921
rect 1210 -1989 1268 -1955
rect 1210 -2023 1222 -1989
rect 1256 -2023 1268 -1989
rect 1210 -2057 1268 -2023
rect 1210 -2091 1222 -2057
rect 1256 -2091 1268 -2057
rect 1210 -2125 1268 -2091
rect 1210 -2159 1222 -2125
rect 1256 -2159 1268 -2125
rect 1210 -2193 1268 -2159
rect 1210 -2227 1222 -2193
rect 1256 -2227 1268 -2193
rect 1210 -2261 1268 -2227
rect 1210 -2295 1222 -2261
rect 1256 -2295 1268 -2261
rect 1210 -2329 1268 -2295
rect 1210 -2363 1222 -2329
rect 1256 -2363 1268 -2329
rect 1210 -2397 1268 -2363
rect 1210 -2431 1222 -2397
rect 1256 -2431 1268 -2397
rect 1210 -2465 1268 -2431
rect 1210 -2499 1222 -2465
rect 1256 -2499 1268 -2465
rect 1210 -2533 1268 -2499
rect 1210 -2567 1222 -2533
rect 1256 -2567 1268 -2533
rect 1210 -2601 1268 -2567
rect 1210 -2635 1222 -2601
rect 1256 -2635 1268 -2601
rect 1210 -2669 1268 -2635
rect 1210 -2703 1222 -2669
rect 1256 -2703 1268 -2669
rect 1210 -2737 1268 -2703
rect 1210 -2771 1222 -2737
rect 1256 -2771 1268 -2737
rect 1210 -2805 1268 -2771
rect 1210 -2839 1222 -2805
rect 1256 -2839 1268 -2805
rect 1210 -2873 1268 -2839
rect 1210 -2907 1222 -2873
rect 1256 -2907 1268 -2873
rect 1210 -2941 1268 -2907
rect 1210 -2975 1222 -2941
rect 1256 -2975 1268 -2941
rect 1210 -3009 1268 -2975
rect 1210 -3043 1222 -3009
rect 1256 -3043 1268 -3009
rect 1210 -3077 1268 -3043
rect 1210 -3111 1222 -3077
rect 1256 -3111 1268 -3077
rect 1210 -3145 1268 -3111
rect 1210 -3179 1222 -3145
rect 1256 -3179 1268 -3145
rect 1210 -3213 1268 -3179
rect 1210 -3247 1222 -3213
rect 1256 -3247 1268 -3213
rect 1210 -3281 1268 -3247
rect 1210 -3315 1222 -3281
rect 1256 -3315 1268 -3281
rect 1210 -3349 1268 -3315
rect 1210 -3383 1222 -3349
rect 1256 -3383 1268 -3349
rect 1210 -3417 1268 -3383
rect 1210 -3451 1222 -3417
rect 1256 -3451 1268 -3417
rect 1210 -3485 1268 -3451
rect 1210 -3519 1222 -3485
rect 1256 -3519 1268 -3485
rect 1210 -3553 1268 -3519
rect 1210 -3587 1222 -3553
rect 1256 -3587 1268 -3553
rect 1210 -3621 1268 -3587
rect 1210 -3655 1222 -3621
rect 1256 -3655 1268 -3621
rect 1210 -3689 1268 -3655
rect 1210 -3723 1222 -3689
rect 1256 -3723 1268 -3689
rect 1210 -3757 1268 -3723
rect 1210 -3791 1222 -3757
rect 1256 -3791 1268 -3757
rect 1210 -3825 1268 -3791
rect 1210 -3859 1222 -3825
rect 1256 -3859 1268 -3825
rect 1210 -3893 1268 -3859
rect 1210 -3927 1222 -3893
rect 1256 -3927 1268 -3893
rect 1210 -3961 1268 -3927
rect 1210 -3995 1222 -3961
rect 1256 -3995 1268 -3961
rect 1210 -4029 1268 -3995
rect 1210 -4063 1222 -4029
rect 1256 -4063 1268 -4029
rect 1210 -4097 1268 -4063
rect 1210 -4131 1222 -4097
rect 1256 -4131 1268 -4097
rect 1210 -4165 1268 -4131
rect 1210 -4199 1222 -4165
rect 1256 -4199 1268 -4165
rect 1210 -4233 1268 -4199
rect 1210 -4267 1222 -4233
rect 1256 -4267 1268 -4233
rect 1210 -4301 1268 -4267
rect 1210 -4335 1222 -4301
rect 1256 -4335 1268 -4301
rect 1210 -4369 1268 -4335
rect 1210 -4403 1222 -4369
rect 1256 -4403 1268 -4369
rect 1210 -4437 1268 -4403
rect 1210 -4471 1222 -4437
rect 1256 -4471 1268 -4437
rect 1210 -4505 1268 -4471
rect 1210 -4539 1222 -4505
rect 1256 -4539 1268 -4505
rect 1210 -4573 1268 -4539
rect 1210 -4607 1222 -4573
rect 1256 -4607 1268 -4573
rect 1210 -4641 1268 -4607
rect 1210 -4675 1222 -4641
rect 1256 -4675 1268 -4641
rect 1210 -4709 1268 -4675
rect 1210 -4743 1222 -4709
rect 1256 -4743 1268 -4709
rect 1210 -4777 1268 -4743
rect 1210 -4811 1222 -4777
rect 1256 -4811 1268 -4777
rect 1210 -4845 1268 -4811
rect 1210 -4879 1222 -4845
rect 1256 -4879 1268 -4845
rect 1210 -4913 1268 -4879
rect 1210 -4947 1222 -4913
rect 1256 -4947 1268 -4913
rect 1210 -4981 1268 -4947
rect 1210 -5015 1222 -4981
rect 1256 -5015 1268 -4981
rect 1210 -5049 1268 -5015
rect 1210 -5083 1222 -5049
rect 1256 -5083 1268 -5049
rect 1210 -5117 1268 -5083
rect 1210 -5151 1222 -5117
rect 1256 -5151 1268 -5117
rect 1210 -5185 1268 -5151
rect 1210 -5219 1222 -5185
rect 1256 -5219 1268 -5185
rect 1210 -5253 1268 -5219
rect 1210 -5287 1222 -5253
rect 1256 -5287 1268 -5253
rect 1210 -5321 1268 -5287
rect 1210 -5355 1222 -5321
rect 1256 -5355 1268 -5321
rect 1210 -5389 1268 -5355
rect 1210 -5423 1222 -5389
rect 1256 -5423 1268 -5389
rect 1210 -5457 1268 -5423
rect 1210 -5491 1222 -5457
rect 1256 -5491 1268 -5457
rect 1210 -5525 1268 -5491
rect 1210 -5559 1222 -5525
rect 1256 -5559 1268 -5525
rect 1210 -5593 1268 -5559
rect 1210 -5627 1222 -5593
rect 1256 -5627 1268 -5593
rect 1210 -5661 1268 -5627
rect 1210 -5695 1222 -5661
rect 1256 -5695 1268 -5661
rect 1210 -5729 1268 -5695
rect 1210 -5763 1222 -5729
rect 1256 -5763 1268 -5729
rect 1210 -5797 1268 -5763
rect 1210 -5831 1222 -5797
rect 1256 -5831 1268 -5797
rect 1210 -5865 1268 -5831
rect 1210 -5899 1222 -5865
rect 1256 -5899 1268 -5865
rect 1210 -5933 1268 -5899
rect 1210 -5967 1222 -5933
rect 1256 -5967 1268 -5933
rect 1210 -6001 1268 -5967
rect 1210 -6035 1222 -6001
rect 1256 -6035 1268 -6001
rect 1210 -6069 1268 -6035
rect 1210 -6103 1222 -6069
rect 1256 -6103 1268 -6069
rect 1210 -6137 1268 -6103
rect 1210 -6171 1222 -6137
rect 1256 -6171 1268 -6137
rect 1210 -6205 1268 -6171
rect 1210 -6239 1222 -6205
rect 1256 -6239 1268 -6205
rect 1210 -6273 1268 -6239
rect 1210 -6307 1222 -6273
rect 1256 -6307 1268 -6273
rect 1210 -6341 1268 -6307
rect 1210 -6375 1222 -6341
rect 1256 -6375 1268 -6341
rect 1210 -6409 1268 -6375
rect 1210 -6443 1222 -6409
rect 1256 -6443 1268 -6409
rect 1210 -6477 1268 -6443
rect 1210 -6511 1222 -6477
rect 1256 -6511 1268 -6477
rect 1210 -6545 1268 -6511
rect 1210 -6579 1222 -6545
rect 1256 -6579 1268 -6545
rect 1210 -6613 1268 -6579
rect 1210 -6647 1222 -6613
rect 1256 -6647 1268 -6613
rect 1210 -6681 1268 -6647
rect 1210 -6715 1222 -6681
rect 1256 -6715 1268 -6681
rect 1210 -6749 1268 -6715
rect 1210 -6783 1222 -6749
rect 1256 -6783 1268 -6749
rect 1210 -6817 1268 -6783
rect 1210 -6851 1222 -6817
rect 1256 -6851 1268 -6817
rect 1210 -6885 1268 -6851
rect 1210 -6919 1222 -6885
rect 1256 -6919 1268 -6885
rect 1210 -6953 1268 -6919
rect 1210 -6987 1222 -6953
rect 1256 -6987 1268 -6953
rect 1210 -7021 1268 -6987
rect 1210 -7055 1222 -7021
rect 1256 -7055 1268 -7021
rect 1210 -7089 1268 -7055
rect 1210 -7123 1222 -7089
rect 1256 -7123 1268 -7089
rect 1210 -7157 1268 -7123
rect 1210 -7191 1222 -7157
rect 1256 -7191 1268 -7157
rect 1210 -7225 1268 -7191
rect 1210 -7259 1222 -7225
rect 1256 -7259 1268 -7225
rect 1210 -7293 1268 -7259
rect 1210 -7327 1222 -7293
rect 1256 -7327 1268 -7293
rect 1210 -7361 1268 -7327
rect 1210 -7395 1222 -7361
rect 1256 -7395 1268 -7361
rect 1210 -7429 1268 -7395
rect 1210 -7463 1222 -7429
rect 1256 -7463 1268 -7429
rect 1210 -7497 1268 -7463
rect 1210 -7531 1222 -7497
rect 1256 -7531 1268 -7497
rect 1210 -7565 1268 -7531
rect 1210 -7599 1222 -7565
rect 1256 -7599 1268 -7565
rect 1210 -7633 1268 -7599
rect 1210 -7667 1222 -7633
rect 1256 -7667 1268 -7633
rect 1210 -7701 1268 -7667
rect 1210 -7735 1222 -7701
rect 1256 -7735 1268 -7701
rect 1210 -7769 1268 -7735
rect 1210 -7803 1222 -7769
rect 1256 -7803 1268 -7769
rect 1210 -7837 1268 -7803
rect 1210 -7871 1222 -7837
rect 1256 -7871 1268 -7837
rect 1210 -7905 1268 -7871
rect 1210 -7939 1222 -7905
rect 1256 -7939 1268 -7905
rect 1210 -7973 1268 -7939
rect 1210 -8007 1222 -7973
rect 1256 -8007 1268 -7973
rect 1210 -8041 1268 -8007
rect 1210 -8075 1222 -8041
rect 1256 -8075 1268 -8041
rect 1210 -8109 1268 -8075
rect 1210 -8143 1222 -8109
rect 1256 -8143 1268 -8109
rect 1210 -8177 1268 -8143
rect 1210 -8211 1222 -8177
rect 1256 -8211 1268 -8177
rect 1210 -8245 1268 -8211
rect 1210 -8279 1222 -8245
rect 1256 -8279 1268 -8245
rect 1210 -8313 1268 -8279
rect 1210 -8347 1222 -8313
rect 1256 -8347 1268 -8313
rect 1210 -8381 1268 -8347
rect 1210 -8415 1222 -8381
rect 1256 -8415 1268 -8381
rect 1210 -8449 1268 -8415
rect 1210 -8483 1222 -8449
rect 1256 -8483 1268 -8449
rect 1210 -8517 1268 -8483
rect 1210 -8551 1222 -8517
rect 1256 -8551 1268 -8517
rect 1210 -8585 1268 -8551
rect 1210 -8619 1222 -8585
rect 1256 -8619 1268 -8585
rect 1210 -8653 1268 -8619
rect 1210 -8687 1222 -8653
rect 1256 -8687 1268 -8653
rect 1210 -8721 1268 -8687
rect 1210 -8755 1222 -8721
rect 1256 -8755 1268 -8721
rect 1210 -8789 1268 -8755
rect 1210 -8823 1222 -8789
rect 1256 -8823 1268 -8789
rect 1210 -8857 1268 -8823
rect 1210 -8891 1222 -8857
rect 1256 -8891 1268 -8857
rect 1210 -8925 1268 -8891
rect 1210 -8959 1222 -8925
rect 1256 -8959 1268 -8925
rect 1210 -8993 1268 -8959
rect 1210 -9027 1222 -8993
rect 1256 -9027 1268 -8993
rect 1210 -9061 1268 -9027
rect 1210 -9095 1222 -9061
rect 1256 -9095 1268 -9061
rect 1210 -9129 1268 -9095
rect 1210 -9163 1222 -9129
rect 1256 -9163 1268 -9129
rect 1210 -9197 1268 -9163
rect 1210 -9231 1222 -9197
rect 1256 -9231 1268 -9197
rect 1210 -9265 1268 -9231
rect 1210 -9299 1222 -9265
rect 1256 -9299 1268 -9265
rect 1210 -9333 1268 -9299
rect 1210 -9367 1222 -9333
rect 1256 -9367 1268 -9333
rect 1210 -9401 1268 -9367
rect 1210 -9435 1222 -9401
rect 1256 -9435 1268 -9401
rect 1210 -9469 1268 -9435
rect 1210 -9503 1222 -9469
rect 1256 -9503 1268 -9469
rect 1210 -9537 1268 -9503
rect 1210 -9571 1222 -9537
rect 1256 -9571 1268 -9537
rect 1210 -9600 1268 -9571
rect 1328 9571 1386 9600
rect 1328 9537 1340 9571
rect 1374 9537 1386 9571
rect 1328 9503 1386 9537
rect 1328 9469 1340 9503
rect 1374 9469 1386 9503
rect 1328 9435 1386 9469
rect 1328 9401 1340 9435
rect 1374 9401 1386 9435
rect 1328 9367 1386 9401
rect 1328 9333 1340 9367
rect 1374 9333 1386 9367
rect 1328 9299 1386 9333
rect 1328 9265 1340 9299
rect 1374 9265 1386 9299
rect 1328 9231 1386 9265
rect 1328 9197 1340 9231
rect 1374 9197 1386 9231
rect 1328 9163 1386 9197
rect 1328 9129 1340 9163
rect 1374 9129 1386 9163
rect 1328 9095 1386 9129
rect 1328 9061 1340 9095
rect 1374 9061 1386 9095
rect 1328 9027 1386 9061
rect 1328 8993 1340 9027
rect 1374 8993 1386 9027
rect 1328 8959 1386 8993
rect 1328 8925 1340 8959
rect 1374 8925 1386 8959
rect 1328 8891 1386 8925
rect 1328 8857 1340 8891
rect 1374 8857 1386 8891
rect 1328 8823 1386 8857
rect 1328 8789 1340 8823
rect 1374 8789 1386 8823
rect 1328 8755 1386 8789
rect 1328 8721 1340 8755
rect 1374 8721 1386 8755
rect 1328 8687 1386 8721
rect 1328 8653 1340 8687
rect 1374 8653 1386 8687
rect 1328 8619 1386 8653
rect 1328 8585 1340 8619
rect 1374 8585 1386 8619
rect 1328 8551 1386 8585
rect 1328 8517 1340 8551
rect 1374 8517 1386 8551
rect 1328 8483 1386 8517
rect 1328 8449 1340 8483
rect 1374 8449 1386 8483
rect 1328 8415 1386 8449
rect 1328 8381 1340 8415
rect 1374 8381 1386 8415
rect 1328 8347 1386 8381
rect 1328 8313 1340 8347
rect 1374 8313 1386 8347
rect 1328 8279 1386 8313
rect 1328 8245 1340 8279
rect 1374 8245 1386 8279
rect 1328 8211 1386 8245
rect 1328 8177 1340 8211
rect 1374 8177 1386 8211
rect 1328 8143 1386 8177
rect 1328 8109 1340 8143
rect 1374 8109 1386 8143
rect 1328 8075 1386 8109
rect 1328 8041 1340 8075
rect 1374 8041 1386 8075
rect 1328 8007 1386 8041
rect 1328 7973 1340 8007
rect 1374 7973 1386 8007
rect 1328 7939 1386 7973
rect 1328 7905 1340 7939
rect 1374 7905 1386 7939
rect 1328 7871 1386 7905
rect 1328 7837 1340 7871
rect 1374 7837 1386 7871
rect 1328 7803 1386 7837
rect 1328 7769 1340 7803
rect 1374 7769 1386 7803
rect 1328 7735 1386 7769
rect 1328 7701 1340 7735
rect 1374 7701 1386 7735
rect 1328 7667 1386 7701
rect 1328 7633 1340 7667
rect 1374 7633 1386 7667
rect 1328 7599 1386 7633
rect 1328 7565 1340 7599
rect 1374 7565 1386 7599
rect 1328 7531 1386 7565
rect 1328 7497 1340 7531
rect 1374 7497 1386 7531
rect 1328 7463 1386 7497
rect 1328 7429 1340 7463
rect 1374 7429 1386 7463
rect 1328 7395 1386 7429
rect 1328 7361 1340 7395
rect 1374 7361 1386 7395
rect 1328 7327 1386 7361
rect 1328 7293 1340 7327
rect 1374 7293 1386 7327
rect 1328 7259 1386 7293
rect 1328 7225 1340 7259
rect 1374 7225 1386 7259
rect 1328 7191 1386 7225
rect 1328 7157 1340 7191
rect 1374 7157 1386 7191
rect 1328 7123 1386 7157
rect 1328 7089 1340 7123
rect 1374 7089 1386 7123
rect 1328 7055 1386 7089
rect 1328 7021 1340 7055
rect 1374 7021 1386 7055
rect 1328 6987 1386 7021
rect 1328 6953 1340 6987
rect 1374 6953 1386 6987
rect 1328 6919 1386 6953
rect 1328 6885 1340 6919
rect 1374 6885 1386 6919
rect 1328 6851 1386 6885
rect 1328 6817 1340 6851
rect 1374 6817 1386 6851
rect 1328 6783 1386 6817
rect 1328 6749 1340 6783
rect 1374 6749 1386 6783
rect 1328 6715 1386 6749
rect 1328 6681 1340 6715
rect 1374 6681 1386 6715
rect 1328 6647 1386 6681
rect 1328 6613 1340 6647
rect 1374 6613 1386 6647
rect 1328 6579 1386 6613
rect 1328 6545 1340 6579
rect 1374 6545 1386 6579
rect 1328 6511 1386 6545
rect 1328 6477 1340 6511
rect 1374 6477 1386 6511
rect 1328 6443 1386 6477
rect 1328 6409 1340 6443
rect 1374 6409 1386 6443
rect 1328 6375 1386 6409
rect 1328 6341 1340 6375
rect 1374 6341 1386 6375
rect 1328 6307 1386 6341
rect 1328 6273 1340 6307
rect 1374 6273 1386 6307
rect 1328 6239 1386 6273
rect 1328 6205 1340 6239
rect 1374 6205 1386 6239
rect 1328 6171 1386 6205
rect 1328 6137 1340 6171
rect 1374 6137 1386 6171
rect 1328 6103 1386 6137
rect 1328 6069 1340 6103
rect 1374 6069 1386 6103
rect 1328 6035 1386 6069
rect 1328 6001 1340 6035
rect 1374 6001 1386 6035
rect 1328 5967 1386 6001
rect 1328 5933 1340 5967
rect 1374 5933 1386 5967
rect 1328 5899 1386 5933
rect 1328 5865 1340 5899
rect 1374 5865 1386 5899
rect 1328 5831 1386 5865
rect 1328 5797 1340 5831
rect 1374 5797 1386 5831
rect 1328 5763 1386 5797
rect 1328 5729 1340 5763
rect 1374 5729 1386 5763
rect 1328 5695 1386 5729
rect 1328 5661 1340 5695
rect 1374 5661 1386 5695
rect 1328 5627 1386 5661
rect 1328 5593 1340 5627
rect 1374 5593 1386 5627
rect 1328 5559 1386 5593
rect 1328 5525 1340 5559
rect 1374 5525 1386 5559
rect 1328 5491 1386 5525
rect 1328 5457 1340 5491
rect 1374 5457 1386 5491
rect 1328 5423 1386 5457
rect 1328 5389 1340 5423
rect 1374 5389 1386 5423
rect 1328 5355 1386 5389
rect 1328 5321 1340 5355
rect 1374 5321 1386 5355
rect 1328 5287 1386 5321
rect 1328 5253 1340 5287
rect 1374 5253 1386 5287
rect 1328 5219 1386 5253
rect 1328 5185 1340 5219
rect 1374 5185 1386 5219
rect 1328 5151 1386 5185
rect 1328 5117 1340 5151
rect 1374 5117 1386 5151
rect 1328 5083 1386 5117
rect 1328 5049 1340 5083
rect 1374 5049 1386 5083
rect 1328 5015 1386 5049
rect 1328 4981 1340 5015
rect 1374 4981 1386 5015
rect 1328 4947 1386 4981
rect 1328 4913 1340 4947
rect 1374 4913 1386 4947
rect 1328 4879 1386 4913
rect 1328 4845 1340 4879
rect 1374 4845 1386 4879
rect 1328 4811 1386 4845
rect 1328 4777 1340 4811
rect 1374 4777 1386 4811
rect 1328 4743 1386 4777
rect 1328 4709 1340 4743
rect 1374 4709 1386 4743
rect 1328 4675 1386 4709
rect 1328 4641 1340 4675
rect 1374 4641 1386 4675
rect 1328 4607 1386 4641
rect 1328 4573 1340 4607
rect 1374 4573 1386 4607
rect 1328 4539 1386 4573
rect 1328 4505 1340 4539
rect 1374 4505 1386 4539
rect 1328 4471 1386 4505
rect 1328 4437 1340 4471
rect 1374 4437 1386 4471
rect 1328 4403 1386 4437
rect 1328 4369 1340 4403
rect 1374 4369 1386 4403
rect 1328 4335 1386 4369
rect 1328 4301 1340 4335
rect 1374 4301 1386 4335
rect 1328 4267 1386 4301
rect 1328 4233 1340 4267
rect 1374 4233 1386 4267
rect 1328 4199 1386 4233
rect 1328 4165 1340 4199
rect 1374 4165 1386 4199
rect 1328 4131 1386 4165
rect 1328 4097 1340 4131
rect 1374 4097 1386 4131
rect 1328 4063 1386 4097
rect 1328 4029 1340 4063
rect 1374 4029 1386 4063
rect 1328 3995 1386 4029
rect 1328 3961 1340 3995
rect 1374 3961 1386 3995
rect 1328 3927 1386 3961
rect 1328 3893 1340 3927
rect 1374 3893 1386 3927
rect 1328 3859 1386 3893
rect 1328 3825 1340 3859
rect 1374 3825 1386 3859
rect 1328 3791 1386 3825
rect 1328 3757 1340 3791
rect 1374 3757 1386 3791
rect 1328 3723 1386 3757
rect 1328 3689 1340 3723
rect 1374 3689 1386 3723
rect 1328 3655 1386 3689
rect 1328 3621 1340 3655
rect 1374 3621 1386 3655
rect 1328 3587 1386 3621
rect 1328 3553 1340 3587
rect 1374 3553 1386 3587
rect 1328 3519 1386 3553
rect 1328 3485 1340 3519
rect 1374 3485 1386 3519
rect 1328 3451 1386 3485
rect 1328 3417 1340 3451
rect 1374 3417 1386 3451
rect 1328 3383 1386 3417
rect 1328 3349 1340 3383
rect 1374 3349 1386 3383
rect 1328 3315 1386 3349
rect 1328 3281 1340 3315
rect 1374 3281 1386 3315
rect 1328 3247 1386 3281
rect 1328 3213 1340 3247
rect 1374 3213 1386 3247
rect 1328 3179 1386 3213
rect 1328 3145 1340 3179
rect 1374 3145 1386 3179
rect 1328 3111 1386 3145
rect 1328 3077 1340 3111
rect 1374 3077 1386 3111
rect 1328 3043 1386 3077
rect 1328 3009 1340 3043
rect 1374 3009 1386 3043
rect 1328 2975 1386 3009
rect 1328 2941 1340 2975
rect 1374 2941 1386 2975
rect 1328 2907 1386 2941
rect 1328 2873 1340 2907
rect 1374 2873 1386 2907
rect 1328 2839 1386 2873
rect 1328 2805 1340 2839
rect 1374 2805 1386 2839
rect 1328 2771 1386 2805
rect 1328 2737 1340 2771
rect 1374 2737 1386 2771
rect 1328 2703 1386 2737
rect 1328 2669 1340 2703
rect 1374 2669 1386 2703
rect 1328 2635 1386 2669
rect 1328 2601 1340 2635
rect 1374 2601 1386 2635
rect 1328 2567 1386 2601
rect 1328 2533 1340 2567
rect 1374 2533 1386 2567
rect 1328 2499 1386 2533
rect 1328 2465 1340 2499
rect 1374 2465 1386 2499
rect 1328 2431 1386 2465
rect 1328 2397 1340 2431
rect 1374 2397 1386 2431
rect 1328 2363 1386 2397
rect 1328 2329 1340 2363
rect 1374 2329 1386 2363
rect 1328 2295 1386 2329
rect 1328 2261 1340 2295
rect 1374 2261 1386 2295
rect 1328 2227 1386 2261
rect 1328 2193 1340 2227
rect 1374 2193 1386 2227
rect 1328 2159 1386 2193
rect 1328 2125 1340 2159
rect 1374 2125 1386 2159
rect 1328 2091 1386 2125
rect 1328 2057 1340 2091
rect 1374 2057 1386 2091
rect 1328 2023 1386 2057
rect 1328 1989 1340 2023
rect 1374 1989 1386 2023
rect 1328 1955 1386 1989
rect 1328 1921 1340 1955
rect 1374 1921 1386 1955
rect 1328 1887 1386 1921
rect 1328 1853 1340 1887
rect 1374 1853 1386 1887
rect 1328 1819 1386 1853
rect 1328 1785 1340 1819
rect 1374 1785 1386 1819
rect 1328 1751 1386 1785
rect 1328 1717 1340 1751
rect 1374 1717 1386 1751
rect 1328 1683 1386 1717
rect 1328 1649 1340 1683
rect 1374 1649 1386 1683
rect 1328 1615 1386 1649
rect 1328 1581 1340 1615
rect 1374 1581 1386 1615
rect 1328 1547 1386 1581
rect 1328 1513 1340 1547
rect 1374 1513 1386 1547
rect 1328 1479 1386 1513
rect 1328 1445 1340 1479
rect 1374 1445 1386 1479
rect 1328 1411 1386 1445
rect 1328 1377 1340 1411
rect 1374 1377 1386 1411
rect 1328 1343 1386 1377
rect 1328 1309 1340 1343
rect 1374 1309 1386 1343
rect 1328 1275 1386 1309
rect 1328 1241 1340 1275
rect 1374 1241 1386 1275
rect 1328 1207 1386 1241
rect 1328 1173 1340 1207
rect 1374 1173 1386 1207
rect 1328 1139 1386 1173
rect 1328 1105 1340 1139
rect 1374 1105 1386 1139
rect 1328 1071 1386 1105
rect 1328 1037 1340 1071
rect 1374 1037 1386 1071
rect 1328 1003 1386 1037
rect 1328 969 1340 1003
rect 1374 969 1386 1003
rect 1328 935 1386 969
rect 1328 901 1340 935
rect 1374 901 1386 935
rect 1328 867 1386 901
rect 1328 833 1340 867
rect 1374 833 1386 867
rect 1328 799 1386 833
rect 1328 765 1340 799
rect 1374 765 1386 799
rect 1328 731 1386 765
rect 1328 697 1340 731
rect 1374 697 1386 731
rect 1328 663 1386 697
rect 1328 629 1340 663
rect 1374 629 1386 663
rect 1328 595 1386 629
rect 1328 561 1340 595
rect 1374 561 1386 595
rect 1328 527 1386 561
rect 1328 493 1340 527
rect 1374 493 1386 527
rect 1328 459 1386 493
rect 1328 425 1340 459
rect 1374 425 1386 459
rect 1328 391 1386 425
rect 1328 357 1340 391
rect 1374 357 1386 391
rect 1328 323 1386 357
rect 1328 289 1340 323
rect 1374 289 1386 323
rect 1328 255 1386 289
rect 1328 221 1340 255
rect 1374 221 1386 255
rect 1328 187 1386 221
rect 1328 153 1340 187
rect 1374 153 1386 187
rect 1328 119 1386 153
rect 1328 85 1340 119
rect 1374 85 1386 119
rect 1328 51 1386 85
rect 1328 17 1340 51
rect 1374 17 1386 51
rect 1328 -17 1386 17
rect 1328 -51 1340 -17
rect 1374 -51 1386 -17
rect 1328 -85 1386 -51
rect 1328 -119 1340 -85
rect 1374 -119 1386 -85
rect 1328 -153 1386 -119
rect 1328 -187 1340 -153
rect 1374 -187 1386 -153
rect 1328 -221 1386 -187
rect 1328 -255 1340 -221
rect 1374 -255 1386 -221
rect 1328 -289 1386 -255
rect 1328 -323 1340 -289
rect 1374 -323 1386 -289
rect 1328 -357 1386 -323
rect 1328 -391 1340 -357
rect 1374 -391 1386 -357
rect 1328 -425 1386 -391
rect 1328 -459 1340 -425
rect 1374 -459 1386 -425
rect 1328 -493 1386 -459
rect 1328 -527 1340 -493
rect 1374 -527 1386 -493
rect 1328 -561 1386 -527
rect 1328 -595 1340 -561
rect 1374 -595 1386 -561
rect 1328 -629 1386 -595
rect 1328 -663 1340 -629
rect 1374 -663 1386 -629
rect 1328 -697 1386 -663
rect 1328 -731 1340 -697
rect 1374 -731 1386 -697
rect 1328 -765 1386 -731
rect 1328 -799 1340 -765
rect 1374 -799 1386 -765
rect 1328 -833 1386 -799
rect 1328 -867 1340 -833
rect 1374 -867 1386 -833
rect 1328 -901 1386 -867
rect 1328 -935 1340 -901
rect 1374 -935 1386 -901
rect 1328 -969 1386 -935
rect 1328 -1003 1340 -969
rect 1374 -1003 1386 -969
rect 1328 -1037 1386 -1003
rect 1328 -1071 1340 -1037
rect 1374 -1071 1386 -1037
rect 1328 -1105 1386 -1071
rect 1328 -1139 1340 -1105
rect 1374 -1139 1386 -1105
rect 1328 -1173 1386 -1139
rect 1328 -1207 1340 -1173
rect 1374 -1207 1386 -1173
rect 1328 -1241 1386 -1207
rect 1328 -1275 1340 -1241
rect 1374 -1275 1386 -1241
rect 1328 -1309 1386 -1275
rect 1328 -1343 1340 -1309
rect 1374 -1343 1386 -1309
rect 1328 -1377 1386 -1343
rect 1328 -1411 1340 -1377
rect 1374 -1411 1386 -1377
rect 1328 -1445 1386 -1411
rect 1328 -1479 1340 -1445
rect 1374 -1479 1386 -1445
rect 1328 -1513 1386 -1479
rect 1328 -1547 1340 -1513
rect 1374 -1547 1386 -1513
rect 1328 -1581 1386 -1547
rect 1328 -1615 1340 -1581
rect 1374 -1615 1386 -1581
rect 1328 -1649 1386 -1615
rect 1328 -1683 1340 -1649
rect 1374 -1683 1386 -1649
rect 1328 -1717 1386 -1683
rect 1328 -1751 1340 -1717
rect 1374 -1751 1386 -1717
rect 1328 -1785 1386 -1751
rect 1328 -1819 1340 -1785
rect 1374 -1819 1386 -1785
rect 1328 -1853 1386 -1819
rect 1328 -1887 1340 -1853
rect 1374 -1887 1386 -1853
rect 1328 -1921 1386 -1887
rect 1328 -1955 1340 -1921
rect 1374 -1955 1386 -1921
rect 1328 -1989 1386 -1955
rect 1328 -2023 1340 -1989
rect 1374 -2023 1386 -1989
rect 1328 -2057 1386 -2023
rect 1328 -2091 1340 -2057
rect 1374 -2091 1386 -2057
rect 1328 -2125 1386 -2091
rect 1328 -2159 1340 -2125
rect 1374 -2159 1386 -2125
rect 1328 -2193 1386 -2159
rect 1328 -2227 1340 -2193
rect 1374 -2227 1386 -2193
rect 1328 -2261 1386 -2227
rect 1328 -2295 1340 -2261
rect 1374 -2295 1386 -2261
rect 1328 -2329 1386 -2295
rect 1328 -2363 1340 -2329
rect 1374 -2363 1386 -2329
rect 1328 -2397 1386 -2363
rect 1328 -2431 1340 -2397
rect 1374 -2431 1386 -2397
rect 1328 -2465 1386 -2431
rect 1328 -2499 1340 -2465
rect 1374 -2499 1386 -2465
rect 1328 -2533 1386 -2499
rect 1328 -2567 1340 -2533
rect 1374 -2567 1386 -2533
rect 1328 -2601 1386 -2567
rect 1328 -2635 1340 -2601
rect 1374 -2635 1386 -2601
rect 1328 -2669 1386 -2635
rect 1328 -2703 1340 -2669
rect 1374 -2703 1386 -2669
rect 1328 -2737 1386 -2703
rect 1328 -2771 1340 -2737
rect 1374 -2771 1386 -2737
rect 1328 -2805 1386 -2771
rect 1328 -2839 1340 -2805
rect 1374 -2839 1386 -2805
rect 1328 -2873 1386 -2839
rect 1328 -2907 1340 -2873
rect 1374 -2907 1386 -2873
rect 1328 -2941 1386 -2907
rect 1328 -2975 1340 -2941
rect 1374 -2975 1386 -2941
rect 1328 -3009 1386 -2975
rect 1328 -3043 1340 -3009
rect 1374 -3043 1386 -3009
rect 1328 -3077 1386 -3043
rect 1328 -3111 1340 -3077
rect 1374 -3111 1386 -3077
rect 1328 -3145 1386 -3111
rect 1328 -3179 1340 -3145
rect 1374 -3179 1386 -3145
rect 1328 -3213 1386 -3179
rect 1328 -3247 1340 -3213
rect 1374 -3247 1386 -3213
rect 1328 -3281 1386 -3247
rect 1328 -3315 1340 -3281
rect 1374 -3315 1386 -3281
rect 1328 -3349 1386 -3315
rect 1328 -3383 1340 -3349
rect 1374 -3383 1386 -3349
rect 1328 -3417 1386 -3383
rect 1328 -3451 1340 -3417
rect 1374 -3451 1386 -3417
rect 1328 -3485 1386 -3451
rect 1328 -3519 1340 -3485
rect 1374 -3519 1386 -3485
rect 1328 -3553 1386 -3519
rect 1328 -3587 1340 -3553
rect 1374 -3587 1386 -3553
rect 1328 -3621 1386 -3587
rect 1328 -3655 1340 -3621
rect 1374 -3655 1386 -3621
rect 1328 -3689 1386 -3655
rect 1328 -3723 1340 -3689
rect 1374 -3723 1386 -3689
rect 1328 -3757 1386 -3723
rect 1328 -3791 1340 -3757
rect 1374 -3791 1386 -3757
rect 1328 -3825 1386 -3791
rect 1328 -3859 1340 -3825
rect 1374 -3859 1386 -3825
rect 1328 -3893 1386 -3859
rect 1328 -3927 1340 -3893
rect 1374 -3927 1386 -3893
rect 1328 -3961 1386 -3927
rect 1328 -3995 1340 -3961
rect 1374 -3995 1386 -3961
rect 1328 -4029 1386 -3995
rect 1328 -4063 1340 -4029
rect 1374 -4063 1386 -4029
rect 1328 -4097 1386 -4063
rect 1328 -4131 1340 -4097
rect 1374 -4131 1386 -4097
rect 1328 -4165 1386 -4131
rect 1328 -4199 1340 -4165
rect 1374 -4199 1386 -4165
rect 1328 -4233 1386 -4199
rect 1328 -4267 1340 -4233
rect 1374 -4267 1386 -4233
rect 1328 -4301 1386 -4267
rect 1328 -4335 1340 -4301
rect 1374 -4335 1386 -4301
rect 1328 -4369 1386 -4335
rect 1328 -4403 1340 -4369
rect 1374 -4403 1386 -4369
rect 1328 -4437 1386 -4403
rect 1328 -4471 1340 -4437
rect 1374 -4471 1386 -4437
rect 1328 -4505 1386 -4471
rect 1328 -4539 1340 -4505
rect 1374 -4539 1386 -4505
rect 1328 -4573 1386 -4539
rect 1328 -4607 1340 -4573
rect 1374 -4607 1386 -4573
rect 1328 -4641 1386 -4607
rect 1328 -4675 1340 -4641
rect 1374 -4675 1386 -4641
rect 1328 -4709 1386 -4675
rect 1328 -4743 1340 -4709
rect 1374 -4743 1386 -4709
rect 1328 -4777 1386 -4743
rect 1328 -4811 1340 -4777
rect 1374 -4811 1386 -4777
rect 1328 -4845 1386 -4811
rect 1328 -4879 1340 -4845
rect 1374 -4879 1386 -4845
rect 1328 -4913 1386 -4879
rect 1328 -4947 1340 -4913
rect 1374 -4947 1386 -4913
rect 1328 -4981 1386 -4947
rect 1328 -5015 1340 -4981
rect 1374 -5015 1386 -4981
rect 1328 -5049 1386 -5015
rect 1328 -5083 1340 -5049
rect 1374 -5083 1386 -5049
rect 1328 -5117 1386 -5083
rect 1328 -5151 1340 -5117
rect 1374 -5151 1386 -5117
rect 1328 -5185 1386 -5151
rect 1328 -5219 1340 -5185
rect 1374 -5219 1386 -5185
rect 1328 -5253 1386 -5219
rect 1328 -5287 1340 -5253
rect 1374 -5287 1386 -5253
rect 1328 -5321 1386 -5287
rect 1328 -5355 1340 -5321
rect 1374 -5355 1386 -5321
rect 1328 -5389 1386 -5355
rect 1328 -5423 1340 -5389
rect 1374 -5423 1386 -5389
rect 1328 -5457 1386 -5423
rect 1328 -5491 1340 -5457
rect 1374 -5491 1386 -5457
rect 1328 -5525 1386 -5491
rect 1328 -5559 1340 -5525
rect 1374 -5559 1386 -5525
rect 1328 -5593 1386 -5559
rect 1328 -5627 1340 -5593
rect 1374 -5627 1386 -5593
rect 1328 -5661 1386 -5627
rect 1328 -5695 1340 -5661
rect 1374 -5695 1386 -5661
rect 1328 -5729 1386 -5695
rect 1328 -5763 1340 -5729
rect 1374 -5763 1386 -5729
rect 1328 -5797 1386 -5763
rect 1328 -5831 1340 -5797
rect 1374 -5831 1386 -5797
rect 1328 -5865 1386 -5831
rect 1328 -5899 1340 -5865
rect 1374 -5899 1386 -5865
rect 1328 -5933 1386 -5899
rect 1328 -5967 1340 -5933
rect 1374 -5967 1386 -5933
rect 1328 -6001 1386 -5967
rect 1328 -6035 1340 -6001
rect 1374 -6035 1386 -6001
rect 1328 -6069 1386 -6035
rect 1328 -6103 1340 -6069
rect 1374 -6103 1386 -6069
rect 1328 -6137 1386 -6103
rect 1328 -6171 1340 -6137
rect 1374 -6171 1386 -6137
rect 1328 -6205 1386 -6171
rect 1328 -6239 1340 -6205
rect 1374 -6239 1386 -6205
rect 1328 -6273 1386 -6239
rect 1328 -6307 1340 -6273
rect 1374 -6307 1386 -6273
rect 1328 -6341 1386 -6307
rect 1328 -6375 1340 -6341
rect 1374 -6375 1386 -6341
rect 1328 -6409 1386 -6375
rect 1328 -6443 1340 -6409
rect 1374 -6443 1386 -6409
rect 1328 -6477 1386 -6443
rect 1328 -6511 1340 -6477
rect 1374 -6511 1386 -6477
rect 1328 -6545 1386 -6511
rect 1328 -6579 1340 -6545
rect 1374 -6579 1386 -6545
rect 1328 -6613 1386 -6579
rect 1328 -6647 1340 -6613
rect 1374 -6647 1386 -6613
rect 1328 -6681 1386 -6647
rect 1328 -6715 1340 -6681
rect 1374 -6715 1386 -6681
rect 1328 -6749 1386 -6715
rect 1328 -6783 1340 -6749
rect 1374 -6783 1386 -6749
rect 1328 -6817 1386 -6783
rect 1328 -6851 1340 -6817
rect 1374 -6851 1386 -6817
rect 1328 -6885 1386 -6851
rect 1328 -6919 1340 -6885
rect 1374 -6919 1386 -6885
rect 1328 -6953 1386 -6919
rect 1328 -6987 1340 -6953
rect 1374 -6987 1386 -6953
rect 1328 -7021 1386 -6987
rect 1328 -7055 1340 -7021
rect 1374 -7055 1386 -7021
rect 1328 -7089 1386 -7055
rect 1328 -7123 1340 -7089
rect 1374 -7123 1386 -7089
rect 1328 -7157 1386 -7123
rect 1328 -7191 1340 -7157
rect 1374 -7191 1386 -7157
rect 1328 -7225 1386 -7191
rect 1328 -7259 1340 -7225
rect 1374 -7259 1386 -7225
rect 1328 -7293 1386 -7259
rect 1328 -7327 1340 -7293
rect 1374 -7327 1386 -7293
rect 1328 -7361 1386 -7327
rect 1328 -7395 1340 -7361
rect 1374 -7395 1386 -7361
rect 1328 -7429 1386 -7395
rect 1328 -7463 1340 -7429
rect 1374 -7463 1386 -7429
rect 1328 -7497 1386 -7463
rect 1328 -7531 1340 -7497
rect 1374 -7531 1386 -7497
rect 1328 -7565 1386 -7531
rect 1328 -7599 1340 -7565
rect 1374 -7599 1386 -7565
rect 1328 -7633 1386 -7599
rect 1328 -7667 1340 -7633
rect 1374 -7667 1386 -7633
rect 1328 -7701 1386 -7667
rect 1328 -7735 1340 -7701
rect 1374 -7735 1386 -7701
rect 1328 -7769 1386 -7735
rect 1328 -7803 1340 -7769
rect 1374 -7803 1386 -7769
rect 1328 -7837 1386 -7803
rect 1328 -7871 1340 -7837
rect 1374 -7871 1386 -7837
rect 1328 -7905 1386 -7871
rect 1328 -7939 1340 -7905
rect 1374 -7939 1386 -7905
rect 1328 -7973 1386 -7939
rect 1328 -8007 1340 -7973
rect 1374 -8007 1386 -7973
rect 1328 -8041 1386 -8007
rect 1328 -8075 1340 -8041
rect 1374 -8075 1386 -8041
rect 1328 -8109 1386 -8075
rect 1328 -8143 1340 -8109
rect 1374 -8143 1386 -8109
rect 1328 -8177 1386 -8143
rect 1328 -8211 1340 -8177
rect 1374 -8211 1386 -8177
rect 1328 -8245 1386 -8211
rect 1328 -8279 1340 -8245
rect 1374 -8279 1386 -8245
rect 1328 -8313 1386 -8279
rect 1328 -8347 1340 -8313
rect 1374 -8347 1386 -8313
rect 1328 -8381 1386 -8347
rect 1328 -8415 1340 -8381
rect 1374 -8415 1386 -8381
rect 1328 -8449 1386 -8415
rect 1328 -8483 1340 -8449
rect 1374 -8483 1386 -8449
rect 1328 -8517 1386 -8483
rect 1328 -8551 1340 -8517
rect 1374 -8551 1386 -8517
rect 1328 -8585 1386 -8551
rect 1328 -8619 1340 -8585
rect 1374 -8619 1386 -8585
rect 1328 -8653 1386 -8619
rect 1328 -8687 1340 -8653
rect 1374 -8687 1386 -8653
rect 1328 -8721 1386 -8687
rect 1328 -8755 1340 -8721
rect 1374 -8755 1386 -8721
rect 1328 -8789 1386 -8755
rect 1328 -8823 1340 -8789
rect 1374 -8823 1386 -8789
rect 1328 -8857 1386 -8823
rect 1328 -8891 1340 -8857
rect 1374 -8891 1386 -8857
rect 1328 -8925 1386 -8891
rect 1328 -8959 1340 -8925
rect 1374 -8959 1386 -8925
rect 1328 -8993 1386 -8959
rect 1328 -9027 1340 -8993
rect 1374 -9027 1386 -8993
rect 1328 -9061 1386 -9027
rect 1328 -9095 1340 -9061
rect 1374 -9095 1386 -9061
rect 1328 -9129 1386 -9095
rect 1328 -9163 1340 -9129
rect 1374 -9163 1386 -9129
rect 1328 -9197 1386 -9163
rect 1328 -9231 1340 -9197
rect 1374 -9231 1386 -9197
rect 1328 -9265 1386 -9231
rect 1328 -9299 1340 -9265
rect 1374 -9299 1386 -9265
rect 1328 -9333 1386 -9299
rect 1328 -9367 1340 -9333
rect 1374 -9367 1386 -9333
rect 1328 -9401 1386 -9367
rect 1328 -9435 1340 -9401
rect 1374 -9435 1386 -9401
rect 1328 -9469 1386 -9435
rect 1328 -9503 1340 -9469
rect 1374 -9503 1386 -9469
rect 1328 -9537 1386 -9503
rect 1328 -9571 1340 -9537
rect 1374 -9571 1386 -9537
rect 1328 -9600 1386 -9571
rect 1446 9571 1504 9600
rect 1446 9537 1458 9571
rect 1492 9537 1504 9571
rect 1446 9503 1504 9537
rect 1446 9469 1458 9503
rect 1492 9469 1504 9503
rect 1446 9435 1504 9469
rect 1446 9401 1458 9435
rect 1492 9401 1504 9435
rect 1446 9367 1504 9401
rect 1446 9333 1458 9367
rect 1492 9333 1504 9367
rect 1446 9299 1504 9333
rect 1446 9265 1458 9299
rect 1492 9265 1504 9299
rect 1446 9231 1504 9265
rect 1446 9197 1458 9231
rect 1492 9197 1504 9231
rect 1446 9163 1504 9197
rect 1446 9129 1458 9163
rect 1492 9129 1504 9163
rect 1446 9095 1504 9129
rect 1446 9061 1458 9095
rect 1492 9061 1504 9095
rect 1446 9027 1504 9061
rect 1446 8993 1458 9027
rect 1492 8993 1504 9027
rect 1446 8959 1504 8993
rect 1446 8925 1458 8959
rect 1492 8925 1504 8959
rect 1446 8891 1504 8925
rect 1446 8857 1458 8891
rect 1492 8857 1504 8891
rect 1446 8823 1504 8857
rect 1446 8789 1458 8823
rect 1492 8789 1504 8823
rect 1446 8755 1504 8789
rect 1446 8721 1458 8755
rect 1492 8721 1504 8755
rect 1446 8687 1504 8721
rect 1446 8653 1458 8687
rect 1492 8653 1504 8687
rect 1446 8619 1504 8653
rect 1446 8585 1458 8619
rect 1492 8585 1504 8619
rect 1446 8551 1504 8585
rect 1446 8517 1458 8551
rect 1492 8517 1504 8551
rect 1446 8483 1504 8517
rect 1446 8449 1458 8483
rect 1492 8449 1504 8483
rect 1446 8415 1504 8449
rect 1446 8381 1458 8415
rect 1492 8381 1504 8415
rect 1446 8347 1504 8381
rect 1446 8313 1458 8347
rect 1492 8313 1504 8347
rect 1446 8279 1504 8313
rect 1446 8245 1458 8279
rect 1492 8245 1504 8279
rect 1446 8211 1504 8245
rect 1446 8177 1458 8211
rect 1492 8177 1504 8211
rect 1446 8143 1504 8177
rect 1446 8109 1458 8143
rect 1492 8109 1504 8143
rect 1446 8075 1504 8109
rect 1446 8041 1458 8075
rect 1492 8041 1504 8075
rect 1446 8007 1504 8041
rect 1446 7973 1458 8007
rect 1492 7973 1504 8007
rect 1446 7939 1504 7973
rect 1446 7905 1458 7939
rect 1492 7905 1504 7939
rect 1446 7871 1504 7905
rect 1446 7837 1458 7871
rect 1492 7837 1504 7871
rect 1446 7803 1504 7837
rect 1446 7769 1458 7803
rect 1492 7769 1504 7803
rect 1446 7735 1504 7769
rect 1446 7701 1458 7735
rect 1492 7701 1504 7735
rect 1446 7667 1504 7701
rect 1446 7633 1458 7667
rect 1492 7633 1504 7667
rect 1446 7599 1504 7633
rect 1446 7565 1458 7599
rect 1492 7565 1504 7599
rect 1446 7531 1504 7565
rect 1446 7497 1458 7531
rect 1492 7497 1504 7531
rect 1446 7463 1504 7497
rect 1446 7429 1458 7463
rect 1492 7429 1504 7463
rect 1446 7395 1504 7429
rect 1446 7361 1458 7395
rect 1492 7361 1504 7395
rect 1446 7327 1504 7361
rect 1446 7293 1458 7327
rect 1492 7293 1504 7327
rect 1446 7259 1504 7293
rect 1446 7225 1458 7259
rect 1492 7225 1504 7259
rect 1446 7191 1504 7225
rect 1446 7157 1458 7191
rect 1492 7157 1504 7191
rect 1446 7123 1504 7157
rect 1446 7089 1458 7123
rect 1492 7089 1504 7123
rect 1446 7055 1504 7089
rect 1446 7021 1458 7055
rect 1492 7021 1504 7055
rect 1446 6987 1504 7021
rect 1446 6953 1458 6987
rect 1492 6953 1504 6987
rect 1446 6919 1504 6953
rect 1446 6885 1458 6919
rect 1492 6885 1504 6919
rect 1446 6851 1504 6885
rect 1446 6817 1458 6851
rect 1492 6817 1504 6851
rect 1446 6783 1504 6817
rect 1446 6749 1458 6783
rect 1492 6749 1504 6783
rect 1446 6715 1504 6749
rect 1446 6681 1458 6715
rect 1492 6681 1504 6715
rect 1446 6647 1504 6681
rect 1446 6613 1458 6647
rect 1492 6613 1504 6647
rect 1446 6579 1504 6613
rect 1446 6545 1458 6579
rect 1492 6545 1504 6579
rect 1446 6511 1504 6545
rect 1446 6477 1458 6511
rect 1492 6477 1504 6511
rect 1446 6443 1504 6477
rect 1446 6409 1458 6443
rect 1492 6409 1504 6443
rect 1446 6375 1504 6409
rect 1446 6341 1458 6375
rect 1492 6341 1504 6375
rect 1446 6307 1504 6341
rect 1446 6273 1458 6307
rect 1492 6273 1504 6307
rect 1446 6239 1504 6273
rect 1446 6205 1458 6239
rect 1492 6205 1504 6239
rect 1446 6171 1504 6205
rect 1446 6137 1458 6171
rect 1492 6137 1504 6171
rect 1446 6103 1504 6137
rect 1446 6069 1458 6103
rect 1492 6069 1504 6103
rect 1446 6035 1504 6069
rect 1446 6001 1458 6035
rect 1492 6001 1504 6035
rect 1446 5967 1504 6001
rect 1446 5933 1458 5967
rect 1492 5933 1504 5967
rect 1446 5899 1504 5933
rect 1446 5865 1458 5899
rect 1492 5865 1504 5899
rect 1446 5831 1504 5865
rect 1446 5797 1458 5831
rect 1492 5797 1504 5831
rect 1446 5763 1504 5797
rect 1446 5729 1458 5763
rect 1492 5729 1504 5763
rect 1446 5695 1504 5729
rect 1446 5661 1458 5695
rect 1492 5661 1504 5695
rect 1446 5627 1504 5661
rect 1446 5593 1458 5627
rect 1492 5593 1504 5627
rect 1446 5559 1504 5593
rect 1446 5525 1458 5559
rect 1492 5525 1504 5559
rect 1446 5491 1504 5525
rect 1446 5457 1458 5491
rect 1492 5457 1504 5491
rect 1446 5423 1504 5457
rect 1446 5389 1458 5423
rect 1492 5389 1504 5423
rect 1446 5355 1504 5389
rect 1446 5321 1458 5355
rect 1492 5321 1504 5355
rect 1446 5287 1504 5321
rect 1446 5253 1458 5287
rect 1492 5253 1504 5287
rect 1446 5219 1504 5253
rect 1446 5185 1458 5219
rect 1492 5185 1504 5219
rect 1446 5151 1504 5185
rect 1446 5117 1458 5151
rect 1492 5117 1504 5151
rect 1446 5083 1504 5117
rect 1446 5049 1458 5083
rect 1492 5049 1504 5083
rect 1446 5015 1504 5049
rect 1446 4981 1458 5015
rect 1492 4981 1504 5015
rect 1446 4947 1504 4981
rect 1446 4913 1458 4947
rect 1492 4913 1504 4947
rect 1446 4879 1504 4913
rect 1446 4845 1458 4879
rect 1492 4845 1504 4879
rect 1446 4811 1504 4845
rect 1446 4777 1458 4811
rect 1492 4777 1504 4811
rect 1446 4743 1504 4777
rect 1446 4709 1458 4743
rect 1492 4709 1504 4743
rect 1446 4675 1504 4709
rect 1446 4641 1458 4675
rect 1492 4641 1504 4675
rect 1446 4607 1504 4641
rect 1446 4573 1458 4607
rect 1492 4573 1504 4607
rect 1446 4539 1504 4573
rect 1446 4505 1458 4539
rect 1492 4505 1504 4539
rect 1446 4471 1504 4505
rect 1446 4437 1458 4471
rect 1492 4437 1504 4471
rect 1446 4403 1504 4437
rect 1446 4369 1458 4403
rect 1492 4369 1504 4403
rect 1446 4335 1504 4369
rect 1446 4301 1458 4335
rect 1492 4301 1504 4335
rect 1446 4267 1504 4301
rect 1446 4233 1458 4267
rect 1492 4233 1504 4267
rect 1446 4199 1504 4233
rect 1446 4165 1458 4199
rect 1492 4165 1504 4199
rect 1446 4131 1504 4165
rect 1446 4097 1458 4131
rect 1492 4097 1504 4131
rect 1446 4063 1504 4097
rect 1446 4029 1458 4063
rect 1492 4029 1504 4063
rect 1446 3995 1504 4029
rect 1446 3961 1458 3995
rect 1492 3961 1504 3995
rect 1446 3927 1504 3961
rect 1446 3893 1458 3927
rect 1492 3893 1504 3927
rect 1446 3859 1504 3893
rect 1446 3825 1458 3859
rect 1492 3825 1504 3859
rect 1446 3791 1504 3825
rect 1446 3757 1458 3791
rect 1492 3757 1504 3791
rect 1446 3723 1504 3757
rect 1446 3689 1458 3723
rect 1492 3689 1504 3723
rect 1446 3655 1504 3689
rect 1446 3621 1458 3655
rect 1492 3621 1504 3655
rect 1446 3587 1504 3621
rect 1446 3553 1458 3587
rect 1492 3553 1504 3587
rect 1446 3519 1504 3553
rect 1446 3485 1458 3519
rect 1492 3485 1504 3519
rect 1446 3451 1504 3485
rect 1446 3417 1458 3451
rect 1492 3417 1504 3451
rect 1446 3383 1504 3417
rect 1446 3349 1458 3383
rect 1492 3349 1504 3383
rect 1446 3315 1504 3349
rect 1446 3281 1458 3315
rect 1492 3281 1504 3315
rect 1446 3247 1504 3281
rect 1446 3213 1458 3247
rect 1492 3213 1504 3247
rect 1446 3179 1504 3213
rect 1446 3145 1458 3179
rect 1492 3145 1504 3179
rect 1446 3111 1504 3145
rect 1446 3077 1458 3111
rect 1492 3077 1504 3111
rect 1446 3043 1504 3077
rect 1446 3009 1458 3043
rect 1492 3009 1504 3043
rect 1446 2975 1504 3009
rect 1446 2941 1458 2975
rect 1492 2941 1504 2975
rect 1446 2907 1504 2941
rect 1446 2873 1458 2907
rect 1492 2873 1504 2907
rect 1446 2839 1504 2873
rect 1446 2805 1458 2839
rect 1492 2805 1504 2839
rect 1446 2771 1504 2805
rect 1446 2737 1458 2771
rect 1492 2737 1504 2771
rect 1446 2703 1504 2737
rect 1446 2669 1458 2703
rect 1492 2669 1504 2703
rect 1446 2635 1504 2669
rect 1446 2601 1458 2635
rect 1492 2601 1504 2635
rect 1446 2567 1504 2601
rect 1446 2533 1458 2567
rect 1492 2533 1504 2567
rect 1446 2499 1504 2533
rect 1446 2465 1458 2499
rect 1492 2465 1504 2499
rect 1446 2431 1504 2465
rect 1446 2397 1458 2431
rect 1492 2397 1504 2431
rect 1446 2363 1504 2397
rect 1446 2329 1458 2363
rect 1492 2329 1504 2363
rect 1446 2295 1504 2329
rect 1446 2261 1458 2295
rect 1492 2261 1504 2295
rect 1446 2227 1504 2261
rect 1446 2193 1458 2227
rect 1492 2193 1504 2227
rect 1446 2159 1504 2193
rect 1446 2125 1458 2159
rect 1492 2125 1504 2159
rect 1446 2091 1504 2125
rect 1446 2057 1458 2091
rect 1492 2057 1504 2091
rect 1446 2023 1504 2057
rect 1446 1989 1458 2023
rect 1492 1989 1504 2023
rect 1446 1955 1504 1989
rect 1446 1921 1458 1955
rect 1492 1921 1504 1955
rect 1446 1887 1504 1921
rect 1446 1853 1458 1887
rect 1492 1853 1504 1887
rect 1446 1819 1504 1853
rect 1446 1785 1458 1819
rect 1492 1785 1504 1819
rect 1446 1751 1504 1785
rect 1446 1717 1458 1751
rect 1492 1717 1504 1751
rect 1446 1683 1504 1717
rect 1446 1649 1458 1683
rect 1492 1649 1504 1683
rect 1446 1615 1504 1649
rect 1446 1581 1458 1615
rect 1492 1581 1504 1615
rect 1446 1547 1504 1581
rect 1446 1513 1458 1547
rect 1492 1513 1504 1547
rect 1446 1479 1504 1513
rect 1446 1445 1458 1479
rect 1492 1445 1504 1479
rect 1446 1411 1504 1445
rect 1446 1377 1458 1411
rect 1492 1377 1504 1411
rect 1446 1343 1504 1377
rect 1446 1309 1458 1343
rect 1492 1309 1504 1343
rect 1446 1275 1504 1309
rect 1446 1241 1458 1275
rect 1492 1241 1504 1275
rect 1446 1207 1504 1241
rect 1446 1173 1458 1207
rect 1492 1173 1504 1207
rect 1446 1139 1504 1173
rect 1446 1105 1458 1139
rect 1492 1105 1504 1139
rect 1446 1071 1504 1105
rect 1446 1037 1458 1071
rect 1492 1037 1504 1071
rect 1446 1003 1504 1037
rect 1446 969 1458 1003
rect 1492 969 1504 1003
rect 1446 935 1504 969
rect 1446 901 1458 935
rect 1492 901 1504 935
rect 1446 867 1504 901
rect 1446 833 1458 867
rect 1492 833 1504 867
rect 1446 799 1504 833
rect 1446 765 1458 799
rect 1492 765 1504 799
rect 1446 731 1504 765
rect 1446 697 1458 731
rect 1492 697 1504 731
rect 1446 663 1504 697
rect 1446 629 1458 663
rect 1492 629 1504 663
rect 1446 595 1504 629
rect 1446 561 1458 595
rect 1492 561 1504 595
rect 1446 527 1504 561
rect 1446 493 1458 527
rect 1492 493 1504 527
rect 1446 459 1504 493
rect 1446 425 1458 459
rect 1492 425 1504 459
rect 1446 391 1504 425
rect 1446 357 1458 391
rect 1492 357 1504 391
rect 1446 323 1504 357
rect 1446 289 1458 323
rect 1492 289 1504 323
rect 1446 255 1504 289
rect 1446 221 1458 255
rect 1492 221 1504 255
rect 1446 187 1504 221
rect 1446 153 1458 187
rect 1492 153 1504 187
rect 1446 119 1504 153
rect 1446 85 1458 119
rect 1492 85 1504 119
rect 1446 51 1504 85
rect 1446 17 1458 51
rect 1492 17 1504 51
rect 1446 -17 1504 17
rect 1446 -51 1458 -17
rect 1492 -51 1504 -17
rect 1446 -85 1504 -51
rect 1446 -119 1458 -85
rect 1492 -119 1504 -85
rect 1446 -153 1504 -119
rect 1446 -187 1458 -153
rect 1492 -187 1504 -153
rect 1446 -221 1504 -187
rect 1446 -255 1458 -221
rect 1492 -255 1504 -221
rect 1446 -289 1504 -255
rect 1446 -323 1458 -289
rect 1492 -323 1504 -289
rect 1446 -357 1504 -323
rect 1446 -391 1458 -357
rect 1492 -391 1504 -357
rect 1446 -425 1504 -391
rect 1446 -459 1458 -425
rect 1492 -459 1504 -425
rect 1446 -493 1504 -459
rect 1446 -527 1458 -493
rect 1492 -527 1504 -493
rect 1446 -561 1504 -527
rect 1446 -595 1458 -561
rect 1492 -595 1504 -561
rect 1446 -629 1504 -595
rect 1446 -663 1458 -629
rect 1492 -663 1504 -629
rect 1446 -697 1504 -663
rect 1446 -731 1458 -697
rect 1492 -731 1504 -697
rect 1446 -765 1504 -731
rect 1446 -799 1458 -765
rect 1492 -799 1504 -765
rect 1446 -833 1504 -799
rect 1446 -867 1458 -833
rect 1492 -867 1504 -833
rect 1446 -901 1504 -867
rect 1446 -935 1458 -901
rect 1492 -935 1504 -901
rect 1446 -969 1504 -935
rect 1446 -1003 1458 -969
rect 1492 -1003 1504 -969
rect 1446 -1037 1504 -1003
rect 1446 -1071 1458 -1037
rect 1492 -1071 1504 -1037
rect 1446 -1105 1504 -1071
rect 1446 -1139 1458 -1105
rect 1492 -1139 1504 -1105
rect 1446 -1173 1504 -1139
rect 1446 -1207 1458 -1173
rect 1492 -1207 1504 -1173
rect 1446 -1241 1504 -1207
rect 1446 -1275 1458 -1241
rect 1492 -1275 1504 -1241
rect 1446 -1309 1504 -1275
rect 1446 -1343 1458 -1309
rect 1492 -1343 1504 -1309
rect 1446 -1377 1504 -1343
rect 1446 -1411 1458 -1377
rect 1492 -1411 1504 -1377
rect 1446 -1445 1504 -1411
rect 1446 -1479 1458 -1445
rect 1492 -1479 1504 -1445
rect 1446 -1513 1504 -1479
rect 1446 -1547 1458 -1513
rect 1492 -1547 1504 -1513
rect 1446 -1581 1504 -1547
rect 1446 -1615 1458 -1581
rect 1492 -1615 1504 -1581
rect 1446 -1649 1504 -1615
rect 1446 -1683 1458 -1649
rect 1492 -1683 1504 -1649
rect 1446 -1717 1504 -1683
rect 1446 -1751 1458 -1717
rect 1492 -1751 1504 -1717
rect 1446 -1785 1504 -1751
rect 1446 -1819 1458 -1785
rect 1492 -1819 1504 -1785
rect 1446 -1853 1504 -1819
rect 1446 -1887 1458 -1853
rect 1492 -1887 1504 -1853
rect 1446 -1921 1504 -1887
rect 1446 -1955 1458 -1921
rect 1492 -1955 1504 -1921
rect 1446 -1989 1504 -1955
rect 1446 -2023 1458 -1989
rect 1492 -2023 1504 -1989
rect 1446 -2057 1504 -2023
rect 1446 -2091 1458 -2057
rect 1492 -2091 1504 -2057
rect 1446 -2125 1504 -2091
rect 1446 -2159 1458 -2125
rect 1492 -2159 1504 -2125
rect 1446 -2193 1504 -2159
rect 1446 -2227 1458 -2193
rect 1492 -2227 1504 -2193
rect 1446 -2261 1504 -2227
rect 1446 -2295 1458 -2261
rect 1492 -2295 1504 -2261
rect 1446 -2329 1504 -2295
rect 1446 -2363 1458 -2329
rect 1492 -2363 1504 -2329
rect 1446 -2397 1504 -2363
rect 1446 -2431 1458 -2397
rect 1492 -2431 1504 -2397
rect 1446 -2465 1504 -2431
rect 1446 -2499 1458 -2465
rect 1492 -2499 1504 -2465
rect 1446 -2533 1504 -2499
rect 1446 -2567 1458 -2533
rect 1492 -2567 1504 -2533
rect 1446 -2601 1504 -2567
rect 1446 -2635 1458 -2601
rect 1492 -2635 1504 -2601
rect 1446 -2669 1504 -2635
rect 1446 -2703 1458 -2669
rect 1492 -2703 1504 -2669
rect 1446 -2737 1504 -2703
rect 1446 -2771 1458 -2737
rect 1492 -2771 1504 -2737
rect 1446 -2805 1504 -2771
rect 1446 -2839 1458 -2805
rect 1492 -2839 1504 -2805
rect 1446 -2873 1504 -2839
rect 1446 -2907 1458 -2873
rect 1492 -2907 1504 -2873
rect 1446 -2941 1504 -2907
rect 1446 -2975 1458 -2941
rect 1492 -2975 1504 -2941
rect 1446 -3009 1504 -2975
rect 1446 -3043 1458 -3009
rect 1492 -3043 1504 -3009
rect 1446 -3077 1504 -3043
rect 1446 -3111 1458 -3077
rect 1492 -3111 1504 -3077
rect 1446 -3145 1504 -3111
rect 1446 -3179 1458 -3145
rect 1492 -3179 1504 -3145
rect 1446 -3213 1504 -3179
rect 1446 -3247 1458 -3213
rect 1492 -3247 1504 -3213
rect 1446 -3281 1504 -3247
rect 1446 -3315 1458 -3281
rect 1492 -3315 1504 -3281
rect 1446 -3349 1504 -3315
rect 1446 -3383 1458 -3349
rect 1492 -3383 1504 -3349
rect 1446 -3417 1504 -3383
rect 1446 -3451 1458 -3417
rect 1492 -3451 1504 -3417
rect 1446 -3485 1504 -3451
rect 1446 -3519 1458 -3485
rect 1492 -3519 1504 -3485
rect 1446 -3553 1504 -3519
rect 1446 -3587 1458 -3553
rect 1492 -3587 1504 -3553
rect 1446 -3621 1504 -3587
rect 1446 -3655 1458 -3621
rect 1492 -3655 1504 -3621
rect 1446 -3689 1504 -3655
rect 1446 -3723 1458 -3689
rect 1492 -3723 1504 -3689
rect 1446 -3757 1504 -3723
rect 1446 -3791 1458 -3757
rect 1492 -3791 1504 -3757
rect 1446 -3825 1504 -3791
rect 1446 -3859 1458 -3825
rect 1492 -3859 1504 -3825
rect 1446 -3893 1504 -3859
rect 1446 -3927 1458 -3893
rect 1492 -3927 1504 -3893
rect 1446 -3961 1504 -3927
rect 1446 -3995 1458 -3961
rect 1492 -3995 1504 -3961
rect 1446 -4029 1504 -3995
rect 1446 -4063 1458 -4029
rect 1492 -4063 1504 -4029
rect 1446 -4097 1504 -4063
rect 1446 -4131 1458 -4097
rect 1492 -4131 1504 -4097
rect 1446 -4165 1504 -4131
rect 1446 -4199 1458 -4165
rect 1492 -4199 1504 -4165
rect 1446 -4233 1504 -4199
rect 1446 -4267 1458 -4233
rect 1492 -4267 1504 -4233
rect 1446 -4301 1504 -4267
rect 1446 -4335 1458 -4301
rect 1492 -4335 1504 -4301
rect 1446 -4369 1504 -4335
rect 1446 -4403 1458 -4369
rect 1492 -4403 1504 -4369
rect 1446 -4437 1504 -4403
rect 1446 -4471 1458 -4437
rect 1492 -4471 1504 -4437
rect 1446 -4505 1504 -4471
rect 1446 -4539 1458 -4505
rect 1492 -4539 1504 -4505
rect 1446 -4573 1504 -4539
rect 1446 -4607 1458 -4573
rect 1492 -4607 1504 -4573
rect 1446 -4641 1504 -4607
rect 1446 -4675 1458 -4641
rect 1492 -4675 1504 -4641
rect 1446 -4709 1504 -4675
rect 1446 -4743 1458 -4709
rect 1492 -4743 1504 -4709
rect 1446 -4777 1504 -4743
rect 1446 -4811 1458 -4777
rect 1492 -4811 1504 -4777
rect 1446 -4845 1504 -4811
rect 1446 -4879 1458 -4845
rect 1492 -4879 1504 -4845
rect 1446 -4913 1504 -4879
rect 1446 -4947 1458 -4913
rect 1492 -4947 1504 -4913
rect 1446 -4981 1504 -4947
rect 1446 -5015 1458 -4981
rect 1492 -5015 1504 -4981
rect 1446 -5049 1504 -5015
rect 1446 -5083 1458 -5049
rect 1492 -5083 1504 -5049
rect 1446 -5117 1504 -5083
rect 1446 -5151 1458 -5117
rect 1492 -5151 1504 -5117
rect 1446 -5185 1504 -5151
rect 1446 -5219 1458 -5185
rect 1492 -5219 1504 -5185
rect 1446 -5253 1504 -5219
rect 1446 -5287 1458 -5253
rect 1492 -5287 1504 -5253
rect 1446 -5321 1504 -5287
rect 1446 -5355 1458 -5321
rect 1492 -5355 1504 -5321
rect 1446 -5389 1504 -5355
rect 1446 -5423 1458 -5389
rect 1492 -5423 1504 -5389
rect 1446 -5457 1504 -5423
rect 1446 -5491 1458 -5457
rect 1492 -5491 1504 -5457
rect 1446 -5525 1504 -5491
rect 1446 -5559 1458 -5525
rect 1492 -5559 1504 -5525
rect 1446 -5593 1504 -5559
rect 1446 -5627 1458 -5593
rect 1492 -5627 1504 -5593
rect 1446 -5661 1504 -5627
rect 1446 -5695 1458 -5661
rect 1492 -5695 1504 -5661
rect 1446 -5729 1504 -5695
rect 1446 -5763 1458 -5729
rect 1492 -5763 1504 -5729
rect 1446 -5797 1504 -5763
rect 1446 -5831 1458 -5797
rect 1492 -5831 1504 -5797
rect 1446 -5865 1504 -5831
rect 1446 -5899 1458 -5865
rect 1492 -5899 1504 -5865
rect 1446 -5933 1504 -5899
rect 1446 -5967 1458 -5933
rect 1492 -5967 1504 -5933
rect 1446 -6001 1504 -5967
rect 1446 -6035 1458 -6001
rect 1492 -6035 1504 -6001
rect 1446 -6069 1504 -6035
rect 1446 -6103 1458 -6069
rect 1492 -6103 1504 -6069
rect 1446 -6137 1504 -6103
rect 1446 -6171 1458 -6137
rect 1492 -6171 1504 -6137
rect 1446 -6205 1504 -6171
rect 1446 -6239 1458 -6205
rect 1492 -6239 1504 -6205
rect 1446 -6273 1504 -6239
rect 1446 -6307 1458 -6273
rect 1492 -6307 1504 -6273
rect 1446 -6341 1504 -6307
rect 1446 -6375 1458 -6341
rect 1492 -6375 1504 -6341
rect 1446 -6409 1504 -6375
rect 1446 -6443 1458 -6409
rect 1492 -6443 1504 -6409
rect 1446 -6477 1504 -6443
rect 1446 -6511 1458 -6477
rect 1492 -6511 1504 -6477
rect 1446 -6545 1504 -6511
rect 1446 -6579 1458 -6545
rect 1492 -6579 1504 -6545
rect 1446 -6613 1504 -6579
rect 1446 -6647 1458 -6613
rect 1492 -6647 1504 -6613
rect 1446 -6681 1504 -6647
rect 1446 -6715 1458 -6681
rect 1492 -6715 1504 -6681
rect 1446 -6749 1504 -6715
rect 1446 -6783 1458 -6749
rect 1492 -6783 1504 -6749
rect 1446 -6817 1504 -6783
rect 1446 -6851 1458 -6817
rect 1492 -6851 1504 -6817
rect 1446 -6885 1504 -6851
rect 1446 -6919 1458 -6885
rect 1492 -6919 1504 -6885
rect 1446 -6953 1504 -6919
rect 1446 -6987 1458 -6953
rect 1492 -6987 1504 -6953
rect 1446 -7021 1504 -6987
rect 1446 -7055 1458 -7021
rect 1492 -7055 1504 -7021
rect 1446 -7089 1504 -7055
rect 1446 -7123 1458 -7089
rect 1492 -7123 1504 -7089
rect 1446 -7157 1504 -7123
rect 1446 -7191 1458 -7157
rect 1492 -7191 1504 -7157
rect 1446 -7225 1504 -7191
rect 1446 -7259 1458 -7225
rect 1492 -7259 1504 -7225
rect 1446 -7293 1504 -7259
rect 1446 -7327 1458 -7293
rect 1492 -7327 1504 -7293
rect 1446 -7361 1504 -7327
rect 1446 -7395 1458 -7361
rect 1492 -7395 1504 -7361
rect 1446 -7429 1504 -7395
rect 1446 -7463 1458 -7429
rect 1492 -7463 1504 -7429
rect 1446 -7497 1504 -7463
rect 1446 -7531 1458 -7497
rect 1492 -7531 1504 -7497
rect 1446 -7565 1504 -7531
rect 1446 -7599 1458 -7565
rect 1492 -7599 1504 -7565
rect 1446 -7633 1504 -7599
rect 1446 -7667 1458 -7633
rect 1492 -7667 1504 -7633
rect 1446 -7701 1504 -7667
rect 1446 -7735 1458 -7701
rect 1492 -7735 1504 -7701
rect 1446 -7769 1504 -7735
rect 1446 -7803 1458 -7769
rect 1492 -7803 1504 -7769
rect 1446 -7837 1504 -7803
rect 1446 -7871 1458 -7837
rect 1492 -7871 1504 -7837
rect 1446 -7905 1504 -7871
rect 1446 -7939 1458 -7905
rect 1492 -7939 1504 -7905
rect 1446 -7973 1504 -7939
rect 1446 -8007 1458 -7973
rect 1492 -8007 1504 -7973
rect 1446 -8041 1504 -8007
rect 1446 -8075 1458 -8041
rect 1492 -8075 1504 -8041
rect 1446 -8109 1504 -8075
rect 1446 -8143 1458 -8109
rect 1492 -8143 1504 -8109
rect 1446 -8177 1504 -8143
rect 1446 -8211 1458 -8177
rect 1492 -8211 1504 -8177
rect 1446 -8245 1504 -8211
rect 1446 -8279 1458 -8245
rect 1492 -8279 1504 -8245
rect 1446 -8313 1504 -8279
rect 1446 -8347 1458 -8313
rect 1492 -8347 1504 -8313
rect 1446 -8381 1504 -8347
rect 1446 -8415 1458 -8381
rect 1492 -8415 1504 -8381
rect 1446 -8449 1504 -8415
rect 1446 -8483 1458 -8449
rect 1492 -8483 1504 -8449
rect 1446 -8517 1504 -8483
rect 1446 -8551 1458 -8517
rect 1492 -8551 1504 -8517
rect 1446 -8585 1504 -8551
rect 1446 -8619 1458 -8585
rect 1492 -8619 1504 -8585
rect 1446 -8653 1504 -8619
rect 1446 -8687 1458 -8653
rect 1492 -8687 1504 -8653
rect 1446 -8721 1504 -8687
rect 1446 -8755 1458 -8721
rect 1492 -8755 1504 -8721
rect 1446 -8789 1504 -8755
rect 1446 -8823 1458 -8789
rect 1492 -8823 1504 -8789
rect 1446 -8857 1504 -8823
rect 1446 -8891 1458 -8857
rect 1492 -8891 1504 -8857
rect 1446 -8925 1504 -8891
rect 1446 -8959 1458 -8925
rect 1492 -8959 1504 -8925
rect 1446 -8993 1504 -8959
rect 1446 -9027 1458 -8993
rect 1492 -9027 1504 -8993
rect 1446 -9061 1504 -9027
rect 1446 -9095 1458 -9061
rect 1492 -9095 1504 -9061
rect 1446 -9129 1504 -9095
rect 1446 -9163 1458 -9129
rect 1492 -9163 1504 -9129
rect 1446 -9197 1504 -9163
rect 1446 -9231 1458 -9197
rect 1492 -9231 1504 -9197
rect 1446 -9265 1504 -9231
rect 1446 -9299 1458 -9265
rect 1492 -9299 1504 -9265
rect 1446 -9333 1504 -9299
rect 1446 -9367 1458 -9333
rect 1492 -9367 1504 -9333
rect 1446 -9401 1504 -9367
rect 1446 -9435 1458 -9401
rect 1492 -9435 1504 -9401
rect 1446 -9469 1504 -9435
rect 1446 -9503 1458 -9469
rect 1492 -9503 1504 -9469
rect 1446 -9537 1504 -9503
rect 1446 -9571 1458 -9537
rect 1492 -9571 1504 -9537
rect 1446 -9600 1504 -9571
<< ndiffc >>
rect -1492 9537 -1458 9571
rect -1492 9469 -1458 9503
rect -1492 9401 -1458 9435
rect -1492 9333 -1458 9367
rect -1492 9265 -1458 9299
rect -1492 9197 -1458 9231
rect -1492 9129 -1458 9163
rect -1492 9061 -1458 9095
rect -1492 8993 -1458 9027
rect -1492 8925 -1458 8959
rect -1492 8857 -1458 8891
rect -1492 8789 -1458 8823
rect -1492 8721 -1458 8755
rect -1492 8653 -1458 8687
rect -1492 8585 -1458 8619
rect -1492 8517 -1458 8551
rect -1492 8449 -1458 8483
rect -1492 8381 -1458 8415
rect -1492 8313 -1458 8347
rect -1492 8245 -1458 8279
rect -1492 8177 -1458 8211
rect -1492 8109 -1458 8143
rect -1492 8041 -1458 8075
rect -1492 7973 -1458 8007
rect -1492 7905 -1458 7939
rect -1492 7837 -1458 7871
rect -1492 7769 -1458 7803
rect -1492 7701 -1458 7735
rect -1492 7633 -1458 7667
rect -1492 7565 -1458 7599
rect -1492 7497 -1458 7531
rect -1492 7429 -1458 7463
rect -1492 7361 -1458 7395
rect -1492 7293 -1458 7327
rect -1492 7225 -1458 7259
rect -1492 7157 -1458 7191
rect -1492 7089 -1458 7123
rect -1492 7021 -1458 7055
rect -1492 6953 -1458 6987
rect -1492 6885 -1458 6919
rect -1492 6817 -1458 6851
rect -1492 6749 -1458 6783
rect -1492 6681 -1458 6715
rect -1492 6613 -1458 6647
rect -1492 6545 -1458 6579
rect -1492 6477 -1458 6511
rect -1492 6409 -1458 6443
rect -1492 6341 -1458 6375
rect -1492 6273 -1458 6307
rect -1492 6205 -1458 6239
rect -1492 6137 -1458 6171
rect -1492 6069 -1458 6103
rect -1492 6001 -1458 6035
rect -1492 5933 -1458 5967
rect -1492 5865 -1458 5899
rect -1492 5797 -1458 5831
rect -1492 5729 -1458 5763
rect -1492 5661 -1458 5695
rect -1492 5593 -1458 5627
rect -1492 5525 -1458 5559
rect -1492 5457 -1458 5491
rect -1492 5389 -1458 5423
rect -1492 5321 -1458 5355
rect -1492 5253 -1458 5287
rect -1492 5185 -1458 5219
rect -1492 5117 -1458 5151
rect -1492 5049 -1458 5083
rect -1492 4981 -1458 5015
rect -1492 4913 -1458 4947
rect -1492 4845 -1458 4879
rect -1492 4777 -1458 4811
rect -1492 4709 -1458 4743
rect -1492 4641 -1458 4675
rect -1492 4573 -1458 4607
rect -1492 4505 -1458 4539
rect -1492 4437 -1458 4471
rect -1492 4369 -1458 4403
rect -1492 4301 -1458 4335
rect -1492 4233 -1458 4267
rect -1492 4165 -1458 4199
rect -1492 4097 -1458 4131
rect -1492 4029 -1458 4063
rect -1492 3961 -1458 3995
rect -1492 3893 -1458 3927
rect -1492 3825 -1458 3859
rect -1492 3757 -1458 3791
rect -1492 3689 -1458 3723
rect -1492 3621 -1458 3655
rect -1492 3553 -1458 3587
rect -1492 3485 -1458 3519
rect -1492 3417 -1458 3451
rect -1492 3349 -1458 3383
rect -1492 3281 -1458 3315
rect -1492 3213 -1458 3247
rect -1492 3145 -1458 3179
rect -1492 3077 -1458 3111
rect -1492 3009 -1458 3043
rect -1492 2941 -1458 2975
rect -1492 2873 -1458 2907
rect -1492 2805 -1458 2839
rect -1492 2737 -1458 2771
rect -1492 2669 -1458 2703
rect -1492 2601 -1458 2635
rect -1492 2533 -1458 2567
rect -1492 2465 -1458 2499
rect -1492 2397 -1458 2431
rect -1492 2329 -1458 2363
rect -1492 2261 -1458 2295
rect -1492 2193 -1458 2227
rect -1492 2125 -1458 2159
rect -1492 2057 -1458 2091
rect -1492 1989 -1458 2023
rect -1492 1921 -1458 1955
rect -1492 1853 -1458 1887
rect -1492 1785 -1458 1819
rect -1492 1717 -1458 1751
rect -1492 1649 -1458 1683
rect -1492 1581 -1458 1615
rect -1492 1513 -1458 1547
rect -1492 1445 -1458 1479
rect -1492 1377 -1458 1411
rect -1492 1309 -1458 1343
rect -1492 1241 -1458 1275
rect -1492 1173 -1458 1207
rect -1492 1105 -1458 1139
rect -1492 1037 -1458 1071
rect -1492 969 -1458 1003
rect -1492 901 -1458 935
rect -1492 833 -1458 867
rect -1492 765 -1458 799
rect -1492 697 -1458 731
rect -1492 629 -1458 663
rect -1492 561 -1458 595
rect -1492 493 -1458 527
rect -1492 425 -1458 459
rect -1492 357 -1458 391
rect -1492 289 -1458 323
rect -1492 221 -1458 255
rect -1492 153 -1458 187
rect -1492 85 -1458 119
rect -1492 17 -1458 51
rect -1492 -51 -1458 -17
rect -1492 -119 -1458 -85
rect -1492 -187 -1458 -153
rect -1492 -255 -1458 -221
rect -1492 -323 -1458 -289
rect -1492 -391 -1458 -357
rect -1492 -459 -1458 -425
rect -1492 -527 -1458 -493
rect -1492 -595 -1458 -561
rect -1492 -663 -1458 -629
rect -1492 -731 -1458 -697
rect -1492 -799 -1458 -765
rect -1492 -867 -1458 -833
rect -1492 -935 -1458 -901
rect -1492 -1003 -1458 -969
rect -1492 -1071 -1458 -1037
rect -1492 -1139 -1458 -1105
rect -1492 -1207 -1458 -1173
rect -1492 -1275 -1458 -1241
rect -1492 -1343 -1458 -1309
rect -1492 -1411 -1458 -1377
rect -1492 -1479 -1458 -1445
rect -1492 -1547 -1458 -1513
rect -1492 -1615 -1458 -1581
rect -1492 -1683 -1458 -1649
rect -1492 -1751 -1458 -1717
rect -1492 -1819 -1458 -1785
rect -1492 -1887 -1458 -1853
rect -1492 -1955 -1458 -1921
rect -1492 -2023 -1458 -1989
rect -1492 -2091 -1458 -2057
rect -1492 -2159 -1458 -2125
rect -1492 -2227 -1458 -2193
rect -1492 -2295 -1458 -2261
rect -1492 -2363 -1458 -2329
rect -1492 -2431 -1458 -2397
rect -1492 -2499 -1458 -2465
rect -1492 -2567 -1458 -2533
rect -1492 -2635 -1458 -2601
rect -1492 -2703 -1458 -2669
rect -1492 -2771 -1458 -2737
rect -1492 -2839 -1458 -2805
rect -1492 -2907 -1458 -2873
rect -1492 -2975 -1458 -2941
rect -1492 -3043 -1458 -3009
rect -1492 -3111 -1458 -3077
rect -1492 -3179 -1458 -3145
rect -1492 -3247 -1458 -3213
rect -1492 -3315 -1458 -3281
rect -1492 -3383 -1458 -3349
rect -1492 -3451 -1458 -3417
rect -1492 -3519 -1458 -3485
rect -1492 -3587 -1458 -3553
rect -1492 -3655 -1458 -3621
rect -1492 -3723 -1458 -3689
rect -1492 -3791 -1458 -3757
rect -1492 -3859 -1458 -3825
rect -1492 -3927 -1458 -3893
rect -1492 -3995 -1458 -3961
rect -1492 -4063 -1458 -4029
rect -1492 -4131 -1458 -4097
rect -1492 -4199 -1458 -4165
rect -1492 -4267 -1458 -4233
rect -1492 -4335 -1458 -4301
rect -1492 -4403 -1458 -4369
rect -1492 -4471 -1458 -4437
rect -1492 -4539 -1458 -4505
rect -1492 -4607 -1458 -4573
rect -1492 -4675 -1458 -4641
rect -1492 -4743 -1458 -4709
rect -1492 -4811 -1458 -4777
rect -1492 -4879 -1458 -4845
rect -1492 -4947 -1458 -4913
rect -1492 -5015 -1458 -4981
rect -1492 -5083 -1458 -5049
rect -1492 -5151 -1458 -5117
rect -1492 -5219 -1458 -5185
rect -1492 -5287 -1458 -5253
rect -1492 -5355 -1458 -5321
rect -1492 -5423 -1458 -5389
rect -1492 -5491 -1458 -5457
rect -1492 -5559 -1458 -5525
rect -1492 -5627 -1458 -5593
rect -1492 -5695 -1458 -5661
rect -1492 -5763 -1458 -5729
rect -1492 -5831 -1458 -5797
rect -1492 -5899 -1458 -5865
rect -1492 -5967 -1458 -5933
rect -1492 -6035 -1458 -6001
rect -1492 -6103 -1458 -6069
rect -1492 -6171 -1458 -6137
rect -1492 -6239 -1458 -6205
rect -1492 -6307 -1458 -6273
rect -1492 -6375 -1458 -6341
rect -1492 -6443 -1458 -6409
rect -1492 -6511 -1458 -6477
rect -1492 -6579 -1458 -6545
rect -1492 -6647 -1458 -6613
rect -1492 -6715 -1458 -6681
rect -1492 -6783 -1458 -6749
rect -1492 -6851 -1458 -6817
rect -1492 -6919 -1458 -6885
rect -1492 -6987 -1458 -6953
rect -1492 -7055 -1458 -7021
rect -1492 -7123 -1458 -7089
rect -1492 -7191 -1458 -7157
rect -1492 -7259 -1458 -7225
rect -1492 -7327 -1458 -7293
rect -1492 -7395 -1458 -7361
rect -1492 -7463 -1458 -7429
rect -1492 -7531 -1458 -7497
rect -1492 -7599 -1458 -7565
rect -1492 -7667 -1458 -7633
rect -1492 -7735 -1458 -7701
rect -1492 -7803 -1458 -7769
rect -1492 -7871 -1458 -7837
rect -1492 -7939 -1458 -7905
rect -1492 -8007 -1458 -7973
rect -1492 -8075 -1458 -8041
rect -1492 -8143 -1458 -8109
rect -1492 -8211 -1458 -8177
rect -1492 -8279 -1458 -8245
rect -1492 -8347 -1458 -8313
rect -1492 -8415 -1458 -8381
rect -1492 -8483 -1458 -8449
rect -1492 -8551 -1458 -8517
rect -1492 -8619 -1458 -8585
rect -1492 -8687 -1458 -8653
rect -1492 -8755 -1458 -8721
rect -1492 -8823 -1458 -8789
rect -1492 -8891 -1458 -8857
rect -1492 -8959 -1458 -8925
rect -1492 -9027 -1458 -8993
rect -1492 -9095 -1458 -9061
rect -1492 -9163 -1458 -9129
rect -1492 -9231 -1458 -9197
rect -1492 -9299 -1458 -9265
rect -1492 -9367 -1458 -9333
rect -1492 -9435 -1458 -9401
rect -1492 -9503 -1458 -9469
rect -1492 -9571 -1458 -9537
rect -1374 9537 -1340 9571
rect -1374 9469 -1340 9503
rect -1374 9401 -1340 9435
rect -1374 9333 -1340 9367
rect -1374 9265 -1340 9299
rect -1374 9197 -1340 9231
rect -1374 9129 -1340 9163
rect -1374 9061 -1340 9095
rect -1374 8993 -1340 9027
rect -1374 8925 -1340 8959
rect -1374 8857 -1340 8891
rect -1374 8789 -1340 8823
rect -1374 8721 -1340 8755
rect -1374 8653 -1340 8687
rect -1374 8585 -1340 8619
rect -1374 8517 -1340 8551
rect -1374 8449 -1340 8483
rect -1374 8381 -1340 8415
rect -1374 8313 -1340 8347
rect -1374 8245 -1340 8279
rect -1374 8177 -1340 8211
rect -1374 8109 -1340 8143
rect -1374 8041 -1340 8075
rect -1374 7973 -1340 8007
rect -1374 7905 -1340 7939
rect -1374 7837 -1340 7871
rect -1374 7769 -1340 7803
rect -1374 7701 -1340 7735
rect -1374 7633 -1340 7667
rect -1374 7565 -1340 7599
rect -1374 7497 -1340 7531
rect -1374 7429 -1340 7463
rect -1374 7361 -1340 7395
rect -1374 7293 -1340 7327
rect -1374 7225 -1340 7259
rect -1374 7157 -1340 7191
rect -1374 7089 -1340 7123
rect -1374 7021 -1340 7055
rect -1374 6953 -1340 6987
rect -1374 6885 -1340 6919
rect -1374 6817 -1340 6851
rect -1374 6749 -1340 6783
rect -1374 6681 -1340 6715
rect -1374 6613 -1340 6647
rect -1374 6545 -1340 6579
rect -1374 6477 -1340 6511
rect -1374 6409 -1340 6443
rect -1374 6341 -1340 6375
rect -1374 6273 -1340 6307
rect -1374 6205 -1340 6239
rect -1374 6137 -1340 6171
rect -1374 6069 -1340 6103
rect -1374 6001 -1340 6035
rect -1374 5933 -1340 5967
rect -1374 5865 -1340 5899
rect -1374 5797 -1340 5831
rect -1374 5729 -1340 5763
rect -1374 5661 -1340 5695
rect -1374 5593 -1340 5627
rect -1374 5525 -1340 5559
rect -1374 5457 -1340 5491
rect -1374 5389 -1340 5423
rect -1374 5321 -1340 5355
rect -1374 5253 -1340 5287
rect -1374 5185 -1340 5219
rect -1374 5117 -1340 5151
rect -1374 5049 -1340 5083
rect -1374 4981 -1340 5015
rect -1374 4913 -1340 4947
rect -1374 4845 -1340 4879
rect -1374 4777 -1340 4811
rect -1374 4709 -1340 4743
rect -1374 4641 -1340 4675
rect -1374 4573 -1340 4607
rect -1374 4505 -1340 4539
rect -1374 4437 -1340 4471
rect -1374 4369 -1340 4403
rect -1374 4301 -1340 4335
rect -1374 4233 -1340 4267
rect -1374 4165 -1340 4199
rect -1374 4097 -1340 4131
rect -1374 4029 -1340 4063
rect -1374 3961 -1340 3995
rect -1374 3893 -1340 3927
rect -1374 3825 -1340 3859
rect -1374 3757 -1340 3791
rect -1374 3689 -1340 3723
rect -1374 3621 -1340 3655
rect -1374 3553 -1340 3587
rect -1374 3485 -1340 3519
rect -1374 3417 -1340 3451
rect -1374 3349 -1340 3383
rect -1374 3281 -1340 3315
rect -1374 3213 -1340 3247
rect -1374 3145 -1340 3179
rect -1374 3077 -1340 3111
rect -1374 3009 -1340 3043
rect -1374 2941 -1340 2975
rect -1374 2873 -1340 2907
rect -1374 2805 -1340 2839
rect -1374 2737 -1340 2771
rect -1374 2669 -1340 2703
rect -1374 2601 -1340 2635
rect -1374 2533 -1340 2567
rect -1374 2465 -1340 2499
rect -1374 2397 -1340 2431
rect -1374 2329 -1340 2363
rect -1374 2261 -1340 2295
rect -1374 2193 -1340 2227
rect -1374 2125 -1340 2159
rect -1374 2057 -1340 2091
rect -1374 1989 -1340 2023
rect -1374 1921 -1340 1955
rect -1374 1853 -1340 1887
rect -1374 1785 -1340 1819
rect -1374 1717 -1340 1751
rect -1374 1649 -1340 1683
rect -1374 1581 -1340 1615
rect -1374 1513 -1340 1547
rect -1374 1445 -1340 1479
rect -1374 1377 -1340 1411
rect -1374 1309 -1340 1343
rect -1374 1241 -1340 1275
rect -1374 1173 -1340 1207
rect -1374 1105 -1340 1139
rect -1374 1037 -1340 1071
rect -1374 969 -1340 1003
rect -1374 901 -1340 935
rect -1374 833 -1340 867
rect -1374 765 -1340 799
rect -1374 697 -1340 731
rect -1374 629 -1340 663
rect -1374 561 -1340 595
rect -1374 493 -1340 527
rect -1374 425 -1340 459
rect -1374 357 -1340 391
rect -1374 289 -1340 323
rect -1374 221 -1340 255
rect -1374 153 -1340 187
rect -1374 85 -1340 119
rect -1374 17 -1340 51
rect -1374 -51 -1340 -17
rect -1374 -119 -1340 -85
rect -1374 -187 -1340 -153
rect -1374 -255 -1340 -221
rect -1374 -323 -1340 -289
rect -1374 -391 -1340 -357
rect -1374 -459 -1340 -425
rect -1374 -527 -1340 -493
rect -1374 -595 -1340 -561
rect -1374 -663 -1340 -629
rect -1374 -731 -1340 -697
rect -1374 -799 -1340 -765
rect -1374 -867 -1340 -833
rect -1374 -935 -1340 -901
rect -1374 -1003 -1340 -969
rect -1374 -1071 -1340 -1037
rect -1374 -1139 -1340 -1105
rect -1374 -1207 -1340 -1173
rect -1374 -1275 -1340 -1241
rect -1374 -1343 -1340 -1309
rect -1374 -1411 -1340 -1377
rect -1374 -1479 -1340 -1445
rect -1374 -1547 -1340 -1513
rect -1374 -1615 -1340 -1581
rect -1374 -1683 -1340 -1649
rect -1374 -1751 -1340 -1717
rect -1374 -1819 -1340 -1785
rect -1374 -1887 -1340 -1853
rect -1374 -1955 -1340 -1921
rect -1374 -2023 -1340 -1989
rect -1374 -2091 -1340 -2057
rect -1374 -2159 -1340 -2125
rect -1374 -2227 -1340 -2193
rect -1374 -2295 -1340 -2261
rect -1374 -2363 -1340 -2329
rect -1374 -2431 -1340 -2397
rect -1374 -2499 -1340 -2465
rect -1374 -2567 -1340 -2533
rect -1374 -2635 -1340 -2601
rect -1374 -2703 -1340 -2669
rect -1374 -2771 -1340 -2737
rect -1374 -2839 -1340 -2805
rect -1374 -2907 -1340 -2873
rect -1374 -2975 -1340 -2941
rect -1374 -3043 -1340 -3009
rect -1374 -3111 -1340 -3077
rect -1374 -3179 -1340 -3145
rect -1374 -3247 -1340 -3213
rect -1374 -3315 -1340 -3281
rect -1374 -3383 -1340 -3349
rect -1374 -3451 -1340 -3417
rect -1374 -3519 -1340 -3485
rect -1374 -3587 -1340 -3553
rect -1374 -3655 -1340 -3621
rect -1374 -3723 -1340 -3689
rect -1374 -3791 -1340 -3757
rect -1374 -3859 -1340 -3825
rect -1374 -3927 -1340 -3893
rect -1374 -3995 -1340 -3961
rect -1374 -4063 -1340 -4029
rect -1374 -4131 -1340 -4097
rect -1374 -4199 -1340 -4165
rect -1374 -4267 -1340 -4233
rect -1374 -4335 -1340 -4301
rect -1374 -4403 -1340 -4369
rect -1374 -4471 -1340 -4437
rect -1374 -4539 -1340 -4505
rect -1374 -4607 -1340 -4573
rect -1374 -4675 -1340 -4641
rect -1374 -4743 -1340 -4709
rect -1374 -4811 -1340 -4777
rect -1374 -4879 -1340 -4845
rect -1374 -4947 -1340 -4913
rect -1374 -5015 -1340 -4981
rect -1374 -5083 -1340 -5049
rect -1374 -5151 -1340 -5117
rect -1374 -5219 -1340 -5185
rect -1374 -5287 -1340 -5253
rect -1374 -5355 -1340 -5321
rect -1374 -5423 -1340 -5389
rect -1374 -5491 -1340 -5457
rect -1374 -5559 -1340 -5525
rect -1374 -5627 -1340 -5593
rect -1374 -5695 -1340 -5661
rect -1374 -5763 -1340 -5729
rect -1374 -5831 -1340 -5797
rect -1374 -5899 -1340 -5865
rect -1374 -5967 -1340 -5933
rect -1374 -6035 -1340 -6001
rect -1374 -6103 -1340 -6069
rect -1374 -6171 -1340 -6137
rect -1374 -6239 -1340 -6205
rect -1374 -6307 -1340 -6273
rect -1374 -6375 -1340 -6341
rect -1374 -6443 -1340 -6409
rect -1374 -6511 -1340 -6477
rect -1374 -6579 -1340 -6545
rect -1374 -6647 -1340 -6613
rect -1374 -6715 -1340 -6681
rect -1374 -6783 -1340 -6749
rect -1374 -6851 -1340 -6817
rect -1374 -6919 -1340 -6885
rect -1374 -6987 -1340 -6953
rect -1374 -7055 -1340 -7021
rect -1374 -7123 -1340 -7089
rect -1374 -7191 -1340 -7157
rect -1374 -7259 -1340 -7225
rect -1374 -7327 -1340 -7293
rect -1374 -7395 -1340 -7361
rect -1374 -7463 -1340 -7429
rect -1374 -7531 -1340 -7497
rect -1374 -7599 -1340 -7565
rect -1374 -7667 -1340 -7633
rect -1374 -7735 -1340 -7701
rect -1374 -7803 -1340 -7769
rect -1374 -7871 -1340 -7837
rect -1374 -7939 -1340 -7905
rect -1374 -8007 -1340 -7973
rect -1374 -8075 -1340 -8041
rect -1374 -8143 -1340 -8109
rect -1374 -8211 -1340 -8177
rect -1374 -8279 -1340 -8245
rect -1374 -8347 -1340 -8313
rect -1374 -8415 -1340 -8381
rect -1374 -8483 -1340 -8449
rect -1374 -8551 -1340 -8517
rect -1374 -8619 -1340 -8585
rect -1374 -8687 -1340 -8653
rect -1374 -8755 -1340 -8721
rect -1374 -8823 -1340 -8789
rect -1374 -8891 -1340 -8857
rect -1374 -8959 -1340 -8925
rect -1374 -9027 -1340 -8993
rect -1374 -9095 -1340 -9061
rect -1374 -9163 -1340 -9129
rect -1374 -9231 -1340 -9197
rect -1374 -9299 -1340 -9265
rect -1374 -9367 -1340 -9333
rect -1374 -9435 -1340 -9401
rect -1374 -9503 -1340 -9469
rect -1374 -9571 -1340 -9537
rect -1256 9537 -1222 9571
rect -1256 9469 -1222 9503
rect -1256 9401 -1222 9435
rect -1256 9333 -1222 9367
rect -1256 9265 -1222 9299
rect -1256 9197 -1222 9231
rect -1256 9129 -1222 9163
rect -1256 9061 -1222 9095
rect -1256 8993 -1222 9027
rect -1256 8925 -1222 8959
rect -1256 8857 -1222 8891
rect -1256 8789 -1222 8823
rect -1256 8721 -1222 8755
rect -1256 8653 -1222 8687
rect -1256 8585 -1222 8619
rect -1256 8517 -1222 8551
rect -1256 8449 -1222 8483
rect -1256 8381 -1222 8415
rect -1256 8313 -1222 8347
rect -1256 8245 -1222 8279
rect -1256 8177 -1222 8211
rect -1256 8109 -1222 8143
rect -1256 8041 -1222 8075
rect -1256 7973 -1222 8007
rect -1256 7905 -1222 7939
rect -1256 7837 -1222 7871
rect -1256 7769 -1222 7803
rect -1256 7701 -1222 7735
rect -1256 7633 -1222 7667
rect -1256 7565 -1222 7599
rect -1256 7497 -1222 7531
rect -1256 7429 -1222 7463
rect -1256 7361 -1222 7395
rect -1256 7293 -1222 7327
rect -1256 7225 -1222 7259
rect -1256 7157 -1222 7191
rect -1256 7089 -1222 7123
rect -1256 7021 -1222 7055
rect -1256 6953 -1222 6987
rect -1256 6885 -1222 6919
rect -1256 6817 -1222 6851
rect -1256 6749 -1222 6783
rect -1256 6681 -1222 6715
rect -1256 6613 -1222 6647
rect -1256 6545 -1222 6579
rect -1256 6477 -1222 6511
rect -1256 6409 -1222 6443
rect -1256 6341 -1222 6375
rect -1256 6273 -1222 6307
rect -1256 6205 -1222 6239
rect -1256 6137 -1222 6171
rect -1256 6069 -1222 6103
rect -1256 6001 -1222 6035
rect -1256 5933 -1222 5967
rect -1256 5865 -1222 5899
rect -1256 5797 -1222 5831
rect -1256 5729 -1222 5763
rect -1256 5661 -1222 5695
rect -1256 5593 -1222 5627
rect -1256 5525 -1222 5559
rect -1256 5457 -1222 5491
rect -1256 5389 -1222 5423
rect -1256 5321 -1222 5355
rect -1256 5253 -1222 5287
rect -1256 5185 -1222 5219
rect -1256 5117 -1222 5151
rect -1256 5049 -1222 5083
rect -1256 4981 -1222 5015
rect -1256 4913 -1222 4947
rect -1256 4845 -1222 4879
rect -1256 4777 -1222 4811
rect -1256 4709 -1222 4743
rect -1256 4641 -1222 4675
rect -1256 4573 -1222 4607
rect -1256 4505 -1222 4539
rect -1256 4437 -1222 4471
rect -1256 4369 -1222 4403
rect -1256 4301 -1222 4335
rect -1256 4233 -1222 4267
rect -1256 4165 -1222 4199
rect -1256 4097 -1222 4131
rect -1256 4029 -1222 4063
rect -1256 3961 -1222 3995
rect -1256 3893 -1222 3927
rect -1256 3825 -1222 3859
rect -1256 3757 -1222 3791
rect -1256 3689 -1222 3723
rect -1256 3621 -1222 3655
rect -1256 3553 -1222 3587
rect -1256 3485 -1222 3519
rect -1256 3417 -1222 3451
rect -1256 3349 -1222 3383
rect -1256 3281 -1222 3315
rect -1256 3213 -1222 3247
rect -1256 3145 -1222 3179
rect -1256 3077 -1222 3111
rect -1256 3009 -1222 3043
rect -1256 2941 -1222 2975
rect -1256 2873 -1222 2907
rect -1256 2805 -1222 2839
rect -1256 2737 -1222 2771
rect -1256 2669 -1222 2703
rect -1256 2601 -1222 2635
rect -1256 2533 -1222 2567
rect -1256 2465 -1222 2499
rect -1256 2397 -1222 2431
rect -1256 2329 -1222 2363
rect -1256 2261 -1222 2295
rect -1256 2193 -1222 2227
rect -1256 2125 -1222 2159
rect -1256 2057 -1222 2091
rect -1256 1989 -1222 2023
rect -1256 1921 -1222 1955
rect -1256 1853 -1222 1887
rect -1256 1785 -1222 1819
rect -1256 1717 -1222 1751
rect -1256 1649 -1222 1683
rect -1256 1581 -1222 1615
rect -1256 1513 -1222 1547
rect -1256 1445 -1222 1479
rect -1256 1377 -1222 1411
rect -1256 1309 -1222 1343
rect -1256 1241 -1222 1275
rect -1256 1173 -1222 1207
rect -1256 1105 -1222 1139
rect -1256 1037 -1222 1071
rect -1256 969 -1222 1003
rect -1256 901 -1222 935
rect -1256 833 -1222 867
rect -1256 765 -1222 799
rect -1256 697 -1222 731
rect -1256 629 -1222 663
rect -1256 561 -1222 595
rect -1256 493 -1222 527
rect -1256 425 -1222 459
rect -1256 357 -1222 391
rect -1256 289 -1222 323
rect -1256 221 -1222 255
rect -1256 153 -1222 187
rect -1256 85 -1222 119
rect -1256 17 -1222 51
rect -1256 -51 -1222 -17
rect -1256 -119 -1222 -85
rect -1256 -187 -1222 -153
rect -1256 -255 -1222 -221
rect -1256 -323 -1222 -289
rect -1256 -391 -1222 -357
rect -1256 -459 -1222 -425
rect -1256 -527 -1222 -493
rect -1256 -595 -1222 -561
rect -1256 -663 -1222 -629
rect -1256 -731 -1222 -697
rect -1256 -799 -1222 -765
rect -1256 -867 -1222 -833
rect -1256 -935 -1222 -901
rect -1256 -1003 -1222 -969
rect -1256 -1071 -1222 -1037
rect -1256 -1139 -1222 -1105
rect -1256 -1207 -1222 -1173
rect -1256 -1275 -1222 -1241
rect -1256 -1343 -1222 -1309
rect -1256 -1411 -1222 -1377
rect -1256 -1479 -1222 -1445
rect -1256 -1547 -1222 -1513
rect -1256 -1615 -1222 -1581
rect -1256 -1683 -1222 -1649
rect -1256 -1751 -1222 -1717
rect -1256 -1819 -1222 -1785
rect -1256 -1887 -1222 -1853
rect -1256 -1955 -1222 -1921
rect -1256 -2023 -1222 -1989
rect -1256 -2091 -1222 -2057
rect -1256 -2159 -1222 -2125
rect -1256 -2227 -1222 -2193
rect -1256 -2295 -1222 -2261
rect -1256 -2363 -1222 -2329
rect -1256 -2431 -1222 -2397
rect -1256 -2499 -1222 -2465
rect -1256 -2567 -1222 -2533
rect -1256 -2635 -1222 -2601
rect -1256 -2703 -1222 -2669
rect -1256 -2771 -1222 -2737
rect -1256 -2839 -1222 -2805
rect -1256 -2907 -1222 -2873
rect -1256 -2975 -1222 -2941
rect -1256 -3043 -1222 -3009
rect -1256 -3111 -1222 -3077
rect -1256 -3179 -1222 -3145
rect -1256 -3247 -1222 -3213
rect -1256 -3315 -1222 -3281
rect -1256 -3383 -1222 -3349
rect -1256 -3451 -1222 -3417
rect -1256 -3519 -1222 -3485
rect -1256 -3587 -1222 -3553
rect -1256 -3655 -1222 -3621
rect -1256 -3723 -1222 -3689
rect -1256 -3791 -1222 -3757
rect -1256 -3859 -1222 -3825
rect -1256 -3927 -1222 -3893
rect -1256 -3995 -1222 -3961
rect -1256 -4063 -1222 -4029
rect -1256 -4131 -1222 -4097
rect -1256 -4199 -1222 -4165
rect -1256 -4267 -1222 -4233
rect -1256 -4335 -1222 -4301
rect -1256 -4403 -1222 -4369
rect -1256 -4471 -1222 -4437
rect -1256 -4539 -1222 -4505
rect -1256 -4607 -1222 -4573
rect -1256 -4675 -1222 -4641
rect -1256 -4743 -1222 -4709
rect -1256 -4811 -1222 -4777
rect -1256 -4879 -1222 -4845
rect -1256 -4947 -1222 -4913
rect -1256 -5015 -1222 -4981
rect -1256 -5083 -1222 -5049
rect -1256 -5151 -1222 -5117
rect -1256 -5219 -1222 -5185
rect -1256 -5287 -1222 -5253
rect -1256 -5355 -1222 -5321
rect -1256 -5423 -1222 -5389
rect -1256 -5491 -1222 -5457
rect -1256 -5559 -1222 -5525
rect -1256 -5627 -1222 -5593
rect -1256 -5695 -1222 -5661
rect -1256 -5763 -1222 -5729
rect -1256 -5831 -1222 -5797
rect -1256 -5899 -1222 -5865
rect -1256 -5967 -1222 -5933
rect -1256 -6035 -1222 -6001
rect -1256 -6103 -1222 -6069
rect -1256 -6171 -1222 -6137
rect -1256 -6239 -1222 -6205
rect -1256 -6307 -1222 -6273
rect -1256 -6375 -1222 -6341
rect -1256 -6443 -1222 -6409
rect -1256 -6511 -1222 -6477
rect -1256 -6579 -1222 -6545
rect -1256 -6647 -1222 -6613
rect -1256 -6715 -1222 -6681
rect -1256 -6783 -1222 -6749
rect -1256 -6851 -1222 -6817
rect -1256 -6919 -1222 -6885
rect -1256 -6987 -1222 -6953
rect -1256 -7055 -1222 -7021
rect -1256 -7123 -1222 -7089
rect -1256 -7191 -1222 -7157
rect -1256 -7259 -1222 -7225
rect -1256 -7327 -1222 -7293
rect -1256 -7395 -1222 -7361
rect -1256 -7463 -1222 -7429
rect -1256 -7531 -1222 -7497
rect -1256 -7599 -1222 -7565
rect -1256 -7667 -1222 -7633
rect -1256 -7735 -1222 -7701
rect -1256 -7803 -1222 -7769
rect -1256 -7871 -1222 -7837
rect -1256 -7939 -1222 -7905
rect -1256 -8007 -1222 -7973
rect -1256 -8075 -1222 -8041
rect -1256 -8143 -1222 -8109
rect -1256 -8211 -1222 -8177
rect -1256 -8279 -1222 -8245
rect -1256 -8347 -1222 -8313
rect -1256 -8415 -1222 -8381
rect -1256 -8483 -1222 -8449
rect -1256 -8551 -1222 -8517
rect -1256 -8619 -1222 -8585
rect -1256 -8687 -1222 -8653
rect -1256 -8755 -1222 -8721
rect -1256 -8823 -1222 -8789
rect -1256 -8891 -1222 -8857
rect -1256 -8959 -1222 -8925
rect -1256 -9027 -1222 -8993
rect -1256 -9095 -1222 -9061
rect -1256 -9163 -1222 -9129
rect -1256 -9231 -1222 -9197
rect -1256 -9299 -1222 -9265
rect -1256 -9367 -1222 -9333
rect -1256 -9435 -1222 -9401
rect -1256 -9503 -1222 -9469
rect -1256 -9571 -1222 -9537
rect -1138 9537 -1104 9571
rect -1138 9469 -1104 9503
rect -1138 9401 -1104 9435
rect -1138 9333 -1104 9367
rect -1138 9265 -1104 9299
rect -1138 9197 -1104 9231
rect -1138 9129 -1104 9163
rect -1138 9061 -1104 9095
rect -1138 8993 -1104 9027
rect -1138 8925 -1104 8959
rect -1138 8857 -1104 8891
rect -1138 8789 -1104 8823
rect -1138 8721 -1104 8755
rect -1138 8653 -1104 8687
rect -1138 8585 -1104 8619
rect -1138 8517 -1104 8551
rect -1138 8449 -1104 8483
rect -1138 8381 -1104 8415
rect -1138 8313 -1104 8347
rect -1138 8245 -1104 8279
rect -1138 8177 -1104 8211
rect -1138 8109 -1104 8143
rect -1138 8041 -1104 8075
rect -1138 7973 -1104 8007
rect -1138 7905 -1104 7939
rect -1138 7837 -1104 7871
rect -1138 7769 -1104 7803
rect -1138 7701 -1104 7735
rect -1138 7633 -1104 7667
rect -1138 7565 -1104 7599
rect -1138 7497 -1104 7531
rect -1138 7429 -1104 7463
rect -1138 7361 -1104 7395
rect -1138 7293 -1104 7327
rect -1138 7225 -1104 7259
rect -1138 7157 -1104 7191
rect -1138 7089 -1104 7123
rect -1138 7021 -1104 7055
rect -1138 6953 -1104 6987
rect -1138 6885 -1104 6919
rect -1138 6817 -1104 6851
rect -1138 6749 -1104 6783
rect -1138 6681 -1104 6715
rect -1138 6613 -1104 6647
rect -1138 6545 -1104 6579
rect -1138 6477 -1104 6511
rect -1138 6409 -1104 6443
rect -1138 6341 -1104 6375
rect -1138 6273 -1104 6307
rect -1138 6205 -1104 6239
rect -1138 6137 -1104 6171
rect -1138 6069 -1104 6103
rect -1138 6001 -1104 6035
rect -1138 5933 -1104 5967
rect -1138 5865 -1104 5899
rect -1138 5797 -1104 5831
rect -1138 5729 -1104 5763
rect -1138 5661 -1104 5695
rect -1138 5593 -1104 5627
rect -1138 5525 -1104 5559
rect -1138 5457 -1104 5491
rect -1138 5389 -1104 5423
rect -1138 5321 -1104 5355
rect -1138 5253 -1104 5287
rect -1138 5185 -1104 5219
rect -1138 5117 -1104 5151
rect -1138 5049 -1104 5083
rect -1138 4981 -1104 5015
rect -1138 4913 -1104 4947
rect -1138 4845 -1104 4879
rect -1138 4777 -1104 4811
rect -1138 4709 -1104 4743
rect -1138 4641 -1104 4675
rect -1138 4573 -1104 4607
rect -1138 4505 -1104 4539
rect -1138 4437 -1104 4471
rect -1138 4369 -1104 4403
rect -1138 4301 -1104 4335
rect -1138 4233 -1104 4267
rect -1138 4165 -1104 4199
rect -1138 4097 -1104 4131
rect -1138 4029 -1104 4063
rect -1138 3961 -1104 3995
rect -1138 3893 -1104 3927
rect -1138 3825 -1104 3859
rect -1138 3757 -1104 3791
rect -1138 3689 -1104 3723
rect -1138 3621 -1104 3655
rect -1138 3553 -1104 3587
rect -1138 3485 -1104 3519
rect -1138 3417 -1104 3451
rect -1138 3349 -1104 3383
rect -1138 3281 -1104 3315
rect -1138 3213 -1104 3247
rect -1138 3145 -1104 3179
rect -1138 3077 -1104 3111
rect -1138 3009 -1104 3043
rect -1138 2941 -1104 2975
rect -1138 2873 -1104 2907
rect -1138 2805 -1104 2839
rect -1138 2737 -1104 2771
rect -1138 2669 -1104 2703
rect -1138 2601 -1104 2635
rect -1138 2533 -1104 2567
rect -1138 2465 -1104 2499
rect -1138 2397 -1104 2431
rect -1138 2329 -1104 2363
rect -1138 2261 -1104 2295
rect -1138 2193 -1104 2227
rect -1138 2125 -1104 2159
rect -1138 2057 -1104 2091
rect -1138 1989 -1104 2023
rect -1138 1921 -1104 1955
rect -1138 1853 -1104 1887
rect -1138 1785 -1104 1819
rect -1138 1717 -1104 1751
rect -1138 1649 -1104 1683
rect -1138 1581 -1104 1615
rect -1138 1513 -1104 1547
rect -1138 1445 -1104 1479
rect -1138 1377 -1104 1411
rect -1138 1309 -1104 1343
rect -1138 1241 -1104 1275
rect -1138 1173 -1104 1207
rect -1138 1105 -1104 1139
rect -1138 1037 -1104 1071
rect -1138 969 -1104 1003
rect -1138 901 -1104 935
rect -1138 833 -1104 867
rect -1138 765 -1104 799
rect -1138 697 -1104 731
rect -1138 629 -1104 663
rect -1138 561 -1104 595
rect -1138 493 -1104 527
rect -1138 425 -1104 459
rect -1138 357 -1104 391
rect -1138 289 -1104 323
rect -1138 221 -1104 255
rect -1138 153 -1104 187
rect -1138 85 -1104 119
rect -1138 17 -1104 51
rect -1138 -51 -1104 -17
rect -1138 -119 -1104 -85
rect -1138 -187 -1104 -153
rect -1138 -255 -1104 -221
rect -1138 -323 -1104 -289
rect -1138 -391 -1104 -357
rect -1138 -459 -1104 -425
rect -1138 -527 -1104 -493
rect -1138 -595 -1104 -561
rect -1138 -663 -1104 -629
rect -1138 -731 -1104 -697
rect -1138 -799 -1104 -765
rect -1138 -867 -1104 -833
rect -1138 -935 -1104 -901
rect -1138 -1003 -1104 -969
rect -1138 -1071 -1104 -1037
rect -1138 -1139 -1104 -1105
rect -1138 -1207 -1104 -1173
rect -1138 -1275 -1104 -1241
rect -1138 -1343 -1104 -1309
rect -1138 -1411 -1104 -1377
rect -1138 -1479 -1104 -1445
rect -1138 -1547 -1104 -1513
rect -1138 -1615 -1104 -1581
rect -1138 -1683 -1104 -1649
rect -1138 -1751 -1104 -1717
rect -1138 -1819 -1104 -1785
rect -1138 -1887 -1104 -1853
rect -1138 -1955 -1104 -1921
rect -1138 -2023 -1104 -1989
rect -1138 -2091 -1104 -2057
rect -1138 -2159 -1104 -2125
rect -1138 -2227 -1104 -2193
rect -1138 -2295 -1104 -2261
rect -1138 -2363 -1104 -2329
rect -1138 -2431 -1104 -2397
rect -1138 -2499 -1104 -2465
rect -1138 -2567 -1104 -2533
rect -1138 -2635 -1104 -2601
rect -1138 -2703 -1104 -2669
rect -1138 -2771 -1104 -2737
rect -1138 -2839 -1104 -2805
rect -1138 -2907 -1104 -2873
rect -1138 -2975 -1104 -2941
rect -1138 -3043 -1104 -3009
rect -1138 -3111 -1104 -3077
rect -1138 -3179 -1104 -3145
rect -1138 -3247 -1104 -3213
rect -1138 -3315 -1104 -3281
rect -1138 -3383 -1104 -3349
rect -1138 -3451 -1104 -3417
rect -1138 -3519 -1104 -3485
rect -1138 -3587 -1104 -3553
rect -1138 -3655 -1104 -3621
rect -1138 -3723 -1104 -3689
rect -1138 -3791 -1104 -3757
rect -1138 -3859 -1104 -3825
rect -1138 -3927 -1104 -3893
rect -1138 -3995 -1104 -3961
rect -1138 -4063 -1104 -4029
rect -1138 -4131 -1104 -4097
rect -1138 -4199 -1104 -4165
rect -1138 -4267 -1104 -4233
rect -1138 -4335 -1104 -4301
rect -1138 -4403 -1104 -4369
rect -1138 -4471 -1104 -4437
rect -1138 -4539 -1104 -4505
rect -1138 -4607 -1104 -4573
rect -1138 -4675 -1104 -4641
rect -1138 -4743 -1104 -4709
rect -1138 -4811 -1104 -4777
rect -1138 -4879 -1104 -4845
rect -1138 -4947 -1104 -4913
rect -1138 -5015 -1104 -4981
rect -1138 -5083 -1104 -5049
rect -1138 -5151 -1104 -5117
rect -1138 -5219 -1104 -5185
rect -1138 -5287 -1104 -5253
rect -1138 -5355 -1104 -5321
rect -1138 -5423 -1104 -5389
rect -1138 -5491 -1104 -5457
rect -1138 -5559 -1104 -5525
rect -1138 -5627 -1104 -5593
rect -1138 -5695 -1104 -5661
rect -1138 -5763 -1104 -5729
rect -1138 -5831 -1104 -5797
rect -1138 -5899 -1104 -5865
rect -1138 -5967 -1104 -5933
rect -1138 -6035 -1104 -6001
rect -1138 -6103 -1104 -6069
rect -1138 -6171 -1104 -6137
rect -1138 -6239 -1104 -6205
rect -1138 -6307 -1104 -6273
rect -1138 -6375 -1104 -6341
rect -1138 -6443 -1104 -6409
rect -1138 -6511 -1104 -6477
rect -1138 -6579 -1104 -6545
rect -1138 -6647 -1104 -6613
rect -1138 -6715 -1104 -6681
rect -1138 -6783 -1104 -6749
rect -1138 -6851 -1104 -6817
rect -1138 -6919 -1104 -6885
rect -1138 -6987 -1104 -6953
rect -1138 -7055 -1104 -7021
rect -1138 -7123 -1104 -7089
rect -1138 -7191 -1104 -7157
rect -1138 -7259 -1104 -7225
rect -1138 -7327 -1104 -7293
rect -1138 -7395 -1104 -7361
rect -1138 -7463 -1104 -7429
rect -1138 -7531 -1104 -7497
rect -1138 -7599 -1104 -7565
rect -1138 -7667 -1104 -7633
rect -1138 -7735 -1104 -7701
rect -1138 -7803 -1104 -7769
rect -1138 -7871 -1104 -7837
rect -1138 -7939 -1104 -7905
rect -1138 -8007 -1104 -7973
rect -1138 -8075 -1104 -8041
rect -1138 -8143 -1104 -8109
rect -1138 -8211 -1104 -8177
rect -1138 -8279 -1104 -8245
rect -1138 -8347 -1104 -8313
rect -1138 -8415 -1104 -8381
rect -1138 -8483 -1104 -8449
rect -1138 -8551 -1104 -8517
rect -1138 -8619 -1104 -8585
rect -1138 -8687 -1104 -8653
rect -1138 -8755 -1104 -8721
rect -1138 -8823 -1104 -8789
rect -1138 -8891 -1104 -8857
rect -1138 -8959 -1104 -8925
rect -1138 -9027 -1104 -8993
rect -1138 -9095 -1104 -9061
rect -1138 -9163 -1104 -9129
rect -1138 -9231 -1104 -9197
rect -1138 -9299 -1104 -9265
rect -1138 -9367 -1104 -9333
rect -1138 -9435 -1104 -9401
rect -1138 -9503 -1104 -9469
rect -1138 -9571 -1104 -9537
rect -1020 9537 -986 9571
rect -1020 9469 -986 9503
rect -1020 9401 -986 9435
rect -1020 9333 -986 9367
rect -1020 9265 -986 9299
rect -1020 9197 -986 9231
rect -1020 9129 -986 9163
rect -1020 9061 -986 9095
rect -1020 8993 -986 9027
rect -1020 8925 -986 8959
rect -1020 8857 -986 8891
rect -1020 8789 -986 8823
rect -1020 8721 -986 8755
rect -1020 8653 -986 8687
rect -1020 8585 -986 8619
rect -1020 8517 -986 8551
rect -1020 8449 -986 8483
rect -1020 8381 -986 8415
rect -1020 8313 -986 8347
rect -1020 8245 -986 8279
rect -1020 8177 -986 8211
rect -1020 8109 -986 8143
rect -1020 8041 -986 8075
rect -1020 7973 -986 8007
rect -1020 7905 -986 7939
rect -1020 7837 -986 7871
rect -1020 7769 -986 7803
rect -1020 7701 -986 7735
rect -1020 7633 -986 7667
rect -1020 7565 -986 7599
rect -1020 7497 -986 7531
rect -1020 7429 -986 7463
rect -1020 7361 -986 7395
rect -1020 7293 -986 7327
rect -1020 7225 -986 7259
rect -1020 7157 -986 7191
rect -1020 7089 -986 7123
rect -1020 7021 -986 7055
rect -1020 6953 -986 6987
rect -1020 6885 -986 6919
rect -1020 6817 -986 6851
rect -1020 6749 -986 6783
rect -1020 6681 -986 6715
rect -1020 6613 -986 6647
rect -1020 6545 -986 6579
rect -1020 6477 -986 6511
rect -1020 6409 -986 6443
rect -1020 6341 -986 6375
rect -1020 6273 -986 6307
rect -1020 6205 -986 6239
rect -1020 6137 -986 6171
rect -1020 6069 -986 6103
rect -1020 6001 -986 6035
rect -1020 5933 -986 5967
rect -1020 5865 -986 5899
rect -1020 5797 -986 5831
rect -1020 5729 -986 5763
rect -1020 5661 -986 5695
rect -1020 5593 -986 5627
rect -1020 5525 -986 5559
rect -1020 5457 -986 5491
rect -1020 5389 -986 5423
rect -1020 5321 -986 5355
rect -1020 5253 -986 5287
rect -1020 5185 -986 5219
rect -1020 5117 -986 5151
rect -1020 5049 -986 5083
rect -1020 4981 -986 5015
rect -1020 4913 -986 4947
rect -1020 4845 -986 4879
rect -1020 4777 -986 4811
rect -1020 4709 -986 4743
rect -1020 4641 -986 4675
rect -1020 4573 -986 4607
rect -1020 4505 -986 4539
rect -1020 4437 -986 4471
rect -1020 4369 -986 4403
rect -1020 4301 -986 4335
rect -1020 4233 -986 4267
rect -1020 4165 -986 4199
rect -1020 4097 -986 4131
rect -1020 4029 -986 4063
rect -1020 3961 -986 3995
rect -1020 3893 -986 3927
rect -1020 3825 -986 3859
rect -1020 3757 -986 3791
rect -1020 3689 -986 3723
rect -1020 3621 -986 3655
rect -1020 3553 -986 3587
rect -1020 3485 -986 3519
rect -1020 3417 -986 3451
rect -1020 3349 -986 3383
rect -1020 3281 -986 3315
rect -1020 3213 -986 3247
rect -1020 3145 -986 3179
rect -1020 3077 -986 3111
rect -1020 3009 -986 3043
rect -1020 2941 -986 2975
rect -1020 2873 -986 2907
rect -1020 2805 -986 2839
rect -1020 2737 -986 2771
rect -1020 2669 -986 2703
rect -1020 2601 -986 2635
rect -1020 2533 -986 2567
rect -1020 2465 -986 2499
rect -1020 2397 -986 2431
rect -1020 2329 -986 2363
rect -1020 2261 -986 2295
rect -1020 2193 -986 2227
rect -1020 2125 -986 2159
rect -1020 2057 -986 2091
rect -1020 1989 -986 2023
rect -1020 1921 -986 1955
rect -1020 1853 -986 1887
rect -1020 1785 -986 1819
rect -1020 1717 -986 1751
rect -1020 1649 -986 1683
rect -1020 1581 -986 1615
rect -1020 1513 -986 1547
rect -1020 1445 -986 1479
rect -1020 1377 -986 1411
rect -1020 1309 -986 1343
rect -1020 1241 -986 1275
rect -1020 1173 -986 1207
rect -1020 1105 -986 1139
rect -1020 1037 -986 1071
rect -1020 969 -986 1003
rect -1020 901 -986 935
rect -1020 833 -986 867
rect -1020 765 -986 799
rect -1020 697 -986 731
rect -1020 629 -986 663
rect -1020 561 -986 595
rect -1020 493 -986 527
rect -1020 425 -986 459
rect -1020 357 -986 391
rect -1020 289 -986 323
rect -1020 221 -986 255
rect -1020 153 -986 187
rect -1020 85 -986 119
rect -1020 17 -986 51
rect -1020 -51 -986 -17
rect -1020 -119 -986 -85
rect -1020 -187 -986 -153
rect -1020 -255 -986 -221
rect -1020 -323 -986 -289
rect -1020 -391 -986 -357
rect -1020 -459 -986 -425
rect -1020 -527 -986 -493
rect -1020 -595 -986 -561
rect -1020 -663 -986 -629
rect -1020 -731 -986 -697
rect -1020 -799 -986 -765
rect -1020 -867 -986 -833
rect -1020 -935 -986 -901
rect -1020 -1003 -986 -969
rect -1020 -1071 -986 -1037
rect -1020 -1139 -986 -1105
rect -1020 -1207 -986 -1173
rect -1020 -1275 -986 -1241
rect -1020 -1343 -986 -1309
rect -1020 -1411 -986 -1377
rect -1020 -1479 -986 -1445
rect -1020 -1547 -986 -1513
rect -1020 -1615 -986 -1581
rect -1020 -1683 -986 -1649
rect -1020 -1751 -986 -1717
rect -1020 -1819 -986 -1785
rect -1020 -1887 -986 -1853
rect -1020 -1955 -986 -1921
rect -1020 -2023 -986 -1989
rect -1020 -2091 -986 -2057
rect -1020 -2159 -986 -2125
rect -1020 -2227 -986 -2193
rect -1020 -2295 -986 -2261
rect -1020 -2363 -986 -2329
rect -1020 -2431 -986 -2397
rect -1020 -2499 -986 -2465
rect -1020 -2567 -986 -2533
rect -1020 -2635 -986 -2601
rect -1020 -2703 -986 -2669
rect -1020 -2771 -986 -2737
rect -1020 -2839 -986 -2805
rect -1020 -2907 -986 -2873
rect -1020 -2975 -986 -2941
rect -1020 -3043 -986 -3009
rect -1020 -3111 -986 -3077
rect -1020 -3179 -986 -3145
rect -1020 -3247 -986 -3213
rect -1020 -3315 -986 -3281
rect -1020 -3383 -986 -3349
rect -1020 -3451 -986 -3417
rect -1020 -3519 -986 -3485
rect -1020 -3587 -986 -3553
rect -1020 -3655 -986 -3621
rect -1020 -3723 -986 -3689
rect -1020 -3791 -986 -3757
rect -1020 -3859 -986 -3825
rect -1020 -3927 -986 -3893
rect -1020 -3995 -986 -3961
rect -1020 -4063 -986 -4029
rect -1020 -4131 -986 -4097
rect -1020 -4199 -986 -4165
rect -1020 -4267 -986 -4233
rect -1020 -4335 -986 -4301
rect -1020 -4403 -986 -4369
rect -1020 -4471 -986 -4437
rect -1020 -4539 -986 -4505
rect -1020 -4607 -986 -4573
rect -1020 -4675 -986 -4641
rect -1020 -4743 -986 -4709
rect -1020 -4811 -986 -4777
rect -1020 -4879 -986 -4845
rect -1020 -4947 -986 -4913
rect -1020 -5015 -986 -4981
rect -1020 -5083 -986 -5049
rect -1020 -5151 -986 -5117
rect -1020 -5219 -986 -5185
rect -1020 -5287 -986 -5253
rect -1020 -5355 -986 -5321
rect -1020 -5423 -986 -5389
rect -1020 -5491 -986 -5457
rect -1020 -5559 -986 -5525
rect -1020 -5627 -986 -5593
rect -1020 -5695 -986 -5661
rect -1020 -5763 -986 -5729
rect -1020 -5831 -986 -5797
rect -1020 -5899 -986 -5865
rect -1020 -5967 -986 -5933
rect -1020 -6035 -986 -6001
rect -1020 -6103 -986 -6069
rect -1020 -6171 -986 -6137
rect -1020 -6239 -986 -6205
rect -1020 -6307 -986 -6273
rect -1020 -6375 -986 -6341
rect -1020 -6443 -986 -6409
rect -1020 -6511 -986 -6477
rect -1020 -6579 -986 -6545
rect -1020 -6647 -986 -6613
rect -1020 -6715 -986 -6681
rect -1020 -6783 -986 -6749
rect -1020 -6851 -986 -6817
rect -1020 -6919 -986 -6885
rect -1020 -6987 -986 -6953
rect -1020 -7055 -986 -7021
rect -1020 -7123 -986 -7089
rect -1020 -7191 -986 -7157
rect -1020 -7259 -986 -7225
rect -1020 -7327 -986 -7293
rect -1020 -7395 -986 -7361
rect -1020 -7463 -986 -7429
rect -1020 -7531 -986 -7497
rect -1020 -7599 -986 -7565
rect -1020 -7667 -986 -7633
rect -1020 -7735 -986 -7701
rect -1020 -7803 -986 -7769
rect -1020 -7871 -986 -7837
rect -1020 -7939 -986 -7905
rect -1020 -8007 -986 -7973
rect -1020 -8075 -986 -8041
rect -1020 -8143 -986 -8109
rect -1020 -8211 -986 -8177
rect -1020 -8279 -986 -8245
rect -1020 -8347 -986 -8313
rect -1020 -8415 -986 -8381
rect -1020 -8483 -986 -8449
rect -1020 -8551 -986 -8517
rect -1020 -8619 -986 -8585
rect -1020 -8687 -986 -8653
rect -1020 -8755 -986 -8721
rect -1020 -8823 -986 -8789
rect -1020 -8891 -986 -8857
rect -1020 -8959 -986 -8925
rect -1020 -9027 -986 -8993
rect -1020 -9095 -986 -9061
rect -1020 -9163 -986 -9129
rect -1020 -9231 -986 -9197
rect -1020 -9299 -986 -9265
rect -1020 -9367 -986 -9333
rect -1020 -9435 -986 -9401
rect -1020 -9503 -986 -9469
rect -1020 -9571 -986 -9537
rect -902 9537 -868 9571
rect -902 9469 -868 9503
rect -902 9401 -868 9435
rect -902 9333 -868 9367
rect -902 9265 -868 9299
rect -902 9197 -868 9231
rect -902 9129 -868 9163
rect -902 9061 -868 9095
rect -902 8993 -868 9027
rect -902 8925 -868 8959
rect -902 8857 -868 8891
rect -902 8789 -868 8823
rect -902 8721 -868 8755
rect -902 8653 -868 8687
rect -902 8585 -868 8619
rect -902 8517 -868 8551
rect -902 8449 -868 8483
rect -902 8381 -868 8415
rect -902 8313 -868 8347
rect -902 8245 -868 8279
rect -902 8177 -868 8211
rect -902 8109 -868 8143
rect -902 8041 -868 8075
rect -902 7973 -868 8007
rect -902 7905 -868 7939
rect -902 7837 -868 7871
rect -902 7769 -868 7803
rect -902 7701 -868 7735
rect -902 7633 -868 7667
rect -902 7565 -868 7599
rect -902 7497 -868 7531
rect -902 7429 -868 7463
rect -902 7361 -868 7395
rect -902 7293 -868 7327
rect -902 7225 -868 7259
rect -902 7157 -868 7191
rect -902 7089 -868 7123
rect -902 7021 -868 7055
rect -902 6953 -868 6987
rect -902 6885 -868 6919
rect -902 6817 -868 6851
rect -902 6749 -868 6783
rect -902 6681 -868 6715
rect -902 6613 -868 6647
rect -902 6545 -868 6579
rect -902 6477 -868 6511
rect -902 6409 -868 6443
rect -902 6341 -868 6375
rect -902 6273 -868 6307
rect -902 6205 -868 6239
rect -902 6137 -868 6171
rect -902 6069 -868 6103
rect -902 6001 -868 6035
rect -902 5933 -868 5967
rect -902 5865 -868 5899
rect -902 5797 -868 5831
rect -902 5729 -868 5763
rect -902 5661 -868 5695
rect -902 5593 -868 5627
rect -902 5525 -868 5559
rect -902 5457 -868 5491
rect -902 5389 -868 5423
rect -902 5321 -868 5355
rect -902 5253 -868 5287
rect -902 5185 -868 5219
rect -902 5117 -868 5151
rect -902 5049 -868 5083
rect -902 4981 -868 5015
rect -902 4913 -868 4947
rect -902 4845 -868 4879
rect -902 4777 -868 4811
rect -902 4709 -868 4743
rect -902 4641 -868 4675
rect -902 4573 -868 4607
rect -902 4505 -868 4539
rect -902 4437 -868 4471
rect -902 4369 -868 4403
rect -902 4301 -868 4335
rect -902 4233 -868 4267
rect -902 4165 -868 4199
rect -902 4097 -868 4131
rect -902 4029 -868 4063
rect -902 3961 -868 3995
rect -902 3893 -868 3927
rect -902 3825 -868 3859
rect -902 3757 -868 3791
rect -902 3689 -868 3723
rect -902 3621 -868 3655
rect -902 3553 -868 3587
rect -902 3485 -868 3519
rect -902 3417 -868 3451
rect -902 3349 -868 3383
rect -902 3281 -868 3315
rect -902 3213 -868 3247
rect -902 3145 -868 3179
rect -902 3077 -868 3111
rect -902 3009 -868 3043
rect -902 2941 -868 2975
rect -902 2873 -868 2907
rect -902 2805 -868 2839
rect -902 2737 -868 2771
rect -902 2669 -868 2703
rect -902 2601 -868 2635
rect -902 2533 -868 2567
rect -902 2465 -868 2499
rect -902 2397 -868 2431
rect -902 2329 -868 2363
rect -902 2261 -868 2295
rect -902 2193 -868 2227
rect -902 2125 -868 2159
rect -902 2057 -868 2091
rect -902 1989 -868 2023
rect -902 1921 -868 1955
rect -902 1853 -868 1887
rect -902 1785 -868 1819
rect -902 1717 -868 1751
rect -902 1649 -868 1683
rect -902 1581 -868 1615
rect -902 1513 -868 1547
rect -902 1445 -868 1479
rect -902 1377 -868 1411
rect -902 1309 -868 1343
rect -902 1241 -868 1275
rect -902 1173 -868 1207
rect -902 1105 -868 1139
rect -902 1037 -868 1071
rect -902 969 -868 1003
rect -902 901 -868 935
rect -902 833 -868 867
rect -902 765 -868 799
rect -902 697 -868 731
rect -902 629 -868 663
rect -902 561 -868 595
rect -902 493 -868 527
rect -902 425 -868 459
rect -902 357 -868 391
rect -902 289 -868 323
rect -902 221 -868 255
rect -902 153 -868 187
rect -902 85 -868 119
rect -902 17 -868 51
rect -902 -51 -868 -17
rect -902 -119 -868 -85
rect -902 -187 -868 -153
rect -902 -255 -868 -221
rect -902 -323 -868 -289
rect -902 -391 -868 -357
rect -902 -459 -868 -425
rect -902 -527 -868 -493
rect -902 -595 -868 -561
rect -902 -663 -868 -629
rect -902 -731 -868 -697
rect -902 -799 -868 -765
rect -902 -867 -868 -833
rect -902 -935 -868 -901
rect -902 -1003 -868 -969
rect -902 -1071 -868 -1037
rect -902 -1139 -868 -1105
rect -902 -1207 -868 -1173
rect -902 -1275 -868 -1241
rect -902 -1343 -868 -1309
rect -902 -1411 -868 -1377
rect -902 -1479 -868 -1445
rect -902 -1547 -868 -1513
rect -902 -1615 -868 -1581
rect -902 -1683 -868 -1649
rect -902 -1751 -868 -1717
rect -902 -1819 -868 -1785
rect -902 -1887 -868 -1853
rect -902 -1955 -868 -1921
rect -902 -2023 -868 -1989
rect -902 -2091 -868 -2057
rect -902 -2159 -868 -2125
rect -902 -2227 -868 -2193
rect -902 -2295 -868 -2261
rect -902 -2363 -868 -2329
rect -902 -2431 -868 -2397
rect -902 -2499 -868 -2465
rect -902 -2567 -868 -2533
rect -902 -2635 -868 -2601
rect -902 -2703 -868 -2669
rect -902 -2771 -868 -2737
rect -902 -2839 -868 -2805
rect -902 -2907 -868 -2873
rect -902 -2975 -868 -2941
rect -902 -3043 -868 -3009
rect -902 -3111 -868 -3077
rect -902 -3179 -868 -3145
rect -902 -3247 -868 -3213
rect -902 -3315 -868 -3281
rect -902 -3383 -868 -3349
rect -902 -3451 -868 -3417
rect -902 -3519 -868 -3485
rect -902 -3587 -868 -3553
rect -902 -3655 -868 -3621
rect -902 -3723 -868 -3689
rect -902 -3791 -868 -3757
rect -902 -3859 -868 -3825
rect -902 -3927 -868 -3893
rect -902 -3995 -868 -3961
rect -902 -4063 -868 -4029
rect -902 -4131 -868 -4097
rect -902 -4199 -868 -4165
rect -902 -4267 -868 -4233
rect -902 -4335 -868 -4301
rect -902 -4403 -868 -4369
rect -902 -4471 -868 -4437
rect -902 -4539 -868 -4505
rect -902 -4607 -868 -4573
rect -902 -4675 -868 -4641
rect -902 -4743 -868 -4709
rect -902 -4811 -868 -4777
rect -902 -4879 -868 -4845
rect -902 -4947 -868 -4913
rect -902 -5015 -868 -4981
rect -902 -5083 -868 -5049
rect -902 -5151 -868 -5117
rect -902 -5219 -868 -5185
rect -902 -5287 -868 -5253
rect -902 -5355 -868 -5321
rect -902 -5423 -868 -5389
rect -902 -5491 -868 -5457
rect -902 -5559 -868 -5525
rect -902 -5627 -868 -5593
rect -902 -5695 -868 -5661
rect -902 -5763 -868 -5729
rect -902 -5831 -868 -5797
rect -902 -5899 -868 -5865
rect -902 -5967 -868 -5933
rect -902 -6035 -868 -6001
rect -902 -6103 -868 -6069
rect -902 -6171 -868 -6137
rect -902 -6239 -868 -6205
rect -902 -6307 -868 -6273
rect -902 -6375 -868 -6341
rect -902 -6443 -868 -6409
rect -902 -6511 -868 -6477
rect -902 -6579 -868 -6545
rect -902 -6647 -868 -6613
rect -902 -6715 -868 -6681
rect -902 -6783 -868 -6749
rect -902 -6851 -868 -6817
rect -902 -6919 -868 -6885
rect -902 -6987 -868 -6953
rect -902 -7055 -868 -7021
rect -902 -7123 -868 -7089
rect -902 -7191 -868 -7157
rect -902 -7259 -868 -7225
rect -902 -7327 -868 -7293
rect -902 -7395 -868 -7361
rect -902 -7463 -868 -7429
rect -902 -7531 -868 -7497
rect -902 -7599 -868 -7565
rect -902 -7667 -868 -7633
rect -902 -7735 -868 -7701
rect -902 -7803 -868 -7769
rect -902 -7871 -868 -7837
rect -902 -7939 -868 -7905
rect -902 -8007 -868 -7973
rect -902 -8075 -868 -8041
rect -902 -8143 -868 -8109
rect -902 -8211 -868 -8177
rect -902 -8279 -868 -8245
rect -902 -8347 -868 -8313
rect -902 -8415 -868 -8381
rect -902 -8483 -868 -8449
rect -902 -8551 -868 -8517
rect -902 -8619 -868 -8585
rect -902 -8687 -868 -8653
rect -902 -8755 -868 -8721
rect -902 -8823 -868 -8789
rect -902 -8891 -868 -8857
rect -902 -8959 -868 -8925
rect -902 -9027 -868 -8993
rect -902 -9095 -868 -9061
rect -902 -9163 -868 -9129
rect -902 -9231 -868 -9197
rect -902 -9299 -868 -9265
rect -902 -9367 -868 -9333
rect -902 -9435 -868 -9401
rect -902 -9503 -868 -9469
rect -902 -9571 -868 -9537
rect -784 9537 -750 9571
rect -784 9469 -750 9503
rect -784 9401 -750 9435
rect -784 9333 -750 9367
rect -784 9265 -750 9299
rect -784 9197 -750 9231
rect -784 9129 -750 9163
rect -784 9061 -750 9095
rect -784 8993 -750 9027
rect -784 8925 -750 8959
rect -784 8857 -750 8891
rect -784 8789 -750 8823
rect -784 8721 -750 8755
rect -784 8653 -750 8687
rect -784 8585 -750 8619
rect -784 8517 -750 8551
rect -784 8449 -750 8483
rect -784 8381 -750 8415
rect -784 8313 -750 8347
rect -784 8245 -750 8279
rect -784 8177 -750 8211
rect -784 8109 -750 8143
rect -784 8041 -750 8075
rect -784 7973 -750 8007
rect -784 7905 -750 7939
rect -784 7837 -750 7871
rect -784 7769 -750 7803
rect -784 7701 -750 7735
rect -784 7633 -750 7667
rect -784 7565 -750 7599
rect -784 7497 -750 7531
rect -784 7429 -750 7463
rect -784 7361 -750 7395
rect -784 7293 -750 7327
rect -784 7225 -750 7259
rect -784 7157 -750 7191
rect -784 7089 -750 7123
rect -784 7021 -750 7055
rect -784 6953 -750 6987
rect -784 6885 -750 6919
rect -784 6817 -750 6851
rect -784 6749 -750 6783
rect -784 6681 -750 6715
rect -784 6613 -750 6647
rect -784 6545 -750 6579
rect -784 6477 -750 6511
rect -784 6409 -750 6443
rect -784 6341 -750 6375
rect -784 6273 -750 6307
rect -784 6205 -750 6239
rect -784 6137 -750 6171
rect -784 6069 -750 6103
rect -784 6001 -750 6035
rect -784 5933 -750 5967
rect -784 5865 -750 5899
rect -784 5797 -750 5831
rect -784 5729 -750 5763
rect -784 5661 -750 5695
rect -784 5593 -750 5627
rect -784 5525 -750 5559
rect -784 5457 -750 5491
rect -784 5389 -750 5423
rect -784 5321 -750 5355
rect -784 5253 -750 5287
rect -784 5185 -750 5219
rect -784 5117 -750 5151
rect -784 5049 -750 5083
rect -784 4981 -750 5015
rect -784 4913 -750 4947
rect -784 4845 -750 4879
rect -784 4777 -750 4811
rect -784 4709 -750 4743
rect -784 4641 -750 4675
rect -784 4573 -750 4607
rect -784 4505 -750 4539
rect -784 4437 -750 4471
rect -784 4369 -750 4403
rect -784 4301 -750 4335
rect -784 4233 -750 4267
rect -784 4165 -750 4199
rect -784 4097 -750 4131
rect -784 4029 -750 4063
rect -784 3961 -750 3995
rect -784 3893 -750 3927
rect -784 3825 -750 3859
rect -784 3757 -750 3791
rect -784 3689 -750 3723
rect -784 3621 -750 3655
rect -784 3553 -750 3587
rect -784 3485 -750 3519
rect -784 3417 -750 3451
rect -784 3349 -750 3383
rect -784 3281 -750 3315
rect -784 3213 -750 3247
rect -784 3145 -750 3179
rect -784 3077 -750 3111
rect -784 3009 -750 3043
rect -784 2941 -750 2975
rect -784 2873 -750 2907
rect -784 2805 -750 2839
rect -784 2737 -750 2771
rect -784 2669 -750 2703
rect -784 2601 -750 2635
rect -784 2533 -750 2567
rect -784 2465 -750 2499
rect -784 2397 -750 2431
rect -784 2329 -750 2363
rect -784 2261 -750 2295
rect -784 2193 -750 2227
rect -784 2125 -750 2159
rect -784 2057 -750 2091
rect -784 1989 -750 2023
rect -784 1921 -750 1955
rect -784 1853 -750 1887
rect -784 1785 -750 1819
rect -784 1717 -750 1751
rect -784 1649 -750 1683
rect -784 1581 -750 1615
rect -784 1513 -750 1547
rect -784 1445 -750 1479
rect -784 1377 -750 1411
rect -784 1309 -750 1343
rect -784 1241 -750 1275
rect -784 1173 -750 1207
rect -784 1105 -750 1139
rect -784 1037 -750 1071
rect -784 969 -750 1003
rect -784 901 -750 935
rect -784 833 -750 867
rect -784 765 -750 799
rect -784 697 -750 731
rect -784 629 -750 663
rect -784 561 -750 595
rect -784 493 -750 527
rect -784 425 -750 459
rect -784 357 -750 391
rect -784 289 -750 323
rect -784 221 -750 255
rect -784 153 -750 187
rect -784 85 -750 119
rect -784 17 -750 51
rect -784 -51 -750 -17
rect -784 -119 -750 -85
rect -784 -187 -750 -153
rect -784 -255 -750 -221
rect -784 -323 -750 -289
rect -784 -391 -750 -357
rect -784 -459 -750 -425
rect -784 -527 -750 -493
rect -784 -595 -750 -561
rect -784 -663 -750 -629
rect -784 -731 -750 -697
rect -784 -799 -750 -765
rect -784 -867 -750 -833
rect -784 -935 -750 -901
rect -784 -1003 -750 -969
rect -784 -1071 -750 -1037
rect -784 -1139 -750 -1105
rect -784 -1207 -750 -1173
rect -784 -1275 -750 -1241
rect -784 -1343 -750 -1309
rect -784 -1411 -750 -1377
rect -784 -1479 -750 -1445
rect -784 -1547 -750 -1513
rect -784 -1615 -750 -1581
rect -784 -1683 -750 -1649
rect -784 -1751 -750 -1717
rect -784 -1819 -750 -1785
rect -784 -1887 -750 -1853
rect -784 -1955 -750 -1921
rect -784 -2023 -750 -1989
rect -784 -2091 -750 -2057
rect -784 -2159 -750 -2125
rect -784 -2227 -750 -2193
rect -784 -2295 -750 -2261
rect -784 -2363 -750 -2329
rect -784 -2431 -750 -2397
rect -784 -2499 -750 -2465
rect -784 -2567 -750 -2533
rect -784 -2635 -750 -2601
rect -784 -2703 -750 -2669
rect -784 -2771 -750 -2737
rect -784 -2839 -750 -2805
rect -784 -2907 -750 -2873
rect -784 -2975 -750 -2941
rect -784 -3043 -750 -3009
rect -784 -3111 -750 -3077
rect -784 -3179 -750 -3145
rect -784 -3247 -750 -3213
rect -784 -3315 -750 -3281
rect -784 -3383 -750 -3349
rect -784 -3451 -750 -3417
rect -784 -3519 -750 -3485
rect -784 -3587 -750 -3553
rect -784 -3655 -750 -3621
rect -784 -3723 -750 -3689
rect -784 -3791 -750 -3757
rect -784 -3859 -750 -3825
rect -784 -3927 -750 -3893
rect -784 -3995 -750 -3961
rect -784 -4063 -750 -4029
rect -784 -4131 -750 -4097
rect -784 -4199 -750 -4165
rect -784 -4267 -750 -4233
rect -784 -4335 -750 -4301
rect -784 -4403 -750 -4369
rect -784 -4471 -750 -4437
rect -784 -4539 -750 -4505
rect -784 -4607 -750 -4573
rect -784 -4675 -750 -4641
rect -784 -4743 -750 -4709
rect -784 -4811 -750 -4777
rect -784 -4879 -750 -4845
rect -784 -4947 -750 -4913
rect -784 -5015 -750 -4981
rect -784 -5083 -750 -5049
rect -784 -5151 -750 -5117
rect -784 -5219 -750 -5185
rect -784 -5287 -750 -5253
rect -784 -5355 -750 -5321
rect -784 -5423 -750 -5389
rect -784 -5491 -750 -5457
rect -784 -5559 -750 -5525
rect -784 -5627 -750 -5593
rect -784 -5695 -750 -5661
rect -784 -5763 -750 -5729
rect -784 -5831 -750 -5797
rect -784 -5899 -750 -5865
rect -784 -5967 -750 -5933
rect -784 -6035 -750 -6001
rect -784 -6103 -750 -6069
rect -784 -6171 -750 -6137
rect -784 -6239 -750 -6205
rect -784 -6307 -750 -6273
rect -784 -6375 -750 -6341
rect -784 -6443 -750 -6409
rect -784 -6511 -750 -6477
rect -784 -6579 -750 -6545
rect -784 -6647 -750 -6613
rect -784 -6715 -750 -6681
rect -784 -6783 -750 -6749
rect -784 -6851 -750 -6817
rect -784 -6919 -750 -6885
rect -784 -6987 -750 -6953
rect -784 -7055 -750 -7021
rect -784 -7123 -750 -7089
rect -784 -7191 -750 -7157
rect -784 -7259 -750 -7225
rect -784 -7327 -750 -7293
rect -784 -7395 -750 -7361
rect -784 -7463 -750 -7429
rect -784 -7531 -750 -7497
rect -784 -7599 -750 -7565
rect -784 -7667 -750 -7633
rect -784 -7735 -750 -7701
rect -784 -7803 -750 -7769
rect -784 -7871 -750 -7837
rect -784 -7939 -750 -7905
rect -784 -8007 -750 -7973
rect -784 -8075 -750 -8041
rect -784 -8143 -750 -8109
rect -784 -8211 -750 -8177
rect -784 -8279 -750 -8245
rect -784 -8347 -750 -8313
rect -784 -8415 -750 -8381
rect -784 -8483 -750 -8449
rect -784 -8551 -750 -8517
rect -784 -8619 -750 -8585
rect -784 -8687 -750 -8653
rect -784 -8755 -750 -8721
rect -784 -8823 -750 -8789
rect -784 -8891 -750 -8857
rect -784 -8959 -750 -8925
rect -784 -9027 -750 -8993
rect -784 -9095 -750 -9061
rect -784 -9163 -750 -9129
rect -784 -9231 -750 -9197
rect -784 -9299 -750 -9265
rect -784 -9367 -750 -9333
rect -784 -9435 -750 -9401
rect -784 -9503 -750 -9469
rect -784 -9571 -750 -9537
rect -666 9537 -632 9571
rect -666 9469 -632 9503
rect -666 9401 -632 9435
rect -666 9333 -632 9367
rect -666 9265 -632 9299
rect -666 9197 -632 9231
rect -666 9129 -632 9163
rect -666 9061 -632 9095
rect -666 8993 -632 9027
rect -666 8925 -632 8959
rect -666 8857 -632 8891
rect -666 8789 -632 8823
rect -666 8721 -632 8755
rect -666 8653 -632 8687
rect -666 8585 -632 8619
rect -666 8517 -632 8551
rect -666 8449 -632 8483
rect -666 8381 -632 8415
rect -666 8313 -632 8347
rect -666 8245 -632 8279
rect -666 8177 -632 8211
rect -666 8109 -632 8143
rect -666 8041 -632 8075
rect -666 7973 -632 8007
rect -666 7905 -632 7939
rect -666 7837 -632 7871
rect -666 7769 -632 7803
rect -666 7701 -632 7735
rect -666 7633 -632 7667
rect -666 7565 -632 7599
rect -666 7497 -632 7531
rect -666 7429 -632 7463
rect -666 7361 -632 7395
rect -666 7293 -632 7327
rect -666 7225 -632 7259
rect -666 7157 -632 7191
rect -666 7089 -632 7123
rect -666 7021 -632 7055
rect -666 6953 -632 6987
rect -666 6885 -632 6919
rect -666 6817 -632 6851
rect -666 6749 -632 6783
rect -666 6681 -632 6715
rect -666 6613 -632 6647
rect -666 6545 -632 6579
rect -666 6477 -632 6511
rect -666 6409 -632 6443
rect -666 6341 -632 6375
rect -666 6273 -632 6307
rect -666 6205 -632 6239
rect -666 6137 -632 6171
rect -666 6069 -632 6103
rect -666 6001 -632 6035
rect -666 5933 -632 5967
rect -666 5865 -632 5899
rect -666 5797 -632 5831
rect -666 5729 -632 5763
rect -666 5661 -632 5695
rect -666 5593 -632 5627
rect -666 5525 -632 5559
rect -666 5457 -632 5491
rect -666 5389 -632 5423
rect -666 5321 -632 5355
rect -666 5253 -632 5287
rect -666 5185 -632 5219
rect -666 5117 -632 5151
rect -666 5049 -632 5083
rect -666 4981 -632 5015
rect -666 4913 -632 4947
rect -666 4845 -632 4879
rect -666 4777 -632 4811
rect -666 4709 -632 4743
rect -666 4641 -632 4675
rect -666 4573 -632 4607
rect -666 4505 -632 4539
rect -666 4437 -632 4471
rect -666 4369 -632 4403
rect -666 4301 -632 4335
rect -666 4233 -632 4267
rect -666 4165 -632 4199
rect -666 4097 -632 4131
rect -666 4029 -632 4063
rect -666 3961 -632 3995
rect -666 3893 -632 3927
rect -666 3825 -632 3859
rect -666 3757 -632 3791
rect -666 3689 -632 3723
rect -666 3621 -632 3655
rect -666 3553 -632 3587
rect -666 3485 -632 3519
rect -666 3417 -632 3451
rect -666 3349 -632 3383
rect -666 3281 -632 3315
rect -666 3213 -632 3247
rect -666 3145 -632 3179
rect -666 3077 -632 3111
rect -666 3009 -632 3043
rect -666 2941 -632 2975
rect -666 2873 -632 2907
rect -666 2805 -632 2839
rect -666 2737 -632 2771
rect -666 2669 -632 2703
rect -666 2601 -632 2635
rect -666 2533 -632 2567
rect -666 2465 -632 2499
rect -666 2397 -632 2431
rect -666 2329 -632 2363
rect -666 2261 -632 2295
rect -666 2193 -632 2227
rect -666 2125 -632 2159
rect -666 2057 -632 2091
rect -666 1989 -632 2023
rect -666 1921 -632 1955
rect -666 1853 -632 1887
rect -666 1785 -632 1819
rect -666 1717 -632 1751
rect -666 1649 -632 1683
rect -666 1581 -632 1615
rect -666 1513 -632 1547
rect -666 1445 -632 1479
rect -666 1377 -632 1411
rect -666 1309 -632 1343
rect -666 1241 -632 1275
rect -666 1173 -632 1207
rect -666 1105 -632 1139
rect -666 1037 -632 1071
rect -666 969 -632 1003
rect -666 901 -632 935
rect -666 833 -632 867
rect -666 765 -632 799
rect -666 697 -632 731
rect -666 629 -632 663
rect -666 561 -632 595
rect -666 493 -632 527
rect -666 425 -632 459
rect -666 357 -632 391
rect -666 289 -632 323
rect -666 221 -632 255
rect -666 153 -632 187
rect -666 85 -632 119
rect -666 17 -632 51
rect -666 -51 -632 -17
rect -666 -119 -632 -85
rect -666 -187 -632 -153
rect -666 -255 -632 -221
rect -666 -323 -632 -289
rect -666 -391 -632 -357
rect -666 -459 -632 -425
rect -666 -527 -632 -493
rect -666 -595 -632 -561
rect -666 -663 -632 -629
rect -666 -731 -632 -697
rect -666 -799 -632 -765
rect -666 -867 -632 -833
rect -666 -935 -632 -901
rect -666 -1003 -632 -969
rect -666 -1071 -632 -1037
rect -666 -1139 -632 -1105
rect -666 -1207 -632 -1173
rect -666 -1275 -632 -1241
rect -666 -1343 -632 -1309
rect -666 -1411 -632 -1377
rect -666 -1479 -632 -1445
rect -666 -1547 -632 -1513
rect -666 -1615 -632 -1581
rect -666 -1683 -632 -1649
rect -666 -1751 -632 -1717
rect -666 -1819 -632 -1785
rect -666 -1887 -632 -1853
rect -666 -1955 -632 -1921
rect -666 -2023 -632 -1989
rect -666 -2091 -632 -2057
rect -666 -2159 -632 -2125
rect -666 -2227 -632 -2193
rect -666 -2295 -632 -2261
rect -666 -2363 -632 -2329
rect -666 -2431 -632 -2397
rect -666 -2499 -632 -2465
rect -666 -2567 -632 -2533
rect -666 -2635 -632 -2601
rect -666 -2703 -632 -2669
rect -666 -2771 -632 -2737
rect -666 -2839 -632 -2805
rect -666 -2907 -632 -2873
rect -666 -2975 -632 -2941
rect -666 -3043 -632 -3009
rect -666 -3111 -632 -3077
rect -666 -3179 -632 -3145
rect -666 -3247 -632 -3213
rect -666 -3315 -632 -3281
rect -666 -3383 -632 -3349
rect -666 -3451 -632 -3417
rect -666 -3519 -632 -3485
rect -666 -3587 -632 -3553
rect -666 -3655 -632 -3621
rect -666 -3723 -632 -3689
rect -666 -3791 -632 -3757
rect -666 -3859 -632 -3825
rect -666 -3927 -632 -3893
rect -666 -3995 -632 -3961
rect -666 -4063 -632 -4029
rect -666 -4131 -632 -4097
rect -666 -4199 -632 -4165
rect -666 -4267 -632 -4233
rect -666 -4335 -632 -4301
rect -666 -4403 -632 -4369
rect -666 -4471 -632 -4437
rect -666 -4539 -632 -4505
rect -666 -4607 -632 -4573
rect -666 -4675 -632 -4641
rect -666 -4743 -632 -4709
rect -666 -4811 -632 -4777
rect -666 -4879 -632 -4845
rect -666 -4947 -632 -4913
rect -666 -5015 -632 -4981
rect -666 -5083 -632 -5049
rect -666 -5151 -632 -5117
rect -666 -5219 -632 -5185
rect -666 -5287 -632 -5253
rect -666 -5355 -632 -5321
rect -666 -5423 -632 -5389
rect -666 -5491 -632 -5457
rect -666 -5559 -632 -5525
rect -666 -5627 -632 -5593
rect -666 -5695 -632 -5661
rect -666 -5763 -632 -5729
rect -666 -5831 -632 -5797
rect -666 -5899 -632 -5865
rect -666 -5967 -632 -5933
rect -666 -6035 -632 -6001
rect -666 -6103 -632 -6069
rect -666 -6171 -632 -6137
rect -666 -6239 -632 -6205
rect -666 -6307 -632 -6273
rect -666 -6375 -632 -6341
rect -666 -6443 -632 -6409
rect -666 -6511 -632 -6477
rect -666 -6579 -632 -6545
rect -666 -6647 -632 -6613
rect -666 -6715 -632 -6681
rect -666 -6783 -632 -6749
rect -666 -6851 -632 -6817
rect -666 -6919 -632 -6885
rect -666 -6987 -632 -6953
rect -666 -7055 -632 -7021
rect -666 -7123 -632 -7089
rect -666 -7191 -632 -7157
rect -666 -7259 -632 -7225
rect -666 -7327 -632 -7293
rect -666 -7395 -632 -7361
rect -666 -7463 -632 -7429
rect -666 -7531 -632 -7497
rect -666 -7599 -632 -7565
rect -666 -7667 -632 -7633
rect -666 -7735 -632 -7701
rect -666 -7803 -632 -7769
rect -666 -7871 -632 -7837
rect -666 -7939 -632 -7905
rect -666 -8007 -632 -7973
rect -666 -8075 -632 -8041
rect -666 -8143 -632 -8109
rect -666 -8211 -632 -8177
rect -666 -8279 -632 -8245
rect -666 -8347 -632 -8313
rect -666 -8415 -632 -8381
rect -666 -8483 -632 -8449
rect -666 -8551 -632 -8517
rect -666 -8619 -632 -8585
rect -666 -8687 -632 -8653
rect -666 -8755 -632 -8721
rect -666 -8823 -632 -8789
rect -666 -8891 -632 -8857
rect -666 -8959 -632 -8925
rect -666 -9027 -632 -8993
rect -666 -9095 -632 -9061
rect -666 -9163 -632 -9129
rect -666 -9231 -632 -9197
rect -666 -9299 -632 -9265
rect -666 -9367 -632 -9333
rect -666 -9435 -632 -9401
rect -666 -9503 -632 -9469
rect -666 -9571 -632 -9537
rect -548 9537 -514 9571
rect -548 9469 -514 9503
rect -548 9401 -514 9435
rect -548 9333 -514 9367
rect -548 9265 -514 9299
rect -548 9197 -514 9231
rect -548 9129 -514 9163
rect -548 9061 -514 9095
rect -548 8993 -514 9027
rect -548 8925 -514 8959
rect -548 8857 -514 8891
rect -548 8789 -514 8823
rect -548 8721 -514 8755
rect -548 8653 -514 8687
rect -548 8585 -514 8619
rect -548 8517 -514 8551
rect -548 8449 -514 8483
rect -548 8381 -514 8415
rect -548 8313 -514 8347
rect -548 8245 -514 8279
rect -548 8177 -514 8211
rect -548 8109 -514 8143
rect -548 8041 -514 8075
rect -548 7973 -514 8007
rect -548 7905 -514 7939
rect -548 7837 -514 7871
rect -548 7769 -514 7803
rect -548 7701 -514 7735
rect -548 7633 -514 7667
rect -548 7565 -514 7599
rect -548 7497 -514 7531
rect -548 7429 -514 7463
rect -548 7361 -514 7395
rect -548 7293 -514 7327
rect -548 7225 -514 7259
rect -548 7157 -514 7191
rect -548 7089 -514 7123
rect -548 7021 -514 7055
rect -548 6953 -514 6987
rect -548 6885 -514 6919
rect -548 6817 -514 6851
rect -548 6749 -514 6783
rect -548 6681 -514 6715
rect -548 6613 -514 6647
rect -548 6545 -514 6579
rect -548 6477 -514 6511
rect -548 6409 -514 6443
rect -548 6341 -514 6375
rect -548 6273 -514 6307
rect -548 6205 -514 6239
rect -548 6137 -514 6171
rect -548 6069 -514 6103
rect -548 6001 -514 6035
rect -548 5933 -514 5967
rect -548 5865 -514 5899
rect -548 5797 -514 5831
rect -548 5729 -514 5763
rect -548 5661 -514 5695
rect -548 5593 -514 5627
rect -548 5525 -514 5559
rect -548 5457 -514 5491
rect -548 5389 -514 5423
rect -548 5321 -514 5355
rect -548 5253 -514 5287
rect -548 5185 -514 5219
rect -548 5117 -514 5151
rect -548 5049 -514 5083
rect -548 4981 -514 5015
rect -548 4913 -514 4947
rect -548 4845 -514 4879
rect -548 4777 -514 4811
rect -548 4709 -514 4743
rect -548 4641 -514 4675
rect -548 4573 -514 4607
rect -548 4505 -514 4539
rect -548 4437 -514 4471
rect -548 4369 -514 4403
rect -548 4301 -514 4335
rect -548 4233 -514 4267
rect -548 4165 -514 4199
rect -548 4097 -514 4131
rect -548 4029 -514 4063
rect -548 3961 -514 3995
rect -548 3893 -514 3927
rect -548 3825 -514 3859
rect -548 3757 -514 3791
rect -548 3689 -514 3723
rect -548 3621 -514 3655
rect -548 3553 -514 3587
rect -548 3485 -514 3519
rect -548 3417 -514 3451
rect -548 3349 -514 3383
rect -548 3281 -514 3315
rect -548 3213 -514 3247
rect -548 3145 -514 3179
rect -548 3077 -514 3111
rect -548 3009 -514 3043
rect -548 2941 -514 2975
rect -548 2873 -514 2907
rect -548 2805 -514 2839
rect -548 2737 -514 2771
rect -548 2669 -514 2703
rect -548 2601 -514 2635
rect -548 2533 -514 2567
rect -548 2465 -514 2499
rect -548 2397 -514 2431
rect -548 2329 -514 2363
rect -548 2261 -514 2295
rect -548 2193 -514 2227
rect -548 2125 -514 2159
rect -548 2057 -514 2091
rect -548 1989 -514 2023
rect -548 1921 -514 1955
rect -548 1853 -514 1887
rect -548 1785 -514 1819
rect -548 1717 -514 1751
rect -548 1649 -514 1683
rect -548 1581 -514 1615
rect -548 1513 -514 1547
rect -548 1445 -514 1479
rect -548 1377 -514 1411
rect -548 1309 -514 1343
rect -548 1241 -514 1275
rect -548 1173 -514 1207
rect -548 1105 -514 1139
rect -548 1037 -514 1071
rect -548 969 -514 1003
rect -548 901 -514 935
rect -548 833 -514 867
rect -548 765 -514 799
rect -548 697 -514 731
rect -548 629 -514 663
rect -548 561 -514 595
rect -548 493 -514 527
rect -548 425 -514 459
rect -548 357 -514 391
rect -548 289 -514 323
rect -548 221 -514 255
rect -548 153 -514 187
rect -548 85 -514 119
rect -548 17 -514 51
rect -548 -51 -514 -17
rect -548 -119 -514 -85
rect -548 -187 -514 -153
rect -548 -255 -514 -221
rect -548 -323 -514 -289
rect -548 -391 -514 -357
rect -548 -459 -514 -425
rect -548 -527 -514 -493
rect -548 -595 -514 -561
rect -548 -663 -514 -629
rect -548 -731 -514 -697
rect -548 -799 -514 -765
rect -548 -867 -514 -833
rect -548 -935 -514 -901
rect -548 -1003 -514 -969
rect -548 -1071 -514 -1037
rect -548 -1139 -514 -1105
rect -548 -1207 -514 -1173
rect -548 -1275 -514 -1241
rect -548 -1343 -514 -1309
rect -548 -1411 -514 -1377
rect -548 -1479 -514 -1445
rect -548 -1547 -514 -1513
rect -548 -1615 -514 -1581
rect -548 -1683 -514 -1649
rect -548 -1751 -514 -1717
rect -548 -1819 -514 -1785
rect -548 -1887 -514 -1853
rect -548 -1955 -514 -1921
rect -548 -2023 -514 -1989
rect -548 -2091 -514 -2057
rect -548 -2159 -514 -2125
rect -548 -2227 -514 -2193
rect -548 -2295 -514 -2261
rect -548 -2363 -514 -2329
rect -548 -2431 -514 -2397
rect -548 -2499 -514 -2465
rect -548 -2567 -514 -2533
rect -548 -2635 -514 -2601
rect -548 -2703 -514 -2669
rect -548 -2771 -514 -2737
rect -548 -2839 -514 -2805
rect -548 -2907 -514 -2873
rect -548 -2975 -514 -2941
rect -548 -3043 -514 -3009
rect -548 -3111 -514 -3077
rect -548 -3179 -514 -3145
rect -548 -3247 -514 -3213
rect -548 -3315 -514 -3281
rect -548 -3383 -514 -3349
rect -548 -3451 -514 -3417
rect -548 -3519 -514 -3485
rect -548 -3587 -514 -3553
rect -548 -3655 -514 -3621
rect -548 -3723 -514 -3689
rect -548 -3791 -514 -3757
rect -548 -3859 -514 -3825
rect -548 -3927 -514 -3893
rect -548 -3995 -514 -3961
rect -548 -4063 -514 -4029
rect -548 -4131 -514 -4097
rect -548 -4199 -514 -4165
rect -548 -4267 -514 -4233
rect -548 -4335 -514 -4301
rect -548 -4403 -514 -4369
rect -548 -4471 -514 -4437
rect -548 -4539 -514 -4505
rect -548 -4607 -514 -4573
rect -548 -4675 -514 -4641
rect -548 -4743 -514 -4709
rect -548 -4811 -514 -4777
rect -548 -4879 -514 -4845
rect -548 -4947 -514 -4913
rect -548 -5015 -514 -4981
rect -548 -5083 -514 -5049
rect -548 -5151 -514 -5117
rect -548 -5219 -514 -5185
rect -548 -5287 -514 -5253
rect -548 -5355 -514 -5321
rect -548 -5423 -514 -5389
rect -548 -5491 -514 -5457
rect -548 -5559 -514 -5525
rect -548 -5627 -514 -5593
rect -548 -5695 -514 -5661
rect -548 -5763 -514 -5729
rect -548 -5831 -514 -5797
rect -548 -5899 -514 -5865
rect -548 -5967 -514 -5933
rect -548 -6035 -514 -6001
rect -548 -6103 -514 -6069
rect -548 -6171 -514 -6137
rect -548 -6239 -514 -6205
rect -548 -6307 -514 -6273
rect -548 -6375 -514 -6341
rect -548 -6443 -514 -6409
rect -548 -6511 -514 -6477
rect -548 -6579 -514 -6545
rect -548 -6647 -514 -6613
rect -548 -6715 -514 -6681
rect -548 -6783 -514 -6749
rect -548 -6851 -514 -6817
rect -548 -6919 -514 -6885
rect -548 -6987 -514 -6953
rect -548 -7055 -514 -7021
rect -548 -7123 -514 -7089
rect -548 -7191 -514 -7157
rect -548 -7259 -514 -7225
rect -548 -7327 -514 -7293
rect -548 -7395 -514 -7361
rect -548 -7463 -514 -7429
rect -548 -7531 -514 -7497
rect -548 -7599 -514 -7565
rect -548 -7667 -514 -7633
rect -548 -7735 -514 -7701
rect -548 -7803 -514 -7769
rect -548 -7871 -514 -7837
rect -548 -7939 -514 -7905
rect -548 -8007 -514 -7973
rect -548 -8075 -514 -8041
rect -548 -8143 -514 -8109
rect -548 -8211 -514 -8177
rect -548 -8279 -514 -8245
rect -548 -8347 -514 -8313
rect -548 -8415 -514 -8381
rect -548 -8483 -514 -8449
rect -548 -8551 -514 -8517
rect -548 -8619 -514 -8585
rect -548 -8687 -514 -8653
rect -548 -8755 -514 -8721
rect -548 -8823 -514 -8789
rect -548 -8891 -514 -8857
rect -548 -8959 -514 -8925
rect -548 -9027 -514 -8993
rect -548 -9095 -514 -9061
rect -548 -9163 -514 -9129
rect -548 -9231 -514 -9197
rect -548 -9299 -514 -9265
rect -548 -9367 -514 -9333
rect -548 -9435 -514 -9401
rect -548 -9503 -514 -9469
rect -548 -9571 -514 -9537
rect -430 9537 -396 9571
rect -430 9469 -396 9503
rect -430 9401 -396 9435
rect -430 9333 -396 9367
rect -430 9265 -396 9299
rect -430 9197 -396 9231
rect -430 9129 -396 9163
rect -430 9061 -396 9095
rect -430 8993 -396 9027
rect -430 8925 -396 8959
rect -430 8857 -396 8891
rect -430 8789 -396 8823
rect -430 8721 -396 8755
rect -430 8653 -396 8687
rect -430 8585 -396 8619
rect -430 8517 -396 8551
rect -430 8449 -396 8483
rect -430 8381 -396 8415
rect -430 8313 -396 8347
rect -430 8245 -396 8279
rect -430 8177 -396 8211
rect -430 8109 -396 8143
rect -430 8041 -396 8075
rect -430 7973 -396 8007
rect -430 7905 -396 7939
rect -430 7837 -396 7871
rect -430 7769 -396 7803
rect -430 7701 -396 7735
rect -430 7633 -396 7667
rect -430 7565 -396 7599
rect -430 7497 -396 7531
rect -430 7429 -396 7463
rect -430 7361 -396 7395
rect -430 7293 -396 7327
rect -430 7225 -396 7259
rect -430 7157 -396 7191
rect -430 7089 -396 7123
rect -430 7021 -396 7055
rect -430 6953 -396 6987
rect -430 6885 -396 6919
rect -430 6817 -396 6851
rect -430 6749 -396 6783
rect -430 6681 -396 6715
rect -430 6613 -396 6647
rect -430 6545 -396 6579
rect -430 6477 -396 6511
rect -430 6409 -396 6443
rect -430 6341 -396 6375
rect -430 6273 -396 6307
rect -430 6205 -396 6239
rect -430 6137 -396 6171
rect -430 6069 -396 6103
rect -430 6001 -396 6035
rect -430 5933 -396 5967
rect -430 5865 -396 5899
rect -430 5797 -396 5831
rect -430 5729 -396 5763
rect -430 5661 -396 5695
rect -430 5593 -396 5627
rect -430 5525 -396 5559
rect -430 5457 -396 5491
rect -430 5389 -396 5423
rect -430 5321 -396 5355
rect -430 5253 -396 5287
rect -430 5185 -396 5219
rect -430 5117 -396 5151
rect -430 5049 -396 5083
rect -430 4981 -396 5015
rect -430 4913 -396 4947
rect -430 4845 -396 4879
rect -430 4777 -396 4811
rect -430 4709 -396 4743
rect -430 4641 -396 4675
rect -430 4573 -396 4607
rect -430 4505 -396 4539
rect -430 4437 -396 4471
rect -430 4369 -396 4403
rect -430 4301 -396 4335
rect -430 4233 -396 4267
rect -430 4165 -396 4199
rect -430 4097 -396 4131
rect -430 4029 -396 4063
rect -430 3961 -396 3995
rect -430 3893 -396 3927
rect -430 3825 -396 3859
rect -430 3757 -396 3791
rect -430 3689 -396 3723
rect -430 3621 -396 3655
rect -430 3553 -396 3587
rect -430 3485 -396 3519
rect -430 3417 -396 3451
rect -430 3349 -396 3383
rect -430 3281 -396 3315
rect -430 3213 -396 3247
rect -430 3145 -396 3179
rect -430 3077 -396 3111
rect -430 3009 -396 3043
rect -430 2941 -396 2975
rect -430 2873 -396 2907
rect -430 2805 -396 2839
rect -430 2737 -396 2771
rect -430 2669 -396 2703
rect -430 2601 -396 2635
rect -430 2533 -396 2567
rect -430 2465 -396 2499
rect -430 2397 -396 2431
rect -430 2329 -396 2363
rect -430 2261 -396 2295
rect -430 2193 -396 2227
rect -430 2125 -396 2159
rect -430 2057 -396 2091
rect -430 1989 -396 2023
rect -430 1921 -396 1955
rect -430 1853 -396 1887
rect -430 1785 -396 1819
rect -430 1717 -396 1751
rect -430 1649 -396 1683
rect -430 1581 -396 1615
rect -430 1513 -396 1547
rect -430 1445 -396 1479
rect -430 1377 -396 1411
rect -430 1309 -396 1343
rect -430 1241 -396 1275
rect -430 1173 -396 1207
rect -430 1105 -396 1139
rect -430 1037 -396 1071
rect -430 969 -396 1003
rect -430 901 -396 935
rect -430 833 -396 867
rect -430 765 -396 799
rect -430 697 -396 731
rect -430 629 -396 663
rect -430 561 -396 595
rect -430 493 -396 527
rect -430 425 -396 459
rect -430 357 -396 391
rect -430 289 -396 323
rect -430 221 -396 255
rect -430 153 -396 187
rect -430 85 -396 119
rect -430 17 -396 51
rect -430 -51 -396 -17
rect -430 -119 -396 -85
rect -430 -187 -396 -153
rect -430 -255 -396 -221
rect -430 -323 -396 -289
rect -430 -391 -396 -357
rect -430 -459 -396 -425
rect -430 -527 -396 -493
rect -430 -595 -396 -561
rect -430 -663 -396 -629
rect -430 -731 -396 -697
rect -430 -799 -396 -765
rect -430 -867 -396 -833
rect -430 -935 -396 -901
rect -430 -1003 -396 -969
rect -430 -1071 -396 -1037
rect -430 -1139 -396 -1105
rect -430 -1207 -396 -1173
rect -430 -1275 -396 -1241
rect -430 -1343 -396 -1309
rect -430 -1411 -396 -1377
rect -430 -1479 -396 -1445
rect -430 -1547 -396 -1513
rect -430 -1615 -396 -1581
rect -430 -1683 -396 -1649
rect -430 -1751 -396 -1717
rect -430 -1819 -396 -1785
rect -430 -1887 -396 -1853
rect -430 -1955 -396 -1921
rect -430 -2023 -396 -1989
rect -430 -2091 -396 -2057
rect -430 -2159 -396 -2125
rect -430 -2227 -396 -2193
rect -430 -2295 -396 -2261
rect -430 -2363 -396 -2329
rect -430 -2431 -396 -2397
rect -430 -2499 -396 -2465
rect -430 -2567 -396 -2533
rect -430 -2635 -396 -2601
rect -430 -2703 -396 -2669
rect -430 -2771 -396 -2737
rect -430 -2839 -396 -2805
rect -430 -2907 -396 -2873
rect -430 -2975 -396 -2941
rect -430 -3043 -396 -3009
rect -430 -3111 -396 -3077
rect -430 -3179 -396 -3145
rect -430 -3247 -396 -3213
rect -430 -3315 -396 -3281
rect -430 -3383 -396 -3349
rect -430 -3451 -396 -3417
rect -430 -3519 -396 -3485
rect -430 -3587 -396 -3553
rect -430 -3655 -396 -3621
rect -430 -3723 -396 -3689
rect -430 -3791 -396 -3757
rect -430 -3859 -396 -3825
rect -430 -3927 -396 -3893
rect -430 -3995 -396 -3961
rect -430 -4063 -396 -4029
rect -430 -4131 -396 -4097
rect -430 -4199 -396 -4165
rect -430 -4267 -396 -4233
rect -430 -4335 -396 -4301
rect -430 -4403 -396 -4369
rect -430 -4471 -396 -4437
rect -430 -4539 -396 -4505
rect -430 -4607 -396 -4573
rect -430 -4675 -396 -4641
rect -430 -4743 -396 -4709
rect -430 -4811 -396 -4777
rect -430 -4879 -396 -4845
rect -430 -4947 -396 -4913
rect -430 -5015 -396 -4981
rect -430 -5083 -396 -5049
rect -430 -5151 -396 -5117
rect -430 -5219 -396 -5185
rect -430 -5287 -396 -5253
rect -430 -5355 -396 -5321
rect -430 -5423 -396 -5389
rect -430 -5491 -396 -5457
rect -430 -5559 -396 -5525
rect -430 -5627 -396 -5593
rect -430 -5695 -396 -5661
rect -430 -5763 -396 -5729
rect -430 -5831 -396 -5797
rect -430 -5899 -396 -5865
rect -430 -5967 -396 -5933
rect -430 -6035 -396 -6001
rect -430 -6103 -396 -6069
rect -430 -6171 -396 -6137
rect -430 -6239 -396 -6205
rect -430 -6307 -396 -6273
rect -430 -6375 -396 -6341
rect -430 -6443 -396 -6409
rect -430 -6511 -396 -6477
rect -430 -6579 -396 -6545
rect -430 -6647 -396 -6613
rect -430 -6715 -396 -6681
rect -430 -6783 -396 -6749
rect -430 -6851 -396 -6817
rect -430 -6919 -396 -6885
rect -430 -6987 -396 -6953
rect -430 -7055 -396 -7021
rect -430 -7123 -396 -7089
rect -430 -7191 -396 -7157
rect -430 -7259 -396 -7225
rect -430 -7327 -396 -7293
rect -430 -7395 -396 -7361
rect -430 -7463 -396 -7429
rect -430 -7531 -396 -7497
rect -430 -7599 -396 -7565
rect -430 -7667 -396 -7633
rect -430 -7735 -396 -7701
rect -430 -7803 -396 -7769
rect -430 -7871 -396 -7837
rect -430 -7939 -396 -7905
rect -430 -8007 -396 -7973
rect -430 -8075 -396 -8041
rect -430 -8143 -396 -8109
rect -430 -8211 -396 -8177
rect -430 -8279 -396 -8245
rect -430 -8347 -396 -8313
rect -430 -8415 -396 -8381
rect -430 -8483 -396 -8449
rect -430 -8551 -396 -8517
rect -430 -8619 -396 -8585
rect -430 -8687 -396 -8653
rect -430 -8755 -396 -8721
rect -430 -8823 -396 -8789
rect -430 -8891 -396 -8857
rect -430 -8959 -396 -8925
rect -430 -9027 -396 -8993
rect -430 -9095 -396 -9061
rect -430 -9163 -396 -9129
rect -430 -9231 -396 -9197
rect -430 -9299 -396 -9265
rect -430 -9367 -396 -9333
rect -430 -9435 -396 -9401
rect -430 -9503 -396 -9469
rect -430 -9571 -396 -9537
rect -312 9537 -278 9571
rect -312 9469 -278 9503
rect -312 9401 -278 9435
rect -312 9333 -278 9367
rect -312 9265 -278 9299
rect -312 9197 -278 9231
rect -312 9129 -278 9163
rect -312 9061 -278 9095
rect -312 8993 -278 9027
rect -312 8925 -278 8959
rect -312 8857 -278 8891
rect -312 8789 -278 8823
rect -312 8721 -278 8755
rect -312 8653 -278 8687
rect -312 8585 -278 8619
rect -312 8517 -278 8551
rect -312 8449 -278 8483
rect -312 8381 -278 8415
rect -312 8313 -278 8347
rect -312 8245 -278 8279
rect -312 8177 -278 8211
rect -312 8109 -278 8143
rect -312 8041 -278 8075
rect -312 7973 -278 8007
rect -312 7905 -278 7939
rect -312 7837 -278 7871
rect -312 7769 -278 7803
rect -312 7701 -278 7735
rect -312 7633 -278 7667
rect -312 7565 -278 7599
rect -312 7497 -278 7531
rect -312 7429 -278 7463
rect -312 7361 -278 7395
rect -312 7293 -278 7327
rect -312 7225 -278 7259
rect -312 7157 -278 7191
rect -312 7089 -278 7123
rect -312 7021 -278 7055
rect -312 6953 -278 6987
rect -312 6885 -278 6919
rect -312 6817 -278 6851
rect -312 6749 -278 6783
rect -312 6681 -278 6715
rect -312 6613 -278 6647
rect -312 6545 -278 6579
rect -312 6477 -278 6511
rect -312 6409 -278 6443
rect -312 6341 -278 6375
rect -312 6273 -278 6307
rect -312 6205 -278 6239
rect -312 6137 -278 6171
rect -312 6069 -278 6103
rect -312 6001 -278 6035
rect -312 5933 -278 5967
rect -312 5865 -278 5899
rect -312 5797 -278 5831
rect -312 5729 -278 5763
rect -312 5661 -278 5695
rect -312 5593 -278 5627
rect -312 5525 -278 5559
rect -312 5457 -278 5491
rect -312 5389 -278 5423
rect -312 5321 -278 5355
rect -312 5253 -278 5287
rect -312 5185 -278 5219
rect -312 5117 -278 5151
rect -312 5049 -278 5083
rect -312 4981 -278 5015
rect -312 4913 -278 4947
rect -312 4845 -278 4879
rect -312 4777 -278 4811
rect -312 4709 -278 4743
rect -312 4641 -278 4675
rect -312 4573 -278 4607
rect -312 4505 -278 4539
rect -312 4437 -278 4471
rect -312 4369 -278 4403
rect -312 4301 -278 4335
rect -312 4233 -278 4267
rect -312 4165 -278 4199
rect -312 4097 -278 4131
rect -312 4029 -278 4063
rect -312 3961 -278 3995
rect -312 3893 -278 3927
rect -312 3825 -278 3859
rect -312 3757 -278 3791
rect -312 3689 -278 3723
rect -312 3621 -278 3655
rect -312 3553 -278 3587
rect -312 3485 -278 3519
rect -312 3417 -278 3451
rect -312 3349 -278 3383
rect -312 3281 -278 3315
rect -312 3213 -278 3247
rect -312 3145 -278 3179
rect -312 3077 -278 3111
rect -312 3009 -278 3043
rect -312 2941 -278 2975
rect -312 2873 -278 2907
rect -312 2805 -278 2839
rect -312 2737 -278 2771
rect -312 2669 -278 2703
rect -312 2601 -278 2635
rect -312 2533 -278 2567
rect -312 2465 -278 2499
rect -312 2397 -278 2431
rect -312 2329 -278 2363
rect -312 2261 -278 2295
rect -312 2193 -278 2227
rect -312 2125 -278 2159
rect -312 2057 -278 2091
rect -312 1989 -278 2023
rect -312 1921 -278 1955
rect -312 1853 -278 1887
rect -312 1785 -278 1819
rect -312 1717 -278 1751
rect -312 1649 -278 1683
rect -312 1581 -278 1615
rect -312 1513 -278 1547
rect -312 1445 -278 1479
rect -312 1377 -278 1411
rect -312 1309 -278 1343
rect -312 1241 -278 1275
rect -312 1173 -278 1207
rect -312 1105 -278 1139
rect -312 1037 -278 1071
rect -312 969 -278 1003
rect -312 901 -278 935
rect -312 833 -278 867
rect -312 765 -278 799
rect -312 697 -278 731
rect -312 629 -278 663
rect -312 561 -278 595
rect -312 493 -278 527
rect -312 425 -278 459
rect -312 357 -278 391
rect -312 289 -278 323
rect -312 221 -278 255
rect -312 153 -278 187
rect -312 85 -278 119
rect -312 17 -278 51
rect -312 -51 -278 -17
rect -312 -119 -278 -85
rect -312 -187 -278 -153
rect -312 -255 -278 -221
rect -312 -323 -278 -289
rect -312 -391 -278 -357
rect -312 -459 -278 -425
rect -312 -527 -278 -493
rect -312 -595 -278 -561
rect -312 -663 -278 -629
rect -312 -731 -278 -697
rect -312 -799 -278 -765
rect -312 -867 -278 -833
rect -312 -935 -278 -901
rect -312 -1003 -278 -969
rect -312 -1071 -278 -1037
rect -312 -1139 -278 -1105
rect -312 -1207 -278 -1173
rect -312 -1275 -278 -1241
rect -312 -1343 -278 -1309
rect -312 -1411 -278 -1377
rect -312 -1479 -278 -1445
rect -312 -1547 -278 -1513
rect -312 -1615 -278 -1581
rect -312 -1683 -278 -1649
rect -312 -1751 -278 -1717
rect -312 -1819 -278 -1785
rect -312 -1887 -278 -1853
rect -312 -1955 -278 -1921
rect -312 -2023 -278 -1989
rect -312 -2091 -278 -2057
rect -312 -2159 -278 -2125
rect -312 -2227 -278 -2193
rect -312 -2295 -278 -2261
rect -312 -2363 -278 -2329
rect -312 -2431 -278 -2397
rect -312 -2499 -278 -2465
rect -312 -2567 -278 -2533
rect -312 -2635 -278 -2601
rect -312 -2703 -278 -2669
rect -312 -2771 -278 -2737
rect -312 -2839 -278 -2805
rect -312 -2907 -278 -2873
rect -312 -2975 -278 -2941
rect -312 -3043 -278 -3009
rect -312 -3111 -278 -3077
rect -312 -3179 -278 -3145
rect -312 -3247 -278 -3213
rect -312 -3315 -278 -3281
rect -312 -3383 -278 -3349
rect -312 -3451 -278 -3417
rect -312 -3519 -278 -3485
rect -312 -3587 -278 -3553
rect -312 -3655 -278 -3621
rect -312 -3723 -278 -3689
rect -312 -3791 -278 -3757
rect -312 -3859 -278 -3825
rect -312 -3927 -278 -3893
rect -312 -3995 -278 -3961
rect -312 -4063 -278 -4029
rect -312 -4131 -278 -4097
rect -312 -4199 -278 -4165
rect -312 -4267 -278 -4233
rect -312 -4335 -278 -4301
rect -312 -4403 -278 -4369
rect -312 -4471 -278 -4437
rect -312 -4539 -278 -4505
rect -312 -4607 -278 -4573
rect -312 -4675 -278 -4641
rect -312 -4743 -278 -4709
rect -312 -4811 -278 -4777
rect -312 -4879 -278 -4845
rect -312 -4947 -278 -4913
rect -312 -5015 -278 -4981
rect -312 -5083 -278 -5049
rect -312 -5151 -278 -5117
rect -312 -5219 -278 -5185
rect -312 -5287 -278 -5253
rect -312 -5355 -278 -5321
rect -312 -5423 -278 -5389
rect -312 -5491 -278 -5457
rect -312 -5559 -278 -5525
rect -312 -5627 -278 -5593
rect -312 -5695 -278 -5661
rect -312 -5763 -278 -5729
rect -312 -5831 -278 -5797
rect -312 -5899 -278 -5865
rect -312 -5967 -278 -5933
rect -312 -6035 -278 -6001
rect -312 -6103 -278 -6069
rect -312 -6171 -278 -6137
rect -312 -6239 -278 -6205
rect -312 -6307 -278 -6273
rect -312 -6375 -278 -6341
rect -312 -6443 -278 -6409
rect -312 -6511 -278 -6477
rect -312 -6579 -278 -6545
rect -312 -6647 -278 -6613
rect -312 -6715 -278 -6681
rect -312 -6783 -278 -6749
rect -312 -6851 -278 -6817
rect -312 -6919 -278 -6885
rect -312 -6987 -278 -6953
rect -312 -7055 -278 -7021
rect -312 -7123 -278 -7089
rect -312 -7191 -278 -7157
rect -312 -7259 -278 -7225
rect -312 -7327 -278 -7293
rect -312 -7395 -278 -7361
rect -312 -7463 -278 -7429
rect -312 -7531 -278 -7497
rect -312 -7599 -278 -7565
rect -312 -7667 -278 -7633
rect -312 -7735 -278 -7701
rect -312 -7803 -278 -7769
rect -312 -7871 -278 -7837
rect -312 -7939 -278 -7905
rect -312 -8007 -278 -7973
rect -312 -8075 -278 -8041
rect -312 -8143 -278 -8109
rect -312 -8211 -278 -8177
rect -312 -8279 -278 -8245
rect -312 -8347 -278 -8313
rect -312 -8415 -278 -8381
rect -312 -8483 -278 -8449
rect -312 -8551 -278 -8517
rect -312 -8619 -278 -8585
rect -312 -8687 -278 -8653
rect -312 -8755 -278 -8721
rect -312 -8823 -278 -8789
rect -312 -8891 -278 -8857
rect -312 -8959 -278 -8925
rect -312 -9027 -278 -8993
rect -312 -9095 -278 -9061
rect -312 -9163 -278 -9129
rect -312 -9231 -278 -9197
rect -312 -9299 -278 -9265
rect -312 -9367 -278 -9333
rect -312 -9435 -278 -9401
rect -312 -9503 -278 -9469
rect -312 -9571 -278 -9537
rect -194 9537 -160 9571
rect -194 9469 -160 9503
rect -194 9401 -160 9435
rect -194 9333 -160 9367
rect -194 9265 -160 9299
rect -194 9197 -160 9231
rect -194 9129 -160 9163
rect -194 9061 -160 9095
rect -194 8993 -160 9027
rect -194 8925 -160 8959
rect -194 8857 -160 8891
rect -194 8789 -160 8823
rect -194 8721 -160 8755
rect -194 8653 -160 8687
rect -194 8585 -160 8619
rect -194 8517 -160 8551
rect -194 8449 -160 8483
rect -194 8381 -160 8415
rect -194 8313 -160 8347
rect -194 8245 -160 8279
rect -194 8177 -160 8211
rect -194 8109 -160 8143
rect -194 8041 -160 8075
rect -194 7973 -160 8007
rect -194 7905 -160 7939
rect -194 7837 -160 7871
rect -194 7769 -160 7803
rect -194 7701 -160 7735
rect -194 7633 -160 7667
rect -194 7565 -160 7599
rect -194 7497 -160 7531
rect -194 7429 -160 7463
rect -194 7361 -160 7395
rect -194 7293 -160 7327
rect -194 7225 -160 7259
rect -194 7157 -160 7191
rect -194 7089 -160 7123
rect -194 7021 -160 7055
rect -194 6953 -160 6987
rect -194 6885 -160 6919
rect -194 6817 -160 6851
rect -194 6749 -160 6783
rect -194 6681 -160 6715
rect -194 6613 -160 6647
rect -194 6545 -160 6579
rect -194 6477 -160 6511
rect -194 6409 -160 6443
rect -194 6341 -160 6375
rect -194 6273 -160 6307
rect -194 6205 -160 6239
rect -194 6137 -160 6171
rect -194 6069 -160 6103
rect -194 6001 -160 6035
rect -194 5933 -160 5967
rect -194 5865 -160 5899
rect -194 5797 -160 5831
rect -194 5729 -160 5763
rect -194 5661 -160 5695
rect -194 5593 -160 5627
rect -194 5525 -160 5559
rect -194 5457 -160 5491
rect -194 5389 -160 5423
rect -194 5321 -160 5355
rect -194 5253 -160 5287
rect -194 5185 -160 5219
rect -194 5117 -160 5151
rect -194 5049 -160 5083
rect -194 4981 -160 5015
rect -194 4913 -160 4947
rect -194 4845 -160 4879
rect -194 4777 -160 4811
rect -194 4709 -160 4743
rect -194 4641 -160 4675
rect -194 4573 -160 4607
rect -194 4505 -160 4539
rect -194 4437 -160 4471
rect -194 4369 -160 4403
rect -194 4301 -160 4335
rect -194 4233 -160 4267
rect -194 4165 -160 4199
rect -194 4097 -160 4131
rect -194 4029 -160 4063
rect -194 3961 -160 3995
rect -194 3893 -160 3927
rect -194 3825 -160 3859
rect -194 3757 -160 3791
rect -194 3689 -160 3723
rect -194 3621 -160 3655
rect -194 3553 -160 3587
rect -194 3485 -160 3519
rect -194 3417 -160 3451
rect -194 3349 -160 3383
rect -194 3281 -160 3315
rect -194 3213 -160 3247
rect -194 3145 -160 3179
rect -194 3077 -160 3111
rect -194 3009 -160 3043
rect -194 2941 -160 2975
rect -194 2873 -160 2907
rect -194 2805 -160 2839
rect -194 2737 -160 2771
rect -194 2669 -160 2703
rect -194 2601 -160 2635
rect -194 2533 -160 2567
rect -194 2465 -160 2499
rect -194 2397 -160 2431
rect -194 2329 -160 2363
rect -194 2261 -160 2295
rect -194 2193 -160 2227
rect -194 2125 -160 2159
rect -194 2057 -160 2091
rect -194 1989 -160 2023
rect -194 1921 -160 1955
rect -194 1853 -160 1887
rect -194 1785 -160 1819
rect -194 1717 -160 1751
rect -194 1649 -160 1683
rect -194 1581 -160 1615
rect -194 1513 -160 1547
rect -194 1445 -160 1479
rect -194 1377 -160 1411
rect -194 1309 -160 1343
rect -194 1241 -160 1275
rect -194 1173 -160 1207
rect -194 1105 -160 1139
rect -194 1037 -160 1071
rect -194 969 -160 1003
rect -194 901 -160 935
rect -194 833 -160 867
rect -194 765 -160 799
rect -194 697 -160 731
rect -194 629 -160 663
rect -194 561 -160 595
rect -194 493 -160 527
rect -194 425 -160 459
rect -194 357 -160 391
rect -194 289 -160 323
rect -194 221 -160 255
rect -194 153 -160 187
rect -194 85 -160 119
rect -194 17 -160 51
rect -194 -51 -160 -17
rect -194 -119 -160 -85
rect -194 -187 -160 -153
rect -194 -255 -160 -221
rect -194 -323 -160 -289
rect -194 -391 -160 -357
rect -194 -459 -160 -425
rect -194 -527 -160 -493
rect -194 -595 -160 -561
rect -194 -663 -160 -629
rect -194 -731 -160 -697
rect -194 -799 -160 -765
rect -194 -867 -160 -833
rect -194 -935 -160 -901
rect -194 -1003 -160 -969
rect -194 -1071 -160 -1037
rect -194 -1139 -160 -1105
rect -194 -1207 -160 -1173
rect -194 -1275 -160 -1241
rect -194 -1343 -160 -1309
rect -194 -1411 -160 -1377
rect -194 -1479 -160 -1445
rect -194 -1547 -160 -1513
rect -194 -1615 -160 -1581
rect -194 -1683 -160 -1649
rect -194 -1751 -160 -1717
rect -194 -1819 -160 -1785
rect -194 -1887 -160 -1853
rect -194 -1955 -160 -1921
rect -194 -2023 -160 -1989
rect -194 -2091 -160 -2057
rect -194 -2159 -160 -2125
rect -194 -2227 -160 -2193
rect -194 -2295 -160 -2261
rect -194 -2363 -160 -2329
rect -194 -2431 -160 -2397
rect -194 -2499 -160 -2465
rect -194 -2567 -160 -2533
rect -194 -2635 -160 -2601
rect -194 -2703 -160 -2669
rect -194 -2771 -160 -2737
rect -194 -2839 -160 -2805
rect -194 -2907 -160 -2873
rect -194 -2975 -160 -2941
rect -194 -3043 -160 -3009
rect -194 -3111 -160 -3077
rect -194 -3179 -160 -3145
rect -194 -3247 -160 -3213
rect -194 -3315 -160 -3281
rect -194 -3383 -160 -3349
rect -194 -3451 -160 -3417
rect -194 -3519 -160 -3485
rect -194 -3587 -160 -3553
rect -194 -3655 -160 -3621
rect -194 -3723 -160 -3689
rect -194 -3791 -160 -3757
rect -194 -3859 -160 -3825
rect -194 -3927 -160 -3893
rect -194 -3995 -160 -3961
rect -194 -4063 -160 -4029
rect -194 -4131 -160 -4097
rect -194 -4199 -160 -4165
rect -194 -4267 -160 -4233
rect -194 -4335 -160 -4301
rect -194 -4403 -160 -4369
rect -194 -4471 -160 -4437
rect -194 -4539 -160 -4505
rect -194 -4607 -160 -4573
rect -194 -4675 -160 -4641
rect -194 -4743 -160 -4709
rect -194 -4811 -160 -4777
rect -194 -4879 -160 -4845
rect -194 -4947 -160 -4913
rect -194 -5015 -160 -4981
rect -194 -5083 -160 -5049
rect -194 -5151 -160 -5117
rect -194 -5219 -160 -5185
rect -194 -5287 -160 -5253
rect -194 -5355 -160 -5321
rect -194 -5423 -160 -5389
rect -194 -5491 -160 -5457
rect -194 -5559 -160 -5525
rect -194 -5627 -160 -5593
rect -194 -5695 -160 -5661
rect -194 -5763 -160 -5729
rect -194 -5831 -160 -5797
rect -194 -5899 -160 -5865
rect -194 -5967 -160 -5933
rect -194 -6035 -160 -6001
rect -194 -6103 -160 -6069
rect -194 -6171 -160 -6137
rect -194 -6239 -160 -6205
rect -194 -6307 -160 -6273
rect -194 -6375 -160 -6341
rect -194 -6443 -160 -6409
rect -194 -6511 -160 -6477
rect -194 -6579 -160 -6545
rect -194 -6647 -160 -6613
rect -194 -6715 -160 -6681
rect -194 -6783 -160 -6749
rect -194 -6851 -160 -6817
rect -194 -6919 -160 -6885
rect -194 -6987 -160 -6953
rect -194 -7055 -160 -7021
rect -194 -7123 -160 -7089
rect -194 -7191 -160 -7157
rect -194 -7259 -160 -7225
rect -194 -7327 -160 -7293
rect -194 -7395 -160 -7361
rect -194 -7463 -160 -7429
rect -194 -7531 -160 -7497
rect -194 -7599 -160 -7565
rect -194 -7667 -160 -7633
rect -194 -7735 -160 -7701
rect -194 -7803 -160 -7769
rect -194 -7871 -160 -7837
rect -194 -7939 -160 -7905
rect -194 -8007 -160 -7973
rect -194 -8075 -160 -8041
rect -194 -8143 -160 -8109
rect -194 -8211 -160 -8177
rect -194 -8279 -160 -8245
rect -194 -8347 -160 -8313
rect -194 -8415 -160 -8381
rect -194 -8483 -160 -8449
rect -194 -8551 -160 -8517
rect -194 -8619 -160 -8585
rect -194 -8687 -160 -8653
rect -194 -8755 -160 -8721
rect -194 -8823 -160 -8789
rect -194 -8891 -160 -8857
rect -194 -8959 -160 -8925
rect -194 -9027 -160 -8993
rect -194 -9095 -160 -9061
rect -194 -9163 -160 -9129
rect -194 -9231 -160 -9197
rect -194 -9299 -160 -9265
rect -194 -9367 -160 -9333
rect -194 -9435 -160 -9401
rect -194 -9503 -160 -9469
rect -194 -9571 -160 -9537
rect -76 9537 -42 9571
rect -76 9469 -42 9503
rect -76 9401 -42 9435
rect -76 9333 -42 9367
rect -76 9265 -42 9299
rect -76 9197 -42 9231
rect -76 9129 -42 9163
rect -76 9061 -42 9095
rect -76 8993 -42 9027
rect -76 8925 -42 8959
rect -76 8857 -42 8891
rect -76 8789 -42 8823
rect -76 8721 -42 8755
rect -76 8653 -42 8687
rect -76 8585 -42 8619
rect -76 8517 -42 8551
rect -76 8449 -42 8483
rect -76 8381 -42 8415
rect -76 8313 -42 8347
rect -76 8245 -42 8279
rect -76 8177 -42 8211
rect -76 8109 -42 8143
rect -76 8041 -42 8075
rect -76 7973 -42 8007
rect -76 7905 -42 7939
rect -76 7837 -42 7871
rect -76 7769 -42 7803
rect -76 7701 -42 7735
rect -76 7633 -42 7667
rect -76 7565 -42 7599
rect -76 7497 -42 7531
rect -76 7429 -42 7463
rect -76 7361 -42 7395
rect -76 7293 -42 7327
rect -76 7225 -42 7259
rect -76 7157 -42 7191
rect -76 7089 -42 7123
rect -76 7021 -42 7055
rect -76 6953 -42 6987
rect -76 6885 -42 6919
rect -76 6817 -42 6851
rect -76 6749 -42 6783
rect -76 6681 -42 6715
rect -76 6613 -42 6647
rect -76 6545 -42 6579
rect -76 6477 -42 6511
rect -76 6409 -42 6443
rect -76 6341 -42 6375
rect -76 6273 -42 6307
rect -76 6205 -42 6239
rect -76 6137 -42 6171
rect -76 6069 -42 6103
rect -76 6001 -42 6035
rect -76 5933 -42 5967
rect -76 5865 -42 5899
rect -76 5797 -42 5831
rect -76 5729 -42 5763
rect -76 5661 -42 5695
rect -76 5593 -42 5627
rect -76 5525 -42 5559
rect -76 5457 -42 5491
rect -76 5389 -42 5423
rect -76 5321 -42 5355
rect -76 5253 -42 5287
rect -76 5185 -42 5219
rect -76 5117 -42 5151
rect -76 5049 -42 5083
rect -76 4981 -42 5015
rect -76 4913 -42 4947
rect -76 4845 -42 4879
rect -76 4777 -42 4811
rect -76 4709 -42 4743
rect -76 4641 -42 4675
rect -76 4573 -42 4607
rect -76 4505 -42 4539
rect -76 4437 -42 4471
rect -76 4369 -42 4403
rect -76 4301 -42 4335
rect -76 4233 -42 4267
rect -76 4165 -42 4199
rect -76 4097 -42 4131
rect -76 4029 -42 4063
rect -76 3961 -42 3995
rect -76 3893 -42 3927
rect -76 3825 -42 3859
rect -76 3757 -42 3791
rect -76 3689 -42 3723
rect -76 3621 -42 3655
rect -76 3553 -42 3587
rect -76 3485 -42 3519
rect -76 3417 -42 3451
rect -76 3349 -42 3383
rect -76 3281 -42 3315
rect -76 3213 -42 3247
rect -76 3145 -42 3179
rect -76 3077 -42 3111
rect -76 3009 -42 3043
rect -76 2941 -42 2975
rect -76 2873 -42 2907
rect -76 2805 -42 2839
rect -76 2737 -42 2771
rect -76 2669 -42 2703
rect -76 2601 -42 2635
rect -76 2533 -42 2567
rect -76 2465 -42 2499
rect -76 2397 -42 2431
rect -76 2329 -42 2363
rect -76 2261 -42 2295
rect -76 2193 -42 2227
rect -76 2125 -42 2159
rect -76 2057 -42 2091
rect -76 1989 -42 2023
rect -76 1921 -42 1955
rect -76 1853 -42 1887
rect -76 1785 -42 1819
rect -76 1717 -42 1751
rect -76 1649 -42 1683
rect -76 1581 -42 1615
rect -76 1513 -42 1547
rect -76 1445 -42 1479
rect -76 1377 -42 1411
rect -76 1309 -42 1343
rect -76 1241 -42 1275
rect -76 1173 -42 1207
rect -76 1105 -42 1139
rect -76 1037 -42 1071
rect -76 969 -42 1003
rect -76 901 -42 935
rect -76 833 -42 867
rect -76 765 -42 799
rect -76 697 -42 731
rect -76 629 -42 663
rect -76 561 -42 595
rect -76 493 -42 527
rect -76 425 -42 459
rect -76 357 -42 391
rect -76 289 -42 323
rect -76 221 -42 255
rect -76 153 -42 187
rect -76 85 -42 119
rect -76 17 -42 51
rect -76 -51 -42 -17
rect -76 -119 -42 -85
rect -76 -187 -42 -153
rect -76 -255 -42 -221
rect -76 -323 -42 -289
rect -76 -391 -42 -357
rect -76 -459 -42 -425
rect -76 -527 -42 -493
rect -76 -595 -42 -561
rect -76 -663 -42 -629
rect -76 -731 -42 -697
rect -76 -799 -42 -765
rect -76 -867 -42 -833
rect -76 -935 -42 -901
rect -76 -1003 -42 -969
rect -76 -1071 -42 -1037
rect -76 -1139 -42 -1105
rect -76 -1207 -42 -1173
rect -76 -1275 -42 -1241
rect -76 -1343 -42 -1309
rect -76 -1411 -42 -1377
rect -76 -1479 -42 -1445
rect -76 -1547 -42 -1513
rect -76 -1615 -42 -1581
rect -76 -1683 -42 -1649
rect -76 -1751 -42 -1717
rect -76 -1819 -42 -1785
rect -76 -1887 -42 -1853
rect -76 -1955 -42 -1921
rect -76 -2023 -42 -1989
rect -76 -2091 -42 -2057
rect -76 -2159 -42 -2125
rect -76 -2227 -42 -2193
rect -76 -2295 -42 -2261
rect -76 -2363 -42 -2329
rect -76 -2431 -42 -2397
rect -76 -2499 -42 -2465
rect -76 -2567 -42 -2533
rect -76 -2635 -42 -2601
rect -76 -2703 -42 -2669
rect -76 -2771 -42 -2737
rect -76 -2839 -42 -2805
rect -76 -2907 -42 -2873
rect -76 -2975 -42 -2941
rect -76 -3043 -42 -3009
rect -76 -3111 -42 -3077
rect -76 -3179 -42 -3145
rect -76 -3247 -42 -3213
rect -76 -3315 -42 -3281
rect -76 -3383 -42 -3349
rect -76 -3451 -42 -3417
rect -76 -3519 -42 -3485
rect -76 -3587 -42 -3553
rect -76 -3655 -42 -3621
rect -76 -3723 -42 -3689
rect -76 -3791 -42 -3757
rect -76 -3859 -42 -3825
rect -76 -3927 -42 -3893
rect -76 -3995 -42 -3961
rect -76 -4063 -42 -4029
rect -76 -4131 -42 -4097
rect -76 -4199 -42 -4165
rect -76 -4267 -42 -4233
rect -76 -4335 -42 -4301
rect -76 -4403 -42 -4369
rect -76 -4471 -42 -4437
rect -76 -4539 -42 -4505
rect -76 -4607 -42 -4573
rect -76 -4675 -42 -4641
rect -76 -4743 -42 -4709
rect -76 -4811 -42 -4777
rect -76 -4879 -42 -4845
rect -76 -4947 -42 -4913
rect -76 -5015 -42 -4981
rect -76 -5083 -42 -5049
rect -76 -5151 -42 -5117
rect -76 -5219 -42 -5185
rect -76 -5287 -42 -5253
rect -76 -5355 -42 -5321
rect -76 -5423 -42 -5389
rect -76 -5491 -42 -5457
rect -76 -5559 -42 -5525
rect -76 -5627 -42 -5593
rect -76 -5695 -42 -5661
rect -76 -5763 -42 -5729
rect -76 -5831 -42 -5797
rect -76 -5899 -42 -5865
rect -76 -5967 -42 -5933
rect -76 -6035 -42 -6001
rect -76 -6103 -42 -6069
rect -76 -6171 -42 -6137
rect -76 -6239 -42 -6205
rect -76 -6307 -42 -6273
rect -76 -6375 -42 -6341
rect -76 -6443 -42 -6409
rect -76 -6511 -42 -6477
rect -76 -6579 -42 -6545
rect -76 -6647 -42 -6613
rect -76 -6715 -42 -6681
rect -76 -6783 -42 -6749
rect -76 -6851 -42 -6817
rect -76 -6919 -42 -6885
rect -76 -6987 -42 -6953
rect -76 -7055 -42 -7021
rect -76 -7123 -42 -7089
rect -76 -7191 -42 -7157
rect -76 -7259 -42 -7225
rect -76 -7327 -42 -7293
rect -76 -7395 -42 -7361
rect -76 -7463 -42 -7429
rect -76 -7531 -42 -7497
rect -76 -7599 -42 -7565
rect -76 -7667 -42 -7633
rect -76 -7735 -42 -7701
rect -76 -7803 -42 -7769
rect -76 -7871 -42 -7837
rect -76 -7939 -42 -7905
rect -76 -8007 -42 -7973
rect -76 -8075 -42 -8041
rect -76 -8143 -42 -8109
rect -76 -8211 -42 -8177
rect -76 -8279 -42 -8245
rect -76 -8347 -42 -8313
rect -76 -8415 -42 -8381
rect -76 -8483 -42 -8449
rect -76 -8551 -42 -8517
rect -76 -8619 -42 -8585
rect -76 -8687 -42 -8653
rect -76 -8755 -42 -8721
rect -76 -8823 -42 -8789
rect -76 -8891 -42 -8857
rect -76 -8959 -42 -8925
rect -76 -9027 -42 -8993
rect -76 -9095 -42 -9061
rect -76 -9163 -42 -9129
rect -76 -9231 -42 -9197
rect -76 -9299 -42 -9265
rect -76 -9367 -42 -9333
rect -76 -9435 -42 -9401
rect -76 -9503 -42 -9469
rect -76 -9571 -42 -9537
rect 42 9537 76 9571
rect 42 9469 76 9503
rect 42 9401 76 9435
rect 42 9333 76 9367
rect 42 9265 76 9299
rect 42 9197 76 9231
rect 42 9129 76 9163
rect 42 9061 76 9095
rect 42 8993 76 9027
rect 42 8925 76 8959
rect 42 8857 76 8891
rect 42 8789 76 8823
rect 42 8721 76 8755
rect 42 8653 76 8687
rect 42 8585 76 8619
rect 42 8517 76 8551
rect 42 8449 76 8483
rect 42 8381 76 8415
rect 42 8313 76 8347
rect 42 8245 76 8279
rect 42 8177 76 8211
rect 42 8109 76 8143
rect 42 8041 76 8075
rect 42 7973 76 8007
rect 42 7905 76 7939
rect 42 7837 76 7871
rect 42 7769 76 7803
rect 42 7701 76 7735
rect 42 7633 76 7667
rect 42 7565 76 7599
rect 42 7497 76 7531
rect 42 7429 76 7463
rect 42 7361 76 7395
rect 42 7293 76 7327
rect 42 7225 76 7259
rect 42 7157 76 7191
rect 42 7089 76 7123
rect 42 7021 76 7055
rect 42 6953 76 6987
rect 42 6885 76 6919
rect 42 6817 76 6851
rect 42 6749 76 6783
rect 42 6681 76 6715
rect 42 6613 76 6647
rect 42 6545 76 6579
rect 42 6477 76 6511
rect 42 6409 76 6443
rect 42 6341 76 6375
rect 42 6273 76 6307
rect 42 6205 76 6239
rect 42 6137 76 6171
rect 42 6069 76 6103
rect 42 6001 76 6035
rect 42 5933 76 5967
rect 42 5865 76 5899
rect 42 5797 76 5831
rect 42 5729 76 5763
rect 42 5661 76 5695
rect 42 5593 76 5627
rect 42 5525 76 5559
rect 42 5457 76 5491
rect 42 5389 76 5423
rect 42 5321 76 5355
rect 42 5253 76 5287
rect 42 5185 76 5219
rect 42 5117 76 5151
rect 42 5049 76 5083
rect 42 4981 76 5015
rect 42 4913 76 4947
rect 42 4845 76 4879
rect 42 4777 76 4811
rect 42 4709 76 4743
rect 42 4641 76 4675
rect 42 4573 76 4607
rect 42 4505 76 4539
rect 42 4437 76 4471
rect 42 4369 76 4403
rect 42 4301 76 4335
rect 42 4233 76 4267
rect 42 4165 76 4199
rect 42 4097 76 4131
rect 42 4029 76 4063
rect 42 3961 76 3995
rect 42 3893 76 3927
rect 42 3825 76 3859
rect 42 3757 76 3791
rect 42 3689 76 3723
rect 42 3621 76 3655
rect 42 3553 76 3587
rect 42 3485 76 3519
rect 42 3417 76 3451
rect 42 3349 76 3383
rect 42 3281 76 3315
rect 42 3213 76 3247
rect 42 3145 76 3179
rect 42 3077 76 3111
rect 42 3009 76 3043
rect 42 2941 76 2975
rect 42 2873 76 2907
rect 42 2805 76 2839
rect 42 2737 76 2771
rect 42 2669 76 2703
rect 42 2601 76 2635
rect 42 2533 76 2567
rect 42 2465 76 2499
rect 42 2397 76 2431
rect 42 2329 76 2363
rect 42 2261 76 2295
rect 42 2193 76 2227
rect 42 2125 76 2159
rect 42 2057 76 2091
rect 42 1989 76 2023
rect 42 1921 76 1955
rect 42 1853 76 1887
rect 42 1785 76 1819
rect 42 1717 76 1751
rect 42 1649 76 1683
rect 42 1581 76 1615
rect 42 1513 76 1547
rect 42 1445 76 1479
rect 42 1377 76 1411
rect 42 1309 76 1343
rect 42 1241 76 1275
rect 42 1173 76 1207
rect 42 1105 76 1139
rect 42 1037 76 1071
rect 42 969 76 1003
rect 42 901 76 935
rect 42 833 76 867
rect 42 765 76 799
rect 42 697 76 731
rect 42 629 76 663
rect 42 561 76 595
rect 42 493 76 527
rect 42 425 76 459
rect 42 357 76 391
rect 42 289 76 323
rect 42 221 76 255
rect 42 153 76 187
rect 42 85 76 119
rect 42 17 76 51
rect 42 -51 76 -17
rect 42 -119 76 -85
rect 42 -187 76 -153
rect 42 -255 76 -221
rect 42 -323 76 -289
rect 42 -391 76 -357
rect 42 -459 76 -425
rect 42 -527 76 -493
rect 42 -595 76 -561
rect 42 -663 76 -629
rect 42 -731 76 -697
rect 42 -799 76 -765
rect 42 -867 76 -833
rect 42 -935 76 -901
rect 42 -1003 76 -969
rect 42 -1071 76 -1037
rect 42 -1139 76 -1105
rect 42 -1207 76 -1173
rect 42 -1275 76 -1241
rect 42 -1343 76 -1309
rect 42 -1411 76 -1377
rect 42 -1479 76 -1445
rect 42 -1547 76 -1513
rect 42 -1615 76 -1581
rect 42 -1683 76 -1649
rect 42 -1751 76 -1717
rect 42 -1819 76 -1785
rect 42 -1887 76 -1853
rect 42 -1955 76 -1921
rect 42 -2023 76 -1989
rect 42 -2091 76 -2057
rect 42 -2159 76 -2125
rect 42 -2227 76 -2193
rect 42 -2295 76 -2261
rect 42 -2363 76 -2329
rect 42 -2431 76 -2397
rect 42 -2499 76 -2465
rect 42 -2567 76 -2533
rect 42 -2635 76 -2601
rect 42 -2703 76 -2669
rect 42 -2771 76 -2737
rect 42 -2839 76 -2805
rect 42 -2907 76 -2873
rect 42 -2975 76 -2941
rect 42 -3043 76 -3009
rect 42 -3111 76 -3077
rect 42 -3179 76 -3145
rect 42 -3247 76 -3213
rect 42 -3315 76 -3281
rect 42 -3383 76 -3349
rect 42 -3451 76 -3417
rect 42 -3519 76 -3485
rect 42 -3587 76 -3553
rect 42 -3655 76 -3621
rect 42 -3723 76 -3689
rect 42 -3791 76 -3757
rect 42 -3859 76 -3825
rect 42 -3927 76 -3893
rect 42 -3995 76 -3961
rect 42 -4063 76 -4029
rect 42 -4131 76 -4097
rect 42 -4199 76 -4165
rect 42 -4267 76 -4233
rect 42 -4335 76 -4301
rect 42 -4403 76 -4369
rect 42 -4471 76 -4437
rect 42 -4539 76 -4505
rect 42 -4607 76 -4573
rect 42 -4675 76 -4641
rect 42 -4743 76 -4709
rect 42 -4811 76 -4777
rect 42 -4879 76 -4845
rect 42 -4947 76 -4913
rect 42 -5015 76 -4981
rect 42 -5083 76 -5049
rect 42 -5151 76 -5117
rect 42 -5219 76 -5185
rect 42 -5287 76 -5253
rect 42 -5355 76 -5321
rect 42 -5423 76 -5389
rect 42 -5491 76 -5457
rect 42 -5559 76 -5525
rect 42 -5627 76 -5593
rect 42 -5695 76 -5661
rect 42 -5763 76 -5729
rect 42 -5831 76 -5797
rect 42 -5899 76 -5865
rect 42 -5967 76 -5933
rect 42 -6035 76 -6001
rect 42 -6103 76 -6069
rect 42 -6171 76 -6137
rect 42 -6239 76 -6205
rect 42 -6307 76 -6273
rect 42 -6375 76 -6341
rect 42 -6443 76 -6409
rect 42 -6511 76 -6477
rect 42 -6579 76 -6545
rect 42 -6647 76 -6613
rect 42 -6715 76 -6681
rect 42 -6783 76 -6749
rect 42 -6851 76 -6817
rect 42 -6919 76 -6885
rect 42 -6987 76 -6953
rect 42 -7055 76 -7021
rect 42 -7123 76 -7089
rect 42 -7191 76 -7157
rect 42 -7259 76 -7225
rect 42 -7327 76 -7293
rect 42 -7395 76 -7361
rect 42 -7463 76 -7429
rect 42 -7531 76 -7497
rect 42 -7599 76 -7565
rect 42 -7667 76 -7633
rect 42 -7735 76 -7701
rect 42 -7803 76 -7769
rect 42 -7871 76 -7837
rect 42 -7939 76 -7905
rect 42 -8007 76 -7973
rect 42 -8075 76 -8041
rect 42 -8143 76 -8109
rect 42 -8211 76 -8177
rect 42 -8279 76 -8245
rect 42 -8347 76 -8313
rect 42 -8415 76 -8381
rect 42 -8483 76 -8449
rect 42 -8551 76 -8517
rect 42 -8619 76 -8585
rect 42 -8687 76 -8653
rect 42 -8755 76 -8721
rect 42 -8823 76 -8789
rect 42 -8891 76 -8857
rect 42 -8959 76 -8925
rect 42 -9027 76 -8993
rect 42 -9095 76 -9061
rect 42 -9163 76 -9129
rect 42 -9231 76 -9197
rect 42 -9299 76 -9265
rect 42 -9367 76 -9333
rect 42 -9435 76 -9401
rect 42 -9503 76 -9469
rect 42 -9571 76 -9537
rect 160 9537 194 9571
rect 160 9469 194 9503
rect 160 9401 194 9435
rect 160 9333 194 9367
rect 160 9265 194 9299
rect 160 9197 194 9231
rect 160 9129 194 9163
rect 160 9061 194 9095
rect 160 8993 194 9027
rect 160 8925 194 8959
rect 160 8857 194 8891
rect 160 8789 194 8823
rect 160 8721 194 8755
rect 160 8653 194 8687
rect 160 8585 194 8619
rect 160 8517 194 8551
rect 160 8449 194 8483
rect 160 8381 194 8415
rect 160 8313 194 8347
rect 160 8245 194 8279
rect 160 8177 194 8211
rect 160 8109 194 8143
rect 160 8041 194 8075
rect 160 7973 194 8007
rect 160 7905 194 7939
rect 160 7837 194 7871
rect 160 7769 194 7803
rect 160 7701 194 7735
rect 160 7633 194 7667
rect 160 7565 194 7599
rect 160 7497 194 7531
rect 160 7429 194 7463
rect 160 7361 194 7395
rect 160 7293 194 7327
rect 160 7225 194 7259
rect 160 7157 194 7191
rect 160 7089 194 7123
rect 160 7021 194 7055
rect 160 6953 194 6987
rect 160 6885 194 6919
rect 160 6817 194 6851
rect 160 6749 194 6783
rect 160 6681 194 6715
rect 160 6613 194 6647
rect 160 6545 194 6579
rect 160 6477 194 6511
rect 160 6409 194 6443
rect 160 6341 194 6375
rect 160 6273 194 6307
rect 160 6205 194 6239
rect 160 6137 194 6171
rect 160 6069 194 6103
rect 160 6001 194 6035
rect 160 5933 194 5967
rect 160 5865 194 5899
rect 160 5797 194 5831
rect 160 5729 194 5763
rect 160 5661 194 5695
rect 160 5593 194 5627
rect 160 5525 194 5559
rect 160 5457 194 5491
rect 160 5389 194 5423
rect 160 5321 194 5355
rect 160 5253 194 5287
rect 160 5185 194 5219
rect 160 5117 194 5151
rect 160 5049 194 5083
rect 160 4981 194 5015
rect 160 4913 194 4947
rect 160 4845 194 4879
rect 160 4777 194 4811
rect 160 4709 194 4743
rect 160 4641 194 4675
rect 160 4573 194 4607
rect 160 4505 194 4539
rect 160 4437 194 4471
rect 160 4369 194 4403
rect 160 4301 194 4335
rect 160 4233 194 4267
rect 160 4165 194 4199
rect 160 4097 194 4131
rect 160 4029 194 4063
rect 160 3961 194 3995
rect 160 3893 194 3927
rect 160 3825 194 3859
rect 160 3757 194 3791
rect 160 3689 194 3723
rect 160 3621 194 3655
rect 160 3553 194 3587
rect 160 3485 194 3519
rect 160 3417 194 3451
rect 160 3349 194 3383
rect 160 3281 194 3315
rect 160 3213 194 3247
rect 160 3145 194 3179
rect 160 3077 194 3111
rect 160 3009 194 3043
rect 160 2941 194 2975
rect 160 2873 194 2907
rect 160 2805 194 2839
rect 160 2737 194 2771
rect 160 2669 194 2703
rect 160 2601 194 2635
rect 160 2533 194 2567
rect 160 2465 194 2499
rect 160 2397 194 2431
rect 160 2329 194 2363
rect 160 2261 194 2295
rect 160 2193 194 2227
rect 160 2125 194 2159
rect 160 2057 194 2091
rect 160 1989 194 2023
rect 160 1921 194 1955
rect 160 1853 194 1887
rect 160 1785 194 1819
rect 160 1717 194 1751
rect 160 1649 194 1683
rect 160 1581 194 1615
rect 160 1513 194 1547
rect 160 1445 194 1479
rect 160 1377 194 1411
rect 160 1309 194 1343
rect 160 1241 194 1275
rect 160 1173 194 1207
rect 160 1105 194 1139
rect 160 1037 194 1071
rect 160 969 194 1003
rect 160 901 194 935
rect 160 833 194 867
rect 160 765 194 799
rect 160 697 194 731
rect 160 629 194 663
rect 160 561 194 595
rect 160 493 194 527
rect 160 425 194 459
rect 160 357 194 391
rect 160 289 194 323
rect 160 221 194 255
rect 160 153 194 187
rect 160 85 194 119
rect 160 17 194 51
rect 160 -51 194 -17
rect 160 -119 194 -85
rect 160 -187 194 -153
rect 160 -255 194 -221
rect 160 -323 194 -289
rect 160 -391 194 -357
rect 160 -459 194 -425
rect 160 -527 194 -493
rect 160 -595 194 -561
rect 160 -663 194 -629
rect 160 -731 194 -697
rect 160 -799 194 -765
rect 160 -867 194 -833
rect 160 -935 194 -901
rect 160 -1003 194 -969
rect 160 -1071 194 -1037
rect 160 -1139 194 -1105
rect 160 -1207 194 -1173
rect 160 -1275 194 -1241
rect 160 -1343 194 -1309
rect 160 -1411 194 -1377
rect 160 -1479 194 -1445
rect 160 -1547 194 -1513
rect 160 -1615 194 -1581
rect 160 -1683 194 -1649
rect 160 -1751 194 -1717
rect 160 -1819 194 -1785
rect 160 -1887 194 -1853
rect 160 -1955 194 -1921
rect 160 -2023 194 -1989
rect 160 -2091 194 -2057
rect 160 -2159 194 -2125
rect 160 -2227 194 -2193
rect 160 -2295 194 -2261
rect 160 -2363 194 -2329
rect 160 -2431 194 -2397
rect 160 -2499 194 -2465
rect 160 -2567 194 -2533
rect 160 -2635 194 -2601
rect 160 -2703 194 -2669
rect 160 -2771 194 -2737
rect 160 -2839 194 -2805
rect 160 -2907 194 -2873
rect 160 -2975 194 -2941
rect 160 -3043 194 -3009
rect 160 -3111 194 -3077
rect 160 -3179 194 -3145
rect 160 -3247 194 -3213
rect 160 -3315 194 -3281
rect 160 -3383 194 -3349
rect 160 -3451 194 -3417
rect 160 -3519 194 -3485
rect 160 -3587 194 -3553
rect 160 -3655 194 -3621
rect 160 -3723 194 -3689
rect 160 -3791 194 -3757
rect 160 -3859 194 -3825
rect 160 -3927 194 -3893
rect 160 -3995 194 -3961
rect 160 -4063 194 -4029
rect 160 -4131 194 -4097
rect 160 -4199 194 -4165
rect 160 -4267 194 -4233
rect 160 -4335 194 -4301
rect 160 -4403 194 -4369
rect 160 -4471 194 -4437
rect 160 -4539 194 -4505
rect 160 -4607 194 -4573
rect 160 -4675 194 -4641
rect 160 -4743 194 -4709
rect 160 -4811 194 -4777
rect 160 -4879 194 -4845
rect 160 -4947 194 -4913
rect 160 -5015 194 -4981
rect 160 -5083 194 -5049
rect 160 -5151 194 -5117
rect 160 -5219 194 -5185
rect 160 -5287 194 -5253
rect 160 -5355 194 -5321
rect 160 -5423 194 -5389
rect 160 -5491 194 -5457
rect 160 -5559 194 -5525
rect 160 -5627 194 -5593
rect 160 -5695 194 -5661
rect 160 -5763 194 -5729
rect 160 -5831 194 -5797
rect 160 -5899 194 -5865
rect 160 -5967 194 -5933
rect 160 -6035 194 -6001
rect 160 -6103 194 -6069
rect 160 -6171 194 -6137
rect 160 -6239 194 -6205
rect 160 -6307 194 -6273
rect 160 -6375 194 -6341
rect 160 -6443 194 -6409
rect 160 -6511 194 -6477
rect 160 -6579 194 -6545
rect 160 -6647 194 -6613
rect 160 -6715 194 -6681
rect 160 -6783 194 -6749
rect 160 -6851 194 -6817
rect 160 -6919 194 -6885
rect 160 -6987 194 -6953
rect 160 -7055 194 -7021
rect 160 -7123 194 -7089
rect 160 -7191 194 -7157
rect 160 -7259 194 -7225
rect 160 -7327 194 -7293
rect 160 -7395 194 -7361
rect 160 -7463 194 -7429
rect 160 -7531 194 -7497
rect 160 -7599 194 -7565
rect 160 -7667 194 -7633
rect 160 -7735 194 -7701
rect 160 -7803 194 -7769
rect 160 -7871 194 -7837
rect 160 -7939 194 -7905
rect 160 -8007 194 -7973
rect 160 -8075 194 -8041
rect 160 -8143 194 -8109
rect 160 -8211 194 -8177
rect 160 -8279 194 -8245
rect 160 -8347 194 -8313
rect 160 -8415 194 -8381
rect 160 -8483 194 -8449
rect 160 -8551 194 -8517
rect 160 -8619 194 -8585
rect 160 -8687 194 -8653
rect 160 -8755 194 -8721
rect 160 -8823 194 -8789
rect 160 -8891 194 -8857
rect 160 -8959 194 -8925
rect 160 -9027 194 -8993
rect 160 -9095 194 -9061
rect 160 -9163 194 -9129
rect 160 -9231 194 -9197
rect 160 -9299 194 -9265
rect 160 -9367 194 -9333
rect 160 -9435 194 -9401
rect 160 -9503 194 -9469
rect 160 -9571 194 -9537
rect 278 9537 312 9571
rect 278 9469 312 9503
rect 278 9401 312 9435
rect 278 9333 312 9367
rect 278 9265 312 9299
rect 278 9197 312 9231
rect 278 9129 312 9163
rect 278 9061 312 9095
rect 278 8993 312 9027
rect 278 8925 312 8959
rect 278 8857 312 8891
rect 278 8789 312 8823
rect 278 8721 312 8755
rect 278 8653 312 8687
rect 278 8585 312 8619
rect 278 8517 312 8551
rect 278 8449 312 8483
rect 278 8381 312 8415
rect 278 8313 312 8347
rect 278 8245 312 8279
rect 278 8177 312 8211
rect 278 8109 312 8143
rect 278 8041 312 8075
rect 278 7973 312 8007
rect 278 7905 312 7939
rect 278 7837 312 7871
rect 278 7769 312 7803
rect 278 7701 312 7735
rect 278 7633 312 7667
rect 278 7565 312 7599
rect 278 7497 312 7531
rect 278 7429 312 7463
rect 278 7361 312 7395
rect 278 7293 312 7327
rect 278 7225 312 7259
rect 278 7157 312 7191
rect 278 7089 312 7123
rect 278 7021 312 7055
rect 278 6953 312 6987
rect 278 6885 312 6919
rect 278 6817 312 6851
rect 278 6749 312 6783
rect 278 6681 312 6715
rect 278 6613 312 6647
rect 278 6545 312 6579
rect 278 6477 312 6511
rect 278 6409 312 6443
rect 278 6341 312 6375
rect 278 6273 312 6307
rect 278 6205 312 6239
rect 278 6137 312 6171
rect 278 6069 312 6103
rect 278 6001 312 6035
rect 278 5933 312 5967
rect 278 5865 312 5899
rect 278 5797 312 5831
rect 278 5729 312 5763
rect 278 5661 312 5695
rect 278 5593 312 5627
rect 278 5525 312 5559
rect 278 5457 312 5491
rect 278 5389 312 5423
rect 278 5321 312 5355
rect 278 5253 312 5287
rect 278 5185 312 5219
rect 278 5117 312 5151
rect 278 5049 312 5083
rect 278 4981 312 5015
rect 278 4913 312 4947
rect 278 4845 312 4879
rect 278 4777 312 4811
rect 278 4709 312 4743
rect 278 4641 312 4675
rect 278 4573 312 4607
rect 278 4505 312 4539
rect 278 4437 312 4471
rect 278 4369 312 4403
rect 278 4301 312 4335
rect 278 4233 312 4267
rect 278 4165 312 4199
rect 278 4097 312 4131
rect 278 4029 312 4063
rect 278 3961 312 3995
rect 278 3893 312 3927
rect 278 3825 312 3859
rect 278 3757 312 3791
rect 278 3689 312 3723
rect 278 3621 312 3655
rect 278 3553 312 3587
rect 278 3485 312 3519
rect 278 3417 312 3451
rect 278 3349 312 3383
rect 278 3281 312 3315
rect 278 3213 312 3247
rect 278 3145 312 3179
rect 278 3077 312 3111
rect 278 3009 312 3043
rect 278 2941 312 2975
rect 278 2873 312 2907
rect 278 2805 312 2839
rect 278 2737 312 2771
rect 278 2669 312 2703
rect 278 2601 312 2635
rect 278 2533 312 2567
rect 278 2465 312 2499
rect 278 2397 312 2431
rect 278 2329 312 2363
rect 278 2261 312 2295
rect 278 2193 312 2227
rect 278 2125 312 2159
rect 278 2057 312 2091
rect 278 1989 312 2023
rect 278 1921 312 1955
rect 278 1853 312 1887
rect 278 1785 312 1819
rect 278 1717 312 1751
rect 278 1649 312 1683
rect 278 1581 312 1615
rect 278 1513 312 1547
rect 278 1445 312 1479
rect 278 1377 312 1411
rect 278 1309 312 1343
rect 278 1241 312 1275
rect 278 1173 312 1207
rect 278 1105 312 1139
rect 278 1037 312 1071
rect 278 969 312 1003
rect 278 901 312 935
rect 278 833 312 867
rect 278 765 312 799
rect 278 697 312 731
rect 278 629 312 663
rect 278 561 312 595
rect 278 493 312 527
rect 278 425 312 459
rect 278 357 312 391
rect 278 289 312 323
rect 278 221 312 255
rect 278 153 312 187
rect 278 85 312 119
rect 278 17 312 51
rect 278 -51 312 -17
rect 278 -119 312 -85
rect 278 -187 312 -153
rect 278 -255 312 -221
rect 278 -323 312 -289
rect 278 -391 312 -357
rect 278 -459 312 -425
rect 278 -527 312 -493
rect 278 -595 312 -561
rect 278 -663 312 -629
rect 278 -731 312 -697
rect 278 -799 312 -765
rect 278 -867 312 -833
rect 278 -935 312 -901
rect 278 -1003 312 -969
rect 278 -1071 312 -1037
rect 278 -1139 312 -1105
rect 278 -1207 312 -1173
rect 278 -1275 312 -1241
rect 278 -1343 312 -1309
rect 278 -1411 312 -1377
rect 278 -1479 312 -1445
rect 278 -1547 312 -1513
rect 278 -1615 312 -1581
rect 278 -1683 312 -1649
rect 278 -1751 312 -1717
rect 278 -1819 312 -1785
rect 278 -1887 312 -1853
rect 278 -1955 312 -1921
rect 278 -2023 312 -1989
rect 278 -2091 312 -2057
rect 278 -2159 312 -2125
rect 278 -2227 312 -2193
rect 278 -2295 312 -2261
rect 278 -2363 312 -2329
rect 278 -2431 312 -2397
rect 278 -2499 312 -2465
rect 278 -2567 312 -2533
rect 278 -2635 312 -2601
rect 278 -2703 312 -2669
rect 278 -2771 312 -2737
rect 278 -2839 312 -2805
rect 278 -2907 312 -2873
rect 278 -2975 312 -2941
rect 278 -3043 312 -3009
rect 278 -3111 312 -3077
rect 278 -3179 312 -3145
rect 278 -3247 312 -3213
rect 278 -3315 312 -3281
rect 278 -3383 312 -3349
rect 278 -3451 312 -3417
rect 278 -3519 312 -3485
rect 278 -3587 312 -3553
rect 278 -3655 312 -3621
rect 278 -3723 312 -3689
rect 278 -3791 312 -3757
rect 278 -3859 312 -3825
rect 278 -3927 312 -3893
rect 278 -3995 312 -3961
rect 278 -4063 312 -4029
rect 278 -4131 312 -4097
rect 278 -4199 312 -4165
rect 278 -4267 312 -4233
rect 278 -4335 312 -4301
rect 278 -4403 312 -4369
rect 278 -4471 312 -4437
rect 278 -4539 312 -4505
rect 278 -4607 312 -4573
rect 278 -4675 312 -4641
rect 278 -4743 312 -4709
rect 278 -4811 312 -4777
rect 278 -4879 312 -4845
rect 278 -4947 312 -4913
rect 278 -5015 312 -4981
rect 278 -5083 312 -5049
rect 278 -5151 312 -5117
rect 278 -5219 312 -5185
rect 278 -5287 312 -5253
rect 278 -5355 312 -5321
rect 278 -5423 312 -5389
rect 278 -5491 312 -5457
rect 278 -5559 312 -5525
rect 278 -5627 312 -5593
rect 278 -5695 312 -5661
rect 278 -5763 312 -5729
rect 278 -5831 312 -5797
rect 278 -5899 312 -5865
rect 278 -5967 312 -5933
rect 278 -6035 312 -6001
rect 278 -6103 312 -6069
rect 278 -6171 312 -6137
rect 278 -6239 312 -6205
rect 278 -6307 312 -6273
rect 278 -6375 312 -6341
rect 278 -6443 312 -6409
rect 278 -6511 312 -6477
rect 278 -6579 312 -6545
rect 278 -6647 312 -6613
rect 278 -6715 312 -6681
rect 278 -6783 312 -6749
rect 278 -6851 312 -6817
rect 278 -6919 312 -6885
rect 278 -6987 312 -6953
rect 278 -7055 312 -7021
rect 278 -7123 312 -7089
rect 278 -7191 312 -7157
rect 278 -7259 312 -7225
rect 278 -7327 312 -7293
rect 278 -7395 312 -7361
rect 278 -7463 312 -7429
rect 278 -7531 312 -7497
rect 278 -7599 312 -7565
rect 278 -7667 312 -7633
rect 278 -7735 312 -7701
rect 278 -7803 312 -7769
rect 278 -7871 312 -7837
rect 278 -7939 312 -7905
rect 278 -8007 312 -7973
rect 278 -8075 312 -8041
rect 278 -8143 312 -8109
rect 278 -8211 312 -8177
rect 278 -8279 312 -8245
rect 278 -8347 312 -8313
rect 278 -8415 312 -8381
rect 278 -8483 312 -8449
rect 278 -8551 312 -8517
rect 278 -8619 312 -8585
rect 278 -8687 312 -8653
rect 278 -8755 312 -8721
rect 278 -8823 312 -8789
rect 278 -8891 312 -8857
rect 278 -8959 312 -8925
rect 278 -9027 312 -8993
rect 278 -9095 312 -9061
rect 278 -9163 312 -9129
rect 278 -9231 312 -9197
rect 278 -9299 312 -9265
rect 278 -9367 312 -9333
rect 278 -9435 312 -9401
rect 278 -9503 312 -9469
rect 278 -9571 312 -9537
rect 396 9537 430 9571
rect 396 9469 430 9503
rect 396 9401 430 9435
rect 396 9333 430 9367
rect 396 9265 430 9299
rect 396 9197 430 9231
rect 396 9129 430 9163
rect 396 9061 430 9095
rect 396 8993 430 9027
rect 396 8925 430 8959
rect 396 8857 430 8891
rect 396 8789 430 8823
rect 396 8721 430 8755
rect 396 8653 430 8687
rect 396 8585 430 8619
rect 396 8517 430 8551
rect 396 8449 430 8483
rect 396 8381 430 8415
rect 396 8313 430 8347
rect 396 8245 430 8279
rect 396 8177 430 8211
rect 396 8109 430 8143
rect 396 8041 430 8075
rect 396 7973 430 8007
rect 396 7905 430 7939
rect 396 7837 430 7871
rect 396 7769 430 7803
rect 396 7701 430 7735
rect 396 7633 430 7667
rect 396 7565 430 7599
rect 396 7497 430 7531
rect 396 7429 430 7463
rect 396 7361 430 7395
rect 396 7293 430 7327
rect 396 7225 430 7259
rect 396 7157 430 7191
rect 396 7089 430 7123
rect 396 7021 430 7055
rect 396 6953 430 6987
rect 396 6885 430 6919
rect 396 6817 430 6851
rect 396 6749 430 6783
rect 396 6681 430 6715
rect 396 6613 430 6647
rect 396 6545 430 6579
rect 396 6477 430 6511
rect 396 6409 430 6443
rect 396 6341 430 6375
rect 396 6273 430 6307
rect 396 6205 430 6239
rect 396 6137 430 6171
rect 396 6069 430 6103
rect 396 6001 430 6035
rect 396 5933 430 5967
rect 396 5865 430 5899
rect 396 5797 430 5831
rect 396 5729 430 5763
rect 396 5661 430 5695
rect 396 5593 430 5627
rect 396 5525 430 5559
rect 396 5457 430 5491
rect 396 5389 430 5423
rect 396 5321 430 5355
rect 396 5253 430 5287
rect 396 5185 430 5219
rect 396 5117 430 5151
rect 396 5049 430 5083
rect 396 4981 430 5015
rect 396 4913 430 4947
rect 396 4845 430 4879
rect 396 4777 430 4811
rect 396 4709 430 4743
rect 396 4641 430 4675
rect 396 4573 430 4607
rect 396 4505 430 4539
rect 396 4437 430 4471
rect 396 4369 430 4403
rect 396 4301 430 4335
rect 396 4233 430 4267
rect 396 4165 430 4199
rect 396 4097 430 4131
rect 396 4029 430 4063
rect 396 3961 430 3995
rect 396 3893 430 3927
rect 396 3825 430 3859
rect 396 3757 430 3791
rect 396 3689 430 3723
rect 396 3621 430 3655
rect 396 3553 430 3587
rect 396 3485 430 3519
rect 396 3417 430 3451
rect 396 3349 430 3383
rect 396 3281 430 3315
rect 396 3213 430 3247
rect 396 3145 430 3179
rect 396 3077 430 3111
rect 396 3009 430 3043
rect 396 2941 430 2975
rect 396 2873 430 2907
rect 396 2805 430 2839
rect 396 2737 430 2771
rect 396 2669 430 2703
rect 396 2601 430 2635
rect 396 2533 430 2567
rect 396 2465 430 2499
rect 396 2397 430 2431
rect 396 2329 430 2363
rect 396 2261 430 2295
rect 396 2193 430 2227
rect 396 2125 430 2159
rect 396 2057 430 2091
rect 396 1989 430 2023
rect 396 1921 430 1955
rect 396 1853 430 1887
rect 396 1785 430 1819
rect 396 1717 430 1751
rect 396 1649 430 1683
rect 396 1581 430 1615
rect 396 1513 430 1547
rect 396 1445 430 1479
rect 396 1377 430 1411
rect 396 1309 430 1343
rect 396 1241 430 1275
rect 396 1173 430 1207
rect 396 1105 430 1139
rect 396 1037 430 1071
rect 396 969 430 1003
rect 396 901 430 935
rect 396 833 430 867
rect 396 765 430 799
rect 396 697 430 731
rect 396 629 430 663
rect 396 561 430 595
rect 396 493 430 527
rect 396 425 430 459
rect 396 357 430 391
rect 396 289 430 323
rect 396 221 430 255
rect 396 153 430 187
rect 396 85 430 119
rect 396 17 430 51
rect 396 -51 430 -17
rect 396 -119 430 -85
rect 396 -187 430 -153
rect 396 -255 430 -221
rect 396 -323 430 -289
rect 396 -391 430 -357
rect 396 -459 430 -425
rect 396 -527 430 -493
rect 396 -595 430 -561
rect 396 -663 430 -629
rect 396 -731 430 -697
rect 396 -799 430 -765
rect 396 -867 430 -833
rect 396 -935 430 -901
rect 396 -1003 430 -969
rect 396 -1071 430 -1037
rect 396 -1139 430 -1105
rect 396 -1207 430 -1173
rect 396 -1275 430 -1241
rect 396 -1343 430 -1309
rect 396 -1411 430 -1377
rect 396 -1479 430 -1445
rect 396 -1547 430 -1513
rect 396 -1615 430 -1581
rect 396 -1683 430 -1649
rect 396 -1751 430 -1717
rect 396 -1819 430 -1785
rect 396 -1887 430 -1853
rect 396 -1955 430 -1921
rect 396 -2023 430 -1989
rect 396 -2091 430 -2057
rect 396 -2159 430 -2125
rect 396 -2227 430 -2193
rect 396 -2295 430 -2261
rect 396 -2363 430 -2329
rect 396 -2431 430 -2397
rect 396 -2499 430 -2465
rect 396 -2567 430 -2533
rect 396 -2635 430 -2601
rect 396 -2703 430 -2669
rect 396 -2771 430 -2737
rect 396 -2839 430 -2805
rect 396 -2907 430 -2873
rect 396 -2975 430 -2941
rect 396 -3043 430 -3009
rect 396 -3111 430 -3077
rect 396 -3179 430 -3145
rect 396 -3247 430 -3213
rect 396 -3315 430 -3281
rect 396 -3383 430 -3349
rect 396 -3451 430 -3417
rect 396 -3519 430 -3485
rect 396 -3587 430 -3553
rect 396 -3655 430 -3621
rect 396 -3723 430 -3689
rect 396 -3791 430 -3757
rect 396 -3859 430 -3825
rect 396 -3927 430 -3893
rect 396 -3995 430 -3961
rect 396 -4063 430 -4029
rect 396 -4131 430 -4097
rect 396 -4199 430 -4165
rect 396 -4267 430 -4233
rect 396 -4335 430 -4301
rect 396 -4403 430 -4369
rect 396 -4471 430 -4437
rect 396 -4539 430 -4505
rect 396 -4607 430 -4573
rect 396 -4675 430 -4641
rect 396 -4743 430 -4709
rect 396 -4811 430 -4777
rect 396 -4879 430 -4845
rect 396 -4947 430 -4913
rect 396 -5015 430 -4981
rect 396 -5083 430 -5049
rect 396 -5151 430 -5117
rect 396 -5219 430 -5185
rect 396 -5287 430 -5253
rect 396 -5355 430 -5321
rect 396 -5423 430 -5389
rect 396 -5491 430 -5457
rect 396 -5559 430 -5525
rect 396 -5627 430 -5593
rect 396 -5695 430 -5661
rect 396 -5763 430 -5729
rect 396 -5831 430 -5797
rect 396 -5899 430 -5865
rect 396 -5967 430 -5933
rect 396 -6035 430 -6001
rect 396 -6103 430 -6069
rect 396 -6171 430 -6137
rect 396 -6239 430 -6205
rect 396 -6307 430 -6273
rect 396 -6375 430 -6341
rect 396 -6443 430 -6409
rect 396 -6511 430 -6477
rect 396 -6579 430 -6545
rect 396 -6647 430 -6613
rect 396 -6715 430 -6681
rect 396 -6783 430 -6749
rect 396 -6851 430 -6817
rect 396 -6919 430 -6885
rect 396 -6987 430 -6953
rect 396 -7055 430 -7021
rect 396 -7123 430 -7089
rect 396 -7191 430 -7157
rect 396 -7259 430 -7225
rect 396 -7327 430 -7293
rect 396 -7395 430 -7361
rect 396 -7463 430 -7429
rect 396 -7531 430 -7497
rect 396 -7599 430 -7565
rect 396 -7667 430 -7633
rect 396 -7735 430 -7701
rect 396 -7803 430 -7769
rect 396 -7871 430 -7837
rect 396 -7939 430 -7905
rect 396 -8007 430 -7973
rect 396 -8075 430 -8041
rect 396 -8143 430 -8109
rect 396 -8211 430 -8177
rect 396 -8279 430 -8245
rect 396 -8347 430 -8313
rect 396 -8415 430 -8381
rect 396 -8483 430 -8449
rect 396 -8551 430 -8517
rect 396 -8619 430 -8585
rect 396 -8687 430 -8653
rect 396 -8755 430 -8721
rect 396 -8823 430 -8789
rect 396 -8891 430 -8857
rect 396 -8959 430 -8925
rect 396 -9027 430 -8993
rect 396 -9095 430 -9061
rect 396 -9163 430 -9129
rect 396 -9231 430 -9197
rect 396 -9299 430 -9265
rect 396 -9367 430 -9333
rect 396 -9435 430 -9401
rect 396 -9503 430 -9469
rect 396 -9571 430 -9537
rect 514 9537 548 9571
rect 514 9469 548 9503
rect 514 9401 548 9435
rect 514 9333 548 9367
rect 514 9265 548 9299
rect 514 9197 548 9231
rect 514 9129 548 9163
rect 514 9061 548 9095
rect 514 8993 548 9027
rect 514 8925 548 8959
rect 514 8857 548 8891
rect 514 8789 548 8823
rect 514 8721 548 8755
rect 514 8653 548 8687
rect 514 8585 548 8619
rect 514 8517 548 8551
rect 514 8449 548 8483
rect 514 8381 548 8415
rect 514 8313 548 8347
rect 514 8245 548 8279
rect 514 8177 548 8211
rect 514 8109 548 8143
rect 514 8041 548 8075
rect 514 7973 548 8007
rect 514 7905 548 7939
rect 514 7837 548 7871
rect 514 7769 548 7803
rect 514 7701 548 7735
rect 514 7633 548 7667
rect 514 7565 548 7599
rect 514 7497 548 7531
rect 514 7429 548 7463
rect 514 7361 548 7395
rect 514 7293 548 7327
rect 514 7225 548 7259
rect 514 7157 548 7191
rect 514 7089 548 7123
rect 514 7021 548 7055
rect 514 6953 548 6987
rect 514 6885 548 6919
rect 514 6817 548 6851
rect 514 6749 548 6783
rect 514 6681 548 6715
rect 514 6613 548 6647
rect 514 6545 548 6579
rect 514 6477 548 6511
rect 514 6409 548 6443
rect 514 6341 548 6375
rect 514 6273 548 6307
rect 514 6205 548 6239
rect 514 6137 548 6171
rect 514 6069 548 6103
rect 514 6001 548 6035
rect 514 5933 548 5967
rect 514 5865 548 5899
rect 514 5797 548 5831
rect 514 5729 548 5763
rect 514 5661 548 5695
rect 514 5593 548 5627
rect 514 5525 548 5559
rect 514 5457 548 5491
rect 514 5389 548 5423
rect 514 5321 548 5355
rect 514 5253 548 5287
rect 514 5185 548 5219
rect 514 5117 548 5151
rect 514 5049 548 5083
rect 514 4981 548 5015
rect 514 4913 548 4947
rect 514 4845 548 4879
rect 514 4777 548 4811
rect 514 4709 548 4743
rect 514 4641 548 4675
rect 514 4573 548 4607
rect 514 4505 548 4539
rect 514 4437 548 4471
rect 514 4369 548 4403
rect 514 4301 548 4335
rect 514 4233 548 4267
rect 514 4165 548 4199
rect 514 4097 548 4131
rect 514 4029 548 4063
rect 514 3961 548 3995
rect 514 3893 548 3927
rect 514 3825 548 3859
rect 514 3757 548 3791
rect 514 3689 548 3723
rect 514 3621 548 3655
rect 514 3553 548 3587
rect 514 3485 548 3519
rect 514 3417 548 3451
rect 514 3349 548 3383
rect 514 3281 548 3315
rect 514 3213 548 3247
rect 514 3145 548 3179
rect 514 3077 548 3111
rect 514 3009 548 3043
rect 514 2941 548 2975
rect 514 2873 548 2907
rect 514 2805 548 2839
rect 514 2737 548 2771
rect 514 2669 548 2703
rect 514 2601 548 2635
rect 514 2533 548 2567
rect 514 2465 548 2499
rect 514 2397 548 2431
rect 514 2329 548 2363
rect 514 2261 548 2295
rect 514 2193 548 2227
rect 514 2125 548 2159
rect 514 2057 548 2091
rect 514 1989 548 2023
rect 514 1921 548 1955
rect 514 1853 548 1887
rect 514 1785 548 1819
rect 514 1717 548 1751
rect 514 1649 548 1683
rect 514 1581 548 1615
rect 514 1513 548 1547
rect 514 1445 548 1479
rect 514 1377 548 1411
rect 514 1309 548 1343
rect 514 1241 548 1275
rect 514 1173 548 1207
rect 514 1105 548 1139
rect 514 1037 548 1071
rect 514 969 548 1003
rect 514 901 548 935
rect 514 833 548 867
rect 514 765 548 799
rect 514 697 548 731
rect 514 629 548 663
rect 514 561 548 595
rect 514 493 548 527
rect 514 425 548 459
rect 514 357 548 391
rect 514 289 548 323
rect 514 221 548 255
rect 514 153 548 187
rect 514 85 548 119
rect 514 17 548 51
rect 514 -51 548 -17
rect 514 -119 548 -85
rect 514 -187 548 -153
rect 514 -255 548 -221
rect 514 -323 548 -289
rect 514 -391 548 -357
rect 514 -459 548 -425
rect 514 -527 548 -493
rect 514 -595 548 -561
rect 514 -663 548 -629
rect 514 -731 548 -697
rect 514 -799 548 -765
rect 514 -867 548 -833
rect 514 -935 548 -901
rect 514 -1003 548 -969
rect 514 -1071 548 -1037
rect 514 -1139 548 -1105
rect 514 -1207 548 -1173
rect 514 -1275 548 -1241
rect 514 -1343 548 -1309
rect 514 -1411 548 -1377
rect 514 -1479 548 -1445
rect 514 -1547 548 -1513
rect 514 -1615 548 -1581
rect 514 -1683 548 -1649
rect 514 -1751 548 -1717
rect 514 -1819 548 -1785
rect 514 -1887 548 -1853
rect 514 -1955 548 -1921
rect 514 -2023 548 -1989
rect 514 -2091 548 -2057
rect 514 -2159 548 -2125
rect 514 -2227 548 -2193
rect 514 -2295 548 -2261
rect 514 -2363 548 -2329
rect 514 -2431 548 -2397
rect 514 -2499 548 -2465
rect 514 -2567 548 -2533
rect 514 -2635 548 -2601
rect 514 -2703 548 -2669
rect 514 -2771 548 -2737
rect 514 -2839 548 -2805
rect 514 -2907 548 -2873
rect 514 -2975 548 -2941
rect 514 -3043 548 -3009
rect 514 -3111 548 -3077
rect 514 -3179 548 -3145
rect 514 -3247 548 -3213
rect 514 -3315 548 -3281
rect 514 -3383 548 -3349
rect 514 -3451 548 -3417
rect 514 -3519 548 -3485
rect 514 -3587 548 -3553
rect 514 -3655 548 -3621
rect 514 -3723 548 -3689
rect 514 -3791 548 -3757
rect 514 -3859 548 -3825
rect 514 -3927 548 -3893
rect 514 -3995 548 -3961
rect 514 -4063 548 -4029
rect 514 -4131 548 -4097
rect 514 -4199 548 -4165
rect 514 -4267 548 -4233
rect 514 -4335 548 -4301
rect 514 -4403 548 -4369
rect 514 -4471 548 -4437
rect 514 -4539 548 -4505
rect 514 -4607 548 -4573
rect 514 -4675 548 -4641
rect 514 -4743 548 -4709
rect 514 -4811 548 -4777
rect 514 -4879 548 -4845
rect 514 -4947 548 -4913
rect 514 -5015 548 -4981
rect 514 -5083 548 -5049
rect 514 -5151 548 -5117
rect 514 -5219 548 -5185
rect 514 -5287 548 -5253
rect 514 -5355 548 -5321
rect 514 -5423 548 -5389
rect 514 -5491 548 -5457
rect 514 -5559 548 -5525
rect 514 -5627 548 -5593
rect 514 -5695 548 -5661
rect 514 -5763 548 -5729
rect 514 -5831 548 -5797
rect 514 -5899 548 -5865
rect 514 -5967 548 -5933
rect 514 -6035 548 -6001
rect 514 -6103 548 -6069
rect 514 -6171 548 -6137
rect 514 -6239 548 -6205
rect 514 -6307 548 -6273
rect 514 -6375 548 -6341
rect 514 -6443 548 -6409
rect 514 -6511 548 -6477
rect 514 -6579 548 -6545
rect 514 -6647 548 -6613
rect 514 -6715 548 -6681
rect 514 -6783 548 -6749
rect 514 -6851 548 -6817
rect 514 -6919 548 -6885
rect 514 -6987 548 -6953
rect 514 -7055 548 -7021
rect 514 -7123 548 -7089
rect 514 -7191 548 -7157
rect 514 -7259 548 -7225
rect 514 -7327 548 -7293
rect 514 -7395 548 -7361
rect 514 -7463 548 -7429
rect 514 -7531 548 -7497
rect 514 -7599 548 -7565
rect 514 -7667 548 -7633
rect 514 -7735 548 -7701
rect 514 -7803 548 -7769
rect 514 -7871 548 -7837
rect 514 -7939 548 -7905
rect 514 -8007 548 -7973
rect 514 -8075 548 -8041
rect 514 -8143 548 -8109
rect 514 -8211 548 -8177
rect 514 -8279 548 -8245
rect 514 -8347 548 -8313
rect 514 -8415 548 -8381
rect 514 -8483 548 -8449
rect 514 -8551 548 -8517
rect 514 -8619 548 -8585
rect 514 -8687 548 -8653
rect 514 -8755 548 -8721
rect 514 -8823 548 -8789
rect 514 -8891 548 -8857
rect 514 -8959 548 -8925
rect 514 -9027 548 -8993
rect 514 -9095 548 -9061
rect 514 -9163 548 -9129
rect 514 -9231 548 -9197
rect 514 -9299 548 -9265
rect 514 -9367 548 -9333
rect 514 -9435 548 -9401
rect 514 -9503 548 -9469
rect 514 -9571 548 -9537
rect 632 9537 666 9571
rect 632 9469 666 9503
rect 632 9401 666 9435
rect 632 9333 666 9367
rect 632 9265 666 9299
rect 632 9197 666 9231
rect 632 9129 666 9163
rect 632 9061 666 9095
rect 632 8993 666 9027
rect 632 8925 666 8959
rect 632 8857 666 8891
rect 632 8789 666 8823
rect 632 8721 666 8755
rect 632 8653 666 8687
rect 632 8585 666 8619
rect 632 8517 666 8551
rect 632 8449 666 8483
rect 632 8381 666 8415
rect 632 8313 666 8347
rect 632 8245 666 8279
rect 632 8177 666 8211
rect 632 8109 666 8143
rect 632 8041 666 8075
rect 632 7973 666 8007
rect 632 7905 666 7939
rect 632 7837 666 7871
rect 632 7769 666 7803
rect 632 7701 666 7735
rect 632 7633 666 7667
rect 632 7565 666 7599
rect 632 7497 666 7531
rect 632 7429 666 7463
rect 632 7361 666 7395
rect 632 7293 666 7327
rect 632 7225 666 7259
rect 632 7157 666 7191
rect 632 7089 666 7123
rect 632 7021 666 7055
rect 632 6953 666 6987
rect 632 6885 666 6919
rect 632 6817 666 6851
rect 632 6749 666 6783
rect 632 6681 666 6715
rect 632 6613 666 6647
rect 632 6545 666 6579
rect 632 6477 666 6511
rect 632 6409 666 6443
rect 632 6341 666 6375
rect 632 6273 666 6307
rect 632 6205 666 6239
rect 632 6137 666 6171
rect 632 6069 666 6103
rect 632 6001 666 6035
rect 632 5933 666 5967
rect 632 5865 666 5899
rect 632 5797 666 5831
rect 632 5729 666 5763
rect 632 5661 666 5695
rect 632 5593 666 5627
rect 632 5525 666 5559
rect 632 5457 666 5491
rect 632 5389 666 5423
rect 632 5321 666 5355
rect 632 5253 666 5287
rect 632 5185 666 5219
rect 632 5117 666 5151
rect 632 5049 666 5083
rect 632 4981 666 5015
rect 632 4913 666 4947
rect 632 4845 666 4879
rect 632 4777 666 4811
rect 632 4709 666 4743
rect 632 4641 666 4675
rect 632 4573 666 4607
rect 632 4505 666 4539
rect 632 4437 666 4471
rect 632 4369 666 4403
rect 632 4301 666 4335
rect 632 4233 666 4267
rect 632 4165 666 4199
rect 632 4097 666 4131
rect 632 4029 666 4063
rect 632 3961 666 3995
rect 632 3893 666 3927
rect 632 3825 666 3859
rect 632 3757 666 3791
rect 632 3689 666 3723
rect 632 3621 666 3655
rect 632 3553 666 3587
rect 632 3485 666 3519
rect 632 3417 666 3451
rect 632 3349 666 3383
rect 632 3281 666 3315
rect 632 3213 666 3247
rect 632 3145 666 3179
rect 632 3077 666 3111
rect 632 3009 666 3043
rect 632 2941 666 2975
rect 632 2873 666 2907
rect 632 2805 666 2839
rect 632 2737 666 2771
rect 632 2669 666 2703
rect 632 2601 666 2635
rect 632 2533 666 2567
rect 632 2465 666 2499
rect 632 2397 666 2431
rect 632 2329 666 2363
rect 632 2261 666 2295
rect 632 2193 666 2227
rect 632 2125 666 2159
rect 632 2057 666 2091
rect 632 1989 666 2023
rect 632 1921 666 1955
rect 632 1853 666 1887
rect 632 1785 666 1819
rect 632 1717 666 1751
rect 632 1649 666 1683
rect 632 1581 666 1615
rect 632 1513 666 1547
rect 632 1445 666 1479
rect 632 1377 666 1411
rect 632 1309 666 1343
rect 632 1241 666 1275
rect 632 1173 666 1207
rect 632 1105 666 1139
rect 632 1037 666 1071
rect 632 969 666 1003
rect 632 901 666 935
rect 632 833 666 867
rect 632 765 666 799
rect 632 697 666 731
rect 632 629 666 663
rect 632 561 666 595
rect 632 493 666 527
rect 632 425 666 459
rect 632 357 666 391
rect 632 289 666 323
rect 632 221 666 255
rect 632 153 666 187
rect 632 85 666 119
rect 632 17 666 51
rect 632 -51 666 -17
rect 632 -119 666 -85
rect 632 -187 666 -153
rect 632 -255 666 -221
rect 632 -323 666 -289
rect 632 -391 666 -357
rect 632 -459 666 -425
rect 632 -527 666 -493
rect 632 -595 666 -561
rect 632 -663 666 -629
rect 632 -731 666 -697
rect 632 -799 666 -765
rect 632 -867 666 -833
rect 632 -935 666 -901
rect 632 -1003 666 -969
rect 632 -1071 666 -1037
rect 632 -1139 666 -1105
rect 632 -1207 666 -1173
rect 632 -1275 666 -1241
rect 632 -1343 666 -1309
rect 632 -1411 666 -1377
rect 632 -1479 666 -1445
rect 632 -1547 666 -1513
rect 632 -1615 666 -1581
rect 632 -1683 666 -1649
rect 632 -1751 666 -1717
rect 632 -1819 666 -1785
rect 632 -1887 666 -1853
rect 632 -1955 666 -1921
rect 632 -2023 666 -1989
rect 632 -2091 666 -2057
rect 632 -2159 666 -2125
rect 632 -2227 666 -2193
rect 632 -2295 666 -2261
rect 632 -2363 666 -2329
rect 632 -2431 666 -2397
rect 632 -2499 666 -2465
rect 632 -2567 666 -2533
rect 632 -2635 666 -2601
rect 632 -2703 666 -2669
rect 632 -2771 666 -2737
rect 632 -2839 666 -2805
rect 632 -2907 666 -2873
rect 632 -2975 666 -2941
rect 632 -3043 666 -3009
rect 632 -3111 666 -3077
rect 632 -3179 666 -3145
rect 632 -3247 666 -3213
rect 632 -3315 666 -3281
rect 632 -3383 666 -3349
rect 632 -3451 666 -3417
rect 632 -3519 666 -3485
rect 632 -3587 666 -3553
rect 632 -3655 666 -3621
rect 632 -3723 666 -3689
rect 632 -3791 666 -3757
rect 632 -3859 666 -3825
rect 632 -3927 666 -3893
rect 632 -3995 666 -3961
rect 632 -4063 666 -4029
rect 632 -4131 666 -4097
rect 632 -4199 666 -4165
rect 632 -4267 666 -4233
rect 632 -4335 666 -4301
rect 632 -4403 666 -4369
rect 632 -4471 666 -4437
rect 632 -4539 666 -4505
rect 632 -4607 666 -4573
rect 632 -4675 666 -4641
rect 632 -4743 666 -4709
rect 632 -4811 666 -4777
rect 632 -4879 666 -4845
rect 632 -4947 666 -4913
rect 632 -5015 666 -4981
rect 632 -5083 666 -5049
rect 632 -5151 666 -5117
rect 632 -5219 666 -5185
rect 632 -5287 666 -5253
rect 632 -5355 666 -5321
rect 632 -5423 666 -5389
rect 632 -5491 666 -5457
rect 632 -5559 666 -5525
rect 632 -5627 666 -5593
rect 632 -5695 666 -5661
rect 632 -5763 666 -5729
rect 632 -5831 666 -5797
rect 632 -5899 666 -5865
rect 632 -5967 666 -5933
rect 632 -6035 666 -6001
rect 632 -6103 666 -6069
rect 632 -6171 666 -6137
rect 632 -6239 666 -6205
rect 632 -6307 666 -6273
rect 632 -6375 666 -6341
rect 632 -6443 666 -6409
rect 632 -6511 666 -6477
rect 632 -6579 666 -6545
rect 632 -6647 666 -6613
rect 632 -6715 666 -6681
rect 632 -6783 666 -6749
rect 632 -6851 666 -6817
rect 632 -6919 666 -6885
rect 632 -6987 666 -6953
rect 632 -7055 666 -7021
rect 632 -7123 666 -7089
rect 632 -7191 666 -7157
rect 632 -7259 666 -7225
rect 632 -7327 666 -7293
rect 632 -7395 666 -7361
rect 632 -7463 666 -7429
rect 632 -7531 666 -7497
rect 632 -7599 666 -7565
rect 632 -7667 666 -7633
rect 632 -7735 666 -7701
rect 632 -7803 666 -7769
rect 632 -7871 666 -7837
rect 632 -7939 666 -7905
rect 632 -8007 666 -7973
rect 632 -8075 666 -8041
rect 632 -8143 666 -8109
rect 632 -8211 666 -8177
rect 632 -8279 666 -8245
rect 632 -8347 666 -8313
rect 632 -8415 666 -8381
rect 632 -8483 666 -8449
rect 632 -8551 666 -8517
rect 632 -8619 666 -8585
rect 632 -8687 666 -8653
rect 632 -8755 666 -8721
rect 632 -8823 666 -8789
rect 632 -8891 666 -8857
rect 632 -8959 666 -8925
rect 632 -9027 666 -8993
rect 632 -9095 666 -9061
rect 632 -9163 666 -9129
rect 632 -9231 666 -9197
rect 632 -9299 666 -9265
rect 632 -9367 666 -9333
rect 632 -9435 666 -9401
rect 632 -9503 666 -9469
rect 632 -9571 666 -9537
rect 750 9537 784 9571
rect 750 9469 784 9503
rect 750 9401 784 9435
rect 750 9333 784 9367
rect 750 9265 784 9299
rect 750 9197 784 9231
rect 750 9129 784 9163
rect 750 9061 784 9095
rect 750 8993 784 9027
rect 750 8925 784 8959
rect 750 8857 784 8891
rect 750 8789 784 8823
rect 750 8721 784 8755
rect 750 8653 784 8687
rect 750 8585 784 8619
rect 750 8517 784 8551
rect 750 8449 784 8483
rect 750 8381 784 8415
rect 750 8313 784 8347
rect 750 8245 784 8279
rect 750 8177 784 8211
rect 750 8109 784 8143
rect 750 8041 784 8075
rect 750 7973 784 8007
rect 750 7905 784 7939
rect 750 7837 784 7871
rect 750 7769 784 7803
rect 750 7701 784 7735
rect 750 7633 784 7667
rect 750 7565 784 7599
rect 750 7497 784 7531
rect 750 7429 784 7463
rect 750 7361 784 7395
rect 750 7293 784 7327
rect 750 7225 784 7259
rect 750 7157 784 7191
rect 750 7089 784 7123
rect 750 7021 784 7055
rect 750 6953 784 6987
rect 750 6885 784 6919
rect 750 6817 784 6851
rect 750 6749 784 6783
rect 750 6681 784 6715
rect 750 6613 784 6647
rect 750 6545 784 6579
rect 750 6477 784 6511
rect 750 6409 784 6443
rect 750 6341 784 6375
rect 750 6273 784 6307
rect 750 6205 784 6239
rect 750 6137 784 6171
rect 750 6069 784 6103
rect 750 6001 784 6035
rect 750 5933 784 5967
rect 750 5865 784 5899
rect 750 5797 784 5831
rect 750 5729 784 5763
rect 750 5661 784 5695
rect 750 5593 784 5627
rect 750 5525 784 5559
rect 750 5457 784 5491
rect 750 5389 784 5423
rect 750 5321 784 5355
rect 750 5253 784 5287
rect 750 5185 784 5219
rect 750 5117 784 5151
rect 750 5049 784 5083
rect 750 4981 784 5015
rect 750 4913 784 4947
rect 750 4845 784 4879
rect 750 4777 784 4811
rect 750 4709 784 4743
rect 750 4641 784 4675
rect 750 4573 784 4607
rect 750 4505 784 4539
rect 750 4437 784 4471
rect 750 4369 784 4403
rect 750 4301 784 4335
rect 750 4233 784 4267
rect 750 4165 784 4199
rect 750 4097 784 4131
rect 750 4029 784 4063
rect 750 3961 784 3995
rect 750 3893 784 3927
rect 750 3825 784 3859
rect 750 3757 784 3791
rect 750 3689 784 3723
rect 750 3621 784 3655
rect 750 3553 784 3587
rect 750 3485 784 3519
rect 750 3417 784 3451
rect 750 3349 784 3383
rect 750 3281 784 3315
rect 750 3213 784 3247
rect 750 3145 784 3179
rect 750 3077 784 3111
rect 750 3009 784 3043
rect 750 2941 784 2975
rect 750 2873 784 2907
rect 750 2805 784 2839
rect 750 2737 784 2771
rect 750 2669 784 2703
rect 750 2601 784 2635
rect 750 2533 784 2567
rect 750 2465 784 2499
rect 750 2397 784 2431
rect 750 2329 784 2363
rect 750 2261 784 2295
rect 750 2193 784 2227
rect 750 2125 784 2159
rect 750 2057 784 2091
rect 750 1989 784 2023
rect 750 1921 784 1955
rect 750 1853 784 1887
rect 750 1785 784 1819
rect 750 1717 784 1751
rect 750 1649 784 1683
rect 750 1581 784 1615
rect 750 1513 784 1547
rect 750 1445 784 1479
rect 750 1377 784 1411
rect 750 1309 784 1343
rect 750 1241 784 1275
rect 750 1173 784 1207
rect 750 1105 784 1139
rect 750 1037 784 1071
rect 750 969 784 1003
rect 750 901 784 935
rect 750 833 784 867
rect 750 765 784 799
rect 750 697 784 731
rect 750 629 784 663
rect 750 561 784 595
rect 750 493 784 527
rect 750 425 784 459
rect 750 357 784 391
rect 750 289 784 323
rect 750 221 784 255
rect 750 153 784 187
rect 750 85 784 119
rect 750 17 784 51
rect 750 -51 784 -17
rect 750 -119 784 -85
rect 750 -187 784 -153
rect 750 -255 784 -221
rect 750 -323 784 -289
rect 750 -391 784 -357
rect 750 -459 784 -425
rect 750 -527 784 -493
rect 750 -595 784 -561
rect 750 -663 784 -629
rect 750 -731 784 -697
rect 750 -799 784 -765
rect 750 -867 784 -833
rect 750 -935 784 -901
rect 750 -1003 784 -969
rect 750 -1071 784 -1037
rect 750 -1139 784 -1105
rect 750 -1207 784 -1173
rect 750 -1275 784 -1241
rect 750 -1343 784 -1309
rect 750 -1411 784 -1377
rect 750 -1479 784 -1445
rect 750 -1547 784 -1513
rect 750 -1615 784 -1581
rect 750 -1683 784 -1649
rect 750 -1751 784 -1717
rect 750 -1819 784 -1785
rect 750 -1887 784 -1853
rect 750 -1955 784 -1921
rect 750 -2023 784 -1989
rect 750 -2091 784 -2057
rect 750 -2159 784 -2125
rect 750 -2227 784 -2193
rect 750 -2295 784 -2261
rect 750 -2363 784 -2329
rect 750 -2431 784 -2397
rect 750 -2499 784 -2465
rect 750 -2567 784 -2533
rect 750 -2635 784 -2601
rect 750 -2703 784 -2669
rect 750 -2771 784 -2737
rect 750 -2839 784 -2805
rect 750 -2907 784 -2873
rect 750 -2975 784 -2941
rect 750 -3043 784 -3009
rect 750 -3111 784 -3077
rect 750 -3179 784 -3145
rect 750 -3247 784 -3213
rect 750 -3315 784 -3281
rect 750 -3383 784 -3349
rect 750 -3451 784 -3417
rect 750 -3519 784 -3485
rect 750 -3587 784 -3553
rect 750 -3655 784 -3621
rect 750 -3723 784 -3689
rect 750 -3791 784 -3757
rect 750 -3859 784 -3825
rect 750 -3927 784 -3893
rect 750 -3995 784 -3961
rect 750 -4063 784 -4029
rect 750 -4131 784 -4097
rect 750 -4199 784 -4165
rect 750 -4267 784 -4233
rect 750 -4335 784 -4301
rect 750 -4403 784 -4369
rect 750 -4471 784 -4437
rect 750 -4539 784 -4505
rect 750 -4607 784 -4573
rect 750 -4675 784 -4641
rect 750 -4743 784 -4709
rect 750 -4811 784 -4777
rect 750 -4879 784 -4845
rect 750 -4947 784 -4913
rect 750 -5015 784 -4981
rect 750 -5083 784 -5049
rect 750 -5151 784 -5117
rect 750 -5219 784 -5185
rect 750 -5287 784 -5253
rect 750 -5355 784 -5321
rect 750 -5423 784 -5389
rect 750 -5491 784 -5457
rect 750 -5559 784 -5525
rect 750 -5627 784 -5593
rect 750 -5695 784 -5661
rect 750 -5763 784 -5729
rect 750 -5831 784 -5797
rect 750 -5899 784 -5865
rect 750 -5967 784 -5933
rect 750 -6035 784 -6001
rect 750 -6103 784 -6069
rect 750 -6171 784 -6137
rect 750 -6239 784 -6205
rect 750 -6307 784 -6273
rect 750 -6375 784 -6341
rect 750 -6443 784 -6409
rect 750 -6511 784 -6477
rect 750 -6579 784 -6545
rect 750 -6647 784 -6613
rect 750 -6715 784 -6681
rect 750 -6783 784 -6749
rect 750 -6851 784 -6817
rect 750 -6919 784 -6885
rect 750 -6987 784 -6953
rect 750 -7055 784 -7021
rect 750 -7123 784 -7089
rect 750 -7191 784 -7157
rect 750 -7259 784 -7225
rect 750 -7327 784 -7293
rect 750 -7395 784 -7361
rect 750 -7463 784 -7429
rect 750 -7531 784 -7497
rect 750 -7599 784 -7565
rect 750 -7667 784 -7633
rect 750 -7735 784 -7701
rect 750 -7803 784 -7769
rect 750 -7871 784 -7837
rect 750 -7939 784 -7905
rect 750 -8007 784 -7973
rect 750 -8075 784 -8041
rect 750 -8143 784 -8109
rect 750 -8211 784 -8177
rect 750 -8279 784 -8245
rect 750 -8347 784 -8313
rect 750 -8415 784 -8381
rect 750 -8483 784 -8449
rect 750 -8551 784 -8517
rect 750 -8619 784 -8585
rect 750 -8687 784 -8653
rect 750 -8755 784 -8721
rect 750 -8823 784 -8789
rect 750 -8891 784 -8857
rect 750 -8959 784 -8925
rect 750 -9027 784 -8993
rect 750 -9095 784 -9061
rect 750 -9163 784 -9129
rect 750 -9231 784 -9197
rect 750 -9299 784 -9265
rect 750 -9367 784 -9333
rect 750 -9435 784 -9401
rect 750 -9503 784 -9469
rect 750 -9571 784 -9537
rect 868 9537 902 9571
rect 868 9469 902 9503
rect 868 9401 902 9435
rect 868 9333 902 9367
rect 868 9265 902 9299
rect 868 9197 902 9231
rect 868 9129 902 9163
rect 868 9061 902 9095
rect 868 8993 902 9027
rect 868 8925 902 8959
rect 868 8857 902 8891
rect 868 8789 902 8823
rect 868 8721 902 8755
rect 868 8653 902 8687
rect 868 8585 902 8619
rect 868 8517 902 8551
rect 868 8449 902 8483
rect 868 8381 902 8415
rect 868 8313 902 8347
rect 868 8245 902 8279
rect 868 8177 902 8211
rect 868 8109 902 8143
rect 868 8041 902 8075
rect 868 7973 902 8007
rect 868 7905 902 7939
rect 868 7837 902 7871
rect 868 7769 902 7803
rect 868 7701 902 7735
rect 868 7633 902 7667
rect 868 7565 902 7599
rect 868 7497 902 7531
rect 868 7429 902 7463
rect 868 7361 902 7395
rect 868 7293 902 7327
rect 868 7225 902 7259
rect 868 7157 902 7191
rect 868 7089 902 7123
rect 868 7021 902 7055
rect 868 6953 902 6987
rect 868 6885 902 6919
rect 868 6817 902 6851
rect 868 6749 902 6783
rect 868 6681 902 6715
rect 868 6613 902 6647
rect 868 6545 902 6579
rect 868 6477 902 6511
rect 868 6409 902 6443
rect 868 6341 902 6375
rect 868 6273 902 6307
rect 868 6205 902 6239
rect 868 6137 902 6171
rect 868 6069 902 6103
rect 868 6001 902 6035
rect 868 5933 902 5967
rect 868 5865 902 5899
rect 868 5797 902 5831
rect 868 5729 902 5763
rect 868 5661 902 5695
rect 868 5593 902 5627
rect 868 5525 902 5559
rect 868 5457 902 5491
rect 868 5389 902 5423
rect 868 5321 902 5355
rect 868 5253 902 5287
rect 868 5185 902 5219
rect 868 5117 902 5151
rect 868 5049 902 5083
rect 868 4981 902 5015
rect 868 4913 902 4947
rect 868 4845 902 4879
rect 868 4777 902 4811
rect 868 4709 902 4743
rect 868 4641 902 4675
rect 868 4573 902 4607
rect 868 4505 902 4539
rect 868 4437 902 4471
rect 868 4369 902 4403
rect 868 4301 902 4335
rect 868 4233 902 4267
rect 868 4165 902 4199
rect 868 4097 902 4131
rect 868 4029 902 4063
rect 868 3961 902 3995
rect 868 3893 902 3927
rect 868 3825 902 3859
rect 868 3757 902 3791
rect 868 3689 902 3723
rect 868 3621 902 3655
rect 868 3553 902 3587
rect 868 3485 902 3519
rect 868 3417 902 3451
rect 868 3349 902 3383
rect 868 3281 902 3315
rect 868 3213 902 3247
rect 868 3145 902 3179
rect 868 3077 902 3111
rect 868 3009 902 3043
rect 868 2941 902 2975
rect 868 2873 902 2907
rect 868 2805 902 2839
rect 868 2737 902 2771
rect 868 2669 902 2703
rect 868 2601 902 2635
rect 868 2533 902 2567
rect 868 2465 902 2499
rect 868 2397 902 2431
rect 868 2329 902 2363
rect 868 2261 902 2295
rect 868 2193 902 2227
rect 868 2125 902 2159
rect 868 2057 902 2091
rect 868 1989 902 2023
rect 868 1921 902 1955
rect 868 1853 902 1887
rect 868 1785 902 1819
rect 868 1717 902 1751
rect 868 1649 902 1683
rect 868 1581 902 1615
rect 868 1513 902 1547
rect 868 1445 902 1479
rect 868 1377 902 1411
rect 868 1309 902 1343
rect 868 1241 902 1275
rect 868 1173 902 1207
rect 868 1105 902 1139
rect 868 1037 902 1071
rect 868 969 902 1003
rect 868 901 902 935
rect 868 833 902 867
rect 868 765 902 799
rect 868 697 902 731
rect 868 629 902 663
rect 868 561 902 595
rect 868 493 902 527
rect 868 425 902 459
rect 868 357 902 391
rect 868 289 902 323
rect 868 221 902 255
rect 868 153 902 187
rect 868 85 902 119
rect 868 17 902 51
rect 868 -51 902 -17
rect 868 -119 902 -85
rect 868 -187 902 -153
rect 868 -255 902 -221
rect 868 -323 902 -289
rect 868 -391 902 -357
rect 868 -459 902 -425
rect 868 -527 902 -493
rect 868 -595 902 -561
rect 868 -663 902 -629
rect 868 -731 902 -697
rect 868 -799 902 -765
rect 868 -867 902 -833
rect 868 -935 902 -901
rect 868 -1003 902 -969
rect 868 -1071 902 -1037
rect 868 -1139 902 -1105
rect 868 -1207 902 -1173
rect 868 -1275 902 -1241
rect 868 -1343 902 -1309
rect 868 -1411 902 -1377
rect 868 -1479 902 -1445
rect 868 -1547 902 -1513
rect 868 -1615 902 -1581
rect 868 -1683 902 -1649
rect 868 -1751 902 -1717
rect 868 -1819 902 -1785
rect 868 -1887 902 -1853
rect 868 -1955 902 -1921
rect 868 -2023 902 -1989
rect 868 -2091 902 -2057
rect 868 -2159 902 -2125
rect 868 -2227 902 -2193
rect 868 -2295 902 -2261
rect 868 -2363 902 -2329
rect 868 -2431 902 -2397
rect 868 -2499 902 -2465
rect 868 -2567 902 -2533
rect 868 -2635 902 -2601
rect 868 -2703 902 -2669
rect 868 -2771 902 -2737
rect 868 -2839 902 -2805
rect 868 -2907 902 -2873
rect 868 -2975 902 -2941
rect 868 -3043 902 -3009
rect 868 -3111 902 -3077
rect 868 -3179 902 -3145
rect 868 -3247 902 -3213
rect 868 -3315 902 -3281
rect 868 -3383 902 -3349
rect 868 -3451 902 -3417
rect 868 -3519 902 -3485
rect 868 -3587 902 -3553
rect 868 -3655 902 -3621
rect 868 -3723 902 -3689
rect 868 -3791 902 -3757
rect 868 -3859 902 -3825
rect 868 -3927 902 -3893
rect 868 -3995 902 -3961
rect 868 -4063 902 -4029
rect 868 -4131 902 -4097
rect 868 -4199 902 -4165
rect 868 -4267 902 -4233
rect 868 -4335 902 -4301
rect 868 -4403 902 -4369
rect 868 -4471 902 -4437
rect 868 -4539 902 -4505
rect 868 -4607 902 -4573
rect 868 -4675 902 -4641
rect 868 -4743 902 -4709
rect 868 -4811 902 -4777
rect 868 -4879 902 -4845
rect 868 -4947 902 -4913
rect 868 -5015 902 -4981
rect 868 -5083 902 -5049
rect 868 -5151 902 -5117
rect 868 -5219 902 -5185
rect 868 -5287 902 -5253
rect 868 -5355 902 -5321
rect 868 -5423 902 -5389
rect 868 -5491 902 -5457
rect 868 -5559 902 -5525
rect 868 -5627 902 -5593
rect 868 -5695 902 -5661
rect 868 -5763 902 -5729
rect 868 -5831 902 -5797
rect 868 -5899 902 -5865
rect 868 -5967 902 -5933
rect 868 -6035 902 -6001
rect 868 -6103 902 -6069
rect 868 -6171 902 -6137
rect 868 -6239 902 -6205
rect 868 -6307 902 -6273
rect 868 -6375 902 -6341
rect 868 -6443 902 -6409
rect 868 -6511 902 -6477
rect 868 -6579 902 -6545
rect 868 -6647 902 -6613
rect 868 -6715 902 -6681
rect 868 -6783 902 -6749
rect 868 -6851 902 -6817
rect 868 -6919 902 -6885
rect 868 -6987 902 -6953
rect 868 -7055 902 -7021
rect 868 -7123 902 -7089
rect 868 -7191 902 -7157
rect 868 -7259 902 -7225
rect 868 -7327 902 -7293
rect 868 -7395 902 -7361
rect 868 -7463 902 -7429
rect 868 -7531 902 -7497
rect 868 -7599 902 -7565
rect 868 -7667 902 -7633
rect 868 -7735 902 -7701
rect 868 -7803 902 -7769
rect 868 -7871 902 -7837
rect 868 -7939 902 -7905
rect 868 -8007 902 -7973
rect 868 -8075 902 -8041
rect 868 -8143 902 -8109
rect 868 -8211 902 -8177
rect 868 -8279 902 -8245
rect 868 -8347 902 -8313
rect 868 -8415 902 -8381
rect 868 -8483 902 -8449
rect 868 -8551 902 -8517
rect 868 -8619 902 -8585
rect 868 -8687 902 -8653
rect 868 -8755 902 -8721
rect 868 -8823 902 -8789
rect 868 -8891 902 -8857
rect 868 -8959 902 -8925
rect 868 -9027 902 -8993
rect 868 -9095 902 -9061
rect 868 -9163 902 -9129
rect 868 -9231 902 -9197
rect 868 -9299 902 -9265
rect 868 -9367 902 -9333
rect 868 -9435 902 -9401
rect 868 -9503 902 -9469
rect 868 -9571 902 -9537
rect 986 9537 1020 9571
rect 986 9469 1020 9503
rect 986 9401 1020 9435
rect 986 9333 1020 9367
rect 986 9265 1020 9299
rect 986 9197 1020 9231
rect 986 9129 1020 9163
rect 986 9061 1020 9095
rect 986 8993 1020 9027
rect 986 8925 1020 8959
rect 986 8857 1020 8891
rect 986 8789 1020 8823
rect 986 8721 1020 8755
rect 986 8653 1020 8687
rect 986 8585 1020 8619
rect 986 8517 1020 8551
rect 986 8449 1020 8483
rect 986 8381 1020 8415
rect 986 8313 1020 8347
rect 986 8245 1020 8279
rect 986 8177 1020 8211
rect 986 8109 1020 8143
rect 986 8041 1020 8075
rect 986 7973 1020 8007
rect 986 7905 1020 7939
rect 986 7837 1020 7871
rect 986 7769 1020 7803
rect 986 7701 1020 7735
rect 986 7633 1020 7667
rect 986 7565 1020 7599
rect 986 7497 1020 7531
rect 986 7429 1020 7463
rect 986 7361 1020 7395
rect 986 7293 1020 7327
rect 986 7225 1020 7259
rect 986 7157 1020 7191
rect 986 7089 1020 7123
rect 986 7021 1020 7055
rect 986 6953 1020 6987
rect 986 6885 1020 6919
rect 986 6817 1020 6851
rect 986 6749 1020 6783
rect 986 6681 1020 6715
rect 986 6613 1020 6647
rect 986 6545 1020 6579
rect 986 6477 1020 6511
rect 986 6409 1020 6443
rect 986 6341 1020 6375
rect 986 6273 1020 6307
rect 986 6205 1020 6239
rect 986 6137 1020 6171
rect 986 6069 1020 6103
rect 986 6001 1020 6035
rect 986 5933 1020 5967
rect 986 5865 1020 5899
rect 986 5797 1020 5831
rect 986 5729 1020 5763
rect 986 5661 1020 5695
rect 986 5593 1020 5627
rect 986 5525 1020 5559
rect 986 5457 1020 5491
rect 986 5389 1020 5423
rect 986 5321 1020 5355
rect 986 5253 1020 5287
rect 986 5185 1020 5219
rect 986 5117 1020 5151
rect 986 5049 1020 5083
rect 986 4981 1020 5015
rect 986 4913 1020 4947
rect 986 4845 1020 4879
rect 986 4777 1020 4811
rect 986 4709 1020 4743
rect 986 4641 1020 4675
rect 986 4573 1020 4607
rect 986 4505 1020 4539
rect 986 4437 1020 4471
rect 986 4369 1020 4403
rect 986 4301 1020 4335
rect 986 4233 1020 4267
rect 986 4165 1020 4199
rect 986 4097 1020 4131
rect 986 4029 1020 4063
rect 986 3961 1020 3995
rect 986 3893 1020 3927
rect 986 3825 1020 3859
rect 986 3757 1020 3791
rect 986 3689 1020 3723
rect 986 3621 1020 3655
rect 986 3553 1020 3587
rect 986 3485 1020 3519
rect 986 3417 1020 3451
rect 986 3349 1020 3383
rect 986 3281 1020 3315
rect 986 3213 1020 3247
rect 986 3145 1020 3179
rect 986 3077 1020 3111
rect 986 3009 1020 3043
rect 986 2941 1020 2975
rect 986 2873 1020 2907
rect 986 2805 1020 2839
rect 986 2737 1020 2771
rect 986 2669 1020 2703
rect 986 2601 1020 2635
rect 986 2533 1020 2567
rect 986 2465 1020 2499
rect 986 2397 1020 2431
rect 986 2329 1020 2363
rect 986 2261 1020 2295
rect 986 2193 1020 2227
rect 986 2125 1020 2159
rect 986 2057 1020 2091
rect 986 1989 1020 2023
rect 986 1921 1020 1955
rect 986 1853 1020 1887
rect 986 1785 1020 1819
rect 986 1717 1020 1751
rect 986 1649 1020 1683
rect 986 1581 1020 1615
rect 986 1513 1020 1547
rect 986 1445 1020 1479
rect 986 1377 1020 1411
rect 986 1309 1020 1343
rect 986 1241 1020 1275
rect 986 1173 1020 1207
rect 986 1105 1020 1139
rect 986 1037 1020 1071
rect 986 969 1020 1003
rect 986 901 1020 935
rect 986 833 1020 867
rect 986 765 1020 799
rect 986 697 1020 731
rect 986 629 1020 663
rect 986 561 1020 595
rect 986 493 1020 527
rect 986 425 1020 459
rect 986 357 1020 391
rect 986 289 1020 323
rect 986 221 1020 255
rect 986 153 1020 187
rect 986 85 1020 119
rect 986 17 1020 51
rect 986 -51 1020 -17
rect 986 -119 1020 -85
rect 986 -187 1020 -153
rect 986 -255 1020 -221
rect 986 -323 1020 -289
rect 986 -391 1020 -357
rect 986 -459 1020 -425
rect 986 -527 1020 -493
rect 986 -595 1020 -561
rect 986 -663 1020 -629
rect 986 -731 1020 -697
rect 986 -799 1020 -765
rect 986 -867 1020 -833
rect 986 -935 1020 -901
rect 986 -1003 1020 -969
rect 986 -1071 1020 -1037
rect 986 -1139 1020 -1105
rect 986 -1207 1020 -1173
rect 986 -1275 1020 -1241
rect 986 -1343 1020 -1309
rect 986 -1411 1020 -1377
rect 986 -1479 1020 -1445
rect 986 -1547 1020 -1513
rect 986 -1615 1020 -1581
rect 986 -1683 1020 -1649
rect 986 -1751 1020 -1717
rect 986 -1819 1020 -1785
rect 986 -1887 1020 -1853
rect 986 -1955 1020 -1921
rect 986 -2023 1020 -1989
rect 986 -2091 1020 -2057
rect 986 -2159 1020 -2125
rect 986 -2227 1020 -2193
rect 986 -2295 1020 -2261
rect 986 -2363 1020 -2329
rect 986 -2431 1020 -2397
rect 986 -2499 1020 -2465
rect 986 -2567 1020 -2533
rect 986 -2635 1020 -2601
rect 986 -2703 1020 -2669
rect 986 -2771 1020 -2737
rect 986 -2839 1020 -2805
rect 986 -2907 1020 -2873
rect 986 -2975 1020 -2941
rect 986 -3043 1020 -3009
rect 986 -3111 1020 -3077
rect 986 -3179 1020 -3145
rect 986 -3247 1020 -3213
rect 986 -3315 1020 -3281
rect 986 -3383 1020 -3349
rect 986 -3451 1020 -3417
rect 986 -3519 1020 -3485
rect 986 -3587 1020 -3553
rect 986 -3655 1020 -3621
rect 986 -3723 1020 -3689
rect 986 -3791 1020 -3757
rect 986 -3859 1020 -3825
rect 986 -3927 1020 -3893
rect 986 -3995 1020 -3961
rect 986 -4063 1020 -4029
rect 986 -4131 1020 -4097
rect 986 -4199 1020 -4165
rect 986 -4267 1020 -4233
rect 986 -4335 1020 -4301
rect 986 -4403 1020 -4369
rect 986 -4471 1020 -4437
rect 986 -4539 1020 -4505
rect 986 -4607 1020 -4573
rect 986 -4675 1020 -4641
rect 986 -4743 1020 -4709
rect 986 -4811 1020 -4777
rect 986 -4879 1020 -4845
rect 986 -4947 1020 -4913
rect 986 -5015 1020 -4981
rect 986 -5083 1020 -5049
rect 986 -5151 1020 -5117
rect 986 -5219 1020 -5185
rect 986 -5287 1020 -5253
rect 986 -5355 1020 -5321
rect 986 -5423 1020 -5389
rect 986 -5491 1020 -5457
rect 986 -5559 1020 -5525
rect 986 -5627 1020 -5593
rect 986 -5695 1020 -5661
rect 986 -5763 1020 -5729
rect 986 -5831 1020 -5797
rect 986 -5899 1020 -5865
rect 986 -5967 1020 -5933
rect 986 -6035 1020 -6001
rect 986 -6103 1020 -6069
rect 986 -6171 1020 -6137
rect 986 -6239 1020 -6205
rect 986 -6307 1020 -6273
rect 986 -6375 1020 -6341
rect 986 -6443 1020 -6409
rect 986 -6511 1020 -6477
rect 986 -6579 1020 -6545
rect 986 -6647 1020 -6613
rect 986 -6715 1020 -6681
rect 986 -6783 1020 -6749
rect 986 -6851 1020 -6817
rect 986 -6919 1020 -6885
rect 986 -6987 1020 -6953
rect 986 -7055 1020 -7021
rect 986 -7123 1020 -7089
rect 986 -7191 1020 -7157
rect 986 -7259 1020 -7225
rect 986 -7327 1020 -7293
rect 986 -7395 1020 -7361
rect 986 -7463 1020 -7429
rect 986 -7531 1020 -7497
rect 986 -7599 1020 -7565
rect 986 -7667 1020 -7633
rect 986 -7735 1020 -7701
rect 986 -7803 1020 -7769
rect 986 -7871 1020 -7837
rect 986 -7939 1020 -7905
rect 986 -8007 1020 -7973
rect 986 -8075 1020 -8041
rect 986 -8143 1020 -8109
rect 986 -8211 1020 -8177
rect 986 -8279 1020 -8245
rect 986 -8347 1020 -8313
rect 986 -8415 1020 -8381
rect 986 -8483 1020 -8449
rect 986 -8551 1020 -8517
rect 986 -8619 1020 -8585
rect 986 -8687 1020 -8653
rect 986 -8755 1020 -8721
rect 986 -8823 1020 -8789
rect 986 -8891 1020 -8857
rect 986 -8959 1020 -8925
rect 986 -9027 1020 -8993
rect 986 -9095 1020 -9061
rect 986 -9163 1020 -9129
rect 986 -9231 1020 -9197
rect 986 -9299 1020 -9265
rect 986 -9367 1020 -9333
rect 986 -9435 1020 -9401
rect 986 -9503 1020 -9469
rect 986 -9571 1020 -9537
rect 1104 9537 1138 9571
rect 1104 9469 1138 9503
rect 1104 9401 1138 9435
rect 1104 9333 1138 9367
rect 1104 9265 1138 9299
rect 1104 9197 1138 9231
rect 1104 9129 1138 9163
rect 1104 9061 1138 9095
rect 1104 8993 1138 9027
rect 1104 8925 1138 8959
rect 1104 8857 1138 8891
rect 1104 8789 1138 8823
rect 1104 8721 1138 8755
rect 1104 8653 1138 8687
rect 1104 8585 1138 8619
rect 1104 8517 1138 8551
rect 1104 8449 1138 8483
rect 1104 8381 1138 8415
rect 1104 8313 1138 8347
rect 1104 8245 1138 8279
rect 1104 8177 1138 8211
rect 1104 8109 1138 8143
rect 1104 8041 1138 8075
rect 1104 7973 1138 8007
rect 1104 7905 1138 7939
rect 1104 7837 1138 7871
rect 1104 7769 1138 7803
rect 1104 7701 1138 7735
rect 1104 7633 1138 7667
rect 1104 7565 1138 7599
rect 1104 7497 1138 7531
rect 1104 7429 1138 7463
rect 1104 7361 1138 7395
rect 1104 7293 1138 7327
rect 1104 7225 1138 7259
rect 1104 7157 1138 7191
rect 1104 7089 1138 7123
rect 1104 7021 1138 7055
rect 1104 6953 1138 6987
rect 1104 6885 1138 6919
rect 1104 6817 1138 6851
rect 1104 6749 1138 6783
rect 1104 6681 1138 6715
rect 1104 6613 1138 6647
rect 1104 6545 1138 6579
rect 1104 6477 1138 6511
rect 1104 6409 1138 6443
rect 1104 6341 1138 6375
rect 1104 6273 1138 6307
rect 1104 6205 1138 6239
rect 1104 6137 1138 6171
rect 1104 6069 1138 6103
rect 1104 6001 1138 6035
rect 1104 5933 1138 5967
rect 1104 5865 1138 5899
rect 1104 5797 1138 5831
rect 1104 5729 1138 5763
rect 1104 5661 1138 5695
rect 1104 5593 1138 5627
rect 1104 5525 1138 5559
rect 1104 5457 1138 5491
rect 1104 5389 1138 5423
rect 1104 5321 1138 5355
rect 1104 5253 1138 5287
rect 1104 5185 1138 5219
rect 1104 5117 1138 5151
rect 1104 5049 1138 5083
rect 1104 4981 1138 5015
rect 1104 4913 1138 4947
rect 1104 4845 1138 4879
rect 1104 4777 1138 4811
rect 1104 4709 1138 4743
rect 1104 4641 1138 4675
rect 1104 4573 1138 4607
rect 1104 4505 1138 4539
rect 1104 4437 1138 4471
rect 1104 4369 1138 4403
rect 1104 4301 1138 4335
rect 1104 4233 1138 4267
rect 1104 4165 1138 4199
rect 1104 4097 1138 4131
rect 1104 4029 1138 4063
rect 1104 3961 1138 3995
rect 1104 3893 1138 3927
rect 1104 3825 1138 3859
rect 1104 3757 1138 3791
rect 1104 3689 1138 3723
rect 1104 3621 1138 3655
rect 1104 3553 1138 3587
rect 1104 3485 1138 3519
rect 1104 3417 1138 3451
rect 1104 3349 1138 3383
rect 1104 3281 1138 3315
rect 1104 3213 1138 3247
rect 1104 3145 1138 3179
rect 1104 3077 1138 3111
rect 1104 3009 1138 3043
rect 1104 2941 1138 2975
rect 1104 2873 1138 2907
rect 1104 2805 1138 2839
rect 1104 2737 1138 2771
rect 1104 2669 1138 2703
rect 1104 2601 1138 2635
rect 1104 2533 1138 2567
rect 1104 2465 1138 2499
rect 1104 2397 1138 2431
rect 1104 2329 1138 2363
rect 1104 2261 1138 2295
rect 1104 2193 1138 2227
rect 1104 2125 1138 2159
rect 1104 2057 1138 2091
rect 1104 1989 1138 2023
rect 1104 1921 1138 1955
rect 1104 1853 1138 1887
rect 1104 1785 1138 1819
rect 1104 1717 1138 1751
rect 1104 1649 1138 1683
rect 1104 1581 1138 1615
rect 1104 1513 1138 1547
rect 1104 1445 1138 1479
rect 1104 1377 1138 1411
rect 1104 1309 1138 1343
rect 1104 1241 1138 1275
rect 1104 1173 1138 1207
rect 1104 1105 1138 1139
rect 1104 1037 1138 1071
rect 1104 969 1138 1003
rect 1104 901 1138 935
rect 1104 833 1138 867
rect 1104 765 1138 799
rect 1104 697 1138 731
rect 1104 629 1138 663
rect 1104 561 1138 595
rect 1104 493 1138 527
rect 1104 425 1138 459
rect 1104 357 1138 391
rect 1104 289 1138 323
rect 1104 221 1138 255
rect 1104 153 1138 187
rect 1104 85 1138 119
rect 1104 17 1138 51
rect 1104 -51 1138 -17
rect 1104 -119 1138 -85
rect 1104 -187 1138 -153
rect 1104 -255 1138 -221
rect 1104 -323 1138 -289
rect 1104 -391 1138 -357
rect 1104 -459 1138 -425
rect 1104 -527 1138 -493
rect 1104 -595 1138 -561
rect 1104 -663 1138 -629
rect 1104 -731 1138 -697
rect 1104 -799 1138 -765
rect 1104 -867 1138 -833
rect 1104 -935 1138 -901
rect 1104 -1003 1138 -969
rect 1104 -1071 1138 -1037
rect 1104 -1139 1138 -1105
rect 1104 -1207 1138 -1173
rect 1104 -1275 1138 -1241
rect 1104 -1343 1138 -1309
rect 1104 -1411 1138 -1377
rect 1104 -1479 1138 -1445
rect 1104 -1547 1138 -1513
rect 1104 -1615 1138 -1581
rect 1104 -1683 1138 -1649
rect 1104 -1751 1138 -1717
rect 1104 -1819 1138 -1785
rect 1104 -1887 1138 -1853
rect 1104 -1955 1138 -1921
rect 1104 -2023 1138 -1989
rect 1104 -2091 1138 -2057
rect 1104 -2159 1138 -2125
rect 1104 -2227 1138 -2193
rect 1104 -2295 1138 -2261
rect 1104 -2363 1138 -2329
rect 1104 -2431 1138 -2397
rect 1104 -2499 1138 -2465
rect 1104 -2567 1138 -2533
rect 1104 -2635 1138 -2601
rect 1104 -2703 1138 -2669
rect 1104 -2771 1138 -2737
rect 1104 -2839 1138 -2805
rect 1104 -2907 1138 -2873
rect 1104 -2975 1138 -2941
rect 1104 -3043 1138 -3009
rect 1104 -3111 1138 -3077
rect 1104 -3179 1138 -3145
rect 1104 -3247 1138 -3213
rect 1104 -3315 1138 -3281
rect 1104 -3383 1138 -3349
rect 1104 -3451 1138 -3417
rect 1104 -3519 1138 -3485
rect 1104 -3587 1138 -3553
rect 1104 -3655 1138 -3621
rect 1104 -3723 1138 -3689
rect 1104 -3791 1138 -3757
rect 1104 -3859 1138 -3825
rect 1104 -3927 1138 -3893
rect 1104 -3995 1138 -3961
rect 1104 -4063 1138 -4029
rect 1104 -4131 1138 -4097
rect 1104 -4199 1138 -4165
rect 1104 -4267 1138 -4233
rect 1104 -4335 1138 -4301
rect 1104 -4403 1138 -4369
rect 1104 -4471 1138 -4437
rect 1104 -4539 1138 -4505
rect 1104 -4607 1138 -4573
rect 1104 -4675 1138 -4641
rect 1104 -4743 1138 -4709
rect 1104 -4811 1138 -4777
rect 1104 -4879 1138 -4845
rect 1104 -4947 1138 -4913
rect 1104 -5015 1138 -4981
rect 1104 -5083 1138 -5049
rect 1104 -5151 1138 -5117
rect 1104 -5219 1138 -5185
rect 1104 -5287 1138 -5253
rect 1104 -5355 1138 -5321
rect 1104 -5423 1138 -5389
rect 1104 -5491 1138 -5457
rect 1104 -5559 1138 -5525
rect 1104 -5627 1138 -5593
rect 1104 -5695 1138 -5661
rect 1104 -5763 1138 -5729
rect 1104 -5831 1138 -5797
rect 1104 -5899 1138 -5865
rect 1104 -5967 1138 -5933
rect 1104 -6035 1138 -6001
rect 1104 -6103 1138 -6069
rect 1104 -6171 1138 -6137
rect 1104 -6239 1138 -6205
rect 1104 -6307 1138 -6273
rect 1104 -6375 1138 -6341
rect 1104 -6443 1138 -6409
rect 1104 -6511 1138 -6477
rect 1104 -6579 1138 -6545
rect 1104 -6647 1138 -6613
rect 1104 -6715 1138 -6681
rect 1104 -6783 1138 -6749
rect 1104 -6851 1138 -6817
rect 1104 -6919 1138 -6885
rect 1104 -6987 1138 -6953
rect 1104 -7055 1138 -7021
rect 1104 -7123 1138 -7089
rect 1104 -7191 1138 -7157
rect 1104 -7259 1138 -7225
rect 1104 -7327 1138 -7293
rect 1104 -7395 1138 -7361
rect 1104 -7463 1138 -7429
rect 1104 -7531 1138 -7497
rect 1104 -7599 1138 -7565
rect 1104 -7667 1138 -7633
rect 1104 -7735 1138 -7701
rect 1104 -7803 1138 -7769
rect 1104 -7871 1138 -7837
rect 1104 -7939 1138 -7905
rect 1104 -8007 1138 -7973
rect 1104 -8075 1138 -8041
rect 1104 -8143 1138 -8109
rect 1104 -8211 1138 -8177
rect 1104 -8279 1138 -8245
rect 1104 -8347 1138 -8313
rect 1104 -8415 1138 -8381
rect 1104 -8483 1138 -8449
rect 1104 -8551 1138 -8517
rect 1104 -8619 1138 -8585
rect 1104 -8687 1138 -8653
rect 1104 -8755 1138 -8721
rect 1104 -8823 1138 -8789
rect 1104 -8891 1138 -8857
rect 1104 -8959 1138 -8925
rect 1104 -9027 1138 -8993
rect 1104 -9095 1138 -9061
rect 1104 -9163 1138 -9129
rect 1104 -9231 1138 -9197
rect 1104 -9299 1138 -9265
rect 1104 -9367 1138 -9333
rect 1104 -9435 1138 -9401
rect 1104 -9503 1138 -9469
rect 1104 -9571 1138 -9537
rect 1222 9537 1256 9571
rect 1222 9469 1256 9503
rect 1222 9401 1256 9435
rect 1222 9333 1256 9367
rect 1222 9265 1256 9299
rect 1222 9197 1256 9231
rect 1222 9129 1256 9163
rect 1222 9061 1256 9095
rect 1222 8993 1256 9027
rect 1222 8925 1256 8959
rect 1222 8857 1256 8891
rect 1222 8789 1256 8823
rect 1222 8721 1256 8755
rect 1222 8653 1256 8687
rect 1222 8585 1256 8619
rect 1222 8517 1256 8551
rect 1222 8449 1256 8483
rect 1222 8381 1256 8415
rect 1222 8313 1256 8347
rect 1222 8245 1256 8279
rect 1222 8177 1256 8211
rect 1222 8109 1256 8143
rect 1222 8041 1256 8075
rect 1222 7973 1256 8007
rect 1222 7905 1256 7939
rect 1222 7837 1256 7871
rect 1222 7769 1256 7803
rect 1222 7701 1256 7735
rect 1222 7633 1256 7667
rect 1222 7565 1256 7599
rect 1222 7497 1256 7531
rect 1222 7429 1256 7463
rect 1222 7361 1256 7395
rect 1222 7293 1256 7327
rect 1222 7225 1256 7259
rect 1222 7157 1256 7191
rect 1222 7089 1256 7123
rect 1222 7021 1256 7055
rect 1222 6953 1256 6987
rect 1222 6885 1256 6919
rect 1222 6817 1256 6851
rect 1222 6749 1256 6783
rect 1222 6681 1256 6715
rect 1222 6613 1256 6647
rect 1222 6545 1256 6579
rect 1222 6477 1256 6511
rect 1222 6409 1256 6443
rect 1222 6341 1256 6375
rect 1222 6273 1256 6307
rect 1222 6205 1256 6239
rect 1222 6137 1256 6171
rect 1222 6069 1256 6103
rect 1222 6001 1256 6035
rect 1222 5933 1256 5967
rect 1222 5865 1256 5899
rect 1222 5797 1256 5831
rect 1222 5729 1256 5763
rect 1222 5661 1256 5695
rect 1222 5593 1256 5627
rect 1222 5525 1256 5559
rect 1222 5457 1256 5491
rect 1222 5389 1256 5423
rect 1222 5321 1256 5355
rect 1222 5253 1256 5287
rect 1222 5185 1256 5219
rect 1222 5117 1256 5151
rect 1222 5049 1256 5083
rect 1222 4981 1256 5015
rect 1222 4913 1256 4947
rect 1222 4845 1256 4879
rect 1222 4777 1256 4811
rect 1222 4709 1256 4743
rect 1222 4641 1256 4675
rect 1222 4573 1256 4607
rect 1222 4505 1256 4539
rect 1222 4437 1256 4471
rect 1222 4369 1256 4403
rect 1222 4301 1256 4335
rect 1222 4233 1256 4267
rect 1222 4165 1256 4199
rect 1222 4097 1256 4131
rect 1222 4029 1256 4063
rect 1222 3961 1256 3995
rect 1222 3893 1256 3927
rect 1222 3825 1256 3859
rect 1222 3757 1256 3791
rect 1222 3689 1256 3723
rect 1222 3621 1256 3655
rect 1222 3553 1256 3587
rect 1222 3485 1256 3519
rect 1222 3417 1256 3451
rect 1222 3349 1256 3383
rect 1222 3281 1256 3315
rect 1222 3213 1256 3247
rect 1222 3145 1256 3179
rect 1222 3077 1256 3111
rect 1222 3009 1256 3043
rect 1222 2941 1256 2975
rect 1222 2873 1256 2907
rect 1222 2805 1256 2839
rect 1222 2737 1256 2771
rect 1222 2669 1256 2703
rect 1222 2601 1256 2635
rect 1222 2533 1256 2567
rect 1222 2465 1256 2499
rect 1222 2397 1256 2431
rect 1222 2329 1256 2363
rect 1222 2261 1256 2295
rect 1222 2193 1256 2227
rect 1222 2125 1256 2159
rect 1222 2057 1256 2091
rect 1222 1989 1256 2023
rect 1222 1921 1256 1955
rect 1222 1853 1256 1887
rect 1222 1785 1256 1819
rect 1222 1717 1256 1751
rect 1222 1649 1256 1683
rect 1222 1581 1256 1615
rect 1222 1513 1256 1547
rect 1222 1445 1256 1479
rect 1222 1377 1256 1411
rect 1222 1309 1256 1343
rect 1222 1241 1256 1275
rect 1222 1173 1256 1207
rect 1222 1105 1256 1139
rect 1222 1037 1256 1071
rect 1222 969 1256 1003
rect 1222 901 1256 935
rect 1222 833 1256 867
rect 1222 765 1256 799
rect 1222 697 1256 731
rect 1222 629 1256 663
rect 1222 561 1256 595
rect 1222 493 1256 527
rect 1222 425 1256 459
rect 1222 357 1256 391
rect 1222 289 1256 323
rect 1222 221 1256 255
rect 1222 153 1256 187
rect 1222 85 1256 119
rect 1222 17 1256 51
rect 1222 -51 1256 -17
rect 1222 -119 1256 -85
rect 1222 -187 1256 -153
rect 1222 -255 1256 -221
rect 1222 -323 1256 -289
rect 1222 -391 1256 -357
rect 1222 -459 1256 -425
rect 1222 -527 1256 -493
rect 1222 -595 1256 -561
rect 1222 -663 1256 -629
rect 1222 -731 1256 -697
rect 1222 -799 1256 -765
rect 1222 -867 1256 -833
rect 1222 -935 1256 -901
rect 1222 -1003 1256 -969
rect 1222 -1071 1256 -1037
rect 1222 -1139 1256 -1105
rect 1222 -1207 1256 -1173
rect 1222 -1275 1256 -1241
rect 1222 -1343 1256 -1309
rect 1222 -1411 1256 -1377
rect 1222 -1479 1256 -1445
rect 1222 -1547 1256 -1513
rect 1222 -1615 1256 -1581
rect 1222 -1683 1256 -1649
rect 1222 -1751 1256 -1717
rect 1222 -1819 1256 -1785
rect 1222 -1887 1256 -1853
rect 1222 -1955 1256 -1921
rect 1222 -2023 1256 -1989
rect 1222 -2091 1256 -2057
rect 1222 -2159 1256 -2125
rect 1222 -2227 1256 -2193
rect 1222 -2295 1256 -2261
rect 1222 -2363 1256 -2329
rect 1222 -2431 1256 -2397
rect 1222 -2499 1256 -2465
rect 1222 -2567 1256 -2533
rect 1222 -2635 1256 -2601
rect 1222 -2703 1256 -2669
rect 1222 -2771 1256 -2737
rect 1222 -2839 1256 -2805
rect 1222 -2907 1256 -2873
rect 1222 -2975 1256 -2941
rect 1222 -3043 1256 -3009
rect 1222 -3111 1256 -3077
rect 1222 -3179 1256 -3145
rect 1222 -3247 1256 -3213
rect 1222 -3315 1256 -3281
rect 1222 -3383 1256 -3349
rect 1222 -3451 1256 -3417
rect 1222 -3519 1256 -3485
rect 1222 -3587 1256 -3553
rect 1222 -3655 1256 -3621
rect 1222 -3723 1256 -3689
rect 1222 -3791 1256 -3757
rect 1222 -3859 1256 -3825
rect 1222 -3927 1256 -3893
rect 1222 -3995 1256 -3961
rect 1222 -4063 1256 -4029
rect 1222 -4131 1256 -4097
rect 1222 -4199 1256 -4165
rect 1222 -4267 1256 -4233
rect 1222 -4335 1256 -4301
rect 1222 -4403 1256 -4369
rect 1222 -4471 1256 -4437
rect 1222 -4539 1256 -4505
rect 1222 -4607 1256 -4573
rect 1222 -4675 1256 -4641
rect 1222 -4743 1256 -4709
rect 1222 -4811 1256 -4777
rect 1222 -4879 1256 -4845
rect 1222 -4947 1256 -4913
rect 1222 -5015 1256 -4981
rect 1222 -5083 1256 -5049
rect 1222 -5151 1256 -5117
rect 1222 -5219 1256 -5185
rect 1222 -5287 1256 -5253
rect 1222 -5355 1256 -5321
rect 1222 -5423 1256 -5389
rect 1222 -5491 1256 -5457
rect 1222 -5559 1256 -5525
rect 1222 -5627 1256 -5593
rect 1222 -5695 1256 -5661
rect 1222 -5763 1256 -5729
rect 1222 -5831 1256 -5797
rect 1222 -5899 1256 -5865
rect 1222 -5967 1256 -5933
rect 1222 -6035 1256 -6001
rect 1222 -6103 1256 -6069
rect 1222 -6171 1256 -6137
rect 1222 -6239 1256 -6205
rect 1222 -6307 1256 -6273
rect 1222 -6375 1256 -6341
rect 1222 -6443 1256 -6409
rect 1222 -6511 1256 -6477
rect 1222 -6579 1256 -6545
rect 1222 -6647 1256 -6613
rect 1222 -6715 1256 -6681
rect 1222 -6783 1256 -6749
rect 1222 -6851 1256 -6817
rect 1222 -6919 1256 -6885
rect 1222 -6987 1256 -6953
rect 1222 -7055 1256 -7021
rect 1222 -7123 1256 -7089
rect 1222 -7191 1256 -7157
rect 1222 -7259 1256 -7225
rect 1222 -7327 1256 -7293
rect 1222 -7395 1256 -7361
rect 1222 -7463 1256 -7429
rect 1222 -7531 1256 -7497
rect 1222 -7599 1256 -7565
rect 1222 -7667 1256 -7633
rect 1222 -7735 1256 -7701
rect 1222 -7803 1256 -7769
rect 1222 -7871 1256 -7837
rect 1222 -7939 1256 -7905
rect 1222 -8007 1256 -7973
rect 1222 -8075 1256 -8041
rect 1222 -8143 1256 -8109
rect 1222 -8211 1256 -8177
rect 1222 -8279 1256 -8245
rect 1222 -8347 1256 -8313
rect 1222 -8415 1256 -8381
rect 1222 -8483 1256 -8449
rect 1222 -8551 1256 -8517
rect 1222 -8619 1256 -8585
rect 1222 -8687 1256 -8653
rect 1222 -8755 1256 -8721
rect 1222 -8823 1256 -8789
rect 1222 -8891 1256 -8857
rect 1222 -8959 1256 -8925
rect 1222 -9027 1256 -8993
rect 1222 -9095 1256 -9061
rect 1222 -9163 1256 -9129
rect 1222 -9231 1256 -9197
rect 1222 -9299 1256 -9265
rect 1222 -9367 1256 -9333
rect 1222 -9435 1256 -9401
rect 1222 -9503 1256 -9469
rect 1222 -9571 1256 -9537
rect 1340 9537 1374 9571
rect 1340 9469 1374 9503
rect 1340 9401 1374 9435
rect 1340 9333 1374 9367
rect 1340 9265 1374 9299
rect 1340 9197 1374 9231
rect 1340 9129 1374 9163
rect 1340 9061 1374 9095
rect 1340 8993 1374 9027
rect 1340 8925 1374 8959
rect 1340 8857 1374 8891
rect 1340 8789 1374 8823
rect 1340 8721 1374 8755
rect 1340 8653 1374 8687
rect 1340 8585 1374 8619
rect 1340 8517 1374 8551
rect 1340 8449 1374 8483
rect 1340 8381 1374 8415
rect 1340 8313 1374 8347
rect 1340 8245 1374 8279
rect 1340 8177 1374 8211
rect 1340 8109 1374 8143
rect 1340 8041 1374 8075
rect 1340 7973 1374 8007
rect 1340 7905 1374 7939
rect 1340 7837 1374 7871
rect 1340 7769 1374 7803
rect 1340 7701 1374 7735
rect 1340 7633 1374 7667
rect 1340 7565 1374 7599
rect 1340 7497 1374 7531
rect 1340 7429 1374 7463
rect 1340 7361 1374 7395
rect 1340 7293 1374 7327
rect 1340 7225 1374 7259
rect 1340 7157 1374 7191
rect 1340 7089 1374 7123
rect 1340 7021 1374 7055
rect 1340 6953 1374 6987
rect 1340 6885 1374 6919
rect 1340 6817 1374 6851
rect 1340 6749 1374 6783
rect 1340 6681 1374 6715
rect 1340 6613 1374 6647
rect 1340 6545 1374 6579
rect 1340 6477 1374 6511
rect 1340 6409 1374 6443
rect 1340 6341 1374 6375
rect 1340 6273 1374 6307
rect 1340 6205 1374 6239
rect 1340 6137 1374 6171
rect 1340 6069 1374 6103
rect 1340 6001 1374 6035
rect 1340 5933 1374 5967
rect 1340 5865 1374 5899
rect 1340 5797 1374 5831
rect 1340 5729 1374 5763
rect 1340 5661 1374 5695
rect 1340 5593 1374 5627
rect 1340 5525 1374 5559
rect 1340 5457 1374 5491
rect 1340 5389 1374 5423
rect 1340 5321 1374 5355
rect 1340 5253 1374 5287
rect 1340 5185 1374 5219
rect 1340 5117 1374 5151
rect 1340 5049 1374 5083
rect 1340 4981 1374 5015
rect 1340 4913 1374 4947
rect 1340 4845 1374 4879
rect 1340 4777 1374 4811
rect 1340 4709 1374 4743
rect 1340 4641 1374 4675
rect 1340 4573 1374 4607
rect 1340 4505 1374 4539
rect 1340 4437 1374 4471
rect 1340 4369 1374 4403
rect 1340 4301 1374 4335
rect 1340 4233 1374 4267
rect 1340 4165 1374 4199
rect 1340 4097 1374 4131
rect 1340 4029 1374 4063
rect 1340 3961 1374 3995
rect 1340 3893 1374 3927
rect 1340 3825 1374 3859
rect 1340 3757 1374 3791
rect 1340 3689 1374 3723
rect 1340 3621 1374 3655
rect 1340 3553 1374 3587
rect 1340 3485 1374 3519
rect 1340 3417 1374 3451
rect 1340 3349 1374 3383
rect 1340 3281 1374 3315
rect 1340 3213 1374 3247
rect 1340 3145 1374 3179
rect 1340 3077 1374 3111
rect 1340 3009 1374 3043
rect 1340 2941 1374 2975
rect 1340 2873 1374 2907
rect 1340 2805 1374 2839
rect 1340 2737 1374 2771
rect 1340 2669 1374 2703
rect 1340 2601 1374 2635
rect 1340 2533 1374 2567
rect 1340 2465 1374 2499
rect 1340 2397 1374 2431
rect 1340 2329 1374 2363
rect 1340 2261 1374 2295
rect 1340 2193 1374 2227
rect 1340 2125 1374 2159
rect 1340 2057 1374 2091
rect 1340 1989 1374 2023
rect 1340 1921 1374 1955
rect 1340 1853 1374 1887
rect 1340 1785 1374 1819
rect 1340 1717 1374 1751
rect 1340 1649 1374 1683
rect 1340 1581 1374 1615
rect 1340 1513 1374 1547
rect 1340 1445 1374 1479
rect 1340 1377 1374 1411
rect 1340 1309 1374 1343
rect 1340 1241 1374 1275
rect 1340 1173 1374 1207
rect 1340 1105 1374 1139
rect 1340 1037 1374 1071
rect 1340 969 1374 1003
rect 1340 901 1374 935
rect 1340 833 1374 867
rect 1340 765 1374 799
rect 1340 697 1374 731
rect 1340 629 1374 663
rect 1340 561 1374 595
rect 1340 493 1374 527
rect 1340 425 1374 459
rect 1340 357 1374 391
rect 1340 289 1374 323
rect 1340 221 1374 255
rect 1340 153 1374 187
rect 1340 85 1374 119
rect 1340 17 1374 51
rect 1340 -51 1374 -17
rect 1340 -119 1374 -85
rect 1340 -187 1374 -153
rect 1340 -255 1374 -221
rect 1340 -323 1374 -289
rect 1340 -391 1374 -357
rect 1340 -459 1374 -425
rect 1340 -527 1374 -493
rect 1340 -595 1374 -561
rect 1340 -663 1374 -629
rect 1340 -731 1374 -697
rect 1340 -799 1374 -765
rect 1340 -867 1374 -833
rect 1340 -935 1374 -901
rect 1340 -1003 1374 -969
rect 1340 -1071 1374 -1037
rect 1340 -1139 1374 -1105
rect 1340 -1207 1374 -1173
rect 1340 -1275 1374 -1241
rect 1340 -1343 1374 -1309
rect 1340 -1411 1374 -1377
rect 1340 -1479 1374 -1445
rect 1340 -1547 1374 -1513
rect 1340 -1615 1374 -1581
rect 1340 -1683 1374 -1649
rect 1340 -1751 1374 -1717
rect 1340 -1819 1374 -1785
rect 1340 -1887 1374 -1853
rect 1340 -1955 1374 -1921
rect 1340 -2023 1374 -1989
rect 1340 -2091 1374 -2057
rect 1340 -2159 1374 -2125
rect 1340 -2227 1374 -2193
rect 1340 -2295 1374 -2261
rect 1340 -2363 1374 -2329
rect 1340 -2431 1374 -2397
rect 1340 -2499 1374 -2465
rect 1340 -2567 1374 -2533
rect 1340 -2635 1374 -2601
rect 1340 -2703 1374 -2669
rect 1340 -2771 1374 -2737
rect 1340 -2839 1374 -2805
rect 1340 -2907 1374 -2873
rect 1340 -2975 1374 -2941
rect 1340 -3043 1374 -3009
rect 1340 -3111 1374 -3077
rect 1340 -3179 1374 -3145
rect 1340 -3247 1374 -3213
rect 1340 -3315 1374 -3281
rect 1340 -3383 1374 -3349
rect 1340 -3451 1374 -3417
rect 1340 -3519 1374 -3485
rect 1340 -3587 1374 -3553
rect 1340 -3655 1374 -3621
rect 1340 -3723 1374 -3689
rect 1340 -3791 1374 -3757
rect 1340 -3859 1374 -3825
rect 1340 -3927 1374 -3893
rect 1340 -3995 1374 -3961
rect 1340 -4063 1374 -4029
rect 1340 -4131 1374 -4097
rect 1340 -4199 1374 -4165
rect 1340 -4267 1374 -4233
rect 1340 -4335 1374 -4301
rect 1340 -4403 1374 -4369
rect 1340 -4471 1374 -4437
rect 1340 -4539 1374 -4505
rect 1340 -4607 1374 -4573
rect 1340 -4675 1374 -4641
rect 1340 -4743 1374 -4709
rect 1340 -4811 1374 -4777
rect 1340 -4879 1374 -4845
rect 1340 -4947 1374 -4913
rect 1340 -5015 1374 -4981
rect 1340 -5083 1374 -5049
rect 1340 -5151 1374 -5117
rect 1340 -5219 1374 -5185
rect 1340 -5287 1374 -5253
rect 1340 -5355 1374 -5321
rect 1340 -5423 1374 -5389
rect 1340 -5491 1374 -5457
rect 1340 -5559 1374 -5525
rect 1340 -5627 1374 -5593
rect 1340 -5695 1374 -5661
rect 1340 -5763 1374 -5729
rect 1340 -5831 1374 -5797
rect 1340 -5899 1374 -5865
rect 1340 -5967 1374 -5933
rect 1340 -6035 1374 -6001
rect 1340 -6103 1374 -6069
rect 1340 -6171 1374 -6137
rect 1340 -6239 1374 -6205
rect 1340 -6307 1374 -6273
rect 1340 -6375 1374 -6341
rect 1340 -6443 1374 -6409
rect 1340 -6511 1374 -6477
rect 1340 -6579 1374 -6545
rect 1340 -6647 1374 -6613
rect 1340 -6715 1374 -6681
rect 1340 -6783 1374 -6749
rect 1340 -6851 1374 -6817
rect 1340 -6919 1374 -6885
rect 1340 -6987 1374 -6953
rect 1340 -7055 1374 -7021
rect 1340 -7123 1374 -7089
rect 1340 -7191 1374 -7157
rect 1340 -7259 1374 -7225
rect 1340 -7327 1374 -7293
rect 1340 -7395 1374 -7361
rect 1340 -7463 1374 -7429
rect 1340 -7531 1374 -7497
rect 1340 -7599 1374 -7565
rect 1340 -7667 1374 -7633
rect 1340 -7735 1374 -7701
rect 1340 -7803 1374 -7769
rect 1340 -7871 1374 -7837
rect 1340 -7939 1374 -7905
rect 1340 -8007 1374 -7973
rect 1340 -8075 1374 -8041
rect 1340 -8143 1374 -8109
rect 1340 -8211 1374 -8177
rect 1340 -8279 1374 -8245
rect 1340 -8347 1374 -8313
rect 1340 -8415 1374 -8381
rect 1340 -8483 1374 -8449
rect 1340 -8551 1374 -8517
rect 1340 -8619 1374 -8585
rect 1340 -8687 1374 -8653
rect 1340 -8755 1374 -8721
rect 1340 -8823 1374 -8789
rect 1340 -8891 1374 -8857
rect 1340 -8959 1374 -8925
rect 1340 -9027 1374 -8993
rect 1340 -9095 1374 -9061
rect 1340 -9163 1374 -9129
rect 1340 -9231 1374 -9197
rect 1340 -9299 1374 -9265
rect 1340 -9367 1374 -9333
rect 1340 -9435 1374 -9401
rect 1340 -9503 1374 -9469
rect 1340 -9571 1374 -9537
rect 1458 9537 1492 9571
rect 1458 9469 1492 9503
rect 1458 9401 1492 9435
rect 1458 9333 1492 9367
rect 1458 9265 1492 9299
rect 1458 9197 1492 9231
rect 1458 9129 1492 9163
rect 1458 9061 1492 9095
rect 1458 8993 1492 9027
rect 1458 8925 1492 8959
rect 1458 8857 1492 8891
rect 1458 8789 1492 8823
rect 1458 8721 1492 8755
rect 1458 8653 1492 8687
rect 1458 8585 1492 8619
rect 1458 8517 1492 8551
rect 1458 8449 1492 8483
rect 1458 8381 1492 8415
rect 1458 8313 1492 8347
rect 1458 8245 1492 8279
rect 1458 8177 1492 8211
rect 1458 8109 1492 8143
rect 1458 8041 1492 8075
rect 1458 7973 1492 8007
rect 1458 7905 1492 7939
rect 1458 7837 1492 7871
rect 1458 7769 1492 7803
rect 1458 7701 1492 7735
rect 1458 7633 1492 7667
rect 1458 7565 1492 7599
rect 1458 7497 1492 7531
rect 1458 7429 1492 7463
rect 1458 7361 1492 7395
rect 1458 7293 1492 7327
rect 1458 7225 1492 7259
rect 1458 7157 1492 7191
rect 1458 7089 1492 7123
rect 1458 7021 1492 7055
rect 1458 6953 1492 6987
rect 1458 6885 1492 6919
rect 1458 6817 1492 6851
rect 1458 6749 1492 6783
rect 1458 6681 1492 6715
rect 1458 6613 1492 6647
rect 1458 6545 1492 6579
rect 1458 6477 1492 6511
rect 1458 6409 1492 6443
rect 1458 6341 1492 6375
rect 1458 6273 1492 6307
rect 1458 6205 1492 6239
rect 1458 6137 1492 6171
rect 1458 6069 1492 6103
rect 1458 6001 1492 6035
rect 1458 5933 1492 5967
rect 1458 5865 1492 5899
rect 1458 5797 1492 5831
rect 1458 5729 1492 5763
rect 1458 5661 1492 5695
rect 1458 5593 1492 5627
rect 1458 5525 1492 5559
rect 1458 5457 1492 5491
rect 1458 5389 1492 5423
rect 1458 5321 1492 5355
rect 1458 5253 1492 5287
rect 1458 5185 1492 5219
rect 1458 5117 1492 5151
rect 1458 5049 1492 5083
rect 1458 4981 1492 5015
rect 1458 4913 1492 4947
rect 1458 4845 1492 4879
rect 1458 4777 1492 4811
rect 1458 4709 1492 4743
rect 1458 4641 1492 4675
rect 1458 4573 1492 4607
rect 1458 4505 1492 4539
rect 1458 4437 1492 4471
rect 1458 4369 1492 4403
rect 1458 4301 1492 4335
rect 1458 4233 1492 4267
rect 1458 4165 1492 4199
rect 1458 4097 1492 4131
rect 1458 4029 1492 4063
rect 1458 3961 1492 3995
rect 1458 3893 1492 3927
rect 1458 3825 1492 3859
rect 1458 3757 1492 3791
rect 1458 3689 1492 3723
rect 1458 3621 1492 3655
rect 1458 3553 1492 3587
rect 1458 3485 1492 3519
rect 1458 3417 1492 3451
rect 1458 3349 1492 3383
rect 1458 3281 1492 3315
rect 1458 3213 1492 3247
rect 1458 3145 1492 3179
rect 1458 3077 1492 3111
rect 1458 3009 1492 3043
rect 1458 2941 1492 2975
rect 1458 2873 1492 2907
rect 1458 2805 1492 2839
rect 1458 2737 1492 2771
rect 1458 2669 1492 2703
rect 1458 2601 1492 2635
rect 1458 2533 1492 2567
rect 1458 2465 1492 2499
rect 1458 2397 1492 2431
rect 1458 2329 1492 2363
rect 1458 2261 1492 2295
rect 1458 2193 1492 2227
rect 1458 2125 1492 2159
rect 1458 2057 1492 2091
rect 1458 1989 1492 2023
rect 1458 1921 1492 1955
rect 1458 1853 1492 1887
rect 1458 1785 1492 1819
rect 1458 1717 1492 1751
rect 1458 1649 1492 1683
rect 1458 1581 1492 1615
rect 1458 1513 1492 1547
rect 1458 1445 1492 1479
rect 1458 1377 1492 1411
rect 1458 1309 1492 1343
rect 1458 1241 1492 1275
rect 1458 1173 1492 1207
rect 1458 1105 1492 1139
rect 1458 1037 1492 1071
rect 1458 969 1492 1003
rect 1458 901 1492 935
rect 1458 833 1492 867
rect 1458 765 1492 799
rect 1458 697 1492 731
rect 1458 629 1492 663
rect 1458 561 1492 595
rect 1458 493 1492 527
rect 1458 425 1492 459
rect 1458 357 1492 391
rect 1458 289 1492 323
rect 1458 221 1492 255
rect 1458 153 1492 187
rect 1458 85 1492 119
rect 1458 17 1492 51
rect 1458 -51 1492 -17
rect 1458 -119 1492 -85
rect 1458 -187 1492 -153
rect 1458 -255 1492 -221
rect 1458 -323 1492 -289
rect 1458 -391 1492 -357
rect 1458 -459 1492 -425
rect 1458 -527 1492 -493
rect 1458 -595 1492 -561
rect 1458 -663 1492 -629
rect 1458 -731 1492 -697
rect 1458 -799 1492 -765
rect 1458 -867 1492 -833
rect 1458 -935 1492 -901
rect 1458 -1003 1492 -969
rect 1458 -1071 1492 -1037
rect 1458 -1139 1492 -1105
rect 1458 -1207 1492 -1173
rect 1458 -1275 1492 -1241
rect 1458 -1343 1492 -1309
rect 1458 -1411 1492 -1377
rect 1458 -1479 1492 -1445
rect 1458 -1547 1492 -1513
rect 1458 -1615 1492 -1581
rect 1458 -1683 1492 -1649
rect 1458 -1751 1492 -1717
rect 1458 -1819 1492 -1785
rect 1458 -1887 1492 -1853
rect 1458 -1955 1492 -1921
rect 1458 -2023 1492 -1989
rect 1458 -2091 1492 -2057
rect 1458 -2159 1492 -2125
rect 1458 -2227 1492 -2193
rect 1458 -2295 1492 -2261
rect 1458 -2363 1492 -2329
rect 1458 -2431 1492 -2397
rect 1458 -2499 1492 -2465
rect 1458 -2567 1492 -2533
rect 1458 -2635 1492 -2601
rect 1458 -2703 1492 -2669
rect 1458 -2771 1492 -2737
rect 1458 -2839 1492 -2805
rect 1458 -2907 1492 -2873
rect 1458 -2975 1492 -2941
rect 1458 -3043 1492 -3009
rect 1458 -3111 1492 -3077
rect 1458 -3179 1492 -3145
rect 1458 -3247 1492 -3213
rect 1458 -3315 1492 -3281
rect 1458 -3383 1492 -3349
rect 1458 -3451 1492 -3417
rect 1458 -3519 1492 -3485
rect 1458 -3587 1492 -3553
rect 1458 -3655 1492 -3621
rect 1458 -3723 1492 -3689
rect 1458 -3791 1492 -3757
rect 1458 -3859 1492 -3825
rect 1458 -3927 1492 -3893
rect 1458 -3995 1492 -3961
rect 1458 -4063 1492 -4029
rect 1458 -4131 1492 -4097
rect 1458 -4199 1492 -4165
rect 1458 -4267 1492 -4233
rect 1458 -4335 1492 -4301
rect 1458 -4403 1492 -4369
rect 1458 -4471 1492 -4437
rect 1458 -4539 1492 -4505
rect 1458 -4607 1492 -4573
rect 1458 -4675 1492 -4641
rect 1458 -4743 1492 -4709
rect 1458 -4811 1492 -4777
rect 1458 -4879 1492 -4845
rect 1458 -4947 1492 -4913
rect 1458 -5015 1492 -4981
rect 1458 -5083 1492 -5049
rect 1458 -5151 1492 -5117
rect 1458 -5219 1492 -5185
rect 1458 -5287 1492 -5253
rect 1458 -5355 1492 -5321
rect 1458 -5423 1492 -5389
rect 1458 -5491 1492 -5457
rect 1458 -5559 1492 -5525
rect 1458 -5627 1492 -5593
rect 1458 -5695 1492 -5661
rect 1458 -5763 1492 -5729
rect 1458 -5831 1492 -5797
rect 1458 -5899 1492 -5865
rect 1458 -5967 1492 -5933
rect 1458 -6035 1492 -6001
rect 1458 -6103 1492 -6069
rect 1458 -6171 1492 -6137
rect 1458 -6239 1492 -6205
rect 1458 -6307 1492 -6273
rect 1458 -6375 1492 -6341
rect 1458 -6443 1492 -6409
rect 1458 -6511 1492 -6477
rect 1458 -6579 1492 -6545
rect 1458 -6647 1492 -6613
rect 1458 -6715 1492 -6681
rect 1458 -6783 1492 -6749
rect 1458 -6851 1492 -6817
rect 1458 -6919 1492 -6885
rect 1458 -6987 1492 -6953
rect 1458 -7055 1492 -7021
rect 1458 -7123 1492 -7089
rect 1458 -7191 1492 -7157
rect 1458 -7259 1492 -7225
rect 1458 -7327 1492 -7293
rect 1458 -7395 1492 -7361
rect 1458 -7463 1492 -7429
rect 1458 -7531 1492 -7497
rect 1458 -7599 1492 -7565
rect 1458 -7667 1492 -7633
rect 1458 -7735 1492 -7701
rect 1458 -7803 1492 -7769
rect 1458 -7871 1492 -7837
rect 1458 -7939 1492 -7905
rect 1458 -8007 1492 -7973
rect 1458 -8075 1492 -8041
rect 1458 -8143 1492 -8109
rect 1458 -8211 1492 -8177
rect 1458 -8279 1492 -8245
rect 1458 -8347 1492 -8313
rect 1458 -8415 1492 -8381
rect 1458 -8483 1492 -8449
rect 1458 -8551 1492 -8517
rect 1458 -8619 1492 -8585
rect 1458 -8687 1492 -8653
rect 1458 -8755 1492 -8721
rect 1458 -8823 1492 -8789
rect 1458 -8891 1492 -8857
rect 1458 -8959 1492 -8925
rect 1458 -9027 1492 -8993
rect 1458 -9095 1492 -9061
rect 1458 -9163 1492 -9129
rect 1458 -9231 1492 -9197
rect 1458 -9299 1492 -9265
rect 1458 -9367 1492 -9333
rect 1458 -9435 1492 -9401
rect 1458 -9503 1492 -9469
rect 1458 -9571 1492 -9537
<< poly >>
rect -1449 9678 -1383 9688
rect -1331 9678 -1265 9688
rect -1449 9632 -1265 9678
rect -1449 9622 -1383 9632
rect -1331 9622 -1265 9632
rect -1213 9678 -1147 9688
rect -1095 9678 -1029 9688
rect -1213 9632 -1029 9678
rect -1213 9622 -1147 9632
rect -1095 9622 -1029 9632
rect -977 9678 -911 9688
rect -859 9678 -793 9688
rect -977 9632 -793 9678
rect -977 9622 -911 9632
rect -859 9622 -793 9632
rect -741 9678 -675 9688
rect -623 9678 -557 9688
rect -741 9632 -557 9678
rect -741 9622 -675 9632
rect -623 9622 -557 9632
rect -505 9678 -439 9688
rect -387 9678 -321 9688
rect -505 9632 -321 9678
rect -505 9622 -439 9632
rect -387 9622 -321 9632
rect -269 9678 -203 9688
rect -151 9678 -85 9688
rect -269 9632 -85 9678
rect -269 9622 -203 9632
rect -151 9622 -85 9632
rect -33 9678 33 9688
rect 85 9678 151 9688
rect -33 9632 151 9678
rect -33 9622 33 9632
rect 85 9622 151 9632
rect 203 9678 269 9688
rect 321 9678 387 9688
rect 203 9632 387 9678
rect 203 9622 269 9632
rect 321 9622 387 9632
rect 439 9678 505 9688
rect 557 9678 623 9688
rect 439 9632 623 9678
rect 439 9622 505 9632
rect 557 9622 623 9632
rect 675 9678 741 9688
rect 793 9678 859 9688
rect 675 9632 859 9678
rect 675 9622 741 9632
rect 793 9622 859 9632
rect 911 9678 977 9688
rect 1029 9678 1095 9688
rect 911 9632 1095 9678
rect 911 9622 977 9632
rect 1029 9622 1095 9632
rect 1147 9678 1213 9688
rect 1265 9678 1331 9688
rect 1147 9632 1331 9678
rect 1147 9622 1213 9632
rect 1265 9622 1331 9632
rect 1383 9622 1449 9688
rect -1446 9600 -1386 9622
rect -1328 9600 -1268 9622
rect -1210 9600 -1150 9622
rect -1092 9600 -1032 9622
rect -974 9600 -914 9622
rect -856 9600 -796 9622
rect -738 9600 -678 9622
rect -620 9600 -560 9622
rect -502 9600 -442 9622
rect -384 9600 -324 9622
rect -266 9600 -206 9622
rect -148 9600 -88 9622
rect -30 9600 30 9622
rect 88 9600 148 9622
rect 206 9600 266 9622
rect 324 9600 384 9622
rect 442 9600 502 9622
rect 560 9600 620 9622
rect 678 9600 738 9622
rect 796 9600 856 9622
rect 914 9600 974 9622
rect 1032 9600 1092 9622
rect 1150 9600 1210 9622
rect 1268 9600 1328 9622
rect 1386 9600 1446 9622
rect -1446 -9622 -1386 -9600
rect -1328 -9622 -1268 -9600
rect -1210 -9622 -1150 -9600
rect -1092 -9622 -1032 -9600
rect -974 -9622 -914 -9600
rect -856 -9622 -796 -9600
rect -738 -9622 -678 -9600
rect -620 -9622 -560 -9600
rect -502 -9622 -442 -9600
rect -384 -9622 -324 -9600
rect -266 -9622 -206 -9600
rect -148 -9622 -88 -9600
rect -30 -9622 30 -9600
rect 88 -9622 148 -9600
rect 206 -9622 266 -9600
rect 324 -9622 384 -9600
rect 442 -9622 502 -9600
rect 560 -9622 620 -9600
rect 678 -9622 738 -9600
rect 796 -9622 856 -9600
rect 914 -9622 974 -9600
rect 1032 -9622 1092 -9600
rect 1150 -9622 1210 -9600
rect 1268 -9622 1328 -9600
rect 1386 -9622 1446 -9600
rect -1449 -9688 -1383 -9622
rect -1331 -9632 -1265 -9622
rect -1213 -9632 -1147 -9622
rect -1331 -9678 -1147 -9632
rect -1331 -9688 -1265 -9678
rect -1213 -9688 -1147 -9678
rect -1095 -9632 -1029 -9622
rect -977 -9632 -911 -9622
rect -1095 -9678 -911 -9632
rect -1095 -9688 -1029 -9678
rect -977 -9688 -911 -9678
rect -859 -9632 -793 -9622
rect -741 -9632 -675 -9622
rect -859 -9678 -675 -9632
rect -859 -9688 -793 -9678
rect -741 -9688 -675 -9678
rect -623 -9632 -557 -9622
rect -505 -9632 -439 -9622
rect -623 -9678 -439 -9632
rect -623 -9688 -557 -9678
rect -505 -9688 -439 -9678
rect -387 -9632 -321 -9622
rect -269 -9632 -203 -9622
rect -387 -9678 -203 -9632
rect -387 -9688 -321 -9678
rect -269 -9688 -203 -9678
rect -151 -9632 -85 -9622
rect -33 -9632 33 -9622
rect -151 -9678 33 -9632
rect -151 -9688 -85 -9678
rect -33 -9688 33 -9678
rect 85 -9632 151 -9622
rect 203 -9632 269 -9622
rect 85 -9678 269 -9632
rect 85 -9688 151 -9678
rect 203 -9688 269 -9678
rect 321 -9632 387 -9622
rect 439 -9632 505 -9622
rect 321 -9678 505 -9632
rect 321 -9688 387 -9678
rect 439 -9688 505 -9678
rect 557 -9632 623 -9622
rect 675 -9632 741 -9622
rect 557 -9678 741 -9632
rect 557 -9688 623 -9678
rect 675 -9688 741 -9678
rect 793 -9632 859 -9622
rect 911 -9632 977 -9622
rect 793 -9678 977 -9632
rect 793 -9688 859 -9678
rect 911 -9688 977 -9678
rect 1029 -9632 1095 -9622
rect 1147 -9632 1213 -9622
rect 1029 -9678 1213 -9632
rect 1029 -9688 1095 -9678
rect 1147 -9688 1213 -9678
rect 1265 -9632 1331 -9622
rect 1383 -9632 1449 -9622
rect 1265 -9678 1449 -9632
rect 1265 -9688 1331 -9678
rect 1383 -9688 1449 -9678
<< locali >>
rect -1492 9571 -1458 9604
rect -1492 9503 -1458 9523
rect -1492 9435 -1458 9451
rect -1492 9367 -1458 9379
rect -1492 9299 -1458 9307
rect -1492 9231 -1458 9235
rect -1492 9125 -1458 9129
rect -1492 9053 -1458 9061
rect -1492 8981 -1458 8993
rect -1492 8909 -1458 8925
rect -1492 8837 -1458 8857
rect -1492 8765 -1458 8789
rect -1492 8693 -1458 8721
rect -1492 8621 -1458 8653
rect -1492 8551 -1458 8585
rect -1492 8483 -1458 8515
rect -1492 8415 -1458 8443
rect -1492 8347 -1458 8371
rect -1492 8279 -1458 8299
rect -1492 8211 -1458 8227
rect -1492 8143 -1458 8155
rect -1492 8075 -1458 8083
rect -1492 8007 -1458 8011
rect -1492 7901 -1458 7905
rect -1492 7829 -1458 7837
rect -1492 7757 -1458 7769
rect -1492 7685 -1458 7701
rect -1492 7613 -1458 7633
rect -1492 7541 -1458 7565
rect -1492 7469 -1458 7497
rect -1492 7397 -1458 7429
rect -1492 7327 -1458 7361
rect -1492 7259 -1458 7291
rect -1492 7191 -1458 7219
rect -1492 7123 -1458 7147
rect -1492 7055 -1458 7075
rect -1492 6987 -1458 7003
rect -1492 6919 -1458 6931
rect -1492 6851 -1458 6859
rect -1492 6783 -1458 6787
rect -1492 6677 -1458 6681
rect -1492 6605 -1458 6613
rect -1492 6533 -1458 6545
rect -1492 6461 -1458 6477
rect -1492 6389 -1458 6409
rect -1492 6317 -1458 6341
rect -1492 6245 -1458 6273
rect -1492 6173 -1458 6205
rect -1492 6103 -1458 6137
rect -1492 6035 -1458 6067
rect -1492 5967 -1458 5995
rect -1492 5899 -1458 5923
rect -1492 5831 -1458 5851
rect -1492 5763 -1458 5779
rect -1492 5695 -1458 5707
rect -1492 5627 -1458 5635
rect -1492 5559 -1458 5563
rect -1492 5453 -1458 5457
rect -1492 5381 -1458 5389
rect -1492 5309 -1458 5321
rect -1492 5237 -1458 5253
rect -1492 5165 -1458 5185
rect -1492 5093 -1458 5117
rect -1492 5021 -1458 5049
rect -1492 4949 -1458 4981
rect -1492 4879 -1458 4913
rect -1492 4811 -1458 4843
rect -1492 4743 -1458 4771
rect -1492 4675 -1458 4699
rect -1492 4607 -1458 4627
rect -1492 4539 -1458 4555
rect -1492 4471 -1458 4483
rect -1492 4403 -1458 4411
rect -1492 4335 -1458 4339
rect -1492 4229 -1458 4233
rect -1492 4157 -1458 4165
rect -1492 4085 -1458 4097
rect -1492 4013 -1458 4029
rect -1492 3941 -1458 3961
rect -1492 3869 -1458 3893
rect -1492 3797 -1458 3825
rect -1492 3725 -1458 3757
rect -1492 3655 -1458 3689
rect -1492 3587 -1458 3619
rect -1492 3519 -1458 3547
rect -1492 3451 -1458 3475
rect -1492 3383 -1458 3403
rect -1492 3315 -1458 3331
rect -1492 3247 -1458 3259
rect -1492 3179 -1458 3187
rect -1492 3111 -1458 3115
rect -1492 3005 -1458 3009
rect -1492 2933 -1458 2941
rect -1492 2861 -1458 2873
rect -1492 2789 -1458 2805
rect -1492 2717 -1458 2737
rect -1492 2645 -1458 2669
rect -1492 2573 -1458 2601
rect -1492 2501 -1458 2533
rect -1492 2431 -1458 2465
rect -1492 2363 -1458 2395
rect -1492 2295 -1458 2323
rect -1492 2227 -1458 2251
rect -1492 2159 -1458 2179
rect -1492 2091 -1458 2107
rect -1492 2023 -1458 2035
rect -1492 1955 -1458 1963
rect -1492 1887 -1458 1891
rect -1492 1781 -1458 1785
rect -1492 1709 -1458 1717
rect -1492 1637 -1458 1649
rect -1492 1565 -1458 1581
rect -1492 1493 -1458 1513
rect -1492 1421 -1458 1445
rect -1492 1349 -1458 1377
rect -1492 1277 -1458 1309
rect -1492 1207 -1458 1241
rect -1492 1139 -1458 1171
rect -1492 1071 -1458 1099
rect -1492 1003 -1458 1027
rect -1492 935 -1458 955
rect -1492 867 -1458 883
rect -1492 799 -1458 811
rect -1492 731 -1458 739
rect -1492 663 -1458 667
rect -1492 557 -1458 561
rect -1492 485 -1458 493
rect -1492 413 -1458 425
rect -1492 341 -1458 357
rect -1492 269 -1458 289
rect -1492 197 -1458 221
rect -1492 125 -1458 153
rect -1492 53 -1458 85
rect -1492 -17 -1458 17
rect -1492 -85 -1458 -53
rect -1492 -153 -1458 -125
rect -1492 -221 -1458 -197
rect -1492 -289 -1458 -269
rect -1492 -357 -1458 -341
rect -1492 -425 -1458 -413
rect -1492 -493 -1458 -485
rect -1492 -561 -1458 -557
rect -1492 -667 -1458 -663
rect -1492 -739 -1458 -731
rect -1492 -811 -1458 -799
rect -1492 -883 -1458 -867
rect -1492 -955 -1458 -935
rect -1492 -1027 -1458 -1003
rect -1492 -1099 -1458 -1071
rect -1492 -1171 -1458 -1139
rect -1492 -1241 -1458 -1207
rect -1492 -1309 -1458 -1277
rect -1492 -1377 -1458 -1349
rect -1492 -1445 -1458 -1421
rect -1492 -1513 -1458 -1493
rect -1492 -1581 -1458 -1565
rect -1492 -1649 -1458 -1637
rect -1492 -1717 -1458 -1709
rect -1492 -1785 -1458 -1781
rect -1492 -1891 -1458 -1887
rect -1492 -1963 -1458 -1955
rect -1492 -2035 -1458 -2023
rect -1492 -2107 -1458 -2091
rect -1492 -2179 -1458 -2159
rect -1492 -2251 -1458 -2227
rect -1492 -2323 -1458 -2295
rect -1492 -2395 -1458 -2363
rect -1492 -2465 -1458 -2431
rect -1492 -2533 -1458 -2501
rect -1492 -2601 -1458 -2573
rect -1492 -2669 -1458 -2645
rect -1492 -2737 -1458 -2717
rect -1492 -2805 -1458 -2789
rect -1492 -2873 -1458 -2861
rect -1492 -2941 -1458 -2933
rect -1492 -3009 -1458 -3005
rect -1492 -3115 -1458 -3111
rect -1492 -3187 -1458 -3179
rect -1492 -3259 -1458 -3247
rect -1492 -3331 -1458 -3315
rect -1492 -3403 -1458 -3383
rect -1492 -3475 -1458 -3451
rect -1492 -3547 -1458 -3519
rect -1492 -3619 -1458 -3587
rect -1492 -3689 -1458 -3655
rect -1492 -3757 -1458 -3725
rect -1492 -3825 -1458 -3797
rect -1492 -3893 -1458 -3869
rect -1492 -3961 -1458 -3941
rect -1492 -4029 -1458 -4013
rect -1492 -4097 -1458 -4085
rect -1492 -4165 -1458 -4157
rect -1492 -4233 -1458 -4229
rect -1492 -4339 -1458 -4335
rect -1492 -4411 -1458 -4403
rect -1492 -4483 -1458 -4471
rect -1492 -4555 -1458 -4539
rect -1492 -4627 -1458 -4607
rect -1492 -4699 -1458 -4675
rect -1492 -4771 -1458 -4743
rect -1492 -4843 -1458 -4811
rect -1492 -4913 -1458 -4879
rect -1492 -4981 -1458 -4949
rect -1492 -5049 -1458 -5021
rect -1492 -5117 -1458 -5093
rect -1492 -5185 -1458 -5165
rect -1492 -5253 -1458 -5237
rect -1492 -5321 -1458 -5309
rect -1492 -5389 -1458 -5381
rect -1492 -5457 -1458 -5453
rect -1492 -5563 -1458 -5559
rect -1492 -5635 -1458 -5627
rect -1492 -5707 -1458 -5695
rect -1492 -5779 -1458 -5763
rect -1492 -5851 -1458 -5831
rect -1492 -5923 -1458 -5899
rect -1492 -5995 -1458 -5967
rect -1492 -6067 -1458 -6035
rect -1492 -6137 -1458 -6103
rect -1492 -6205 -1458 -6173
rect -1492 -6273 -1458 -6245
rect -1492 -6341 -1458 -6317
rect -1492 -6409 -1458 -6389
rect -1492 -6477 -1458 -6461
rect -1492 -6545 -1458 -6533
rect -1492 -6613 -1458 -6605
rect -1492 -6681 -1458 -6677
rect -1492 -6787 -1458 -6783
rect -1492 -6859 -1458 -6851
rect -1492 -6931 -1458 -6919
rect -1492 -7003 -1458 -6987
rect -1492 -7075 -1458 -7055
rect -1492 -7147 -1458 -7123
rect -1492 -7219 -1458 -7191
rect -1492 -7291 -1458 -7259
rect -1492 -7361 -1458 -7327
rect -1492 -7429 -1458 -7397
rect -1492 -7497 -1458 -7469
rect -1492 -7565 -1458 -7541
rect -1492 -7633 -1458 -7613
rect -1492 -7701 -1458 -7685
rect -1492 -7769 -1458 -7757
rect -1492 -7837 -1458 -7829
rect -1492 -7905 -1458 -7901
rect -1492 -8011 -1458 -8007
rect -1492 -8083 -1458 -8075
rect -1492 -8155 -1458 -8143
rect -1492 -8227 -1458 -8211
rect -1492 -8299 -1458 -8279
rect -1492 -8371 -1458 -8347
rect -1492 -8443 -1458 -8415
rect -1492 -8515 -1458 -8483
rect -1492 -8585 -1458 -8551
rect -1492 -8653 -1458 -8621
rect -1492 -8721 -1458 -8693
rect -1492 -8789 -1458 -8765
rect -1492 -8857 -1458 -8837
rect -1492 -8925 -1458 -8909
rect -1492 -8993 -1458 -8981
rect -1492 -9061 -1458 -9053
rect -1492 -9129 -1458 -9125
rect -1492 -9235 -1458 -9231
rect -1492 -9307 -1458 -9299
rect -1492 -9379 -1458 -9367
rect -1492 -9451 -1458 -9435
rect -1492 -9523 -1458 -9503
rect -1492 -9604 -1458 -9571
rect -1374 9571 -1340 9604
rect -1374 9503 -1340 9523
rect -1374 9435 -1340 9451
rect -1374 9367 -1340 9379
rect -1374 9299 -1340 9307
rect -1374 9231 -1340 9235
rect -1374 9125 -1340 9129
rect -1374 9053 -1340 9061
rect -1374 8981 -1340 8993
rect -1374 8909 -1340 8925
rect -1374 8837 -1340 8857
rect -1374 8765 -1340 8789
rect -1374 8693 -1340 8721
rect -1374 8621 -1340 8653
rect -1374 8551 -1340 8585
rect -1374 8483 -1340 8515
rect -1374 8415 -1340 8443
rect -1374 8347 -1340 8371
rect -1374 8279 -1340 8299
rect -1374 8211 -1340 8227
rect -1374 8143 -1340 8155
rect -1374 8075 -1340 8083
rect -1374 8007 -1340 8011
rect -1374 7901 -1340 7905
rect -1374 7829 -1340 7837
rect -1374 7757 -1340 7769
rect -1374 7685 -1340 7701
rect -1374 7613 -1340 7633
rect -1374 7541 -1340 7565
rect -1374 7469 -1340 7497
rect -1374 7397 -1340 7429
rect -1374 7327 -1340 7361
rect -1374 7259 -1340 7291
rect -1374 7191 -1340 7219
rect -1374 7123 -1340 7147
rect -1374 7055 -1340 7075
rect -1374 6987 -1340 7003
rect -1374 6919 -1340 6931
rect -1374 6851 -1340 6859
rect -1374 6783 -1340 6787
rect -1374 6677 -1340 6681
rect -1374 6605 -1340 6613
rect -1374 6533 -1340 6545
rect -1374 6461 -1340 6477
rect -1374 6389 -1340 6409
rect -1374 6317 -1340 6341
rect -1374 6245 -1340 6273
rect -1374 6173 -1340 6205
rect -1374 6103 -1340 6137
rect -1374 6035 -1340 6067
rect -1374 5967 -1340 5995
rect -1374 5899 -1340 5923
rect -1374 5831 -1340 5851
rect -1374 5763 -1340 5779
rect -1374 5695 -1340 5707
rect -1374 5627 -1340 5635
rect -1374 5559 -1340 5563
rect -1374 5453 -1340 5457
rect -1374 5381 -1340 5389
rect -1374 5309 -1340 5321
rect -1374 5237 -1340 5253
rect -1374 5165 -1340 5185
rect -1374 5093 -1340 5117
rect -1374 5021 -1340 5049
rect -1374 4949 -1340 4981
rect -1374 4879 -1340 4913
rect -1374 4811 -1340 4843
rect -1374 4743 -1340 4771
rect -1374 4675 -1340 4699
rect -1374 4607 -1340 4627
rect -1374 4539 -1340 4555
rect -1374 4471 -1340 4483
rect -1374 4403 -1340 4411
rect -1374 4335 -1340 4339
rect -1374 4229 -1340 4233
rect -1374 4157 -1340 4165
rect -1374 4085 -1340 4097
rect -1374 4013 -1340 4029
rect -1374 3941 -1340 3961
rect -1374 3869 -1340 3893
rect -1374 3797 -1340 3825
rect -1374 3725 -1340 3757
rect -1374 3655 -1340 3689
rect -1374 3587 -1340 3619
rect -1374 3519 -1340 3547
rect -1374 3451 -1340 3475
rect -1374 3383 -1340 3403
rect -1374 3315 -1340 3331
rect -1374 3247 -1340 3259
rect -1374 3179 -1340 3187
rect -1374 3111 -1340 3115
rect -1374 3005 -1340 3009
rect -1374 2933 -1340 2941
rect -1374 2861 -1340 2873
rect -1374 2789 -1340 2805
rect -1374 2717 -1340 2737
rect -1374 2645 -1340 2669
rect -1374 2573 -1340 2601
rect -1374 2501 -1340 2533
rect -1374 2431 -1340 2465
rect -1374 2363 -1340 2395
rect -1374 2295 -1340 2323
rect -1374 2227 -1340 2251
rect -1374 2159 -1340 2179
rect -1374 2091 -1340 2107
rect -1374 2023 -1340 2035
rect -1374 1955 -1340 1963
rect -1374 1887 -1340 1891
rect -1374 1781 -1340 1785
rect -1374 1709 -1340 1717
rect -1374 1637 -1340 1649
rect -1374 1565 -1340 1581
rect -1374 1493 -1340 1513
rect -1374 1421 -1340 1445
rect -1374 1349 -1340 1377
rect -1374 1277 -1340 1309
rect -1374 1207 -1340 1241
rect -1374 1139 -1340 1171
rect -1374 1071 -1340 1099
rect -1374 1003 -1340 1027
rect -1374 935 -1340 955
rect -1374 867 -1340 883
rect -1374 799 -1340 811
rect -1374 731 -1340 739
rect -1374 663 -1340 667
rect -1374 557 -1340 561
rect -1374 485 -1340 493
rect -1374 413 -1340 425
rect -1374 341 -1340 357
rect -1374 269 -1340 289
rect -1374 197 -1340 221
rect -1374 125 -1340 153
rect -1374 53 -1340 85
rect -1374 -17 -1340 17
rect -1374 -85 -1340 -53
rect -1374 -153 -1340 -125
rect -1374 -221 -1340 -197
rect -1374 -289 -1340 -269
rect -1374 -357 -1340 -341
rect -1374 -425 -1340 -413
rect -1374 -493 -1340 -485
rect -1374 -561 -1340 -557
rect -1374 -667 -1340 -663
rect -1374 -739 -1340 -731
rect -1374 -811 -1340 -799
rect -1374 -883 -1340 -867
rect -1374 -955 -1340 -935
rect -1374 -1027 -1340 -1003
rect -1374 -1099 -1340 -1071
rect -1374 -1171 -1340 -1139
rect -1374 -1241 -1340 -1207
rect -1374 -1309 -1340 -1277
rect -1374 -1377 -1340 -1349
rect -1374 -1445 -1340 -1421
rect -1374 -1513 -1340 -1493
rect -1374 -1581 -1340 -1565
rect -1374 -1649 -1340 -1637
rect -1374 -1717 -1340 -1709
rect -1374 -1785 -1340 -1781
rect -1374 -1891 -1340 -1887
rect -1374 -1963 -1340 -1955
rect -1374 -2035 -1340 -2023
rect -1374 -2107 -1340 -2091
rect -1374 -2179 -1340 -2159
rect -1374 -2251 -1340 -2227
rect -1374 -2323 -1340 -2295
rect -1374 -2395 -1340 -2363
rect -1374 -2465 -1340 -2431
rect -1374 -2533 -1340 -2501
rect -1374 -2601 -1340 -2573
rect -1374 -2669 -1340 -2645
rect -1374 -2737 -1340 -2717
rect -1374 -2805 -1340 -2789
rect -1374 -2873 -1340 -2861
rect -1374 -2941 -1340 -2933
rect -1374 -3009 -1340 -3005
rect -1374 -3115 -1340 -3111
rect -1374 -3187 -1340 -3179
rect -1374 -3259 -1340 -3247
rect -1374 -3331 -1340 -3315
rect -1374 -3403 -1340 -3383
rect -1374 -3475 -1340 -3451
rect -1374 -3547 -1340 -3519
rect -1374 -3619 -1340 -3587
rect -1374 -3689 -1340 -3655
rect -1374 -3757 -1340 -3725
rect -1374 -3825 -1340 -3797
rect -1374 -3893 -1340 -3869
rect -1374 -3961 -1340 -3941
rect -1374 -4029 -1340 -4013
rect -1374 -4097 -1340 -4085
rect -1374 -4165 -1340 -4157
rect -1374 -4233 -1340 -4229
rect -1374 -4339 -1340 -4335
rect -1374 -4411 -1340 -4403
rect -1374 -4483 -1340 -4471
rect -1374 -4555 -1340 -4539
rect -1374 -4627 -1340 -4607
rect -1374 -4699 -1340 -4675
rect -1374 -4771 -1340 -4743
rect -1374 -4843 -1340 -4811
rect -1374 -4913 -1340 -4879
rect -1374 -4981 -1340 -4949
rect -1374 -5049 -1340 -5021
rect -1374 -5117 -1340 -5093
rect -1374 -5185 -1340 -5165
rect -1374 -5253 -1340 -5237
rect -1374 -5321 -1340 -5309
rect -1374 -5389 -1340 -5381
rect -1374 -5457 -1340 -5453
rect -1374 -5563 -1340 -5559
rect -1374 -5635 -1340 -5627
rect -1374 -5707 -1340 -5695
rect -1374 -5779 -1340 -5763
rect -1374 -5851 -1340 -5831
rect -1374 -5923 -1340 -5899
rect -1374 -5995 -1340 -5967
rect -1374 -6067 -1340 -6035
rect -1374 -6137 -1340 -6103
rect -1374 -6205 -1340 -6173
rect -1374 -6273 -1340 -6245
rect -1374 -6341 -1340 -6317
rect -1374 -6409 -1340 -6389
rect -1374 -6477 -1340 -6461
rect -1374 -6545 -1340 -6533
rect -1374 -6613 -1340 -6605
rect -1374 -6681 -1340 -6677
rect -1374 -6787 -1340 -6783
rect -1374 -6859 -1340 -6851
rect -1374 -6931 -1340 -6919
rect -1374 -7003 -1340 -6987
rect -1374 -7075 -1340 -7055
rect -1374 -7147 -1340 -7123
rect -1374 -7219 -1340 -7191
rect -1374 -7291 -1340 -7259
rect -1374 -7361 -1340 -7327
rect -1374 -7429 -1340 -7397
rect -1374 -7497 -1340 -7469
rect -1374 -7565 -1340 -7541
rect -1374 -7633 -1340 -7613
rect -1374 -7701 -1340 -7685
rect -1374 -7769 -1340 -7757
rect -1374 -7837 -1340 -7829
rect -1374 -7905 -1340 -7901
rect -1374 -8011 -1340 -8007
rect -1374 -8083 -1340 -8075
rect -1374 -8155 -1340 -8143
rect -1374 -8227 -1340 -8211
rect -1374 -8299 -1340 -8279
rect -1374 -8371 -1340 -8347
rect -1374 -8443 -1340 -8415
rect -1374 -8515 -1340 -8483
rect -1374 -8585 -1340 -8551
rect -1374 -8653 -1340 -8621
rect -1374 -8721 -1340 -8693
rect -1374 -8789 -1340 -8765
rect -1374 -8857 -1340 -8837
rect -1374 -8925 -1340 -8909
rect -1374 -8993 -1340 -8981
rect -1374 -9061 -1340 -9053
rect -1374 -9129 -1340 -9125
rect -1374 -9235 -1340 -9231
rect -1374 -9307 -1340 -9299
rect -1374 -9379 -1340 -9367
rect -1374 -9451 -1340 -9435
rect -1374 -9523 -1340 -9503
rect -1374 -9604 -1340 -9571
rect -1256 9571 -1222 9604
rect -1256 9503 -1222 9523
rect -1256 9435 -1222 9451
rect -1256 9367 -1222 9379
rect -1256 9299 -1222 9307
rect -1256 9231 -1222 9235
rect -1256 9125 -1222 9129
rect -1256 9053 -1222 9061
rect -1256 8981 -1222 8993
rect -1256 8909 -1222 8925
rect -1256 8837 -1222 8857
rect -1256 8765 -1222 8789
rect -1256 8693 -1222 8721
rect -1256 8621 -1222 8653
rect -1256 8551 -1222 8585
rect -1256 8483 -1222 8515
rect -1256 8415 -1222 8443
rect -1256 8347 -1222 8371
rect -1256 8279 -1222 8299
rect -1256 8211 -1222 8227
rect -1256 8143 -1222 8155
rect -1256 8075 -1222 8083
rect -1256 8007 -1222 8011
rect -1256 7901 -1222 7905
rect -1256 7829 -1222 7837
rect -1256 7757 -1222 7769
rect -1256 7685 -1222 7701
rect -1256 7613 -1222 7633
rect -1256 7541 -1222 7565
rect -1256 7469 -1222 7497
rect -1256 7397 -1222 7429
rect -1256 7327 -1222 7361
rect -1256 7259 -1222 7291
rect -1256 7191 -1222 7219
rect -1256 7123 -1222 7147
rect -1256 7055 -1222 7075
rect -1256 6987 -1222 7003
rect -1256 6919 -1222 6931
rect -1256 6851 -1222 6859
rect -1256 6783 -1222 6787
rect -1256 6677 -1222 6681
rect -1256 6605 -1222 6613
rect -1256 6533 -1222 6545
rect -1256 6461 -1222 6477
rect -1256 6389 -1222 6409
rect -1256 6317 -1222 6341
rect -1256 6245 -1222 6273
rect -1256 6173 -1222 6205
rect -1256 6103 -1222 6137
rect -1256 6035 -1222 6067
rect -1256 5967 -1222 5995
rect -1256 5899 -1222 5923
rect -1256 5831 -1222 5851
rect -1256 5763 -1222 5779
rect -1256 5695 -1222 5707
rect -1256 5627 -1222 5635
rect -1256 5559 -1222 5563
rect -1256 5453 -1222 5457
rect -1256 5381 -1222 5389
rect -1256 5309 -1222 5321
rect -1256 5237 -1222 5253
rect -1256 5165 -1222 5185
rect -1256 5093 -1222 5117
rect -1256 5021 -1222 5049
rect -1256 4949 -1222 4981
rect -1256 4879 -1222 4913
rect -1256 4811 -1222 4843
rect -1256 4743 -1222 4771
rect -1256 4675 -1222 4699
rect -1256 4607 -1222 4627
rect -1256 4539 -1222 4555
rect -1256 4471 -1222 4483
rect -1256 4403 -1222 4411
rect -1256 4335 -1222 4339
rect -1256 4229 -1222 4233
rect -1256 4157 -1222 4165
rect -1256 4085 -1222 4097
rect -1256 4013 -1222 4029
rect -1256 3941 -1222 3961
rect -1256 3869 -1222 3893
rect -1256 3797 -1222 3825
rect -1256 3725 -1222 3757
rect -1256 3655 -1222 3689
rect -1256 3587 -1222 3619
rect -1256 3519 -1222 3547
rect -1256 3451 -1222 3475
rect -1256 3383 -1222 3403
rect -1256 3315 -1222 3331
rect -1256 3247 -1222 3259
rect -1256 3179 -1222 3187
rect -1256 3111 -1222 3115
rect -1256 3005 -1222 3009
rect -1256 2933 -1222 2941
rect -1256 2861 -1222 2873
rect -1256 2789 -1222 2805
rect -1256 2717 -1222 2737
rect -1256 2645 -1222 2669
rect -1256 2573 -1222 2601
rect -1256 2501 -1222 2533
rect -1256 2431 -1222 2465
rect -1256 2363 -1222 2395
rect -1256 2295 -1222 2323
rect -1256 2227 -1222 2251
rect -1256 2159 -1222 2179
rect -1256 2091 -1222 2107
rect -1256 2023 -1222 2035
rect -1256 1955 -1222 1963
rect -1256 1887 -1222 1891
rect -1256 1781 -1222 1785
rect -1256 1709 -1222 1717
rect -1256 1637 -1222 1649
rect -1256 1565 -1222 1581
rect -1256 1493 -1222 1513
rect -1256 1421 -1222 1445
rect -1256 1349 -1222 1377
rect -1256 1277 -1222 1309
rect -1256 1207 -1222 1241
rect -1256 1139 -1222 1171
rect -1256 1071 -1222 1099
rect -1256 1003 -1222 1027
rect -1256 935 -1222 955
rect -1256 867 -1222 883
rect -1256 799 -1222 811
rect -1256 731 -1222 739
rect -1256 663 -1222 667
rect -1256 557 -1222 561
rect -1256 485 -1222 493
rect -1256 413 -1222 425
rect -1256 341 -1222 357
rect -1256 269 -1222 289
rect -1256 197 -1222 221
rect -1256 125 -1222 153
rect -1256 53 -1222 85
rect -1256 -17 -1222 17
rect -1256 -85 -1222 -53
rect -1256 -153 -1222 -125
rect -1256 -221 -1222 -197
rect -1256 -289 -1222 -269
rect -1256 -357 -1222 -341
rect -1256 -425 -1222 -413
rect -1256 -493 -1222 -485
rect -1256 -561 -1222 -557
rect -1256 -667 -1222 -663
rect -1256 -739 -1222 -731
rect -1256 -811 -1222 -799
rect -1256 -883 -1222 -867
rect -1256 -955 -1222 -935
rect -1256 -1027 -1222 -1003
rect -1256 -1099 -1222 -1071
rect -1256 -1171 -1222 -1139
rect -1256 -1241 -1222 -1207
rect -1256 -1309 -1222 -1277
rect -1256 -1377 -1222 -1349
rect -1256 -1445 -1222 -1421
rect -1256 -1513 -1222 -1493
rect -1256 -1581 -1222 -1565
rect -1256 -1649 -1222 -1637
rect -1256 -1717 -1222 -1709
rect -1256 -1785 -1222 -1781
rect -1256 -1891 -1222 -1887
rect -1256 -1963 -1222 -1955
rect -1256 -2035 -1222 -2023
rect -1256 -2107 -1222 -2091
rect -1256 -2179 -1222 -2159
rect -1256 -2251 -1222 -2227
rect -1256 -2323 -1222 -2295
rect -1256 -2395 -1222 -2363
rect -1256 -2465 -1222 -2431
rect -1256 -2533 -1222 -2501
rect -1256 -2601 -1222 -2573
rect -1256 -2669 -1222 -2645
rect -1256 -2737 -1222 -2717
rect -1256 -2805 -1222 -2789
rect -1256 -2873 -1222 -2861
rect -1256 -2941 -1222 -2933
rect -1256 -3009 -1222 -3005
rect -1256 -3115 -1222 -3111
rect -1256 -3187 -1222 -3179
rect -1256 -3259 -1222 -3247
rect -1256 -3331 -1222 -3315
rect -1256 -3403 -1222 -3383
rect -1256 -3475 -1222 -3451
rect -1256 -3547 -1222 -3519
rect -1256 -3619 -1222 -3587
rect -1256 -3689 -1222 -3655
rect -1256 -3757 -1222 -3725
rect -1256 -3825 -1222 -3797
rect -1256 -3893 -1222 -3869
rect -1256 -3961 -1222 -3941
rect -1256 -4029 -1222 -4013
rect -1256 -4097 -1222 -4085
rect -1256 -4165 -1222 -4157
rect -1256 -4233 -1222 -4229
rect -1256 -4339 -1222 -4335
rect -1256 -4411 -1222 -4403
rect -1256 -4483 -1222 -4471
rect -1256 -4555 -1222 -4539
rect -1256 -4627 -1222 -4607
rect -1256 -4699 -1222 -4675
rect -1256 -4771 -1222 -4743
rect -1256 -4843 -1222 -4811
rect -1256 -4913 -1222 -4879
rect -1256 -4981 -1222 -4949
rect -1256 -5049 -1222 -5021
rect -1256 -5117 -1222 -5093
rect -1256 -5185 -1222 -5165
rect -1256 -5253 -1222 -5237
rect -1256 -5321 -1222 -5309
rect -1256 -5389 -1222 -5381
rect -1256 -5457 -1222 -5453
rect -1256 -5563 -1222 -5559
rect -1256 -5635 -1222 -5627
rect -1256 -5707 -1222 -5695
rect -1256 -5779 -1222 -5763
rect -1256 -5851 -1222 -5831
rect -1256 -5923 -1222 -5899
rect -1256 -5995 -1222 -5967
rect -1256 -6067 -1222 -6035
rect -1256 -6137 -1222 -6103
rect -1256 -6205 -1222 -6173
rect -1256 -6273 -1222 -6245
rect -1256 -6341 -1222 -6317
rect -1256 -6409 -1222 -6389
rect -1256 -6477 -1222 -6461
rect -1256 -6545 -1222 -6533
rect -1256 -6613 -1222 -6605
rect -1256 -6681 -1222 -6677
rect -1256 -6787 -1222 -6783
rect -1256 -6859 -1222 -6851
rect -1256 -6931 -1222 -6919
rect -1256 -7003 -1222 -6987
rect -1256 -7075 -1222 -7055
rect -1256 -7147 -1222 -7123
rect -1256 -7219 -1222 -7191
rect -1256 -7291 -1222 -7259
rect -1256 -7361 -1222 -7327
rect -1256 -7429 -1222 -7397
rect -1256 -7497 -1222 -7469
rect -1256 -7565 -1222 -7541
rect -1256 -7633 -1222 -7613
rect -1256 -7701 -1222 -7685
rect -1256 -7769 -1222 -7757
rect -1256 -7837 -1222 -7829
rect -1256 -7905 -1222 -7901
rect -1256 -8011 -1222 -8007
rect -1256 -8083 -1222 -8075
rect -1256 -8155 -1222 -8143
rect -1256 -8227 -1222 -8211
rect -1256 -8299 -1222 -8279
rect -1256 -8371 -1222 -8347
rect -1256 -8443 -1222 -8415
rect -1256 -8515 -1222 -8483
rect -1256 -8585 -1222 -8551
rect -1256 -8653 -1222 -8621
rect -1256 -8721 -1222 -8693
rect -1256 -8789 -1222 -8765
rect -1256 -8857 -1222 -8837
rect -1256 -8925 -1222 -8909
rect -1256 -8993 -1222 -8981
rect -1256 -9061 -1222 -9053
rect -1256 -9129 -1222 -9125
rect -1256 -9235 -1222 -9231
rect -1256 -9307 -1222 -9299
rect -1256 -9379 -1222 -9367
rect -1256 -9451 -1222 -9435
rect -1256 -9523 -1222 -9503
rect -1256 -9604 -1222 -9571
rect -1138 9571 -1104 9604
rect -1138 9503 -1104 9523
rect -1138 9435 -1104 9451
rect -1138 9367 -1104 9379
rect -1138 9299 -1104 9307
rect -1138 9231 -1104 9235
rect -1138 9125 -1104 9129
rect -1138 9053 -1104 9061
rect -1138 8981 -1104 8993
rect -1138 8909 -1104 8925
rect -1138 8837 -1104 8857
rect -1138 8765 -1104 8789
rect -1138 8693 -1104 8721
rect -1138 8621 -1104 8653
rect -1138 8551 -1104 8585
rect -1138 8483 -1104 8515
rect -1138 8415 -1104 8443
rect -1138 8347 -1104 8371
rect -1138 8279 -1104 8299
rect -1138 8211 -1104 8227
rect -1138 8143 -1104 8155
rect -1138 8075 -1104 8083
rect -1138 8007 -1104 8011
rect -1138 7901 -1104 7905
rect -1138 7829 -1104 7837
rect -1138 7757 -1104 7769
rect -1138 7685 -1104 7701
rect -1138 7613 -1104 7633
rect -1138 7541 -1104 7565
rect -1138 7469 -1104 7497
rect -1138 7397 -1104 7429
rect -1138 7327 -1104 7361
rect -1138 7259 -1104 7291
rect -1138 7191 -1104 7219
rect -1138 7123 -1104 7147
rect -1138 7055 -1104 7075
rect -1138 6987 -1104 7003
rect -1138 6919 -1104 6931
rect -1138 6851 -1104 6859
rect -1138 6783 -1104 6787
rect -1138 6677 -1104 6681
rect -1138 6605 -1104 6613
rect -1138 6533 -1104 6545
rect -1138 6461 -1104 6477
rect -1138 6389 -1104 6409
rect -1138 6317 -1104 6341
rect -1138 6245 -1104 6273
rect -1138 6173 -1104 6205
rect -1138 6103 -1104 6137
rect -1138 6035 -1104 6067
rect -1138 5967 -1104 5995
rect -1138 5899 -1104 5923
rect -1138 5831 -1104 5851
rect -1138 5763 -1104 5779
rect -1138 5695 -1104 5707
rect -1138 5627 -1104 5635
rect -1138 5559 -1104 5563
rect -1138 5453 -1104 5457
rect -1138 5381 -1104 5389
rect -1138 5309 -1104 5321
rect -1138 5237 -1104 5253
rect -1138 5165 -1104 5185
rect -1138 5093 -1104 5117
rect -1138 5021 -1104 5049
rect -1138 4949 -1104 4981
rect -1138 4879 -1104 4913
rect -1138 4811 -1104 4843
rect -1138 4743 -1104 4771
rect -1138 4675 -1104 4699
rect -1138 4607 -1104 4627
rect -1138 4539 -1104 4555
rect -1138 4471 -1104 4483
rect -1138 4403 -1104 4411
rect -1138 4335 -1104 4339
rect -1138 4229 -1104 4233
rect -1138 4157 -1104 4165
rect -1138 4085 -1104 4097
rect -1138 4013 -1104 4029
rect -1138 3941 -1104 3961
rect -1138 3869 -1104 3893
rect -1138 3797 -1104 3825
rect -1138 3725 -1104 3757
rect -1138 3655 -1104 3689
rect -1138 3587 -1104 3619
rect -1138 3519 -1104 3547
rect -1138 3451 -1104 3475
rect -1138 3383 -1104 3403
rect -1138 3315 -1104 3331
rect -1138 3247 -1104 3259
rect -1138 3179 -1104 3187
rect -1138 3111 -1104 3115
rect -1138 3005 -1104 3009
rect -1138 2933 -1104 2941
rect -1138 2861 -1104 2873
rect -1138 2789 -1104 2805
rect -1138 2717 -1104 2737
rect -1138 2645 -1104 2669
rect -1138 2573 -1104 2601
rect -1138 2501 -1104 2533
rect -1138 2431 -1104 2465
rect -1138 2363 -1104 2395
rect -1138 2295 -1104 2323
rect -1138 2227 -1104 2251
rect -1138 2159 -1104 2179
rect -1138 2091 -1104 2107
rect -1138 2023 -1104 2035
rect -1138 1955 -1104 1963
rect -1138 1887 -1104 1891
rect -1138 1781 -1104 1785
rect -1138 1709 -1104 1717
rect -1138 1637 -1104 1649
rect -1138 1565 -1104 1581
rect -1138 1493 -1104 1513
rect -1138 1421 -1104 1445
rect -1138 1349 -1104 1377
rect -1138 1277 -1104 1309
rect -1138 1207 -1104 1241
rect -1138 1139 -1104 1171
rect -1138 1071 -1104 1099
rect -1138 1003 -1104 1027
rect -1138 935 -1104 955
rect -1138 867 -1104 883
rect -1138 799 -1104 811
rect -1138 731 -1104 739
rect -1138 663 -1104 667
rect -1138 557 -1104 561
rect -1138 485 -1104 493
rect -1138 413 -1104 425
rect -1138 341 -1104 357
rect -1138 269 -1104 289
rect -1138 197 -1104 221
rect -1138 125 -1104 153
rect -1138 53 -1104 85
rect -1138 -17 -1104 17
rect -1138 -85 -1104 -53
rect -1138 -153 -1104 -125
rect -1138 -221 -1104 -197
rect -1138 -289 -1104 -269
rect -1138 -357 -1104 -341
rect -1138 -425 -1104 -413
rect -1138 -493 -1104 -485
rect -1138 -561 -1104 -557
rect -1138 -667 -1104 -663
rect -1138 -739 -1104 -731
rect -1138 -811 -1104 -799
rect -1138 -883 -1104 -867
rect -1138 -955 -1104 -935
rect -1138 -1027 -1104 -1003
rect -1138 -1099 -1104 -1071
rect -1138 -1171 -1104 -1139
rect -1138 -1241 -1104 -1207
rect -1138 -1309 -1104 -1277
rect -1138 -1377 -1104 -1349
rect -1138 -1445 -1104 -1421
rect -1138 -1513 -1104 -1493
rect -1138 -1581 -1104 -1565
rect -1138 -1649 -1104 -1637
rect -1138 -1717 -1104 -1709
rect -1138 -1785 -1104 -1781
rect -1138 -1891 -1104 -1887
rect -1138 -1963 -1104 -1955
rect -1138 -2035 -1104 -2023
rect -1138 -2107 -1104 -2091
rect -1138 -2179 -1104 -2159
rect -1138 -2251 -1104 -2227
rect -1138 -2323 -1104 -2295
rect -1138 -2395 -1104 -2363
rect -1138 -2465 -1104 -2431
rect -1138 -2533 -1104 -2501
rect -1138 -2601 -1104 -2573
rect -1138 -2669 -1104 -2645
rect -1138 -2737 -1104 -2717
rect -1138 -2805 -1104 -2789
rect -1138 -2873 -1104 -2861
rect -1138 -2941 -1104 -2933
rect -1138 -3009 -1104 -3005
rect -1138 -3115 -1104 -3111
rect -1138 -3187 -1104 -3179
rect -1138 -3259 -1104 -3247
rect -1138 -3331 -1104 -3315
rect -1138 -3403 -1104 -3383
rect -1138 -3475 -1104 -3451
rect -1138 -3547 -1104 -3519
rect -1138 -3619 -1104 -3587
rect -1138 -3689 -1104 -3655
rect -1138 -3757 -1104 -3725
rect -1138 -3825 -1104 -3797
rect -1138 -3893 -1104 -3869
rect -1138 -3961 -1104 -3941
rect -1138 -4029 -1104 -4013
rect -1138 -4097 -1104 -4085
rect -1138 -4165 -1104 -4157
rect -1138 -4233 -1104 -4229
rect -1138 -4339 -1104 -4335
rect -1138 -4411 -1104 -4403
rect -1138 -4483 -1104 -4471
rect -1138 -4555 -1104 -4539
rect -1138 -4627 -1104 -4607
rect -1138 -4699 -1104 -4675
rect -1138 -4771 -1104 -4743
rect -1138 -4843 -1104 -4811
rect -1138 -4913 -1104 -4879
rect -1138 -4981 -1104 -4949
rect -1138 -5049 -1104 -5021
rect -1138 -5117 -1104 -5093
rect -1138 -5185 -1104 -5165
rect -1138 -5253 -1104 -5237
rect -1138 -5321 -1104 -5309
rect -1138 -5389 -1104 -5381
rect -1138 -5457 -1104 -5453
rect -1138 -5563 -1104 -5559
rect -1138 -5635 -1104 -5627
rect -1138 -5707 -1104 -5695
rect -1138 -5779 -1104 -5763
rect -1138 -5851 -1104 -5831
rect -1138 -5923 -1104 -5899
rect -1138 -5995 -1104 -5967
rect -1138 -6067 -1104 -6035
rect -1138 -6137 -1104 -6103
rect -1138 -6205 -1104 -6173
rect -1138 -6273 -1104 -6245
rect -1138 -6341 -1104 -6317
rect -1138 -6409 -1104 -6389
rect -1138 -6477 -1104 -6461
rect -1138 -6545 -1104 -6533
rect -1138 -6613 -1104 -6605
rect -1138 -6681 -1104 -6677
rect -1138 -6787 -1104 -6783
rect -1138 -6859 -1104 -6851
rect -1138 -6931 -1104 -6919
rect -1138 -7003 -1104 -6987
rect -1138 -7075 -1104 -7055
rect -1138 -7147 -1104 -7123
rect -1138 -7219 -1104 -7191
rect -1138 -7291 -1104 -7259
rect -1138 -7361 -1104 -7327
rect -1138 -7429 -1104 -7397
rect -1138 -7497 -1104 -7469
rect -1138 -7565 -1104 -7541
rect -1138 -7633 -1104 -7613
rect -1138 -7701 -1104 -7685
rect -1138 -7769 -1104 -7757
rect -1138 -7837 -1104 -7829
rect -1138 -7905 -1104 -7901
rect -1138 -8011 -1104 -8007
rect -1138 -8083 -1104 -8075
rect -1138 -8155 -1104 -8143
rect -1138 -8227 -1104 -8211
rect -1138 -8299 -1104 -8279
rect -1138 -8371 -1104 -8347
rect -1138 -8443 -1104 -8415
rect -1138 -8515 -1104 -8483
rect -1138 -8585 -1104 -8551
rect -1138 -8653 -1104 -8621
rect -1138 -8721 -1104 -8693
rect -1138 -8789 -1104 -8765
rect -1138 -8857 -1104 -8837
rect -1138 -8925 -1104 -8909
rect -1138 -8993 -1104 -8981
rect -1138 -9061 -1104 -9053
rect -1138 -9129 -1104 -9125
rect -1138 -9235 -1104 -9231
rect -1138 -9307 -1104 -9299
rect -1138 -9379 -1104 -9367
rect -1138 -9451 -1104 -9435
rect -1138 -9523 -1104 -9503
rect -1138 -9604 -1104 -9571
rect -1020 9571 -986 9604
rect -1020 9503 -986 9523
rect -1020 9435 -986 9451
rect -1020 9367 -986 9379
rect -1020 9299 -986 9307
rect -1020 9231 -986 9235
rect -1020 9125 -986 9129
rect -1020 9053 -986 9061
rect -1020 8981 -986 8993
rect -1020 8909 -986 8925
rect -1020 8837 -986 8857
rect -1020 8765 -986 8789
rect -1020 8693 -986 8721
rect -1020 8621 -986 8653
rect -1020 8551 -986 8585
rect -1020 8483 -986 8515
rect -1020 8415 -986 8443
rect -1020 8347 -986 8371
rect -1020 8279 -986 8299
rect -1020 8211 -986 8227
rect -1020 8143 -986 8155
rect -1020 8075 -986 8083
rect -1020 8007 -986 8011
rect -1020 7901 -986 7905
rect -1020 7829 -986 7837
rect -1020 7757 -986 7769
rect -1020 7685 -986 7701
rect -1020 7613 -986 7633
rect -1020 7541 -986 7565
rect -1020 7469 -986 7497
rect -1020 7397 -986 7429
rect -1020 7327 -986 7361
rect -1020 7259 -986 7291
rect -1020 7191 -986 7219
rect -1020 7123 -986 7147
rect -1020 7055 -986 7075
rect -1020 6987 -986 7003
rect -1020 6919 -986 6931
rect -1020 6851 -986 6859
rect -1020 6783 -986 6787
rect -1020 6677 -986 6681
rect -1020 6605 -986 6613
rect -1020 6533 -986 6545
rect -1020 6461 -986 6477
rect -1020 6389 -986 6409
rect -1020 6317 -986 6341
rect -1020 6245 -986 6273
rect -1020 6173 -986 6205
rect -1020 6103 -986 6137
rect -1020 6035 -986 6067
rect -1020 5967 -986 5995
rect -1020 5899 -986 5923
rect -1020 5831 -986 5851
rect -1020 5763 -986 5779
rect -1020 5695 -986 5707
rect -1020 5627 -986 5635
rect -1020 5559 -986 5563
rect -1020 5453 -986 5457
rect -1020 5381 -986 5389
rect -1020 5309 -986 5321
rect -1020 5237 -986 5253
rect -1020 5165 -986 5185
rect -1020 5093 -986 5117
rect -1020 5021 -986 5049
rect -1020 4949 -986 4981
rect -1020 4879 -986 4913
rect -1020 4811 -986 4843
rect -1020 4743 -986 4771
rect -1020 4675 -986 4699
rect -1020 4607 -986 4627
rect -1020 4539 -986 4555
rect -1020 4471 -986 4483
rect -1020 4403 -986 4411
rect -1020 4335 -986 4339
rect -1020 4229 -986 4233
rect -1020 4157 -986 4165
rect -1020 4085 -986 4097
rect -1020 4013 -986 4029
rect -1020 3941 -986 3961
rect -1020 3869 -986 3893
rect -1020 3797 -986 3825
rect -1020 3725 -986 3757
rect -1020 3655 -986 3689
rect -1020 3587 -986 3619
rect -1020 3519 -986 3547
rect -1020 3451 -986 3475
rect -1020 3383 -986 3403
rect -1020 3315 -986 3331
rect -1020 3247 -986 3259
rect -1020 3179 -986 3187
rect -1020 3111 -986 3115
rect -1020 3005 -986 3009
rect -1020 2933 -986 2941
rect -1020 2861 -986 2873
rect -1020 2789 -986 2805
rect -1020 2717 -986 2737
rect -1020 2645 -986 2669
rect -1020 2573 -986 2601
rect -1020 2501 -986 2533
rect -1020 2431 -986 2465
rect -1020 2363 -986 2395
rect -1020 2295 -986 2323
rect -1020 2227 -986 2251
rect -1020 2159 -986 2179
rect -1020 2091 -986 2107
rect -1020 2023 -986 2035
rect -1020 1955 -986 1963
rect -1020 1887 -986 1891
rect -1020 1781 -986 1785
rect -1020 1709 -986 1717
rect -1020 1637 -986 1649
rect -1020 1565 -986 1581
rect -1020 1493 -986 1513
rect -1020 1421 -986 1445
rect -1020 1349 -986 1377
rect -1020 1277 -986 1309
rect -1020 1207 -986 1241
rect -1020 1139 -986 1171
rect -1020 1071 -986 1099
rect -1020 1003 -986 1027
rect -1020 935 -986 955
rect -1020 867 -986 883
rect -1020 799 -986 811
rect -1020 731 -986 739
rect -1020 663 -986 667
rect -1020 557 -986 561
rect -1020 485 -986 493
rect -1020 413 -986 425
rect -1020 341 -986 357
rect -1020 269 -986 289
rect -1020 197 -986 221
rect -1020 125 -986 153
rect -1020 53 -986 85
rect -1020 -17 -986 17
rect -1020 -85 -986 -53
rect -1020 -153 -986 -125
rect -1020 -221 -986 -197
rect -1020 -289 -986 -269
rect -1020 -357 -986 -341
rect -1020 -425 -986 -413
rect -1020 -493 -986 -485
rect -1020 -561 -986 -557
rect -1020 -667 -986 -663
rect -1020 -739 -986 -731
rect -1020 -811 -986 -799
rect -1020 -883 -986 -867
rect -1020 -955 -986 -935
rect -1020 -1027 -986 -1003
rect -1020 -1099 -986 -1071
rect -1020 -1171 -986 -1139
rect -1020 -1241 -986 -1207
rect -1020 -1309 -986 -1277
rect -1020 -1377 -986 -1349
rect -1020 -1445 -986 -1421
rect -1020 -1513 -986 -1493
rect -1020 -1581 -986 -1565
rect -1020 -1649 -986 -1637
rect -1020 -1717 -986 -1709
rect -1020 -1785 -986 -1781
rect -1020 -1891 -986 -1887
rect -1020 -1963 -986 -1955
rect -1020 -2035 -986 -2023
rect -1020 -2107 -986 -2091
rect -1020 -2179 -986 -2159
rect -1020 -2251 -986 -2227
rect -1020 -2323 -986 -2295
rect -1020 -2395 -986 -2363
rect -1020 -2465 -986 -2431
rect -1020 -2533 -986 -2501
rect -1020 -2601 -986 -2573
rect -1020 -2669 -986 -2645
rect -1020 -2737 -986 -2717
rect -1020 -2805 -986 -2789
rect -1020 -2873 -986 -2861
rect -1020 -2941 -986 -2933
rect -1020 -3009 -986 -3005
rect -1020 -3115 -986 -3111
rect -1020 -3187 -986 -3179
rect -1020 -3259 -986 -3247
rect -1020 -3331 -986 -3315
rect -1020 -3403 -986 -3383
rect -1020 -3475 -986 -3451
rect -1020 -3547 -986 -3519
rect -1020 -3619 -986 -3587
rect -1020 -3689 -986 -3655
rect -1020 -3757 -986 -3725
rect -1020 -3825 -986 -3797
rect -1020 -3893 -986 -3869
rect -1020 -3961 -986 -3941
rect -1020 -4029 -986 -4013
rect -1020 -4097 -986 -4085
rect -1020 -4165 -986 -4157
rect -1020 -4233 -986 -4229
rect -1020 -4339 -986 -4335
rect -1020 -4411 -986 -4403
rect -1020 -4483 -986 -4471
rect -1020 -4555 -986 -4539
rect -1020 -4627 -986 -4607
rect -1020 -4699 -986 -4675
rect -1020 -4771 -986 -4743
rect -1020 -4843 -986 -4811
rect -1020 -4913 -986 -4879
rect -1020 -4981 -986 -4949
rect -1020 -5049 -986 -5021
rect -1020 -5117 -986 -5093
rect -1020 -5185 -986 -5165
rect -1020 -5253 -986 -5237
rect -1020 -5321 -986 -5309
rect -1020 -5389 -986 -5381
rect -1020 -5457 -986 -5453
rect -1020 -5563 -986 -5559
rect -1020 -5635 -986 -5627
rect -1020 -5707 -986 -5695
rect -1020 -5779 -986 -5763
rect -1020 -5851 -986 -5831
rect -1020 -5923 -986 -5899
rect -1020 -5995 -986 -5967
rect -1020 -6067 -986 -6035
rect -1020 -6137 -986 -6103
rect -1020 -6205 -986 -6173
rect -1020 -6273 -986 -6245
rect -1020 -6341 -986 -6317
rect -1020 -6409 -986 -6389
rect -1020 -6477 -986 -6461
rect -1020 -6545 -986 -6533
rect -1020 -6613 -986 -6605
rect -1020 -6681 -986 -6677
rect -1020 -6787 -986 -6783
rect -1020 -6859 -986 -6851
rect -1020 -6931 -986 -6919
rect -1020 -7003 -986 -6987
rect -1020 -7075 -986 -7055
rect -1020 -7147 -986 -7123
rect -1020 -7219 -986 -7191
rect -1020 -7291 -986 -7259
rect -1020 -7361 -986 -7327
rect -1020 -7429 -986 -7397
rect -1020 -7497 -986 -7469
rect -1020 -7565 -986 -7541
rect -1020 -7633 -986 -7613
rect -1020 -7701 -986 -7685
rect -1020 -7769 -986 -7757
rect -1020 -7837 -986 -7829
rect -1020 -7905 -986 -7901
rect -1020 -8011 -986 -8007
rect -1020 -8083 -986 -8075
rect -1020 -8155 -986 -8143
rect -1020 -8227 -986 -8211
rect -1020 -8299 -986 -8279
rect -1020 -8371 -986 -8347
rect -1020 -8443 -986 -8415
rect -1020 -8515 -986 -8483
rect -1020 -8585 -986 -8551
rect -1020 -8653 -986 -8621
rect -1020 -8721 -986 -8693
rect -1020 -8789 -986 -8765
rect -1020 -8857 -986 -8837
rect -1020 -8925 -986 -8909
rect -1020 -8993 -986 -8981
rect -1020 -9061 -986 -9053
rect -1020 -9129 -986 -9125
rect -1020 -9235 -986 -9231
rect -1020 -9307 -986 -9299
rect -1020 -9379 -986 -9367
rect -1020 -9451 -986 -9435
rect -1020 -9523 -986 -9503
rect -1020 -9604 -986 -9571
rect -902 9571 -868 9604
rect -902 9503 -868 9523
rect -902 9435 -868 9451
rect -902 9367 -868 9379
rect -902 9299 -868 9307
rect -902 9231 -868 9235
rect -902 9125 -868 9129
rect -902 9053 -868 9061
rect -902 8981 -868 8993
rect -902 8909 -868 8925
rect -902 8837 -868 8857
rect -902 8765 -868 8789
rect -902 8693 -868 8721
rect -902 8621 -868 8653
rect -902 8551 -868 8585
rect -902 8483 -868 8515
rect -902 8415 -868 8443
rect -902 8347 -868 8371
rect -902 8279 -868 8299
rect -902 8211 -868 8227
rect -902 8143 -868 8155
rect -902 8075 -868 8083
rect -902 8007 -868 8011
rect -902 7901 -868 7905
rect -902 7829 -868 7837
rect -902 7757 -868 7769
rect -902 7685 -868 7701
rect -902 7613 -868 7633
rect -902 7541 -868 7565
rect -902 7469 -868 7497
rect -902 7397 -868 7429
rect -902 7327 -868 7361
rect -902 7259 -868 7291
rect -902 7191 -868 7219
rect -902 7123 -868 7147
rect -902 7055 -868 7075
rect -902 6987 -868 7003
rect -902 6919 -868 6931
rect -902 6851 -868 6859
rect -902 6783 -868 6787
rect -902 6677 -868 6681
rect -902 6605 -868 6613
rect -902 6533 -868 6545
rect -902 6461 -868 6477
rect -902 6389 -868 6409
rect -902 6317 -868 6341
rect -902 6245 -868 6273
rect -902 6173 -868 6205
rect -902 6103 -868 6137
rect -902 6035 -868 6067
rect -902 5967 -868 5995
rect -902 5899 -868 5923
rect -902 5831 -868 5851
rect -902 5763 -868 5779
rect -902 5695 -868 5707
rect -902 5627 -868 5635
rect -902 5559 -868 5563
rect -902 5453 -868 5457
rect -902 5381 -868 5389
rect -902 5309 -868 5321
rect -902 5237 -868 5253
rect -902 5165 -868 5185
rect -902 5093 -868 5117
rect -902 5021 -868 5049
rect -902 4949 -868 4981
rect -902 4879 -868 4913
rect -902 4811 -868 4843
rect -902 4743 -868 4771
rect -902 4675 -868 4699
rect -902 4607 -868 4627
rect -902 4539 -868 4555
rect -902 4471 -868 4483
rect -902 4403 -868 4411
rect -902 4335 -868 4339
rect -902 4229 -868 4233
rect -902 4157 -868 4165
rect -902 4085 -868 4097
rect -902 4013 -868 4029
rect -902 3941 -868 3961
rect -902 3869 -868 3893
rect -902 3797 -868 3825
rect -902 3725 -868 3757
rect -902 3655 -868 3689
rect -902 3587 -868 3619
rect -902 3519 -868 3547
rect -902 3451 -868 3475
rect -902 3383 -868 3403
rect -902 3315 -868 3331
rect -902 3247 -868 3259
rect -902 3179 -868 3187
rect -902 3111 -868 3115
rect -902 3005 -868 3009
rect -902 2933 -868 2941
rect -902 2861 -868 2873
rect -902 2789 -868 2805
rect -902 2717 -868 2737
rect -902 2645 -868 2669
rect -902 2573 -868 2601
rect -902 2501 -868 2533
rect -902 2431 -868 2465
rect -902 2363 -868 2395
rect -902 2295 -868 2323
rect -902 2227 -868 2251
rect -902 2159 -868 2179
rect -902 2091 -868 2107
rect -902 2023 -868 2035
rect -902 1955 -868 1963
rect -902 1887 -868 1891
rect -902 1781 -868 1785
rect -902 1709 -868 1717
rect -902 1637 -868 1649
rect -902 1565 -868 1581
rect -902 1493 -868 1513
rect -902 1421 -868 1445
rect -902 1349 -868 1377
rect -902 1277 -868 1309
rect -902 1207 -868 1241
rect -902 1139 -868 1171
rect -902 1071 -868 1099
rect -902 1003 -868 1027
rect -902 935 -868 955
rect -902 867 -868 883
rect -902 799 -868 811
rect -902 731 -868 739
rect -902 663 -868 667
rect -902 557 -868 561
rect -902 485 -868 493
rect -902 413 -868 425
rect -902 341 -868 357
rect -902 269 -868 289
rect -902 197 -868 221
rect -902 125 -868 153
rect -902 53 -868 85
rect -902 -17 -868 17
rect -902 -85 -868 -53
rect -902 -153 -868 -125
rect -902 -221 -868 -197
rect -902 -289 -868 -269
rect -902 -357 -868 -341
rect -902 -425 -868 -413
rect -902 -493 -868 -485
rect -902 -561 -868 -557
rect -902 -667 -868 -663
rect -902 -739 -868 -731
rect -902 -811 -868 -799
rect -902 -883 -868 -867
rect -902 -955 -868 -935
rect -902 -1027 -868 -1003
rect -902 -1099 -868 -1071
rect -902 -1171 -868 -1139
rect -902 -1241 -868 -1207
rect -902 -1309 -868 -1277
rect -902 -1377 -868 -1349
rect -902 -1445 -868 -1421
rect -902 -1513 -868 -1493
rect -902 -1581 -868 -1565
rect -902 -1649 -868 -1637
rect -902 -1717 -868 -1709
rect -902 -1785 -868 -1781
rect -902 -1891 -868 -1887
rect -902 -1963 -868 -1955
rect -902 -2035 -868 -2023
rect -902 -2107 -868 -2091
rect -902 -2179 -868 -2159
rect -902 -2251 -868 -2227
rect -902 -2323 -868 -2295
rect -902 -2395 -868 -2363
rect -902 -2465 -868 -2431
rect -902 -2533 -868 -2501
rect -902 -2601 -868 -2573
rect -902 -2669 -868 -2645
rect -902 -2737 -868 -2717
rect -902 -2805 -868 -2789
rect -902 -2873 -868 -2861
rect -902 -2941 -868 -2933
rect -902 -3009 -868 -3005
rect -902 -3115 -868 -3111
rect -902 -3187 -868 -3179
rect -902 -3259 -868 -3247
rect -902 -3331 -868 -3315
rect -902 -3403 -868 -3383
rect -902 -3475 -868 -3451
rect -902 -3547 -868 -3519
rect -902 -3619 -868 -3587
rect -902 -3689 -868 -3655
rect -902 -3757 -868 -3725
rect -902 -3825 -868 -3797
rect -902 -3893 -868 -3869
rect -902 -3961 -868 -3941
rect -902 -4029 -868 -4013
rect -902 -4097 -868 -4085
rect -902 -4165 -868 -4157
rect -902 -4233 -868 -4229
rect -902 -4339 -868 -4335
rect -902 -4411 -868 -4403
rect -902 -4483 -868 -4471
rect -902 -4555 -868 -4539
rect -902 -4627 -868 -4607
rect -902 -4699 -868 -4675
rect -902 -4771 -868 -4743
rect -902 -4843 -868 -4811
rect -902 -4913 -868 -4879
rect -902 -4981 -868 -4949
rect -902 -5049 -868 -5021
rect -902 -5117 -868 -5093
rect -902 -5185 -868 -5165
rect -902 -5253 -868 -5237
rect -902 -5321 -868 -5309
rect -902 -5389 -868 -5381
rect -902 -5457 -868 -5453
rect -902 -5563 -868 -5559
rect -902 -5635 -868 -5627
rect -902 -5707 -868 -5695
rect -902 -5779 -868 -5763
rect -902 -5851 -868 -5831
rect -902 -5923 -868 -5899
rect -902 -5995 -868 -5967
rect -902 -6067 -868 -6035
rect -902 -6137 -868 -6103
rect -902 -6205 -868 -6173
rect -902 -6273 -868 -6245
rect -902 -6341 -868 -6317
rect -902 -6409 -868 -6389
rect -902 -6477 -868 -6461
rect -902 -6545 -868 -6533
rect -902 -6613 -868 -6605
rect -902 -6681 -868 -6677
rect -902 -6787 -868 -6783
rect -902 -6859 -868 -6851
rect -902 -6931 -868 -6919
rect -902 -7003 -868 -6987
rect -902 -7075 -868 -7055
rect -902 -7147 -868 -7123
rect -902 -7219 -868 -7191
rect -902 -7291 -868 -7259
rect -902 -7361 -868 -7327
rect -902 -7429 -868 -7397
rect -902 -7497 -868 -7469
rect -902 -7565 -868 -7541
rect -902 -7633 -868 -7613
rect -902 -7701 -868 -7685
rect -902 -7769 -868 -7757
rect -902 -7837 -868 -7829
rect -902 -7905 -868 -7901
rect -902 -8011 -868 -8007
rect -902 -8083 -868 -8075
rect -902 -8155 -868 -8143
rect -902 -8227 -868 -8211
rect -902 -8299 -868 -8279
rect -902 -8371 -868 -8347
rect -902 -8443 -868 -8415
rect -902 -8515 -868 -8483
rect -902 -8585 -868 -8551
rect -902 -8653 -868 -8621
rect -902 -8721 -868 -8693
rect -902 -8789 -868 -8765
rect -902 -8857 -868 -8837
rect -902 -8925 -868 -8909
rect -902 -8993 -868 -8981
rect -902 -9061 -868 -9053
rect -902 -9129 -868 -9125
rect -902 -9235 -868 -9231
rect -902 -9307 -868 -9299
rect -902 -9379 -868 -9367
rect -902 -9451 -868 -9435
rect -902 -9523 -868 -9503
rect -902 -9604 -868 -9571
rect -784 9571 -750 9604
rect -784 9503 -750 9523
rect -784 9435 -750 9451
rect -784 9367 -750 9379
rect -784 9299 -750 9307
rect -784 9231 -750 9235
rect -784 9125 -750 9129
rect -784 9053 -750 9061
rect -784 8981 -750 8993
rect -784 8909 -750 8925
rect -784 8837 -750 8857
rect -784 8765 -750 8789
rect -784 8693 -750 8721
rect -784 8621 -750 8653
rect -784 8551 -750 8585
rect -784 8483 -750 8515
rect -784 8415 -750 8443
rect -784 8347 -750 8371
rect -784 8279 -750 8299
rect -784 8211 -750 8227
rect -784 8143 -750 8155
rect -784 8075 -750 8083
rect -784 8007 -750 8011
rect -784 7901 -750 7905
rect -784 7829 -750 7837
rect -784 7757 -750 7769
rect -784 7685 -750 7701
rect -784 7613 -750 7633
rect -784 7541 -750 7565
rect -784 7469 -750 7497
rect -784 7397 -750 7429
rect -784 7327 -750 7361
rect -784 7259 -750 7291
rect -784 7191 -750 7219
rect -784 7123 -750 7147
rect -784 7055 -750 7075
rect -784 6987 -750 7003
rect -784 6919 -750 6931
rect -784 6851 -750 6859
rect -784 6783 -750 6787
rect -784 6677 -750 6681
rect -784 6605 -750 6613
rect -784 6533 -750 6545
rect -784 6461 -750 6477
rect -784 6389 -750 6409
rect -784 6317 -750 6341
rect -784 6245 -750 6273
rect -784 6173 -750 6205
rect -784 6103 -750 6137
rect -784 6035 -750 6067
rect -784 5967 -750 5995
rect -784 5899 -750 5923
rect -784 5831 -750 5851
rect -784 5763 -750 5779
rect -784 5695 -750 5707
rect -784 5627 -750 5635
rect -784 5559 -750 5563
rect -784 5453 -750 5457
rect -784 5381 -750 5389
rect -784 5309 -750 5321
rect -784 5237 -750 5253
rect -784 5165 -750 5185
rect -784 5093 -750 5117
rect -784 5021 -750 5049
rect -784 4949 -750 4981
rect -784 4879 -750 4913
rect -784 4811 -750 4843
rect -784 4743 -750 4771
rect -784 4675 -750 4699
rect -784 4607 -750 4627
rect -784 4539 -750 4555
rect -784 4471 -750 4483
rect -784 4403 -750 4411
rect -784 4335 -750 4339
rect -784 4229 -750 4233
rect -784 4157 -750 4165
rect -784 4085 -750 4097
rect -784 4013 -750 4029
rect -784 3941 -750 3961
rect -784 3869 -750 3893
rect -784 3797 -750 3825
rect -784 3725 -750 3757
rect -784 3655 -750 3689
rect -784 3587 -750 3619
rect -784 3519 -750 3547
rect -784 3451 -750 3475
rect -784 3383 -750 3403
rect -784 3315 -750 3331
rect -784 3247 -750 3259
rect -784 3179 -750 3187
rect -784 3111 -750 3115
rect -784 3005 -750 3009
rect -784 2933 -750 2941
rect -784 2861 -750 2873
rect -784 2789 -750 2805
rect -784 2717 -750 2737
rect -784 2645 -750 2669
rect -784 2573 -750 2601
rect -784 2501 -750 2533
rect -784 2431 -750 2465
rect -784 2363 -750 2395
rect -784 2295 -750 2323
rect -784 2227 -750 2251
rect -784 2159 -750 2179
rect -784 2091 -750 2107
rect -784 2023 -750 2035
rect -784 1955 -750 1963
rect -784 1887 -750 1891
rect -784 1781 -750 1785
rect -784 1709 -750 1717
rect -784 1637 -750 1649
rect -784 1565 -750 1581
rect -784 1493 -750 1513
rect -784 1421 -750 1445
rect -784 1349 -750 1377
rect -784 1277 -750 1309
rect -784 1207 -750 1241
rect -784 1139 -750 1171
rect -784 1071 -750 1099
rect -784 1003 -750 1027
rect -784 935 -750 955
rect -784 867 -750 883
rect -784 799 -750 811
rect -784 731 -750 739
rect -784 663 -750 667
rect -784 557 -750 561
rect -784 485 -750 493
rect -784 413 -750 425
rect -784 341 -750 357
rect -784 269 -750 289
rect -784 197 -750 221
rect -784 125 -750 153
rect -784 53 -750 85
rect -784 -17 -750 17
rect -784 -85 -750 -53
rect -784 -153 -750 -125
rect -784 -221 -750 -197
rect -784 -289 -750 -269
rect -784 -357 -750 -341
rect -784 -425 -750 -413
rect -784 -493 -750 -485
rect -784 -561 -750 -557
rect -784 -667 -750 -663
rect -784 -739 -750 -731
rect -784 -811 -750 -799
rect -784 -883 -750 -867
rect -784 -955 -750 -935
rect -784 -1027 -750 -1003
rect -784 -1099 -750 -1071
rect -784 -1171 -750 -1139
rect -784 -1241 -750 -1207
rect -784 -1309 -750 -1277
rect -784 -1377 -750 -1349
rect -784 -1445 -750 -1421
rect -784 -1513 -750 -1493
rect -784 -1581 -750 -1565
rect -784 -1649 -750 -1637
rect -784 -1717 -750 -1709
rect -784 -1785 -750 -1781
rect -784 -1891 -750 -1887
rect -784 -1963 -750 -1955
rect -784 -2035 -750 -2023
rect -784 -2107 -750 -2091
rect -784 -2179 -750 -2159
rect -784 -2251 -750 -2227
rect -784 -2323 -750 -2295
rect -784 -2395 -750 -2363
rect -784 -2465 -750 -2431
rect -784 -2533 -750 -2501
rect -784 -2601 -750 -2573
rect -784 -2669 -750 -2645
rect -784 -2737 -750 -2717
rect -784 -2805 -750 -2789
rect -784 -2873 -750 -2861
rect -784 -2941 -750 -2933
rect -784 -3009 -750 -3005
rect -784 -3115 -750 -3111
rect -784 -3187 -750 -3179
rect -784 -3259 -750 -3247
rect -784 -3331 -750 -3315
rect -784 -3403 -750 -3383
rect -784 -3475 -750 -3451
rect -784 -3547 -750 -3519
rect -784 -3619 -750 -3587
rect -784 -3689 -750 -3655
rect -784 -3757 -750 -3725
rect -784 -3825 -750 -3797
rect -784 -3893 -750 -3869
rect -784 -3961 -750 -3941
rect -784 -4029 -750 -4013
rect -784 -4097 -750 -4085
rect -784 -4165 -750 -4157
rect -784 -4233 -750 -4229
rect -784 -4339 -750 -4335
rect -784 -4411 -750 -4403
rect -784 -4483 -750 -4471
rect -784 -4555 -750 -4539
rect -784 -4627 -750 -4607
rect -784 -4699 -750 -4675
rect -784 -4771 -750 -4743
rect -784 -4843 -750 -4811
rect -784 -4913 -750 -4879
rect -784 -4981 -750 -4949
rect -784 -5049 -750 -5021
rect -784 -5117 -750 -5093
rect -784 -5185 -750 -5165
rect -784 -5253 -750 -5237
rect -784 -5321 -750 -5309
rect -784 -5389 -750 -5381
rect -784 -5457 -750 -5453
rect -784 -5563 -750 -5559
rect -784 -5635 -750 -5627
rect -784 -5707 -750 -5695
rect -784 -5779 -750 -5763
rect -784 -5851 -750 -5831
rect -784 -5923 -750 -5899
rect -784 -5995 -750 -5967
rect -784 -6067 -750 -6035
rect -784 -6137 -750 -6103
rect -784 -6205 -750 -6173
rect -784 -6273 -750 -6245
rect -784 -6341 -750 -6317
rect -784 -6409 -750 -6389
rect -784 -6477 -750 -6461
rect -784 -6545 -750 -6533
rect -784 -6613 -750 -6605
rect -784 -6681 -750 -6677
rect -784 -6787 -750 -6783
rect -784 -6859 -750 -6851
rect -784 -6931 -750 -6919
rect -784 -7003 -750 -6987
rect -784 -7075 -750 -7055
rect -784 -7147 -750 -7123
rect -784 -7219 -750 -7191
rect -784 -7291 -750 -7259
rect -784 -7361 -750 -7327
rect -784 -7429 -750 -7397
rect -784 -7497 -750 -7469
rect -784 -7565 -750 -7541
rect -784 -7633 -750 -7613
rect -784 -7701 -750 -7685
rect -784 -7769 -750 -7757
rect -784 -7837 -750 -7829
rect -784 -7905 -750 -7901
rect -784 -8011 -750 -8007
rect -784 -8083 -750 -8075
rect -784 -8155 -750 -8143
rect -784 -8227 -750 -8211
rect -784 -8299 -750 -8279
rect -784 -8371 -750 -8347
rect -784 -8443 -750 -8415
rect -784 -8515 -750 -8483
rect -784 -8585 -750 -8551
rect -784 -8653 -750 -8621
rect -784 -8721 -750 -8693
rect -784 -8789 -750 -8765
rect -784 -8857 -750 -8837
rect -784 -8925 -750 -8909
rect -784 -8993 -750 -8981
rect -784 -9061 -750 -9053
rect -784 -9129 -750 -9125
rect -784 -9235 -750 -9231
rect -784 -9307 -750 -9299
rect -784 -9379 -750 -9367
rect -784 -9451 -750 -9435
rect -784 -9523 -750 -9503
rect -784 -9604 -750 -9571
rect -666 9571 -632 9604
rect -666 9503 -632 9523
rect -666 9435 -632 9451
rect -666 9367 -632 9379
rect -666 9299 -632 9307
rect -666 9231 -632 9235
rect -666 9125 -632 9129
rect -666 9053 -632 9061
rect -666 8981 -632 8993
rect -666 8909 -632 8925
rect -666 8837 -632 8857
rect -666 8765 -632 8789
rect -666 8693 -632 8721
rect -666 8621 -632 8653
rect -666 8551 -632 8585
rect -666 8483 -632 8515
rect -666 8415 -632 8443
rect -666 8347 -632 8371
rect -666 8279 -632 8299
rect -666 8211 -632 8227
rect -666 8143 -632 8155
rect -666 8075 -632 8083
rect -666 8007 -632 8011
rect -666 7901 -632 7905
rect -666 7829 -632 7837
rect -666 7757 -632 7769
rect -666 7685 -632 7701
rect -666 7613 -632 7633
rect -666 7541 -632 7565
rect -666 7469 -632 7497
rect -666 7397 -632 7429
rect -666 7327 -632 7361
rect -666 7259 -632 7291
rect -666 7191 -632 7219
rect -666 7123 -632 7147
rect -666 7055 -632 7075
rect -666 6987 -632 7003
rect -666 6919 -632 6931
rect -666 6851 -632 6859
rect -666 6783 -632 6787
rect -666 6677 -632 6681
rect -666 6605 -632 6613
rect -666 6533 -632 6545
rect -666 6461 -632 6477
rect -666 6389 -632 6409
rect -666 6317 -632 6341
rect -666 6245 -632 6273
rect -666 6173 -632 6205
rect -666 6103 -632 6137
rect -666 6035 -632 6067
rect -666 5967 -632 5995
rect -666 5899 -632 5923
rect -666 5831 -632 5851
rect -666 5763 -632 5779
rect -666 5695 -632 5707
rect -666 5627 -632 5635
rect -666 5559 -632 5563
rect -666 5453 -632 5457
rect -666 5381 -632 5389
rect -666 5309 -632 5321
rect -666 5237 -632 5253
rect -666 5165 -632 5185
rect -666 5093 -632 5117
rect -666 5021 -632 5049
rect -666 4949 -632 4981
rect -666 4879 -632 4913
rect -666 4811 -632 4843
rect -666 4743 -632 4771
rect -666 4675 -632 4699
rect -666 4607 -632 4627
rect -666 4539 -632 4555
rect -666 4471 -632 4483
rect -666 4403 -632 4411
rect -666 4335 -632 4339
rect -666 4229 -632 4233
rect -666 4157 -632 4165
rect -666 4085 -632 4097
rect -666 4013 -632 4029
rect -666 3941 -632 3961
rect -666 3869 -632 3893
rect -666 3797 -632 3825
rect -666 3725 -632 3757
rect -666 3655 -632 3689
rect -666 3587 -632 3619
rect -666 3519 -632 3547
rect -666 3451 -632 3475
rect -666 3383 -632 3403
rect -666 3315 -632 3331
rect -666 3247 -632 3259
rect -666 3179 -632 3187
rect -666 3111 -632 3115
rect -666 3005 -632 3009
rect -666 2933 -632 2941
rect -666 2861 -632 2873
rect -666 2789 -632 2805
rect -666 2717 -632 2737
rect -666 2645 -632 2669
rect -666 2573 -632 2601
rect -666 2501 -632 2533
rect -666 2431 -632 2465
rect -666 2363 -632 2395
rect -666 2295 -632 2323
rect -666 2227 -632 2251
rect -666 2159 -632 2179
rect -666 2091 -632 2107
rect -666 2023 -632 2035
rect -666 1955 -632 1963
rect -666 1887 -632 1891
rect -666 1781 -632 1785
rect -666 1709 -632 1717
rect -666 1637 -632 1649
rect -666 1565 -632 1581
rect -666 1493 -632 1513
rect -666 1421 -632 1445
rect -666 1349 -632 1377
rect -666 1277 -632 1309
rect -666 1207 -632 1241
rect -666 1139 -632 1171
rect -666 1071 -632 1099
rect -666 1003 -632 1027
rect -666 935 -632 955
rect -666 867 -632 883
rect -666 799 -632 811
rect -666 731 -632 739
rect -666 663 -632 667
rect -666 557 -632 561
rect -666 485 -632 493
rect -666 413 -632 425
rect -666 341 -632 357
rect -666 269 -632 289
rect -666 197 -632 221
rect -666 125 -632 153
rect -666 53 -632 85
rect -666 -17 -632 17
rect -666 -85 -632 -53
rect -666 -153 -632 -125
rect -666 -221 -632 -197
rect -666 -289 -632 -269
rect -666 -357 -632 -341
rect -666 -425 -632 -413
rect -666 -493 -632 -485
rect -666 -561 -632 -557
rect -666 -667 -632 -663
rect -666 -739 -632 -731
rect -666 -811 -632 -799
rect -666 -883 -632 -867
rect -666 -955 -632 -935
rect -666 -1027 -632 -1003
rect -666 -1099 -632 -1071
rect -666 -1171 -632 -1139
rect -666 -1241 -632 -1207
rect -666 -1309 -632 -1277
rect -666 -1377 -632 -1349
rect -666 -1445 -632 -1421
rect -666 -1513 -632 -1493
rect -666 -1581 -632 -1565
rect -666 -1649 -632 -1637
rect -666 -1717 -632 -1709
rect -666 -1785 -632 -1781
rect -666 -1891 -632 -1887
rect -666 -1963 -632 -1955
rect -666 -2035 -632 -2023
rect -666 -2107 -632 -2091
rect -666 -2179 -632 -2159
rect -666 -2251 -632 -2227
rect -666 -2323 -632 -2295
rect -666 -2395 -632 -2363
rect -666 -2465 -632 -2431
rect -666 -2533 -632 -2501
rect -666 -2601 -632 -2573
rect -666 -2669 -632 -2645
rect -666 -2737 -632 -2717
rect -666 -2805 -632 -2789
rect -666 -2873 -632 -2861
rect -666 -2941 -632 -2933
rect -666 -3009 -632 -3005
rect -666 -3115 -632 -3111
rect -666 -3187 -632 -3179
rect -666 -3259 -632 -3247
rect -666 -3331 -632 -3315
rect -666 -3403 -632 -3383
rect -666 -3475 -632 -3451
rect -666 -3547 -632 -3519
rect -666 -3619 -632 -3587
rect -666 -3689 -632 -3655
rect -666 -3757 -632 -3725
rect -666 -3825 -632 -3797
rect -666 -3893 -632 -3869
rect -666 -3961 -632 -3941
rect -666 -4029 -632 -4013
rect -666 -4097 -632 -4085
rect -666 -4165 -632 -4157
rect -666 -4233 -632 -4229
rect -666 -4339 -632 -4335
rect -666 -4411 -632 -4403
rect -666 -4483 -632 -4471
rect -666 -4555 -632 -4539
rect -666 -4627 -632 -4607
rect -666 -4699 -632 -4675
rect -666 -4771 -632 -4743
rect -666 -4843 -632 -4811
rect -666 -4913 -632 -4879
rect -666 -4981 -632 -4949
rect -666 -5049 -632 -5021
rect -666 -5117 -632 -5093
rect -666 -5185 -632 -5165
rect -666 -5253 -632 -5237
rect -666 -5321 -632 -5309
rect -666 -5389 -632 -5381
rect -666 -5457 -632 -5453
rect -666 -5563 -632 -5559
rect -666 -5635 -632 -5627
rect -666 -5707 -632 -5695
rect -666 -5779 -632 -5763
rect -666 -5851 -632 -5831
rect -666 -5923 -632 -5899
rect -666 -5995 -632 -5967
rect -666 -6067 -632 -6035
rect -666 -6137 -632 -6103
rect -666 -6205 -632 -6173
rect -666 -6273 -632 -6245
rect -666 -6341 -632 -6317
rect -666 -6409 -632 -6389
rect -666 -6477 -632 -6461
rect -666 -6545 -632 -6533
rect -666 -6613 -632 -6605
rect -666 -6681 -632 -6677
rect -666 -6787 -632 -6783
rect -666 -6859 -632 -6851
rect -666 -6931 -632 -6919
rect -666 -7003 -632 -6987
rect -666 -7075 -632 -7055
rect -666 -7147 -632 -7123
rect -666 -7219 -632 -7191
rect -666 -7291 -632 -7259
rect -666 -7361 -632 -7327
rect -666 -7429 -632 -7397
rect -666 -7497 -632 -7469
rect -666 -7565 -632 -7541
rect -666 -7633 -632 -7613
rect -666 -7701 -632 -7685
rect -666 -7769 -632 -7757
rect -666 -7837 -632 -7829
rect -666 -7905 -632 -7901
rect -666 -8011 -632 -8007
rect -666 -8083 -632 -8075
rect -666 -8155 -632 -8143
rect -666 -8227 -632 -8211
rect -666 -8299 -632 -8279
rect -666 -8371 -632 -8347
rect -666 -8443 -632 -8415
rect -666 -8515 -632 -8483
rect -666 -8585 -632 -8551
rect -666 -8653 -632 -8621
rect -666 -8721 -632 -8693
rect -666 -8789 -632 -8765
rect -666 -8857 -632 -8837
rect -666 -8925 -632 -8909
rect -666 -8993 -632 -8981
rect -666 -9061 -632 -9053
rect -666 -9129 -632 -9125
rect -666 -9235 -632 -9231
rect -666 -9307 -632 -9299
rect -666 -9379 -632 -9367
rect -666 -9451 -632 -9435
rect -666 -9523 -632 -9503
rect -666 -9604 -632 -9571
rect -548 9571 -514 9604
rect -548 9503 -514 9523
rect -548 9435 -514 9451
rect -548 9367 -514 9379
rect -548 9299 -514 9307
rect -548 9231 -514 9235
rect -548 9125 -514 9129
rect -548 9053 -514 9061
rect -548 8981 -514 8993
rect -548 8909 -514 8925
rect -548 8837 -514 8857
rect -548 8765 -514 8789
rect -548 8693 -514 8721
rect -548 8621 -514 8653
rect -548 8551 -514 8585
rect -548 8483 -514 8515
rect -548 8415 -514 8443
rect -548 8347 -514 8371
rect -548 8279 -514 8299
rect -548 8211 -514 8227
rect -548 8143 -514 8155
rect -548 8075 -514 8083
rect -548 8007 -514 8011
rect -548 7901 -514 7905
rect -548 7829 -514 7837
rect -548 7757 -514 7769
rect -548 7685 -514 7701
rect -548 7613 -514 7633
rect -548 7541 -514 7565
rect -548 7469 -514 7497
rect -548 7397 -514 7429
rect -548 7327 -514 7361
rect -548 7259 -514 7291
rect -548 7191 -514 7219
rect -548 7123 -514 7147
rect -548 7055 -514 7075
rect -548 6987 -514 7003
rect -548 6919 -514 6931
rect -548 6851 -514 6859
rect -548 6783 -514 6787
rect -548 6677 -514 6681
rect -548 6605 -514 6613
rect -548 6533 -514 6545
rect -548 6461 -514 6477
rect -548 6389 -514 6409
rect -548 6317 -514 6341
rect -548 6245 -514 6273
rect -548 6173 -514 6205
rect -548 6103 -514 6137
rect -548 6035 -514 6067
rect -548 5967 -514 5995
rect -548 5899 -514 5923
rect -548 5831 -514 5851
rect -548 5763 -514 5779
rect -548 5695 -514 5707
rect -548 5627 -514 5635
rect -548 5559 -514 5563
rect -548 5453 -514 5457
rect -548 5381 -514 5389
rect -548 5309 -514 5321
rect -548 5237 -514 5253
rect -548 5165 -514 5185
rect -548 5093 -514 5117
rect -548 5021 -514 5049
rect -548 4949 -514 4981
rect -548 4879 -514 4913
rect -548 4811 -514 4843
rect -548 4743 -514 4771
rect -548 4675 -514 4699
rect -548 4607 -514 4627
rect -548 4539 -514 4555
rect -548 4471 -514 4483
rect -548 4403 -514 4411
rect -548 4335 -514 4339
rect -548 4229 -514 4233
rect -548 4157 -514 4165
rect -548 4085 -514 4097
rect -548 4013 -514 4029
rect -548 3941 -514 3961
rect -548 3869 -514 3893
rect -548 3797 -514 3825
rect -548 3725 -514 3757
rect -548 3655 -514 3689
rect -548 3587 -514 3619
rect -548 3519 -514 3547
rect -548 3451 -514 3475
rect -548 3383 -514 3403
rect -548 3315 -514 3331
rect -548 3247 -514 3259
rect -548 3179 -514 3187
rect -548 3111 -514 3115
rect -548 3005 -514 3009
rect -548 2933 -514 2941
rect -548 2861 -514 2873
rect -548 2789 -514 2805
rect -548 2717 -514 2737
rect -548 2645 -514 2669
rect -548 2573 -514 2601
rect -548 2501 -514 2533
rect -548 2431 -514 2465
rect -548 2363 -514 2395
rect -548 2295 -514 2323
rect -548 2227 -514 2251
rect -548 2159 -514 2179
rect -548 2091 -514 2107
rect -548 2023 -514 2035
rect -548 1955 -514 1963
rect -548 1887 -514 1891
rect -548 1781 -514 1785
rect -548 1709 -514 1717
rect -548 1637 -514 1649
rect -548 1565 -514 1581
rect -548 1493 -514 1513
rect -548 1421 -514 1445
rect -548 1349 -514 1377
rect -548 1277 -514 1309
rect -548 1207 -514 1241
rect -548 1139 -514 1171
rect -548 1071 -514 1099
rect -548 1003 -514 1027
rect -548 935 -514 955
rect -548 867 -514 883
rect -548 799 -514 811
rect -548 731 -514 739
rect -548 663 -514 667
rect -548 557 -514 561
rect -548 485 -514 493
rect -548 413 -514 425
rect -548 341 -514 357
rect -548 269 -514 289
rect -548 197 -514 221
rect -548 125 -514 153
rect -548 53 -514 85
rect -548 -17 -514 17
rect -548 -85 -514 -53
rect -548 -153 -514 -125
rect -548 -221 -514 -197
rect -548 -289 -514 -269
rect -548 -357 -514 -341
rect -548 -425 -514 -413
rect -548 -493 -514 -485
rect -548 -561 -514 -557
rect -548 -667 -514 -663
rect -548 -739 -514 -731
rect -548 -811 -514 -799
rect -548 -883 -514 -867
rect -548 -955 -514 -935
rect -548 -1027 -514 -1003
rect -548 -1099 -514 -1071
rect -548 -1171 -514 -1139
rect -548 -1241 -514 -1207
rect -548 -1309 -514 -1277
rect -548 -1377 -514 -1349
rect -548 -1445 -514 -1421
rect -548 -1513 -514 -1493
rect -548 -1581 -514 -1565
rect -548 -1649 -514 -1637
rect -548 -1717 -514 -1709
rect -548 -1785 -514 -1781
rect -548 -1891 -514 -1887
rect -548 -1963 -514 -1955
rect -548 -2035 -514 -2023
rect -548 -2107 -514 -2091
rect -548 -2179 -514 -2159
rect -548 -2251 -514 -2227
rect -548 -2323 -514 -2295
rect -548 -2395 -514 -2363
rect -548 -2465 -514 -2431
rect -548 -2533 -514 -2501
rect -548 -2601 -514 -2573
rect -548 -2669 -514 -2645
rect -548 -2737 -514 -2717
rect -548 -2805 -514 -2789
rect -548 -2873 -514 -2861
rect -548 -2941 -514 -2933
rect -548 -3009 -514 -3005
rect -548 -3115 -514 -3111
rect -548 -3187 -514 -3179
rect -548 -3259 -514 -3247
rect -548 -3331 -514 -3315
rect -548 -3403 -514 -3383
rect -548 -3475 -514 -3451
rect -548 -3547 -514 -3519
rect -548 -3619 -514 -3587
rect -548 -3689 -514 -3655
rect -548 -3757 -514 -3725
rect -548 -3825 -514 -3797
rect -548 -3893 -514 -3869
rect -548 -3961 -514 -3941
rect -548 -4029 -514 -4013
rect -548 -4097 -514 -4085
rect -548 -4165 -514 -4157
rect -548 -4233 -514 -4229
rect -548 -4339 -514 -4335
rect -548 -4411 -514 -4403
rect -548 -4483 -514 -4471
rect -548 -4555 -514 -4539
rect -548 -4627 -514 -4607
rect -548 -4699 -514 -4675
rect -548 -4771 -514 -4743
rect -548 -4843 -514 -4811
rect -548 -4913 -514 -4879
rect -548 -4981 -514 -4949
rect -548 -5049 -514 -5021
rect -548 -5117 -514 -5093
rect -548 -5185 -514 -5165
rect -548 -5253 -514 -5237
rect -548 -5321 -514 -5309
rect -548 -5389 -514 -5381
rect -548 -5457 -514 -5453
rect -548 -5563 -514 -5559
rect -548 -5635 -514 -5627
rect -548 -5707 -514 -5695
rect -548 -5779 -514 -5763
rect -548 -5851 -514 -5831
rect -548 -5923 -514 -5899
rect -548 -5995 -514 -5967
rect -548 -6067 -514 -6035
rect -548 -6137 -514 -6103
rect -548 -6205 -514 -6173
rect -548 -6273 -514 -6245
rect -548 -6341 -514 -6317
rect -548 -6409 -514 -6389
rect -548 -6477 -514 -6461
rect -548 -6545 -514 -6533
rect -548 -6613 -514 -6605
rect -548 -6681 -514 -6677
rect -548 -6787 -514 -6783
rect -548 -6859 -514 -6851
rect -548 -6931 -514 -6919
rect -548 -7003 -514 -6987
rect -548 -7075 -514 -7055
rect -548 -7147 -514 -7123
rect -548 -7219 -514 -7191
rect -548 -7291 -514 -7259
rect -548 -7361 -514 -7327
rect -548 -7429 -514 -7397
rect -548 -7497 -514 -7469
rect -548 -7565 -514 -7541
rect -548 -7633 -514 -7613
rect -548 -7701 -514 -7685
rect -548 -7769 -514 -7757
rect -548 -7837 -514 -7829
rect -548 -7905 -514 -7901
rect -548 -8011 -514 -8007
rect -548 -8083 -514 -8075
rect -548 -8155 -514 -8143
rect -548 -8227 -514 -8211
rect -548 -8299 -514 -8279
rect -548 -8371 -514 -8347
rect -548 -8443 -514 -8415
rect -548 -8515 -514 -8483
rect -548 -8585 -514 -8551
rect -548 -8653 -514 -8621
rect -548 -8721 -514 -8693
rect -548 -8789 -514 -8765
rect -548 -8857 -514 -8837
rect -548 -8925 -514 -8909
rect -548 -8993 -514 -8981
rect -548 -9061 -514 -9053
rect -548 -9129 -514 -9125
rect -548 -9235 -514 -9231
rect -548 -9307 -514 -9299
rect -548 -9379 -514 -9367
rect -548 -9451 -514 -9435
rect -548 -9523 -514 -9503
rect -548 -9604 -514 -9571
rect -430 9571 -396 9604
rect -430 9503 -396 9523
rect -430 9435 -396 9451
rect -430 9367 -396 9379
rect -430 9299 -396 9307
rect -430 9231 -396 9235
rect -430 9125 -396 9129
rect -430 9053 -396 9061
rect -430 8981 -396 8993
rect -430 8909 -396 8925
rect -430 8837 -396 8857
rect -430 8765 -396 8789
rect -430 8693 -396 8721
rect -430 8621 -396 8653
rect -430 8551 -396 8585
rect -430 8483 -396 8515
rect -430 8415 -396 8443
rect -430 8347 -396 8371
rect -430 8279 -396 8299
rect -430 8211 -396 8227
rect -430 8143 -396 8155
rect -430 8075 -396 8083
rect -430 8007 -396 8011
rect -430 7901 -396 7905
rect -430 7829 -396 7837
rect -430 7757 -396 7769
rect -430 7685 -396 7701
rect -430 7613 -396 7633
rect -430 7541 -396 7565
rect -430 7469 -396 7497
rect -430 7397 -396 7429
rect -430 7327 -396 7361
rect -430 7259 -396 7291
rect -430 7191 -396 7219
rect -430 7123 -396 7147
rect -430 7055 -396 7075
rect -430 6987 -396 7003
rect -430 6919 -396 6931
rect -430 6851 -396 6859
rect -430 6783 -396 6787
rect -430 6677 -396 6681
rect -430 6605 -396 6613
rect -430 6533 -396 6545
rect -430 6461 -396 6477
rect -430 6389 -396 6409
rect -430 6317 -396 6341
rect -430 6245 -396 6273
rect -430 6173 -396 6205
rect -430 6103 -396 6137
rect -430 6035 -396 6067
rect -430 5967 -396 5995
rect -430 5899 -396 5923
rect -430 5831 -396 5851
rect -430 5763 -396 5779
rect -430 5695 -396 5707
rect -430 5627 -396 5635
rect -430 5559 -396 5563
rect -430 5453 -396 5457
rect -430 5381 -396 5389
rect -430 5309 -396 5321
rect -430 5237 -396 5253
rect -430 5165 -396 5185
rect -430 5093 -396 5117
rect -430 5021 -396 5049
rect -430 4949 -396 4981
rect -430 4879 -396 4913
rect -430 4811 -396 4843
rect -430 4743 -396 4771
rect -430 4675 -396 4699
rect -430 4607 -396 4627
rect -430 4539 -396 4555
rect -430 4471 -396 4483
rect -430 4403 -396 4411
rect -430 4335 -396 4339
rect -430 4229 -396 4233
rect -430 4157 -396 4165
rect -430 4085 -396 4097
rect -430 4013 -396 4029
rect -430 3941 -396 3961
rect -430 3869 -396 3893
rect -430 3797 -396 3825
rect -430 3725 -396 3757
rect -430 3655 -396 3689
rect -430 3587 -396 3619
rect -430 3519 -396 3547
rect -430 3451 -396 3475
rect -430 3383 -396 3403
rect -430 3315 -396 3331
rect -430 3247 -396 3259
rect -430 3179 -396 3187
rect -430 3111 -396 3115
rect -430 3005 -396 3009
rect -430 2933 -396 2941
rect -430 2861 -396 2873
rect -430 2789 -396 2805
rect -430 2717 -396 2737
rect -430 2645 -396 2669
rect -430 2573 -396 2601
rect -430 2501 -396 2533
rect -430 2431 -396 2465
rect -430 2363 -396 2395
rect -430 2295 -396 2323
rect -430 2227 -396 2251
rect -430 2159 -396 2179
rect -430 2091 -396 2107
rect -430 2023 -396 2035
rect -430 1955 -396 1963
rect -430 1887 -396 1891
rect -430 1781 -396 1785
rect -430 1709 -396 1717
rect -430 1637 -396 1649
rect -430 1565 -396 1581
rect -430 1493 -396 1513
rect -430 1421 -396 1445
rect -430 1349 -396 1377
rect -430 1277 -396 1309
rect -430 1207 -396 1241
rect -430 1139 -396 1171
rect -430 1071 -396 1099
rect -430 1003 -396 1027
rect -430 935 -396 955
rect -430 867 -396 883
rect -430 799 -396 811
rect -430 731 -396 739
rect -430 663 -396 667
rect -430 557 -396 561
rect -430 485 -396 493
rect -430 413 -396 425
rect -430 341 -396 357
rect -430 269 -396 289
rect -430 197 -396 221
rect -430 125 -396 153
rect -430 53 -396 85
rect -430 -17 -396 17
rect -430 -85 -396 -53
rect -430 -153 -396 -125
rect -430 -221 -396 -197
rect -430 -289 -396 -269
rect -430 -357 -396 -341
rect -430 -425 -396 -413
rect -430 -493 -396 -485
rect -430 -561 -396 -557
rect -430 -667 -396 -663
rect -430 -739 -396 -731
rect -430 -811 -396 -799
rect -430 -883 -396 -867
rect -430 -955 -396 -935
rect -430 -1027 -396 -1003
rect -430 -1099 -396 -1071
rect -430 -1171 -396 -1139
rect -430 -1241 -396 -1207
rect -430 -1309 -396 -1277
rect -430 -1377 -396 -1349
rect -430 -1445 -396 -1421
rect -430 -1513 -396 -1493
rect -430 -1581 -396 -1565
rect -430 -1649 -396 -1637
rect -430 -1717 -396 -1709
rect -430 -1785 -396 -1781
rect -430 -1891 -396 -1887
rect -430 -1963 -396 -1955
rect -430 -2035 -396 -2023
rect -430 -2107 -396 -2091
rect -430 -2179 -396 -2159
rect -430 -2251 -396 -2227
rect -430 -2323 -396 -2295
rect -430 -2395 -396 -2363
rect -430 -2465 -396 -2431
rect -430 -2533 -396 -2501
rect -430 -2601 -396 -2573
rect -430 -2669 -396 -2645
rect -430 -2737 -396 -2717
rect -430 -2805 -396 -2789
rect -430 -2873 -396 -2861
rect -430 -2941 -396 -2933
rect -430 -3009 -396 -3005
rect -430 -3115 -396 -3111
rect -430 -3187 -396 -3179
rect -430 -3259 -396 -3247
rect -430 -3331 -396 -3315
rect -430 -3403 -396 -3383
rect -430 -3475 -396 -3451
rect -430 -3547 -396 -3519
rect -430 -3619 -396 -3587
rect -430 -3689 -396 -3655
rect -430 -3757 -396 -3725
rect -430 -3825 -396 -3797
rect -430 -3893 -396 -3869
rect -430 -3961 -396 -3941
rect -430 -4029 -396 -4013
rect -430 -4097 -396 -4085
rect -430 -4165 -396 -4157
rect -430 -4233 -396 -4229
rect -430 -4339 -396 -4335
rect -430 -4411 -396 -4403
rect -430 -4483 -396 -4471
rect -430 -4555 -396 -4539
rect -430 -4627 -396 -4607
rect -430 -4699 -396 -4675
rect -430 -4771 -396 -4743
rect -430 -4843 -396 -4811
rect -430 -4913 -396 -4879
rect -430 -4981 -396 -4949
rect -430 -5049 -396 -5021
rect -430 -5117 -396 -5093
rect -430 -5185 -396 -5165
rect -430 -5253 -396 -5237
rect -430 -5321 -396 -5309
rect -430 -5389 -396 -5381
rect -430 -5457 -396 -5453
rect -430 -5563 -396 -5559
rect -430 -5635 -396 -5627
rect -430 -5707 -396 -5695
rect -430 -5779 -396 -5763
rect -430 -5851 -396 -5831
rect -430 -5923 -396 -5899
rect -430 -5995 -396 -5967
rect -430 -6067 -396 -6035
rect -430 -6137 -396 -6103
rect -430 -6205 -396 -6173
rect -430 -6273 -396 -6245
rect -430 -6341 -396 -6317
rect -430 -6409 -396 -6389
rect -430 -6477 -396 -6461
rect -430 -6545 -396 -6533
rect -430 -6613 -396 -6605
rect -430 -6681 -396 -6677
rect -430 -6787 -396 -6783
rect -430 -6859 -396 -6851
rect -430 -6931 -396 -6919
rect -430 -7003 -396 -6987
rect -430 -7075 -396 -7055
rect -430 -7147 -396 -7123
rect -430 -7219 -396 -7191
rect -430 -7291 -396 -7259
rect -430 -7361 -396 -7327
rect -430 -7429 -396 -7397
rect -430 -7497 -396 -7469
rect -430 -7565 -396 -7541
rect -430 -7633 -396 -7613
rect -430 -7701 -396 -7685
rect -430 -7769 -396 -7757
rect -430 -7837 -396 -7829
rect -430 -7905 -396 -7901
rect -430 -8011 -396 -8007
rect -430 -8083 -396 -8075
rect -430 -8155 -396 -8143
rect -430 -8227 -396 -8211
rect -430 -8299 -396 -8279
rect -430 -8371 -396 -8347
rect -430 -8443 -396 -8415
rect -430 -8515 -396 -8483
rect -430 -8585 -396 -8551
rect -430 -8653 -396 -8621
rect -430 -8721 -396 -8693
rect -430 -8789 -396 -8765
rect -430 -8857 -396 -8837
rect -430 -8925 -396 -8909
rect -430 -8993 -396 -8981
rect -430 -9061 -396 -9053
rect -430 -9129 -396 -9125
rect -430 -9235 -396 -9231
rect -430 -9307 -396 -9299
rect -430 -9379 -396 -9367
rect -430 -9451 -396 -9435
rect -430 -9523 -396 -9503
rect -430 -9604 -396 -9571
rect -312 9571 -278 9604
rect -312 9503 -278 9523
rect -312 9435 -278 9451
rect -312 9367 -278 9379
rect -312 9299 -278 9307
rect -312 9231 -278 9235
rect -312 9125 -278 9129
rect -312 9053 -278 9061
rect -312 8981 -278 8993
rect -312 8909 -278 8925
rect -312 8837 -278 8857
rect -312 8765 -278 8789
rect -312 8693 -278 8721
rect -312 8621 -278 8653
rect -312 8551 -278 8585
rect -312 8483 -278 8515
rect -312 8415 -278 8443
rect -312 8347 -278 8371
rect -312 8279 -278 8299
rect -312 8211 -278 8227
rect -312 8143 -278 8155
rect -312 8075 -278 8083
rect -312 8007 -278 8011
rect -312 7901 -278 7905
rect -312 7829 -278 7837
rect -312 7757 -278 7769
rect -312 7685 -278 7701
rect -312 7613 -278 7633
rect -312 7541 -278 7565
rect -312 7469 -278 7497
rect -312 7397 -278 7429
rect -312 7327 -278 7361
rect -312 7259 -278 7291
rect -312 7191 -278 7219
rect -312 7123 -278 7147
rect -312 7055 -278 7075
rect -312 6987 -278 7003
rect -312 6919 -278 6931
rect -312 6851 -278 6859
rect -312 6783 -278 6787
rect -312 6677 -278 6681
rect -312 6605 -278 6613
rect -312 6533 -278 6545
rect -312 6461 -278 6477
rect -312 6389 -278 6409
rect -312 6317 -278 6341
rect -312 6245 -278 6273
rect -312 6173 -278 6205
rect -312 6103 -278 6137
rect -312 6035 -278 6067
rect -312 5967 -278 5995
rect -312 5899 -278 5923
rect -312 5831 -278 5851
rect -312 5763 -278 5779
rect -312 5695 -278 5707
rect -312 5627 -278 5635
rect -312 5559 -278 5563
rect -312 5453 -278 5457
rect -312 5381 -278 5389
rect -312 5309 -278 5321
rect -312 5237 -278 5253
rect -312 5165 -278 5185
rect -312 5093 -278 5117
rect -312 5021 -278 5049
rect -312 4949 -278 4981
rect -312 4879 -278 4913
rect -312 4811 -278 4843
rect -312 4743 -278 4771
rect -312 4675 -278 4699
rect -312 4607 -278 4627
rect -312 4539 -278 4555
rect -312 4471 -278 4483
rect -312 4403 -278 4411
rect -312 4335 -278 4339
rect -312 4229 -278 4233
rect -312 4157 -278 4165
rect -312 4085 -278 4097
rect -312 4013 -278 4029
rect -312 3941 -278 3961
rect -312 3869 -278 3893
rect -312 3797 -278 3825
rect -312 3725 -278 3757
rect -312 3655 -278 3689
rect -312 3587 -278 3619
rect -312 3519 -278 3547
rect -312 3451 -278 3475
rect -312 3383 -278 3403
rect -312 3315 -278 3331
rect -312 3247 -278 3259
rect -312 3179 -278 3187
rect -312 3111 -278 3115
rect -312 3005 -278 3009
rect -312 2933 -278 2941
rect -312 2861 -278 2873
rect -312 2789 -278 2805
rect -312 2717 -278 2737
rect -312 2645 -278 2669
rect -312 2573 -278 2601
rect -312 2501 -278 2533
rect -312 2431 -278 2465
rect -312 2363 -278 2395
rect -312 2295 -278 2323
rect -312 2227 -278 2251
rect -312 2159 -278 2179
rect -312 2091 -278 2107
rect -312 2023 -278 2035
rect -312 1955 -278 1963
rect -312 1887 -278 1891
rect -312 1781 -278 1785
rect -312 1709 -278 1717
rect -312 1637 -278 1649
rect -312 1565 -278 1581
rect -312 1493 -278 1513
rect -312 1421 -278 1445
rect -312 1349 -278 1377
rect -312 1277 -278 1309
rect -312 1207 -278 1241
rect -312 1139 -278 1171
rect -312 1071 -278 1099
rect -312 1003 -278 1027
rect -312 935 -278 955
rect -312 867 -278 883
rect -312 799 -278 811
rect -312 731 -278 739
rect -312 663 -278 667
rect -312 557 -278 561
rect -312 485 -278 493
rect -312 413 -278 425
rect -312 341 -278 357
rect -312 269 -278 289
rect -312 197 -278 221
rect -312 125 -278 153
rect -312 53 -278 85
rect -312 -17 -278 17
rect -312 -85 -278 -53
rect -312 -153 -278 -125
rect -312 -221 -278 -197
rect -312 -289 -278 -269
rect -312 -357 -278 -341
rect -312 -425 -278 -413
rect -312 -493 -278 -485
rect -312 -561 -278 -557
rect -312 -667 -278 -663
rect -312 -739 -278 -731
rect -312 -811 -278 -799
rect -312 -883 -278 -867
rect -312 -955 -278 -935
rect -312 -1027 -278 -1003
rect -312 -1099 -278 -1071
rect -312 -1171 -278 -1139
rect -312 -1241 -278 -1207
rect -312 -1309 -278 -1277
rect -312 -1377 -278 -1349
rect -312 -1445 -278 -1421
rect -312 -1513 -278 -1493
rect -312 -1581 -278 -1565
rect -312 -1649 -278 -1637
rect -312 -1717 -278 -1709
rect -312 -1785 -278 -1781
rect -312 -1891 -278 -1887
rect -312 -1963 -278 -1955
rect -312 -2035 -278 -2023
rect -312 -2107 -278 -2091
rect -312 -2179 -278 -2159
rect -312 -2251 -278 -2227
rect -312 -2323 -278 -2295
rect -312 -2395 -278 -2363
rect -312 -2465 -278 -2431
rect -312 -2533 -278 -2501
rect -312 -2601 -278 -2573
rect -312 -2669 -278 -2645
rect -312 -2737 -278 -2717
rect -312 -2805 -278 -2789
rect -312 -2873 -278 -2861
rect -312 -2941 -278 -2933
rect -312 -3009 -278 -3005
rect -312 -3115 -278 -3111
rect -312 -3187 -278 -3179
rect -312 -3259 -278 -3247
rect -312 -3331 -278 -3315
rect -312 -3403 -278 -3383
rect -312 -3475 -278 -3451
rect -312 -3547 -278 -3519
rect -312 -3619 -278 -3587
rect -312 -3689 -278 -3655
rect -312 -3757 -278 -3725
rect -312 -3825 -278 -3797
rect -312 -3893 -278 -3869
rect -312 -3961 -278 -3941
rect -312 -4029 -278 -4013
rect -312 -4097 -278 -4085
rect -312 -4165 -278 -4157
rect -312 -4233 -278 -4229
rect -312 -4339 -278 -4335
rect -312 -4411 -278 -4403
rect -312 -4483 -278 -4471
rect -312 -4555 -278 -4539
rect -312 -4627 -278 -4607
rect -312 -4699 -278 -4675
rect -312 -4771 -278 -4743
rect -312 -4843 -278 -4811
rect -312 -4913 -278 -4879
rect -312 -4981 -278 -4949
rect -312 -5049 -278 -5021
rect -312 -5117 -278 -5093
rect -312 -5185 -278 -5165
rect -312 -5253 -278 -5237
rect -312 -5321 -278 -5309
rect -312 -5389 -278 -5381
rect -312 -5457 -278 -5453
rect -312 -5563 -278 -5559
rect -312 -5635 -278 -5627
rect -312 -5707 -278 -5695
rect -312 -5779 -278 -5763
rect -312 -5851 -278 -5831
rect -312 -5923 -278 -5899
rect -312 -5995 -278 -5967
rect -312 -6067 -278 -6035
rect -312 -6137 -278 -6103
rect -312 -6205 -278 -6173
rect -312 -6273 -278 -6245
rect -312 -6341 -278 -6317
rect -312 -6409 -278 -6389
rect -312 -6477 -278 -6461
rect -312 -6545 -278 -6533
rect -312 -6613 -278 -6605
rect -312 -6681 -278 -6677
rect -312 -6787 -278 -6783
rect -312 -6859 -278 -6851
rect -312 -6931 -278 -6919
rect -312 -7003 -278 -6987
rect -312 -7075 -278 -7055
rect -312 -7147 -278 -7123
rect -312 -7219 -278 -7191
rect -312 -7291 -278 -7259
rect -312 -7361 -278 -7327
rect -312 -7429 -278 -7397
rect -312 -7497 -278 -7469
rect -312 -7565 -278 -7541
rect -312 -7633 -278 -7613
rect -312 -7701 -278 -7685
rect -312 -7769 -278 -7757
rect -312 -7837 -278 -7829
rect -312 -7905 -278 -7901
rect -312 -8011 -278 -8007
rect -312 -8083 -278 -8075
rect -312 -8155 -278 -8143
rect -312 -8227 -278 -8211
rect -312 -8299 -278 -8279
rect -312 -8371 -278 -8347
rect -312 -8443 -278 -8415
rect -312 -8515 -278 -8483
rect -312 -8585 -278 -8551
rect -312 -8653 -278 -8621
rect -312 -8721 -278 -8693
rect -312 -8789 -278 -8765
rect -312 -8857 -278 -8837
rect -312 -8925 -278 -8909
rect -312 -8993 -278 -8981
rect -312 -9061 -278 -9053
rect -312 -9129 -278 -9125
rect -312 -9235 -278 -9231
rect -312 -9307 -278 -9299
rect -312 -9379 -278 -9367
rect -312 -9451 -278 -9435
rect -312 -9523 -278 -9503
rect -312 -9604 -278 -9571
rect -194 9571 -160 9604
rect -194 9503 -160 9523
rect -194 9435 -160 9451
rect -194 9367 -160 9379
rect -194 9299 -160 9307
rect -194 9231 -160 9235
rect -194 9125 -160 9129
rect -194 9053 -160 9061
rect -194 8981 -160 8993
rect -194 8909 -160 8925
rect -194 8837 -160 8857
rect -194 8765 -160 8789
rect -194 8693 -160 8721
rect -194 8621 -160 8653
rect -194 8551 -160 8585
rect -194 8483 -160 8515
rect -194 8415 -160 8443
rect -194 8347 -160 8371
rect -194 8279 -160 8299
rect -194 8211 -160 8227
rect -194 8143 -160 8155
rect -194 8075 -160 8083
rect -194 8007 -160 8011
rect -194 7901 -160 7905
rect -194 7829 -160 7837
rect -194 7757 -160 7769
rect -194 7685 -160 7701
rect -194 7613 -160 7633
rect -194 7541 -160 7565
rect -194 7469 -160 7497
rect -194 7397 -160 7429
rect -194 7327 -160 7361
rect -194 7259 -160 7291
rect -194 7191 -160 7219
rect -194 7123 -160 7147
rect -194 7055 -160 7075
rect -194 6987 -160 7003
rect -194 6919 -160 6931
rect -194 6851 -160 6859
rect -194 6783 -160 6787
rect -194 6677 -160 6681
rect -194 6605 -160 6613
rect -194 6533 -160 6545
rect -194 6461 -160 6477
rect -194 6389 -160 6409
rect -194 6317 -160 6341
rect -194 6245 -160 6273
rect -194 6173 -160 6205
rect -194 6103 -160 6137
rect -194 6035 -160 6067
rect -194 5967 -160 5995
rect -194 5899 -160 5923
rect -194 5831 -160 5851
rect -194 5763 -160 5779
rect -194 5695 -160 5707
rect -194 5627 -160 5635
rect -194 5559 -160 5563
rect -194 5453 -160 5457
rect -194 5381 -160 5389
rect -194 5309 -160 5321
rect -194 5237 -160 5253
rect -194 5165 -160 5185
rect -194 5093 -160 5117
rect -194 5021 -160 5049
rect -194 4949 -160 4981
rect -194 4879 -160 4913
rect -194 4811 -160 4843
rect -194 4743 -160 4771
rect -194 4675 -160 4699
rect -194 4607 -160 4627
rect -194 4539 -160 4555
rect -194 4471 -160 4483
rect -194 4403 -160 4411
rect -194 4335 -160 4339
rect -194 4229 -160 4233
rect -194 4157 -160 4165
rect -194 4085 -160 4097
rect -194 4013 -160 4029
rect -194 3941 -160 3961
rect -194 3869 -160 3893
rect -194 3797 -160 3825
rect -194 3725 -160 3757
rect -194 3655 -160 3689
rect -194 3587 -160 3619
rect -194 3519 -160 3547
rect -194 3451 -160 3475
rect -194 3383 -160 3403
rect -194 3315 -160 3331
rect -194 3247 -160 3259
rect -194 3179 -160 3187
rect -194 3111 -160 3115
rect -194 3005 -160 3009
rect -194 2933 -160 2941
rect -194 2861 -160 2873
rect -194 2789 -160 2805
rect -194 2717 -160 2737
rect -194 2645 -160 2669
rect -194 2573 -160 2601
rect -194 2501 -160 2533
rect -194 2431 -160 2465
rect -194 2363 -160 2395
rect -194 2295 -160 2323
rect -194 2227 -160 2251
rect -194 2159 -160 2179
rect -194 2091 -160 2107
rect -194 2023 -160 2035
rect -194 1955 -160 1963
rect -194 1887 -160 1891
rect -194 1781 -160 1785
rect -194 1709 -160 1717
rect -194 1637 -160 1649
rect -194 1565 -160 1581
rect -194 1493 -160 1513
rect -194 1421 -160 1445
rect -194 1349 -160 1377
rect -194 1277 -160 1309
rect -194 1207 -160 1241
rect -194 1139 -160 1171
rect -194 1071 -160 1099
rect -194 1003 -160 1027
rect -194 935 -160 955
rect -194 867 -160 883
rect -194 799 -160 811
rect -194 731 -160 739
rect -194 663 -160 667
rect -194 557 -160 561
rect -194 485 -160 493
rect -194 413 -160 425
rect -194 341 -160 357
rect -194 269 -160 289
rect -194 197 -160 221
rect -194 125 -160 153
rect -194 53 -160 85
rect -194 -17 -160 17
rect -194 -85 -160 -53
rect -194 -153 -160 -125
rect -194 -221 -160 -197
rect -194 -289 -160 -269
rect -194 -357 -160 -341
rect -194 -425 -160 -413
rect -194 -493 -160 -485
rect -194 -561 -160 -557
rect -194 -667 -160 -663
rect -194 -739 -160 -731
rect -194 -811 -160 -799
rect -194 -883 -160 -867
rect -194 -955 -160 -935
rect -194 -1027 -160 -1003
rect -194 -1099 -160 -1071
rect -194 -1171 -160 -1139
rect -194 -1241 -160 -1207
rect -194 -1309 -160 -1277
rect -194 -1377 -160 -1349
rect -194 -1445 -160 -1421
rect -194 -1513 -160 -1493
rect -194 -1581 -160 -1565
rect -194 -1649 -160 -1637
rect -194 -1717 -160 -1709
rect -194 -1785 -160 -1781
rect -194 -1891 -160 -1887
rect -194 -1963 -160 -1955
rect -194 -2035 -160 -2023
rect -194 -2107 -160 -2091
rect -194 -2179 -160 -2159
rect -194 -2251 -160 -2227
rect -194 -2323 -160 -2295
rect -194 -2395 -160 -2363
rect -194 -2465 -160 -2431
rect -194 -2533 -160 -2501
rect -194 -2601 -160 -2573
rect -194 -2669 -160 -2645
rect -194 -2737 -160 -2717
rect -194 -2805 -160 -2789
rect -194 -2873 -160 -2861
rect -194 -2941 -160 -2933
rect -194 -3009 -160 -3005
rect -194 -3115 -160 -3111
rect -194 -3187 -160 -3179
rect -194 -3259 -160 -3247
rect -194 -3331 -160 -3315
rect -194 -3403 -160 -3383
rect -194 -3475 -160 -3451
rect -194 -3547 -160 -3519
rect -194 -3619 -160 -3587
rect -194 -3689 -160 -3655
rect -194 -3757 -160 -3725
rect -194 -3825 -160 -3797
rect -194 -3893 -160 -3869
rect -194 -3961 -160 -3941
rect -194 -4029 -160 -4013
rect -194 -4097 -160 -4085
rect -194 -4165 -160 -4157
rect -194 -4233 -160 -4229
rect -194 -4339 -160 -4335
rect -194 -4411 -160 -4403
rect -194 -4483 -160 -4471
rect -194 -4555 -160 -4539
rect -194 -4627 -160 -4607
rect -194 -4699 -160 -4675
rect -194 -4771 -160 -4743
rect -194 -4843 -160 -4811
rect -194 -4913 -160 -4879
rect -194 -4981 -160 -4949
rect -194 -5049 -160 -5021
rect -194 -5117 -160 -5093
rect -194 -5185 -160 -5165
rect -194 -5253 -160 -5237
rect -194 -5321 -160 -5309
rect -194 -5389 -160 -5381
rect -194 -5457 -160 -5453
rect -194 -5563 -160 -5559
rect -194 -5635 -160 -5627
rect -194 -5707 -160 -5695
rect -194 -5779 -160 -5763
rect -194 -5851 -160 -5831
rect -194 -5923 -160 -5899
rect -194 -5995 -160 -5967
rect -194 -6067 -160 -6035
rect -194 -6137 -160 -6103
rect -194 -6205 -160 -6173
rect -194 -6273 -160 -6245
rect -194 -6341 -160 -6317
rect -194 -6409 -160 -6389
rect -194 -6477 -160 -6461
rect -194 -6545 -160 -6533
rect -194 -6613 -160 -6605
rect -194 -6681 -160 -6677
rect -194 -6787 -160 -6783
rect -194 -6859 -160 -6851
rect -194 -6931 -160 -6919
rect -194 -7003 -160 -6987
rect -194 -7075 -160 -7055
rect -194 -7147 -160 -7123
rect -194 -7219 -160 -7191
rect -194 -7291 -160 -7259
rect -194 -7361 -160 -7327
rect -194 -7429 -160 -7397
rect -194 -7497 -160 -7469
rect -194 -7565 -160 -7541
rect -194 -7633 -160 -7613
rect -194 -7701 -160 -7685
rect -194 -7769 -160 -7757
rect -194 -7837 -160 -7829
rect -194 -7905 -160 -7901
rect -194 -8011 -160 -8007
rect -194 -8083 -160 -8075
rect -194 -8155 -160 -8143
rect -194 -8227 -160 -8211
rect -194 -8299 -160 -8279
rect -194 -8371 -160 -8347
rect -194 -8443 -160 -8415
rect -194 -8515 -160 -8483
rect -194 -8585 -160 -8551
rect -194 -8653 -160 -8621
rect -194 -8721 -160 -8693
rect -194 -8789 -160 -8765
rect -194 -8857 -160 -8837
rect -194 -8925 -160 -8909
rect -194 -8993 -160 -8981
rect -194 -9061 -160 -9053
rect -194 -9129 -160 -9125
rect -194 -9235 -160 -9231
rect -194 -9307 -160 -9299
rect -194 -9379 -160 -9367
rect -194 -9451 -160 -9435
rect -194 -9523 -160 -9503
rect -194 -9604 -160 -9571
rect -76 9571 -42 9604
rect -76 9503 -42 9523
rect -76 9435 -42 9451
rect -76 9367 -42 9379
rect -76 9299 -42 9307
rect -76 9231 -42 9235
rect -76 9125 -42 9129
rect -76 9053 -42 9061
rect -76 8981 -42 8993
rect -76 8909 -42 8925
rect -76 8837 -42 8857
rect -76 8765 -42 8789
rect -76 8693 -42 8721
rect -76 8621 -42 8653
rect -76 8551 -42 8585
rect -76 8483 -42 8515
rect -76 8415 -42 8443
rect -76 8347 -42 8371
rect -76 8279 -42 8299
rect -76 8211 -42 8227
rect -76 8143 -42 8155
rect -76 8075 -42 8083
rect -76 8007 -42 8011
rect -76 7901 -42 7905
rect -76 7829 -42 7837
rect -76 7757 -42 7769
rect -76 7685 -42 7701
rect -76 7613 -42 7633
rect -76 7541 -42 7565
rect -76 7469 -42 7497
rect -76 7397 -42 7429
rect -76 7327 -42 7361
rect -76 7259 -42 7291
rect -76 7191 -42 7219
rect -76 7123 -42 7147
rect -76 7055 -42 7075
rect -76 6987 -42 7003
rect -76 6919 -42 6931
rect -76 6851 -42 6859
rect -76 6783 -42 6787
rect -76 6677 -42 6681
rect -76 6605 -42 6613
rect -76 6533 -42 6545
rect -76 6461 -42 6477
rect -76 6389 -42 6409
rect -76 6317 -42 6341
rect -76 6245 -42 6273
rect -76 6173 -42 6205
rect -76 6103 -42 6137
rect -76 6035 -42 6067
rect -76 5967 -42 5995
rect -76 5899 -42 5923
rect -76 5831 -42 5851
rect -76 5763 -42 5779
rect -76 5695 -42 5707
rect -76 5627 -42 5635
rect -76 5559 -42 5563
rect -76 5453 -42 5457
rect -76 5381 -42 5389
rect -76 5309 -42 5321
rect -76 5237 -42 5253
rect -76 5165 -42 5185
rect -76 5093 -42 5117
rect -76 5021 -42 5049
rect -76 4949 -42 4981
rect -76 4879 -42 4913
rect -76 4811 -42 4843
rect -76 4743 -42 4771
rect -76 4675 -42 4699
rect -76 4607 -42 4627
rect -76 4539 -42 4555
rect -76 4471 -42 4483
rect -76 4403 -42 4411
rect -76 4335 -42 4339
rect -76 4229 -42 4233
rect -76 4157 -42 4165
rect -76 4085 -42 4097
rect -76 4013 -42 4029
rect -76 3941 -42 3961
rect -76 3869 -42 3893
rect -76 3797 -42 3825
rect -76 3725 -42 3757
rect -76 3655 -42 3689
rect -76 3587 -42 3619
rect -76 3519 -42 3547
rect -76 3451 -42 3475
rect -76 3383 -42 3403
rect -76 3315 -42 3331
rect -76 3247 -42 3259
rect -76 3179 -42 3187
rect -76 3111 -42 3115
rect -76 3005 -42 3009
rect -76 2933 -42 2941
rect -76 2861 -42 2873
rect -76 2789 -42 2805
rect -76 2717 -42 2737
rect -76 2645 -42 2669
rect -76 2573 -42 2601
rect -76 2501 -42 2533
rect -76 2431 -42 2465
rect -76 2363 -42 2395
rect -76 2295 -42 2323
rect -76 2227 -42 2251
rect -76 2159 -42 2179
rect -76 2091 -42 2107
rect -76 2023 -42 2035
rect -76 1955 -42 1963
rect -76 1887 -42 1891
rect -76 1781 -42 1785
rect -76 1709 -42 1717
rect -76 1637 -42 1649
rect -76 1565 -42 1581
rect -76 1493 -42 1513
rect -76 1421 -42 1445
rect -76 1349 -42 1377
rect -76 1277 -42 1309
rect -76 1207 -42 1241
rect -76 1139 -42 1171
rect -76 1071 -42 1099
rect -76 1003 -42 1027
rect -76 935 -42 955
rect -76 867 -42 883
rect -76 799 -42 811
rect -76 731 -42 739
rect -76 663 -42 667
rect -76 557 -42 561
rect -76 485 -42 493
rect -76 413 -42 425
rect -76 341 -42 357
rect -76 269 -42 289
rect -76 197 -42 221
rect -76 125 -42 153
rect -76 53 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -53
rect -76 -153 -42 -125
rect -76 -221 -42 -197
rect -76 -289 -42 -269
rect -76 -357 -42 -341
rect -76 -425 -42 -413
rect -76 -493 -42 -485
rect -76 -561 -42 -557
rect -76 -667 -42 -663
rect -76 -739 -42 -731
rect -76 -811 -42 -799
rect -76 -883 -42 -867
rect -76 -955 -42 -935
rect -76 -1027 -42 -1003
rect -76 -1099 -42 -1071
rect -76 -1171 -42 -1139
rect -76 -1241 -42 -1207
rect -76 -1309 -42 -1277
rect -76 -1377 -42 -1349
rect -76 -1445 -42 -1421
rect -76 -1513 -42 -1493
rect -76 -1581 -42 -1565
rect -76 -1649 -42 -1637
rect -76 -1717 -42 -1709
rect -76 -1785 -42 -1781
rect -76 -1891 -42 -1887
rect -76 -1963 -42 -1955
rect -76 -2035 -42 -2023
rect -76 -2107 -42 -2091
rect -76 -2179 -42 -2159
rect -76 -2251 -42 -2227
rect -76 -2323 -42 -2295
rect -76 -2395 -42 -2363
rect -76 -2465 -42 -2431
rect -76 -2533 -42 -2501
rect -76 -2601 -42 -2573
rect -76 -2669 -42 -2645
rect -76 -2737 -42 -2717
rect -76 -2805 -42 -2789
rect -76 -2873 -42 -2861
rect -76 -2941 -42 -2933
rect -76 -3009 -42 -3005
rect -76 -3115 -42 -3111
rect -76 -3187 -42 -3179
rect -76 -3259 -42 -3247
rect -76 -3331 -42 -3315
rect -76 -3403 -42 -3383
rect -76 -3475 -42 -3451
rect -76 -3547 -42 -3519
rect -76 -3619 -42 -3587
rect -76 -3689 -42 -3655
rect -76 -3757 -42 -3725
rect -76 -3825 -42 -3797
rect -76 -3893 -42 -3869
rect -76 -3961 -42 -3941
rect -76 -4029 -42 -4013
rect -76 -4097 -42 -4085
rect -76 -4165 -42 -4157
rect -76 -4233 -42 -4229
rect -76 -4339 -42 -4335
rect -76 -4411 -42 -4403
rect -76 -4483 -42 -4471
rect -76 -4555 -42 -4539
rect -76 -4627 -42 -4607
rect -76 -4699 -42 -4675
rect -76 -4771 -42 -4743
rect -76 -4843 -42 -4811
rect -76 -4913 -42 -4879
rect -76 -4981 -42 -4949
rect -76 -5049 -42 -5021
rect -76 -5117 -42 -5093
rect -76 -5185 -42 -5165
rect -76 -5253 -42 -5237
rect -76 -5321 -42 -5309
rect -76 -5389 -42 -5381
rect -76 -5457 -42 -5453
rect -76 -5563 -42 -5559
rect -76 -5635 -42 -5627
rect -76 -5707 -42 -5695
rect -76 -5779 -42 -5763
rect -76 -5851 -42 -5831
rect -76 -5923 -42 -5899
rect -76 -5995 -42 -5967
rect -76 -6067 -42 -6035
rect -76 -6137 -42 -6103
rect -76 -6205 -42 -6173
rect -76 -6273 -42 -6245
rect -76 -6341 -42 -6317
rect -76 -6409 -42 -6389
rect -76 -6477 -42 -6461
rect -76 -6545 -42 -6533
rect -76 -6613 -42 -6605
rect -76 -6681 -42 -6677
rect -76 -6787 -42 -6783
rect -76 -6859 -42 -6851
rect -76 -6931 -42 -6919
rect -76 -7003 -42 -6987
rect -76 -7075 -42 -7055
rect -76 -7147 -42 -7123
rect -76 -7219 -42 -7191
rect -76 -7291 -42 -7259
rect -76 -7361 -42 -7327
rect -76 -7429 -42 -7397
rect -76 -7497 -42 -7469
rect -76 -7565 -42 -7541
rect -76 -7633 -42 -7613
rect -76 -7701 -42 -7685
rect -76 -7769 -42 -7757
rect -76 -7837 -42 -7829
rect -76 -7905 -42 -7901
rect -76 -8011 -42 -8007
rect -76 -8083 -42 -8075
rect -76 -8155 -42 -8143
rect -76 -8227 -42 -8211
rect -76 -8299 -42 -8279
rect -76 -8371 -42 -8347
rect -76 -8443 -42 -8415
rect -76 -8515 -42 -8483
rect -76 -8585 -42 -8551
rect -76 -8653 -42 -8621
rect -76 -8721 -42 -8693
rect -76 -8789 -42 -8765
rect -76 -8857 -42 -8837
rect -76 -8925 -42 -8909
rect -76 -8993 -42 -8981
rect -76 -9061 -42 -9053
rect -76 -9129 -42 -9125
rect -76 -9235 -42 -9231
rect -76 -9307 -42 -9299
rect -76 -9379 -42 -9367
rect -76 -9451 -42 -9435
rect -76 -9523 -42 -9503
rect -76 -9604 -42 -9571
rect 42 9571 76 9604
rect 42 9503 76 9523
rect 42 9435 76 9451
rect 42 9367 76 9379
rect 42 9299 76 9307
rect 42 9231 76 9235
rect 42 9125 76 9129
rect 42 9053 76 9061
rect 42 8981 76 8993
rect 42 8909 76 8925
rect 42 8837 76 8857
rect 42 8765 76 8789
rect 42 8693 76 8721
rect 42 8621 76 8653
rect 42 8551 76 8585
rect 42 8483 76 8515
rect 42 8415 76 8443
rect 42 8347 76 8371
rect 42 8279 76 8299
rect 42 8211 76 8227
rect 42 8143 76 8155
rect 42 8075 76 8083
rect 42 8007 76 8011
rect 42 7901 76 7905
rect 42 7829 76 7837
rect 42 7757 76 7769
rect 42 7685 76 7701
rect 42 7613 76 7633
rect 42 7541 76 7565
rect 42 7469 76 7497
rect 42 7397 76 7429
rect 42 7327 76 7361
rect 42 7259 76 7291
rect 42 7191 76 7219
rect 42 7123 76 7147
rect 42 7055 76 7075
rect 42 6987 76 7003
rect 42 6919 76 6931
rect 42 6851 76 6859
rect 42 6783 76 6787
rect 42 6677 76 6681
rect 42 6605 76 6613
rect 42 6533 76 6545
rect 42 6461 76 6477
rect 42 6389 76 6409
rect 42 6317 76 6341
rect 42 6245 76 6273
rect 42 6173 76 6205
rect 42 6103 76 6137
rect 42 6035 76 6067
rect 42 5967 76 5995
rect 42 5899 76 5923
rect 42 5831 76 5851
rect 42 5763 76 5779
rect 42 5695 76 5707
rect 42 5627 76 5635
rect 42 5559 76 5563
rect 42 5453 76 5457
rect 42 5381 76 5389
rect 42 5309 76 5321
rect 42 5237 76 5253
rect 42 5165 76 5185
rect 42 5093 76 5117
rect 42 5021 76 5049
rect 42 4949 76 4981
rect 42 4879 76 4913
rect 42 4811 76 4843
rect 42 4743 76 4771
rect 42 4675 76 4699
rect 42 4607 76 4627
rect 42 4539 76 4555
rect 42 4471 76 4483
rect 42 4403 76 4411
rect 42 4335 76 4339
rect 42 4229 76 4233
rect 42 4157 76 4165
rect 42 4085 76 4097
rect 42 4013 76 4029
rect 42 3941 76 3961
rect 42 3869 76 3893
rect 42 3797 76 3825
rect 42 3725 76 3757
rect 42 3655 76 3689
rect 42 3587 76 3619
rect 42 3519 76 3547
rect 42 3451 76 3475
rect 42 3383 76 3403
rect 42 3315 76 3331
rect 42 3247 76 3259
rect 42 3179 76 3187
rect 42 3111 76 3115
rect 42 3005 76 3009
rect 42 2933 76 2941
rect 42 2861 76 2873
rect 42 2789 76 2805
rect 42 2717 76 2737
rect 42 2645 76 2669
rect 42 2573 76 2601
rect 42 2501 76 2533
rect 42 2431 76 2465
rect 42 2363 76 2395
rect 42 2295 76 2323
rect 42 2227 76 2251
rect 42 2159 76 2179
rect 42 2091 76 2107
rect 42 2023 76 2035
rect 42 1955 76 1963
rect 42 1887 76 1891
rect 42 1781 76 1785
rect 42 1709 76 1717
rect 42 1637 76 1649
rect 42 1565 76 1581
rect 42 1493 76 1513
rect 42 1421 76 1445
rect 42 1349 76 1377
rect 42 1277 76 1309
rect 42 1207 76 1241
rect 42 1139 76 1171
rect 42 1071 76 1099
rect 42 1003 76 1027
rect 42 935 76 955
rect 42 867 76 883
rect 42 799 76 811
rect 42 731 76 739
rect 42 663 76 667
rect 42 557 76 561
rect 42 485 76 493
rect 42 413 76 425
rect 42 341 76 357
rect 42 269 76 289
rect 42 197 76 221
rect 42 125 76 153
rect 42 53 76 85
rect 42 -17 76 17
rect 42 -85 76 -53
rect 42 -153 76 -125
rect 42 -221 76 -197
rect 42 -289 76 -269
rect 42 -357 76 -341
rect 42 -425 76 -413
rect 42 -493 76 -485
rect 42 -561 76 -557
rect 42 -667 76 -663
rect 42 -739 76 -731
rect 42 -811 76 -799
rect 42 -883 76 -867
rect 42 -955 76 -935
rect 42 -1027 76 -1003
rect 42 -1099 76 -1071
rect 42 -1171 76 -1139
rect 42 -1241 76 -1207
rect 42 -1309 76 -1277
rect 42 -1377 76 -1349
rect 42 -1445 76 -1421
rect 42 -1513 76 -1493
rect 42 -1581 76 -1565
rect 42 -1649 76 -1637
rect 42 -1717 76 -1709
rect 42 -1785 76 -1781
rect 42 -1891 76 -1887
rect 42 -1963 76 -1955
rect 42 -2035 76 -2023
rect 42 -2107 76 -2091
rect 42 -2179 76 -2159
rect 42 -2251 76 -2227
rect 42 -2323 76 -2295
rect 42 -2395 76 -2363
rect 42 -2465 76 -2431
rect 42 -2533 76 -2501
rect 42 -2601 76 -2573
rect 42 -2669 76 -2645
rect 42 -2737 76 -2717
rect 42 -2805 76 -2789
rect 42 -2873 76 -2861
rect 42 -2941 76 -2933
rect 42 -3009 76 -3005
rect 42 -3115 76 -3111
rect 42 -3187 76 -3179
rect 42 -3259 76 -3247
rect 42 -3331 76 -3315
rect 42 -3403 76 -3383
rect 42 -3475 76 -3451
rect 42 -3547 76 -3519
rect 42 -3619 76 -3587
rect 42 -3689 76 -3655
rect 42 -3757 76 -3725
rect 42 -3825 76 -3797
rect 42 -3893 76 -3869
rect 42 -3961 76 -3941
rect 42 -4029 76 -4013
rect 42 -4097 76 -4085
rect 42 -4165 76 -4157
rect 42 -4233 76 -4229
rect 42 -4339 76 -4335
rect 42 -4411 76 -4403
rect 42 -4483 76 -4471
rect 42 -4555 76 -4539
rect 42 -4627 76 -4607
rect 42 -4699 76 -4675
rect 42 -4771 76 -4743
rect 42 -4843 76 -4811
rect 42 -4913 76 -4879
rect 42 -4981 76 -4949
rect 42 -5049 76 -5021
rect 42 -5117 76 -5093
rect 42 -5185 76 -5165
rect 42 -5253 76 -5237
rect 42 -5321 76 -5309
rect 42 -5389 76 -5381
rect 42 -5457 76 -5453
rect 42 -5563 76 -5559
rect 42 -5635 76 -5627
rect 42 -5707 76 -5695
rect 42 -5779 76 -5763
rect 42 -5851 76 -5831
rect 42 -5923 76 -5899
rect 42 -5995 76 -5967
rect 42 -6067 76 -6035
rect 42 -6137 76 -6103
rect 42 -6205 76 -6173
rect 42 -6273 76 -6245
rect 42 -6341 76 -6317
rect 42 -6409 76 -6389
rect 42 -6477 76 -6461
rect 42 -6545 76 -6533
rect 42 -6613 76 -6605
rect 42 -6681 76 -6677
rect 42 -6787 76 -6783
rect 42 -6859 76 -6851
rect 42 -6931 76 -6919
rect 42 -7003 76 -6987
rect 42 -7075 76 -7055
rect 42 -7147 76 -7123
rect 42 -7219 76 -7191
rect 42 -7291 76 -7259
rect 42 -7361 76 -7327
rect 42 -7429 76 -7397
rect 42 -7497 76 -7469
rect 42 -7565 76 -7541
rect 42 -7633 76 -7613
rect 42 -7701 76 -7685
rect 42 -7769 76 -7757
rect 42 -7837 76 -7829
rect 42 -7905 76 -7901
rect 42 -8011 76 -8007
rect 42 -8083 76 -8075
rect 42 -8155 76 -8143
rect 42 -8227 76 -8211
rect 42 -8299 76 -8279
rect 42 -8371 76 -8347
rect 42 -8443 76 -8415
rect 42 -8515 76 -8483
rect 42 -8585 76 -8551
rect 42 -8653 76 -8621
rect 42 -8721 76 -8693
rect 42 -8789 76 -8765
rect 42 -8857 76 -8837
rect 42 -8925 76 -8909
rect 42 -8993 76 -8981
rect 42 -9061 76 -9053
rect 42 -9129 76 -9125
rect 42 -9235 76 -9231
rect 42 -9307 76 -9299
rect 42 -9379 76 -9367
rect 42 -9451 76 -9435
rect 42 -9523 76 -9503
rect 42 -9604 76 -9571
rect 160 9571 194 9604
rect 160 9503 194 9523
rect 160 9435 194 9451
rect 160 9367 194 9379
rect 160 9299 194 9307
rect 160 9231 194 9235
rect 160 9125 194 9129
rect 160 9053 194 9061
rect 160 8981 194 8993
rect 160 8909 194 8925
rect 160 8837 194 8857
rect 160 8765 194 8789
rect 160 8693 194 8721
rect 160 8621 194 8653
rect 160 8551 194 8585
rect 160 8483 194 8515
rect 160 8415 194 8443
rect 160 8347 194 8371
rect 160 8279 194 8299
rect 160 8211 194 8227
rect 160 8143 194 8155
rect 160 8075 194 8083
rect 160 8007 194 8011
rect 160 7901 194 7905
rect 160 7829 194 7837
rect 160 7757 194 7769
rect 160 7685 194 7701
rect 160 7613 194 7633
rect 160 7541 194 7565
rect 160 7469 194 7497
rect 160 7397 194 7429
rect 160 7327 194 7361
rect 160 7259 194 7291
rect 160 7191 194 7219
rect 160 7123 194 7147
rect 160 7055 194 7075
rect 160 6987 194 7003
rect 160 6919 194 6931
rect 160 6851 194 6859
rect 160 6783 194 6787
rect 160 6677 194 6681
rect 160 6605 194 6613
rect 160 6533 194 6545
rect 160 6461 194 6477
rect 160 6389 194 6409
rect 160 6317 194 6341
rect 160 6245 194 6273
rect 160 6173 194 6205
rect 160 6103 194 6137
rect 160 6035 194 6067
rect 160 5967 194 5995
rect 160 5899 194 5923
rect 160 5831 194 5851
rect 160 5763 194 5779
rect 160 5695 194 5707
rect 160 5627 194 5635
rect 160 5559 194 5563
rect 160 5453 194 5457
rect 160 5381 194 5389
rect 160 5309 194 5321
rect 160 5237 194 5253
rect 160 5165 194 5185
rect 160 5093 194 5117
rect 160 5021 194 5049
rect 160 4949 194 4981
rect 160 4879 194 4913
rect 160 4811 194 4843
rect 160 4743 194 4771
rect 160 4675 194 4699
rect 160 4607 194 4627
rect 160 4539 194 4555
rect 160 4471 194 4483
rect 160 4403 194 4411
rect 160 4335 194 4339
rect 160 4229 194 4233
rect 160 4157 194 4165
rect 160 4085 194 4097
rect 160 4013 194 4029
rect 160 3941 194 3961
rect 160 3869 194 3893
rect 160 3797 194 3825
rect 160 3725 194 3757
rect 160 3655 194 3689
rect 160 3587 194 3619
rect 160 3519 194 3547
rect 160 3451 194 3475
rect 160 3383 194 3403
rect 160 3315 194 3331
rect 160 3247 194 3259
rect 160 3179 194 3187
rect 160 3111 194 3115
rect 160 3005 194 3009
rect 160 2933 194 2941
rect 160 2861 194 2873
rect 160 2789 194 2805
rect 160 2717 194 2737
rect 160 2645 194 2669
rect 160 2573 194 2601
rect 160 2501 194 2533
rect 160 2431 194 2465
rect 160 2363 194 2395
rect 160 2295 194 2323
rect 160 2227 194 2251
rect 160 2159 194 2179
rect 160 2091 194 2107
rect 160 2023 194 2035
rect 160 1955 194 1963
rect 160 1887 194 1891
rect 160 1781 194 1785
rect 160 1709 194 1717
rect 160 1637 194 1649
rect 160 1565 194 1581
rect 160 1493 194 1513
rect 160 1421 194 1445
rect 160 1349 194 1377
rect 160 1277 194 1309
rect 160 1207 194 1241
rect 160 1139 194 1171
rect 160 1071 194 1099
rect 160 1003 194 1027
rect 160 935 194 955
rect 160 867 194 883
rect 160 799 194 811
rect 160 731 194 739
rect 160 663 194 667
rect 160 557 194 561
rect 160 485 194 493
rect 160 413 194 425
rect 160 341 194 357
rect 160 269 194 289
rect 160 197 194 221
rect 160 125 194 153
rect 160 53 194 85
rect 160 -17 194 17
rect 160 -85 194 -53
rect 160 -153 194 -125
rect 160 -221 194 -197
rect 160 -289 194 -269
rect 160 -357 194 -341
rect 160 -425 194 -413
rect 160 -493 194 -485
rect 160 -561 194 -557
rect 160 -667 194 -663
rect 160 -739 194 -731
rect 160 -811 194 -799
rect 160 -883 194 -867
rect 160 -955 194 -935
rect 160 -1027 194 -1003
rect 160 -1099 194 -1071
rect 160 -1171 194 -1139
rect 160 -1241 194 -1207
rect 160 -1309 194 -1277
rect 160 -1377 194 -1349
rect 160 -1445 194 -1421
rect 160 -1513 194 -1493
rect 160 -1581 194 -1565
rect 160 -1649 194 -1637
rect 160 -1717 194 -1709
rect 160 -1785 194 -1781
rect 160 -1891 194 -1887
rect 160 -1963 194 -1955
rect 160 -2035 194 -2023
rect 160 -2107 194 -2091
rect 160 -2179 194 -2159
rect 160 -2251 194 -2227
rect 160 -2323 194 -2295
rect 160 -2395 194 -2363
rect 160 -2465 194 -2431
rect 160 -2533 194 -2501
rect 160 -2601 194 -2573
rect 160 -2669 194 -2645
rect 160 -2737 194 -2717
rect 160 -2805 194 -2789
rect 160 -2873 194 -2861
rect 160 -2941 194 -2933
rect 160 -3009 194 -3005
rect 160 -3115 194 -3111
rect 160 -3187 194 -3179
rect 160 -3259 194 -3247
rect 160 -3331 194 -3315
rect 160 -3403 194 -3383
rect 160 -3475 194 -3451
rect 160 -3547 194 -3519
rect 160 -3619 194 -3587
rect 160 -3689 194 -3655
rect 160 -3757 194 -3725
rect 160 -3825 194 -3797
rect 160 -3893 194 -3869
rect 160 -3961 194 -3941
rect 160 -4029 194 -4013
rect 160 -4097 194 -4085
rect 160 -4165 194 -4157
rect 160 -4233 194 -4229
rect 160 -4339 194 -4335
rect 160 -4411 194 -4403
rect 160 -4483 194 -4471
rect 160 -4555 194 -4539
rect 160 -4627 194 -4607
rect 160 -4699 194 -4675
rect 160 -4771 194 -4743
rect 160 -4843 194 -4811
rect 160 -4913 194 -4879
rect 160 -4981 194 -4949
rect 160 -5049 194 -5021
rect 160 -5117 194 -5093
rect 160 -5185 194 -5165
rect 160 -5253 194 -5237
rect 160 -5321 194 -5309
rect 160 -5389 194 -5381
rect 160 -5457 194 -5453
rect 160 -5563 194 -5559
rect 160 -5635 194 -5627
rect 160 -5707 194 -5695
rect 160 -5779 194 -5763
rect 160 -5851 194 -5831
rect 160 -5923 194 -5899
rect 160 -5995 194 -5967
rect 160 -6067 194 -6035
rect 160 -6137 194 -6103
rect 160 -6205 194 -6173
rect 160 -6273 194 -6245
rect 160 -6341 194 -6317
rect 160 -6409 194 -6389
rect 160 -6477 194 -6461
rect 160 -6545 194 -6533
rect 160 -6613 194 -6605
rect 160 -6681 194 -6677
rect 160 -6787 194 -6783
rect 160 -6859 194 -6851
rect 160 -6931 194 -6919
rect 160 -7003 194 -6987
rect 160 -7075 194 -7055
rect 160 -7147 194 -7123
rect 160 -7219 194 -7191
rect 160 -7291 194 -7259
rect 160 -7361 194 -7327
rect 160 -7429 194 -7397
rect 160 -7497 194 -7469
rect 160 -7565 194 -7541
rect 160 -7633 194 -7613
rect 160 -7701 194 -7685
rect 160 -7769 194 -7757
rect 160 -7837 194 -7829
rect 160 -7905 194 -7901
rect 160 -8011 194 -8007
rect 160 -8083 194 -8075
rect 160 -8155 194 -8143
rect 160 -8227 194 -8211
rect 160 -8299 194 -8279
rect 160 -8371 194 -8347
rect 160 -8443 194 -8415
rect 160 -8515 194 -8483
rect 160 -8585 194 -8551
rect 160 -8653 194 -8621
rect 160 -8721 194 -8693
rect 160 -8789 194 -8765
rect 160 -8857 194 -8837
rect 160 -8925 194 -8909
rect 160 -8993 194 -8981
rect 160 -9061 194 -9053
rect 160 -9129 194 -9125
rect 160 -9235 194 -9231
rect 160 -9307 194 -9299
rect 160 -9379 194 -9367
rect 160 -9451 194 -9435
rect 160 -9523 194 -9503
rect 160 -9604 194 -9571
rect 278 9571 312 9604
rect 278 9503 312 9523
rect 278 9435 312 9451
rect 278 9367 312 9379
rect 278 9299 312 9307
rect 278 9231 312 9235
rect 278 9125 312 9129
rect 278 9053 312 9061
rect 278 8981 312 8993
rect 278 8909 312 8925
rect 278 8837 312 8857
rect 278 8765 312 8789
rect 278 8693 312 8721
rect 278 8621 312 8653
rect 278 8551 312 8585
rect 278 8483 312 8515
rect 278 8415 312 8443
rect 278 8347 312 8371
rect 278 8279 312 8299
rect 278 8211 312 8227
rect 278 8143 312 8155
rect 278 8075 312 8083
rect 278 8007 312 8011
rect 278 7901 312 7905
rect 278 7829 312 7837
rect 278 7757 312 7769
rect 278 7685 312 7701
rect 278 7613 312 7633
rect 278 7541 312 7565
rect 278 7469 312 7497
rect 278 7397 312 7429
rect 278 7327 312 7361
rect 278 7259 312 7291
rect 278 7191 312 7219
rect 278 7123 312 7147
rect 278 7055 312 7075
rect 278 6987 312 7003
rect 278 6919 312 6931
rect 278 6851 312 6859
rect 278 6783 312 6787
rect 278 6677 312 6681
rect 278 6605 312 6613
rect 278 6533 312 6545
rect 278 6461 312 6477
rect 278 6389 312 6409
rect 278 6317 312 6341
rect 278 6245 312 6273
rect 278 6173 312 6205
rect 278 6103 312 6137
rect 278 6035 312 6067
rect 278 5967 312 5995
rect 278 5899 312 5923
rect 278 5831 312 5851
rect 278 5763 312 5779
rect 278 5695 312 5707
rect 278 5627 312 5635
rect 278 5559 312 5563
rect 278 5453 312 5457
rect 278 5381 312 5389
rect 278 5309 312 5321
rect 278 5237 312 5253
rect 278 5165 312 5185
rect 278 5093 312 5117
rect 278 5021 312 5049
rect 278 4949 312 4981
rect 278 4879 312 4913
rect 278 4811 312 4843
rect 278 4743 312 4771
rect 278 4675 312 4699
rect 278 4607 312 4627
rect 278 4539 312 4555
rect 278 4471 312 4483
rect 278 4403 312 4411
rect 278 4335 312 4339
rect 278 4229 312 4233
rect 278 4157 312 4165
rect 278 4085 312 4097
rect 278 4013 312 4029
rect 278 3941 312 3961
rect 278 3869 312 3893
rect 278 3797 312 3825
rect 278 3725 312 3757
rect 278 3655 312 3689
rect 278 3587 312 3619
rect 278 3519 312 3547
rect 278 3451 312 3475
rect 278 3383 312 3403
rect 278 3315 312 3331
rect 278 3247 312 3259
rect 278 3179 312 3187
rect 278 3111 312 3115
rect 278 3005 312 3009
rect 278 2933 312 2941
rect 278 2861 312 2873
rect 278 2789 312 2805
rect 278 2717 312 2737
rect 278 2645 312 2669
rect 278 2573 312 2601
rect 278 2501 312 2533
rect 278 2431 312 2465
rect 278 2363 312 2395
rect 278 2295 312 2323
rect 278 2227 312 2251
rect 278 2159 312 2179
rect 278 2091 312 2107
rect 278 2023 312 2035
rect 278 1955 312 1963
rect 278 1887 312 1891
rect 278 1781 312 1785
rect 278 1709 312 1717
rect 278 1637 312 1649
rect 278 1565 312 1581
rect 278 1493 312 1513
rect 278 1421 312 1445
rect 278 1349 312 1377
rect 278 1277 312 1309
rect 278 1207 312 1241
rect 278 1139 312 1171
rect 278 1071 312 1099
rect 278 1003 312 1027
rect 278 935 312 955
rect 278 867 312 883
rect 278 799 312 811
rect 278 731 312 739
rect 278 663 312 667
rect 278 557 312 561
rect 278 485 312 493
rect 278 413 312 425
rect 278 341 312 357
rect 278 269 312 289
rect 278 197 312 221
rect 278 125 312 153
rect 278 53 312 85
rect 278 -17 312 17
rect 278 -85 312 -53
rect 278 -153 312 -125
rect 278 -221 312 -197
rect 278 -289 312 -269
rect 278 -357 312 -341
rect 278 -425 312 -413
rect 278 -493 312 -485
rect 278 -561 312 -557
rect 278 -667 312 -663
rect 278 -739 312 -731
rect 278 -811 312 -799
rect 278 -883 312 -867
rect 278 -955 312 -935
rect 278 -1027 312 -1003
rect 278 -1099 312 -1071
rect 278 -1171 312 -1139
rect 278 -1241 312 -1207
rect 278 -1309 312 -1277
rect 278 -1377 312 -1349
rect 278 -1445 312 -1421
rect 278 -1513 312 -1493
rect 278 -1581 312 -1565
rect 278 -1649 312 -1637
rect 278 -1717 312 -1709
rect 278 -1785 312 -1781
rect 278 -1891 312 -1887
rect 278 -1963 312 -1955
rect 278 -2035 312 -2023
rect 278 -2107 312 -2091
rect 278 -2179 312 -2159
rect 278 -2251 312 -2227
rect 278 -2323 312 -2295
rect 278 -2395 312 -2363
rect 278 -2465 312 -2431
rect 278 -2533 312 -2501
rect 278 -2601 312 -2573
rect 278 -2669 312 -2645
rect 278 -2737 312 -2717
rect 278 -2805 312 -2789
rect 278 -2873 312 -2861
rect 278 -2941 312 -2933
rect 278 -3009 312 -3005
rect 278 -3115 312 -3111
rect 278 -3187 312 -3179
rect 278 -3259 312 -3247
rect 278 -3331 312 -3315
rect 278 -3403 312 -3383
rect 278 -3475 312 -3451
rect 278 -3547 312 -3519
rect 278 -3619 312 -3587
rect 278 -3689 312 -3655
rect 278 -3757 312 -3725
rect 278 -3825 312 -3797
rect 278 -3893 312 -3869
rect 278 -3961 312 -3941
rect 278 -4029 312 -4013
rect 278 -4097 312 -4085
rect 278 -4165 312 -4157
rect 278 -4233 312 -4229
rect 278 -4339 312 -4335
rect 278 -4411 312 -4403
rect 278 -4483 312 -4471
rect 278 -4555 312 -4539
rect 278 -4627 312 -4607
rect 278 -4699 312 -4675
rect 278 -4771 312 -4743
rect 278 -4843 312 -4811
rect 278 -4913 312 -4879
rect 278 -4981 312 -4949
rect 278 -5049 312 -5021
rect 278 -5117 312 -5093
rect 278 -5185 312 -5165
rect 278 -5253 312 -5237
rect 278 -5321 312 -5309
rect 278 -5389 312 -5381
rect 278 -5457 312 -5453
rect 278 -5563 312 -5559
rect 278 -5635 312 -5627
rect 278 -5707 312 -5695
rect 278 -5779 312 -5763
rect 278 -5851 312 -5831
rect 278 -5923 312 -5899
rect 278 -5995 312 -5967
rect 278 -6067 312 -6035
rect 278 -6137 312 -6103
rect 278 -6205 312 -6173
rect 278 -6273 312 -6245
rect 278 -6341 312 -6317
rect 278 -6409 312 -6389
rect 278 -6477 312 -6461
rect 278 -6545 312 -6533
rect 278 -6613 312 -6605
rect 278 -6681 312 -6677
rect 278 -6787 312 -6783
rect 278 -6859 312 -6851
rect 278 -6931 312 -6919
rect 278 -7003 312 -6987
rect 278 -7075 312 -7055
rect 278 -7147 312 -7123
rect 278 -7219 312 -7191
rect 278 -7291 312 -7259
rect 278 -7361 312 -7327
rect 278 -7429 312 -7397
rect 278 -7497 312 -7469
rect 278 -7565 312 -7541
rect 278 -7633 312 -7613
rect 278 -7701 312 -7685
rect 278 -7769 312 -7757
rect 278 -7837 312 -7829
rect 278 -7905 312 -7901
rect 278 -8011 312 -8007
rect 278 -8083 312 -8075
rect 278 -8155 312 -8143
rect 278 -8227 312 -8211
rect 278 -8299 312 -8279
rect 278 -8371 312 -8347
rect 278 -8443 312 -8415
rect 278 -8515 312 -8483
rect 278 -8585 312 -8551
rect 278 -8653 312 -8621
rect 278 -8721 312 -8693
rect 278 -8789 312 -8765
rect 278 -8857 312 -8837
rect 278 -8925 312 -8909
rect 278 -8993 312 -8981
rect 278 -9061 312 -9053
rect 278 -9129 312 -9125
rect 278 -9235 312 -9231
rect 278 -9307 312 -9299
rect 278 -9379 312 -9367
rect 278 -9451 312 -9435
rect 278 -9523 312 -9503
rect 278 -9604 312 -9571
rect 396 9571 430 9604
rect 396 9503 430 9523
rect 396 9435 430 9451
rect 396 9367 430 9379
rect 396 9299 430 9307
rect 396 9231 430 9235
rect 396 9125 430 9129
rect 396 9053 430 9061
rect 396 8981 430 8993
rect 396 8909 430 8925
rect 396 8837 430 8857
rect 396 8765 430 8789
rect 396 8693 430 8721
rect 396 8621 430 8653
rect 396 8551 430 8585
rect 396 8483 430 8515
rect 396 8415 430 8443
rect 396 8347 430 8371
rect 396 8279 430 8299
rect 396 8211 430 8227
rect 396 8143 430 8155
rect 396 8075 430 8083
rect 396 8007 430 8011
rect 396 7901 430 7905
rect 396 7829 430 7837
rect 396 7757 430 7769
rect 396 7685 430 7701
rect 396 7613 430 7633
rect 396 7541 430 7565
rect 396 7469 430 7497
rect 396 7397 430 7429
rect 396 7327 430 7361
rect 396 7259 430 7291
rect 396 7191 430 7219
rect 396 7123 430 7147
rect 396 7055 430 7075
rect 396 6987 430 7003
rect 396 6919 430 6931
rect 396 6851 430 6859
rect 396 6783 430 6787
rect 396 6677 430 6681
rect 396 6605 430 6613
rect 396 6533 430 6545
rect 396 6461 430 6477
rect 396 6389 430 6409
rect 396 6317 430 6341
rect 396 6245 430 6273
rect 396 6173 430 6205
rect 396 6103 430 6137
rect 396 6035 430 6067
rect 396 5967 430 5995
rect 396 5899 430 5923
rect 396 5831 430 5851
rect 396 5763 430 5779
rect 396 5695 430 5707
rect 396 5627 430 5635
rect 396 5559 430 5563
rect 396 5453 430 5457
rect 396 5381 430 5389
rect 396 5309 430 5321
rect 396 5237 430 5253
rect 396 5165 430 5185
rect 396 5093 430 5117
rect 396 5021 430 5049
rect 396 4949 430 4981
rect 396 4879 430 4913
rect 396 4811 430 4843
rect 396 4743 430 4771
rect 396 4675 430 4699
rect 396 4607 430 4627
rect 396 4539 430 4555
rect 396 4471 430 4483
rect 396 4403 430 4411
rect 396 4335 430 4339
rect 396 4229 430 4233
rect 396 4157 430 4165
rect 396 4085 430 4097
rect 396 4013 430 4029
rect 396 3941 430 3961
rect 396 3869 430 3893
rect 396 3797 430 3825
rect 396 3725 430 3757
rect 396 3655 430 3689
rect 396 3587 430 3619
rect 396 3519 430 3547
rect 396 3451 430 3475
rect 396 3383 430 3403
rect 396 3315 430 3331
rect 396 3247 430 3259
rect 396 3179 430 3187
rect 396 3111 430 3115
rect 396 3005 430 3009
rect 396 2933 430 2941
rect 396 2861 430 2873
rect 396 2789 430 2805
rect 396 2717 430 2737
rect 396 2645 430 2669
rect 396 2573 430 2601
rect 396 2501 430 2533
rect 396 2431 430 2465
rect 396 2363 430 2395
rect 396 2295 430 2323
rect 396 2227 430 2251
rect 396 2159 430 2179
rect 396 2091 430 2107
rect 396 2023 430 2035
rect 396 1955 430 1963
rect 396 1887 430 1891
rect 396 1781 430 1785
rect 396 1709 430 1717
rect 396 1637 430 1649
rect 396 1565 430 1581
rect 396 1493 430 1513
rect 396 1421 430 1445
rect 396 1349 430 1377
rect 396 1277 430 1309
rect 396 1207 430 1241
rect 396 1139 430 1171
rect 396 1071 430 1099
rect 396 1003 430 1027
rect 396 935 430 955
rect 396 867 430 883
rect 396 799 430 811
rect 396 731 430 739
rect 396 663 430 667
rect 396 557 430 561
rect 396 485 430 493
rect 396 413 430 425
rect 396 341 430 357
rect 396 269 430 289
rect 396 197 430 221
rect 396 125 430 153
rect 396 53 430 85
rect 396 -17 430 17
rect 396 -85 430 -53
rect 396 -153 430 -125
rect 396 -221 430 -197
rect 396 -289 430 -269
rect 396 -357 430 -341
rect 396 -425 430 -413
rect 396 -493 430 -485
rect 396 -561 430 -557
rect 396 -667 430 -663
rect 396 -739 430 -731
rect 396 -811 430 -799
rect 396 -883 430 -867
rect 396 -955 430 -935
rect 396 -1027 430 -1003
rect 396 -1099 430 -1071
rect 396 -1171 430 -1139
rect 396 -1241 430 -1207
rect 396 -1309 430 -1277
rect 396 -1377 430 -1349
rect 396 -1445 430 -1421
rect 396 -1513 430 -1493
rect 396 -1581 430 -1565
rect 396 -1649 430 -1637
rect 396 -1717 430 -1709
rect 396 -1785 430 -1781
rect 396 -1891 430 -1887
rect 396 -1963 430 -1955
rect 396 -2035 430 -2023
rect 396 -2107 430 -2091
rect 396 -2179 430 -2159
rect 396 -2251 430 -2227
rect 396 -2323 430 -2295
rect 396 -2395 430 -2363
rect 396 -2465 430 -2431
rect 396 -2533 430 -2501
rect 396 -2601 430 -2573
rect 396 -2669 430 -2645
rect 396 -2737 430 -2717
rect 396 -2805 430 -2789
rect 396 -2873 430 -2861
rect 396 -2941 430 -2933
rect 396 -3009 430 -3005
rect 396 -3115 430 -3111
rect 396 -3187 430 -3179
rect 396 -3259 430 -3247
rect 396 -3331 430 -3315
rect 396 -3403 430 -3383
rect 396 -3475 430 -3451
rect 396 -3547 430 -3519
rect 396 -3619 430 -3587
rect 396 -3689 430 -3655
rect 396 -3757 430 -3725
rect 396 -3825 430 -3797
rect 396 -3893 430 -3869
rect 396 -3961 430 -3941
rect 396 -4029 430 -4013
rect 396 -4097 430 -4085
rect 396 -4165 430 -4157
rect 396 -4233 430 -4229
rect 396 -4339 430 -4335
rect 396 -4411 430 -4403
rect 396 -4483 430 -4471
rect 396 -4555 430 -4539
rect 396 -4627 430 -4607
rect 396 -4699 430 -4675
rect 396 -4771 430 -4743
rect 396 -4843 430 -4811
rect 396 -4913 430 -4879
rect 396 -4981 430 -4949
rect 396 -5049 430 -5021
rect 396 -5117 430 -5093
rect 396 -5185 430 -5165
rect 396 -5253 430 -5237
rect 396 -5321 430 -5309
rect 396 -5389 430 -5381
rect 396 -5457 430 -5453
rect 396 -5563 430 -5559
rect 396 -5635 430 -5627
rect 396 -5707 430 -5695
rect 396 -5779 430 -5763
rect 396 -5851 430 -5831
rect 396 -5923 430 -5899
rect 396 -5995 430 -5967
rect 396 -6067 430 -6035
rect 396 -6137 430 -6103
rect 396 -6205 430 -6173
rect 396 -6273 430 -6245
rect 396 -6341 430 -6317
rect 396 -6409 430 -6389
rect 396 -6477 430 -6461
rect 396 -6545 430 -6533
rect 396 -6613 430 -6605
rect 396 -6681 430 -6677
rect 396 -6787 430 -6783
rect 396 -6859 430 -6851
rect 396 -6931 430 -6919
rect 396 -7003 430 -6987
rect 396 -7075 430 -7055
rect 396 -7147 430 -7123
rect 396 -7219 430 -7191
rect 396 -7291 430 -7259
rect 396 -7361 430 -7327
rect 396 -7429 430 -7397
rect 396 -7497 430 -7469
rect 396 -7565 430 -7541
rect 396 -7633 430 -7613
rect 396 -7701 430 -7685
rect 396 -7769 430 -7757
rect 396 -7837 430 -7829
rect 396 -7905 430 -7901
rect 396 -8011 430 -8007
rect 396 -8083 430 -8075
rect 396 -8155 430 -8143
rect 396 -8227 430 -8211
rect 396 -8299 430 -8279
rect 396 -8371 430 -8347
rect 396 -8443 430 -8415
rect 396 -8515 430 -8483
rect 396 -8585 430 -8551
rect 396 -8653 430 -8621
rect 396 -8721 430 -8693
rect 396 -8789 430 -8765
rect 396 -8857 430 -8837
rect 396 -8925 430 -8909
rect 396 -8993 430 -8981
rect 396 -9061 430 -9053
rect 396 -9129 430 -9125
rect 396 -9235 430 -9231
rect 396 -9307 430 -9299
rect 396 -9379 430 -9367
rect 396 -9451 430 -9435
rect 396 -9523 430 -9503
rect 396 -9604 430 -9571
rect 514 9571 548 9604
rect 514 9503 548 9523
rect 514 9435 548 9451
rect 514 9367 548 9379
rect 514 9299 548 9307
rect 514 9231 548 9235
rect 514 9125 548 9129
rect 514 9053 548 9061
rect 514 8981 548 8993
rect 514 8909 548 8925
rect 514 8837 548 8857
rect 514 8765 548 8789
rect 514 8693 548 8721
rect 514 8621 548 8653
rect 514 8551 548 8585
rect 514 8483 548 8515
rect 514 8415 548 8443
rect 514 8347 548 8371
rect 514 8279 548 8299
rect 514 8211 548 8227
rect 514 8143 548 8155
rect 514 8075 548 8083
rect 514 8007 548 8011
rect 514 7901 548 7905
rect 514 7829 548 7837
rect 514 7757 548 7769
rect 514 7685 548 7701
rect 514 7613 548 7633
rect 514 7541 548 7565
rect 514 7469 548 7497
rect 514 7397 548 7429
rect 514 7327 548 7361
rect 514 7259 548 7291
rect 514 7191 548 7219
rect 514 7123 548 7147
rect 514 7055 548 7075
rect 514 6987 548 7003
rect 514 6919 548 6931
rect 514 6851 548 6859
rect 514 6783 548 6787
rect 514 6677 548 6681
rect 514 6605 548 6613
rect 514 6533 548 6545
rect 514 6461 548 6477
rect 514 6389 548 6409
rect 514 6317 548 6341
rect 514 6245 548 6273
rect 514 6173 548 6205
rect 514 6103 548 6137
rect 514 6035 548 6067
rect 514 5967 548 5995
rect 514 5899 548 5923
rect 514 5831 548 5851
rect 514 5763 548 5779
rect 514 5695 548 5707
rect 514 5627 548 5635
rect 514 5559 548 5563
rect 514 5453 548 5457
rect 514 5381 548 5389
rect 514 5309 548 5321
rect 514 5237 548 5253
rect 514 5165 548 5185
rect 514 5093 548 5117
rect 514 5021 548 5049
rect 514 4949 548 4981
rect 514 4879 548 4913
rect 514 4811 548 4843
rect 514 4743 548 4771
rect 514 4675 548 4699
rect 514 4607 548 4627
rect 514 4539 548 4555
rect 514 4471 548 4483
rect 514 4403 548 4411
rect 514 4335 548 4339
rect 514 4229 548 4233
rect 514 4157 548 4165
rect 514 4085 548 4097
rect 514 4013 548 4029
rect 514 3941 548 3961
rect 514 3869 548 3893
rect 514 3797 548 3825
rect 514 3725 548 3757
rect 514 3655 548 3689
rect 514 3587 548 3619
rect 514 3519 548 3547
rect 514 3451 548 3475
rect 514 3383 548 3403
rect 514 3315 548 3331
rect 514 3247 548 3259
rect 514 3179 548 3187
rect 514 3111 548 3115
rect 514 3005 548 3009
rect 514 2933 548 2941
rect 514 2861 548 2873
rect 514 2789 548 2805
rect 514 2717 548 2737
rect 514 2645 548 2669
rect 514 2573 548 2601
rect 514 2501 548 2533
rect 514 2431 548 2465
rect 514 2363 548 2395
rect 514 2295 548 2323
rect 514 2227 548 2251
rect 514 2159 548 2179
rect 514 2091 548 2107
rect 514 2023 548 2035
rect 514 1955 548 1963
rect 514 1887 548 1891
rect 514 1781 548 1785
rect 514 1709 548 1717
rect 514 1637 548 1649
rect 514 1565 548 1581
rect 514 1493 548 1513
rect 514 1421 548 1445
rect 514 1349 548 1377
rect 514 1277 548 1309
rect 514 1207 548 1241
rect 514 1139 548 1171
rect 514 1071 548 1099
rect 514 1003 548 1027
rect 514 935 548 955
rect 514 867 548 883
rect 514 799 548 811
rect 514 731 548 739
rect 514 663 548 667
rect 514 557 548 561
rect 514 485 548 493
rect 514 413 548 425
rect 514 341 548 357
rect 514 269 548 289
rect 514 197 548 221
rect 514 125 548 153
rect 514 53 548 85
rect 514 -17 548 17
rect 514 -85 548 -53
rect 514 -153 548 -125
rect 514 -221 548 -197
rect 514 -289 548 -269
rect 514 -357 548 -341
rect 514 -425 548 -413
rect 514 -493 548 -485
rect 514 -561 548 -557
rect 514 -667 548 -663
rect 514 -739 548 -731
rect 514 -811 548 -799
rect 514 -883 548 -867
rect 514 -955 548 -935
rect 514 -1027 548 -1003
rect 514 -1099 548 -1071
rect 514 -1171 548 -1139
rect 514 -1241 548 -1207
rect 514 -1309 548 -1277
rect 514 -1377 548 -1349
rect 514 -1445 548 -1421
rect 514 -1513 548 -1493
rect 514 -1581 548 -1565
rect 514 -1649 548 -1637
rect 514 -1717 548 -1709
rect 514 -1785 548 -1781
rect 514 -1891 548 -1887
rect 514 -1963 548 -1955
rect 514 -2035 548 -2023
rect 514 -2107 548 -2091
rect 514 -2179 548 -2159
rect 514 -2251 548 -2227
rect 514 -2323 548 -2295
rect 514 -2395 548 -2363
rect 514 -2465 548 -2431
rect 514 -2533 548 -2501
rect 514 -2601 548 -2573
rect 514 -2669 548 -2645
rect 514 -2737 548 -2717
rect 514 -2805 548 -2789
rect 514 -2873 548 -2861
rect 514 -2941 548 -2933
rect 514 -3009 548 -3005
rect 514 -3115 548 -3111
rect 514 -3187 548 -3179
rect 514 -3259 548 -3247
rect 514 -3331 548 -3315
rect 514 -3403 548 -3383
rect 514 -3475 548 -3451
rect 514 -3547 548 -3519
rect 514 -3619 548 -3587
rect 514 -3689 548 -3655
rect 514 -3757 548 -3725
rect 514 -3825 548 -3797
rect 514 -3893 548 -3869
rect 514 -3961 548 -3941
rect 514 -4029 548 -4013
rect 514 -4097 548 -4085
rect 514 -4165 548 -4157
rect 514 -4233 548 -4229
rect 514 -4339 548 -4335
rect 514 -4411 548 -4403
rect 514 -4483 548 -4471
rect 514 -4555 548 -4539
rect 514 -4627 548 -4607
rect 514 -4699 548 -4675
rect 514 -4771 548 -4743
rect 514 -4843 548 -4811
rect 514 -4913 548 -4879
rect 514 -4981 548 -4949
rect 514 -5049 548 -5021
rect 514 -5117 548 -5093
rect 514 -5185 548 -5165
rect 514 -5253 548 -5237
rect 514 -5321 548 -5309
rect 514 -5389 548 -5381
rect 514 -5457 548 -5453
rect 514 -5563 548 -5559
rect 514 -5635 548 -5627
rect 514 -5707 548 -5695
rect 514 -5779 548 -5763
rect 514 -5851 548 -5831
rect 514 -5923 548 -5899
rect 514 -5995 548 -5967
rect 514 -6067 548 -6035
rect 514 -6137 548 -6103
rect 514 -6205 548 -6173
rect 514 -6273 548 -6245
rect 514 -6341 548 -6317
rect 514 -6409 548 -6389
rect 514 -6477 548 -6461
rect 514 -6545 548 -6533
rect 514 -6613 548 -6605
rect 514 -6681 548 -6677
rect 514 -6787 548 -6783
rect 514 -6859 548 -6851
rect 514 -6931 548 -6919
rect 514 -7003 548 -6987
rect 514 -7075 548 -7055
rect 514 -7147 548 -7123
rect 514 -7219 548 -7191
rect 514 -7291 548 -7259
rect 514 -7361 548 -7327
rect 514 -7429 548 -7397
rect 514 -7497 548 -7469
rect 514 -7565 548 -7541
rect 514 -7633 548 -7613
rect 514 -7701 548 -7685
rect 514 -7769 548 -7757
rect 514 -7837 548 -7829
rect 514 -7905 548 -7901
rect 514 -8011 548 -8007
rect 514 -8083 548 -8075
rect 514 -8155 548 -8143
rect 514 -8227 548 -8211
rect 514 -8299 548 -8279
rect 514 -8371 548 -8347
rect 514 -8443 548 -8415
rect 514 -8515 548 -8483
rect 514 -8585 548 -8551
rect 514 -8653 548 -8621
rect 514 -8721 548 -8693
rect 514 -8789 548 -8765
rect 514 -8857 548 -8837
rect 514 -8925 548 -8909
rect 514 -8993 548 -8981
rect 514 -9061 548 -9053
rect 514 -9129 548 -9125
rect 514 -9235 548 -9231
rect 514 -9307 548 -9299
rect 514 -9379 548 -9367
rect 514 -9451 548 -9435
rect 514 -9523 548 -9503
rect 514 -9604 548 -9571
rect 632 9571 666 9604
rect 632 9503 666 9523
rect 632 9435 666 9451
rect 632 9367 666 9379
rect 632 9299 666 9307
rect 632 9231 666 9235
rect 632 9125 666 9129
rect 632 9053 666 9061
rect 632 8981 666 8993
rect 632 8909 666 8925
rect 632 8837 666 8857
rect 632 8765 666 8789
rect 632 8693 666 8721
rect 632 8621 666 8653
rect 632 8551 666 8585
rect 632 8483 666 8515
rect 632 8415 666 8443
rect 632 8347 666 8371
rect 632 8279 666 8299
rect 632 8211 666 8227
rect 632 8143 666 8155
rect 632 8075 666 8083
rect 632 8007 666 8011
rect 632 7901 666 7905
rect 632 7829 666 7837
rect 632 7757 666 7769
rect 632 7685 666 7701
rect 632 7613 666 7633
rect 632 7541 666 7565
rect 632 7469 666 7497
rect 632 7397 666 7429
rect 632 7327 666 7361
rect 632 7259 666 7291
rect 632 7191 666 7219
rect 632 7123 666 7147
rect 632 7055 666 7075
rect 632 6987 666 7003
rect 632 6919 666 6931
rect 632 6851 666 6859
rect 632 6783 666 6787
rect 632 6677 666 6681
rect 632 6605 666 6613
rect 632 6533 666 6545
rect 632 6461 666 6477
rect 632 6389 666 6409
rect 632 6317 666 6341
rect 632 6245 666 6273
rect 632 6173 666 6205
rect 632 6103 666 6137
rect 632 6035 666 6067
rect 632 5967 666 5995
rect 632 5899 666 5923
rect 632 5831 666 5851
rect 632 5763 666 5779
rect 632 5695 666 5707
rect 632 5627 666 5635
rect 632 5559 666 5563
rect 632 5453 666 5457
rect 632 5381 666 5389
rect 632 5309 666 5321
rect 632 5237 666 5253
rect 632 5165 666 5185
rect 632 5093 666 5117
rect 632 5021 666 5049
rect 632 4949 666 4981
rect 632 4879 666 4913
rect 632 4811 666 4843
rect 632 4743 666 4771
rect 632 4675 666 4699
rect 632 4607 666 4627
rect 632 4539 666 4555
rect 632 4471 666 4483
rect 632 4403 666 4411
rect 632 4335 666 4339
rect 632 4229 666 4233
rect 632 4157 666 4165
rect 632 4085 666 4097
rect 632 4013 666 4029
rect 632 3941 666 3961
rect 632 3869 666 3893
rect 632 3797 666 3825
rect 632 3725 666 3757
rect 632 3655 666 3689
rect 632 3587 666 3619
rect 632 3519 666 3547
rect 632 3451 666 3475
rect 632 3383 666 3403
rect 632 3315 666 3331
rect 632 3247 666 3259
rect 632 3179 666 3187
rect 632 3111 666 3115
rect 632 3005 666 3009
rect 632 2933 666 2941
rect 632 2861 666 2873
rect 632 2789 666 2805
rect 632 2717 666 2737
rect 632 2645 666 2669
rect 632 2573 666 2601
rect 632 2501 666 2533
rect 632 2431 666 2465
rect 632 2363 666 2395
rect 632 2295 666 2323
rect 632 2227 666 2251
rect 632 2159 666 2179
rect 632 2091 666 2107
rect 632 2023 666 2035
rect 632 1955 666 1963
rect 632 1887 666 1891
rect 632 1781 666 1785
rect 632 1709 666 1717
rect 632 1637 666 1649
rect 632 1565 666 1581
rect 632 1493 666 1513
rect 632 1421 666 1445
rect 632 1349 666 1377
rect 632 1277 666 1309
rect 632 1207 666 1241
rect 632 1139 666 1171
rect 632 1071 666 1099
rect 632 1003 666 1027
rect 632 935 666 955
rect 632 867 666 883
rect 632 799 666 811
rect 632 731 666 739
rect 632 663 666 667
rect 632 557 666 561
rect 632 485 666 493
rect 632 413 666 425
rect 632 341 666 357
rect 632 269 666 289
rect 632 197 666 221
rect 632 125 666 153
rect 632 53 666 85
rect 632 -17 666 17
rect 632 -85 666 -53
rect 632 -153 666 -125
rect 632 -221 666 -197
rect 632 -289 666 -269
rect 632 -357 666 -341
rect 632 -425 666 -413
rect 632 -493 666 -485
rect 632 -561 666 -557
rect 632 -667 666 -663
rect 632 -739 666 -731
rect 632 -811 666 -799
rect 632 -883 666 -867
rect 632 -955 666 -935
rect 632 -1027 666 -1003
rect 632 -1099 666 -1071
rect 632 -1171 666 -1139
rect 632 -1241 666 -1207
rect 632 -1309 666 -1277
rect 632 -1377 666 -1349
rect 632 -1445 666 -1421
rect 632 -1513 666 -1493
rect 632 -1581 666 -1565
rect 632 -1649 666 -1637
rect 632 -1717 666 -1709
rect 632 -1785 666 -1781
rect 632 -1891 666 -1887
rect 632 -1963 666 -1955
rect 632 -2035 666 -2023
rect 632 -2107 666 -2091
rect 632 -2179 666 -2159
rect 632 -2251 666 -2227
rect 632 -2323 666 -2295
rect 632 -2395 666 -2363
rect 632 -2465 666 -2431
rect 632 -2533 666 -2501
rect 632 -2601 666 -2573
rect 632 -2669 666 -2645
rect 632 -2737 666 -2717
rect 632 -2805 666 -2789
rect 632 -2873 666 -2861
rect 632 -2941 666 -2933
rect 632 -3009 666 -3005
rect 632 -3115 666 -3111
rect 632 -3187 666 -3179
rect 632 -3259 666 -3247
rect 632 -3331 666 -3315
rect 632 -3403 666 -3383
rect 632 -3475 666 -3451
rect 632 -3547 666 -3519
rect 632 -3619 666 -3587
rect 632 -3689 666 -3655
rect 632 -3757 666 -3725
rect 632 -3825 666 -3797
rect 632 -3893 666 -3869
rect 632 -3961 666 -3941
rect 632 -4029 666 -4013
rect 632 -4097 666 -4085
rect 632 -4165 666 -4157
rect 632 -4233 666 -4229
rect 632 -4339 666 -4335
rect 632 -4411 666 -4403
rect 632 -4483 666 -4471
rect 632 -4555 666 -4539
rect 632 -4627 666 -4607
rect 632 -4699 666 -4675
rect 632 -4771 666 -4743
rect 632 -4843 666 -4811
rect 632 -4913 666 -4879
rect 632 -4981 666 -4949
rect 632 -5049 666 -5021
rect 632 -5117 666 -5093
rect 632 -5185 666 -5165
rect 632 -5253 666 -5237
rect 632 -5321 666 -5309
rect 632 -5389 666 -5381
rect 632 -5457 666 -5453
rect 632 -5563 666 -5559
rect 632 -5635 666 -5627
rect 632 -5707 666 -5695
rect 632 -5779 666 -5763
rect 632 -5851 666 -5831
rect 632 -5923 666 -5899
rect 632 -5995 666 -5967
rect 632 -6067 666 -6035
rect 632 -6137 666 -6103
rect 632 -6205 666 -6173
rect 632 -6273 666 -6245
rect 632 -6341 666 -6317
rect 632 -6409 666 -6389
rect 632 -6477 666 -6461
rect 632 -6545 666 -6533
rect 632 -6613 666 -6605
rect 632 -6681 666 -6677
rect 632 -6787 666 -6783
rect 632 -6859 666 -6851
rect 632 -6931 666 -6919
rect 632 -7003 666 -6987
rect 632 -7075 666 -7055
rect 632 -7147 666 -7123
rect 632 -7219 666 -7191
rect 632 -7291 666 -7259
rect 632 -7361 666 -7327
rect 632 -7429 666 -7397
rect 632 -7497 666 -7469
rect 632 -7565 666 -7541
rect 632 -7633 666 -7613
rect 632 -7701 666 -7685
rect 632 -7769 666 -7757
rect 632 -7837 666 -7829
rect 632 -7905 666 -7901
rect 632 -8011 666 -8007
rect 632 -8083 666 -8075
rect 632 -8155 666 -8143
rect 632 -8227 666 -8211
rect 632 -8299 666 -8279
rect 632 -8371 666 -8347
rect 632 -8443 666 -8415
rect 632 -8515 666 -8483
rect 632 -8585 666 -8551
rect 632 -8653 666 -8621
rect 632 -8721 666 -8693
rect 632 -8789 666 -8765
rect 632 -8857 666 -8837
rect 632 -8925 666 -8909
rect 632 -8993 666 -8981
rect 632 -9061 666 -9053
rect 632 -9129 666 -9125
rect 632 -9235 666 -9231
rect 632 -9307 666 -9299
rect 632 -9379 666 -9367
rect 632 -9451 666 -9435
rect 632 -9523 666 -9503
rect 632 -9604 666 -9571
rect 750 9571 784 9604
rect 750 9503 784 9523
rect 750 9435 784 9451
rect 750 9367 784 9379
rect 750 9299 784 9307
rect 750 9231 784 9235
rect 750 9125 784 9129
rect 750 9053 784 9061
rect 750 8981 784 8993
rect 750 8909 784 8925
rect 750 8837 784 8857
rect 750 8765 784 8789
rect 750 8693 784 8721
rect 750 8621 784 8653
rect 750 8551 784 8585
rect 750 8483 784 8515
rect 750 8415 784 8443
rect 750 8347 784 8371
rect 750 8279 784 8299
rect 750 8211 784 8227
rect 750 8143 784 8155
rect 750 8075 784 8083
rect 750 8007 784 8011
rect 750 7901 784 7905
rect 750 7829 784 7837
rect 750 7757 784 7769
rect 750 7685 784 7701
rect 750 7613 784 7633
rect 750 7541 784 7565
rect 750 7469 784 7497
rect 750 7397 784 7429
rect 750 7327 784 7361
rect 750 7259 784 7291
rect 750 7191 784 7219
rect 750 7123 784 7147
rect 750 7055 784 7075
rect 750 6987 784 7003
rect 750 6919 784 6931
rect 750 6851 784 6859
rect 750 6783 784 6787
rect 750 6677 784 6681
rect 750 6605 784 6613
rect 750 6533 784 6545
rect 750 6461 784 6477
rect 750 6389 784 6409
rect 750 6317 784 6341
rect 750 6245 784 6273
rect 750 6173 784 6205
rect 750 6103 784 6137
rect 750 6035 784 6067
rect 750 5967 784 5995
rect 750 5899 784 5923
rect 750 5831 784 5851
rect 750 5763 784 5779
rect 750 5695 784 5707
rect 750 5627 784 5635
rect 750 5559 784 5563
rect 750 5453 784 5457
rect 750 5381 784 5389
rect 750 5309 784 5321
rect 750 5237 784 5253
rect 750 5165 784 5185
rect 750 5093 784 5117
rect 750 5021 784 5049
rect 750 4949 784 4981
rect 750 4879 784 4913
rect 750 4811 784 4843
rect 750 4743 784 4771
rect 750 4675 784 4699
rect 750 4607 784 4627
rect 750 4539 784 4555
rect 750 4471 784 4483
rect 750 4403 784 4411
rect 750 4335 784 4339
rect 750 4229 784 4233
rect 750 4157 784 4165
rect 750 4085 784 4097
rect 750 4013 784 4029
rect 750 3941 784 3961
rect 750 3869 784 3893
rect 750 3797 784 3825
rect 750 3725 784 3757
rect 750 3655 784 3689
rect 750 3587 784 3619
rect 750 3519 784 3547
rect 750 3451 784 3475
rect 750 3383 784 3403
rect 750 3315 784 3331
rect 750 3247 784 3259
rect 750 3179 784 3187
rect 750 3111 784 3115
rect 750 3005 784 3009
rect 750 2933 784 2941
rect 750 2861 784 2873
rect 750 2789 784 2805
rect 750 2717 784 2737
rect 750 2645 784 2669
rect 750 2573 784 2601
rect 750 2501 784 2533
rect 750 2431 784 2465
rect 750 2363 784 2395
rect 750 2295 784 2323
rect 750 2227 784 2251
rect 750 2159 784 2179
rect 750 2091 784 2107
rect 750 2023 784 2035
rect 750 1955 784 1963
rect 750 1887 784 1891
rect 750 1781 784 1785
rect 750 1709 784 1717
rect 750 1637 784 1649
rect 750 1565 784 1581
rect 750 1493 784 1513
rect 750 1421 784 1445
rect 750 1349 784 1377
rect 750 1277 784 1309
rect 750 1207 784 1241
rect 750 1139 784 1171
rect 750 1071 784 1099
rect 750 1003 784 1027
rect 750 935 784 955
rect 750 867 784 883
rect 750 799 784 811
rect 750 731 784 739
rect 750 663 784 667
rect 750 557 784 561
rect 750 485 784 493
rect 750 413 784 425
rect 750 341 784 357
rect 750 269 784 289
rect 750 197 784 221
rect 750 125 784 153
rect 750 53 784 85
rect 750 -17 784 17
rect 750 -85 784 -53
rect 750 -153 784 -125
rect 750 -221 784 -197
rect 750 -289 784 -269
rect 750 -357 784 -341
rect 750 -425 784 -413
rect 750 -493 784 -485
rect 750 -561 784 -557
rect 750 -667 784 -663
rect 750 -739 784 -731
rect 750 -811 784 -799
rect 750 -883 784 -867
rect 750 -955 784 -935
rect 750 -1027 784 -1003
rect 750 -1099 784 -1071
rect 750 -1171 784 -1139
rect 750 -1241 784 -1207
rect 750 -1309 784 -1277
rect 750 -1377 784 -1349
rect 750 -1445 784 -1421
rect 750 -1513 784 -1493
rect 750 -1581 784 -1565
rect 750 -1649 784 -1637
rect 750 -1717 784 -1709
rect 750 -1785 784 -1781
rect 750 -1891 784 -1887
rect 750 -1963 784 -1955
rect 750 -2035 784 -2023
rect 750 -2107 784 -2091
rect 750 -2179 784 -2159
rect 750 -2251 784 -2227
rect 750 -2323 784 -2295
rect 750 -2395 784 -2363
rect 750 -2465 784 -2431
rect 750 -2533 784 -2501
rect 750 -2601 784 -2573
rect 750 -2669 784 -2645
rect 750 -2737 784 -2717
rect 750 -2805 784 -2789
rect 750 -2873 784 -2861
rect 750 -2941 784 -2933
rect 750 -3009 784 -3005
rect 750 -3115 784 -3111
rect 750 -3187 784 -3179
rect 750 -3259 784 -3247
rect 750 -3331 784 -3315
rect 750 -3403 784 -3383
rect 750 -3475 784 -3451
rect 750 -3547 784 -3519
rect 750 -3619 784 -3587
rect 750 -3689 784 -3655
rect 750 -3757 784 -3725
rect 750 -3825 784 -3797
rect 750 -3893 784 -3869
rect 750 -3961 784 -3941
rect 750 -4029 784 -4013
rect 750 -4097 784 -4085
rect 750 -4165 784 -4157
rect 750 -4233 784 -4229
rect 750 -4339 784 -4335
rect 750 -4411 784 -4403
rect 750 -4483 784 -4471
rect 750 -4555 784 -4539
rect 750 -4627 784 -4607
rect 750 -4699 784 -4675
rect 750 -4771 784 -4743
rect 750 -4843 784 -4811
rect 750 -4913 784 -4879
rect 750 -4981 784 -4949
rect 750 -5049 784 -5021
rect 750 -5117 784 -5093
rect 750 -5185 784 -5165
rect 750 -5253 784 -5237
rect 750 -5321 784 -5309
rect 750 -5389 784 -5381
rect 750 -5457 784 -5453
rect 750 -5563 784 -5559
rect 750 -5635 784 -5627
rect 750 -5707 784 -5695
rect 750 -5779 784 -5763
rect 750 -5851 784 -5831
rect 750 -5923 784 -5899
rect 750 -5995 784 -5967
rect 750 -6067 784 -6035
rect 750 -6137 784 -6103
rect 750 -6205 784 -6173
rect 750 -6273 784 -6245
rect 750 -6341 784 -6317
rect 750 -6409 784 -6389
rect 750 -6477 784 -6461
rect 750 -6545 784 -6533
rect 750 -6613 784 -6605
rect 750 -6681 784 -6677
rect 750 -6787 784 -6783
rect 750 -6859 784 -6851
rect 750 -6931 784 -6919
rect 750 -7003 784 -6987
rect 750 -7075 784 -7055
rect 750 -7147 784 -7123
rect 750 -7219 784 -7191
rect 750 -7291 784 -7259
rect 750 -7361 784 -7327
rect 750 -7429 784 -7397
rect 750 -7497 784 -7469
rect 750 -7565 784 -7541
rect 750 -7633 784 -7613
rect 750 -7701 784 -7685
rect 750 -7769 784 -7757
rect 750 -7837 784 -7829
rect 750 -7905 784 -7901
rect 750 -8011 784 -8007
rect 750 -8083 784 -8075
rect 750 -8155 784 -8143
rect 750 -8227 784 -8211
rect 750 -8299 784 -8279
rect 750 -8371 784 -8347
rect 750 -8443 784 -8415
rect 750 -8515 784 -8483
rect 750 -8585 784 -8551
rect 750 -8653 784 -8621
rect 750 -8721 784 -8693
rect 750 -8789 784 -8765
rect 750 -8857 784 -8837
rect 750 -8925 784 -8909
rect 750 -8993 784 -8981
rect 750 -9061 784 -9053
rect 750 -9129 784 -9125
rect 750 -9235 784 -9231
rect 750 -9307 784 -9299
rect 750 -9379 784 -9367
rect 750 -9451 784 -9435
rect 750 -9523 784 -9503
rect 750 -9604 784 -9571
rect 868 9571 902 9604
rect 868 9503 902 9523
rect 868 9435 902 9451
rect 868 9367 902 9379
rect 868 9299 902 9307
rect 868 9231 902 9235
rect 868 9125 902 9129
rect 868 9053 902 9061
rect 868 8981 902 8993
rect 868 8909 902 8925
rect 868 8837 902 8857
rect 868 8765 902 8789
rect 868 8693 902 8721
rect 868 8621 902 8653
rect 868 8551 902 8585
rect 868 8483 902 8515
rect 868 8415 902 8443
rect 868 8347 902 8371
rect 868 8279 902 8299
rect 868 8211 902 8227
rect 868 8143 902 8155
rect 868 8075 902 8083
rect 868 8007 902 8011
rect 868 7901 902 7905
rect 868 7829 902 7837
rect 868 7757 902 7769
rect 868 7685 902 7701
rect 868 7613 902 7633
rect 868 7541 902 7565
rect 868 7469 902 7497
rect 868 7397 902 7429
rect 868 7327 902 7361
rect 868 7259 902 7291
rect 868 7191 902 7219
rect 868 7123 902 7147
rect 868 7055 902 7075
rect 868 6987 902 7003
rect 868 6919 902 6931
rect 868 6851 902 6859
rect 868 6783 902 6787
rect 868 6677 902 6681
rect 868 6605 902 6613
rect 868 6533 902 6545
rect 868 6461 902 6477
rect 868 6389 902 6409
rect 868 6317 902 6341
rect 868 6245 902 6273
rect 868 6173 902 6205
rect 868 6103 902 6137
rect 868 6035 902 6067
rect 868 5967 902 5995
rect 868 5899 902 5923
rect 868 5831 902 5851
rect 868 5763 902 5779
rect 868 5695 902 5707
rect 868 5627 902 5635
rect 868 5559 902 5563
rect 868 5453 902 5457
rect 868 5381 902 5389
rect 868 5309 902 5321
rect 868 5237 902 5253
rect 868 5165 902 5185
rect 868 5093 902 5117
rect 868 5021 902 5049
rect 868 4949 902 4981
rect 868 4879 902 4913
rect 868 4811 902 4843
rect 868 4743 902 4771
rect 868 4675 902 4699
rect 868 4607 902 4627
rect 868 4539 902 4555
rect 868 4471 902 4483
rect 868 4403 902 4411
rect 868 4335 902 4339
rect 868 4229 902 4233
rect 868 4157 902 4165
rect 868 4085 902 4097
rect 868 4013 902 4029
rect 868 3941 902 3961
rect 868 3869 902 3893
rect 868 3797 902 3825
rect 868 3725 902 3757
rect 868 3655 902 3689
rect 868 3587 902 3619
rect 868 3519 902 3547
rect 868 3451 902 3475
rect 868 3383 902 3403
rect 868 3315 902 3331
rect 868 3247 902 3259
rect 868 3179 902 3187
rect 868 3111 902 3115
rect 868 3005 902 3009
rect 868 2933 902 2941
rect 868 2861 902 2873
rect 868 2789 902 2805
rect 868 2717 902 2737
rect 868 2645 902 2669
rect 868 2573 902 2601
rect 868 2501 902 2533
rect 868 2431 902 2465
rect 868 2363 902 2395
rect 868 2295 902 2323
rect 868 2227 902 2251
rect 868 2159 902 2179
rect 868 2091 902 2107
rect 868 2023 902 2035
rect 868 1955 902 1963
rect 868 1887 902 1891
rect 868 1781 902 1785
rect 868 1709 902 1717
rect 868 1637 902 1649
rect 868 1565 902 1581
rect 868 1493 902 1513
rect 868 1421 902 1445
rect 868 1349 902 1377
rect 868 1277 902 1309
rect 868 1207 902 1241
rect 868 1139 902 1171
rect 868 1071 902 1099
rect 868 1003 902 1027
rect 868 935 902 955
rect 868 867 902 883
rect 868 799 902 811
rect 868 731 902 739
rect 868 663 902 667
rect 868 557 902 561
rect 868 485 902 493
rect 868 413 902 425
rect 868 341 902 357
rect 868 269 902 289
rect 868 197 902 221
rect 868 125 902 153
rect 868 53 902 85
rect 868 -17 902 17
rect 868 -85 902 -53
rect 868 -153 902 -125
rect 868 -221 902 -197
rect 868 -289 902 -269
rect 868 -357 902 -341
rect 868 -425 902 -413
rect 868 -493 902 -485
rect 868 -561 902 -557
rect 868 -667 902 -663
rect 868 -739 902 -731
rect 868 -811 902 -799
rect 868 -883 902 -867
rect 868 -955 902 -935
rect 868 -1027 902 -1003
rect 868 -1099 902 -1071
rect 868 -1171 902 -1139
rect 868 -1241 902 -1207
rect 868 -1309 902 -1277
rect 868 -1377 902 -1349
rect 868 -1445 902 -1421
rect 868 -1513 902 -1493
rect 868 -1581 902 -1565
rect 868 -1649 902 -1637
rect 868 -1717 902 -1709
rect 868 -1785 902 -1781
rect 868 -1891 902 -1887
rect 868 -1963 902 -1955
rect 868 -2035 902 -2023
rect 868 -2107 902 -2091
rect 868 -2179 902 -2159
rect 868 -2251 902 -2227
rect 868 -2323 902 -2295
rect 868 -2395 902 -2363
rect 868 -2465 902 -2431
rect 868 -2533 902 -2501
rect 868 -2601 902 -2573
rect 868 -2669 902 -2645
rect 868 -2737 902 -2717
rect 868 -2805 902 -2789
rect 868 -2873 902 -2861
rect 868 -2941 902 -2933
rect 868 -3009 902 -3005
rect 868 -3115 902 -3111
rect 868 -3187 902 -3179
rect 868 -3259 902 -3247
rect 868 -3331 902 -3315
rect 868 -3403 902 -3383
rect 868 -3475 902 -3451
rect 868 -3547 902 -3519
rect 868 -3619 902 -3587
rect 868 -3689 902 -3655
rect 868 -3757 902 -3725
rect 868 -3825 902 -3797
rect 868 -3893 902 -3869
rect 868 -3961 902 -3941
rect 868 -4029 902 -4013
rect 868 -4097 902 -4085
rect 868 -4165 902 -4157
rect 868 -4233 902 -4229
rect 868 -4339 902 -4335
rect 868 -4411 902 -4403
rect 868 -4483 902 -4471
rect 868 -4555 902 -4539
rect 868 -4627 902 -4607
rect 868 -4699 902 -4675
rect 868 -4771 902 -4743
rect 868 -4843 902 -4811
rect 868 -4913 902 -4879
rect 868 -4981 902 -4949
rect 868 -5049 902 -5021
rect 868 -5117 902 -5093
rect 868 -5185 902 -5165
rect 868 -5253 902 -5237
rect 868 -5321 902 -5309
rect 868 -5389 902 -5381
rect 868 -5457 902 -5453
rect 868 -5563 902 -5559
rect 868 -5635 902 -5627
rect 868 -5707 902 -5695
rect 868 -5779 902 -5763
rect 868 -5851 902 -5831
rect 868 -5923 902 -5899
rect 868 -5995 902 -5967
rect 868 -6067 902 -6035
rect 868 -6137 902 -6103
rect 868 -6205 902 -6173
rect 868 -6273 902 -6245
rect 868 -6341 902 -6317
rect 868 -6409 902 -6389
rect 868 -6477 902 -6461
rect 868 -6545 902 -6533
rect 868 -6613 902 -6605
rect 868 -6681 902 -6677
rect 868 -6787 902 -6783
rect 868 -6859 902 -6851
rect 868 -6931 902 -6919
rect 868 -7003 902 -6987
rect 868 -7075 902 -7055
rect 868 -7147 902 -7123
rect 868 -7219 902 -7191
rect 868 -7291 902 -7259
rect 868 -7361 902 -7327
rect 868 -7429 902 -7397
rect 868 -7497 902 -7469
rect 868 -7565 902 -7541
rect 868 -7633 902 -7613
rect 868 -7701 902 -7685
rect 868 -7769 902 -7757
rect 868 -7837 902 -7829
rect 868 -7905 902 -7901
rect 868 -8011 902 -8007
rect 868 -8083 902 -8075
rect 868 -8155 902 -8143
rect 868 -8227 902 -8211
rect 868 -8299 902 -8279
rect 868 -8371 902 -8347
rect 868 -8443 902 -8415
rect 868 -8515 902 -8483
rect 868 -8585 902 -8551
rect 868 -8653 902 -8621
rect 868 -8721 902 -8693
rect 868 -8789 902 -8765
rect 868 -8857 902 -8837
rect 868 -8925 902 -8909
rect 868 -8993 902 -8981
rect 868 -9061 902 -9053
rect 868 -9129 902 -9125
rect 868 -9235 902 -9231
rect 868 -9307 902 -9299
rect 868 -9379 902 -9367
rect 868 -9451 902 -9435
rect 868 -9523 902 -9503
rect 868 -9604 902 -9571
rect 986 9571 1020 9604
rect 986 9503 1020 9523
rect 986 9435 1020 9451
rect 986 9367 1020 9379
rect 986 9299 1020 9307
rect 986 9231 1020 9235
rect 986 9125 1020 9129
rect 986 9053 1020 9061
rect 986 8981 1020 8993
rect 986 8909 1020 8925
rect 986 8837 1020 8857
rect 986 8765 1020 8789
rect 986 8693 1020 8721
rect 986 8621 1020 8653
rect 986 8551 1020 8585
rect 986 8483 1020 8515
rect 986 8415 1020 8443
rect 986 8347 1020 8371
rect 986 8279 1020 8299
rect 986 8211 1020 8227
rect 986 8143 1020 8155
rect 986 8075 1020 8083
rect 986 8007 1020 8011
rect 986 7901 1020 7905
rect 986 7829 1020 7837
rect 986 7757 1020 7769
rect 986 7685 1020 7701
rect 986 7613 1020 7633
rect 986 7541 1020 7565
rect 986 7469 1020 7497
rect 986 7397 1020 7429
rect 986 7327 1020 7361
rect 986 7259 1020 7291
rect 986 7191 1020 7219
rect 986 7123 1020 7147
rect 986 7055 1020 7075
rect 986 6987 1020 7003
rect 986 6919 1020 6931
rect 986 6851 1020 6859
rect 986 6783 1020 6787
rect 986 6677 1020 6681
rect 986 6605 1020 6613
rect 986 6533 1020 6545
rect 986 6461 1020 6477
rect 986 6389 1020 6409
rect 986 6317 1020 6341
rect 986 6245 1020 6273
rect 986 6173 1020 6205
rect 986 6103 1020 6137
rect 986 6035 1020 6067
rect 986 5967 1020 5995
rect 986 5899 1020 5923
rect 986 5831 1020 5851
rect 986 5763 1020 5779
rect 986 5695 1020 5707
rect 986 5627 1020 5635
rect 986 5559 1020 5563
rect 986 5453 1020 5457
rect 986 5381 1020 5389
rect 986 5309 1020 5321
rect 986 5237 1020 5253
rect 986 5165 1020 5185
rect 986 5093 1020 5117
rect 986 5021 1020 5049
rect 986 4949 1020 4981
rect 986 4879 1020 4913
rect 986 4811 1020 4843
rect 986 4743 1020 4771
rect 986 4675 1020 4699
rect 986 4607 1020 4627
rect 986 4539 1020 4555
rect 986 4471 1020 4483
rect 986 4403 1020 4411
rect 986 4335 1020 4339
rect 986 4229 1020 4233
rect 986 4157 1020 4165
rect 986 4085 1020 4097
rect 986 4013 1020 4029
rect 986 3941 1020 3961
rect 986 3869 1020 3893
rect 986 3797 1020 3825
rect 986 3725 1020 3757
rect 986 3655 1020 3689
rect 986 3587 1020 3619
rect 986 3519 1020 3547
rect 986 3451 1020 3475
rect 986 3383 1020 3403
rect 986 3315 1020 3331
rect 986 3247 1020 3259
rect 986 3179 1020 3187
rect 986 3111 1020 3115
rect 986 3005 1020 3009
rect 986 2933 1020 2941
rect 986 2861 1020 2873
rect 986 2789 1020 2805
rect 986 2717 1020 2737
rect 986 2645 1020 2669
rect 986 2573 1020 2601
rect 986 2501 1020 2533
rect 986 2431 1020 2465
rect 986 2363 1020 2395
rect 986 2295 1020 2323
rect 986 2227 1020 2251
rect 986 2159 1020 2179
rect 986 2091 1020 2107
rect 986 2023 1020 2035
rect 986 1955 1020 1963
rect 986 1887 1020 1891
rect 986 1781 1020 1785
rect 986 1709 1020 1717
rect 986 1637 1020 1649
rect 986 1565 1020 1581
rect 986 1493 1020 1513
rect 986 1421 1020 1445
rect 986 1349 1020 1377
rect 986 1277 1020 1309
rect 986 1207 1020 1241
rect 986 1139 1020 1171
rect 986 1071 1020 1099
rect 986 1003 1020 1027
rect 986 935 1020 955
rect 986 867 1020 883
rect 986 799 1020 811
rect 986 731 1020 739
rect 986 663 1020 667
rect 986 557 1020 561
rect 986 485 1020 493
rect 986 413 1020 425
rect 986 341 1020 357
rect 986 269 1020 289
rect 986 197 1020 221
rect 986 125 1020 153
rect 986 53 1020 85
rect 986 -17 1020 17
rect 986 -85 1020 -53
rect 986 -153 1020 -125
rect 986 -221 1020 -197
rect 986 -289 1020 -269
rect 986 -357 1020 -341
rect 986 -425 1020 -413
rect 986 -493 1020 -485
rect 986 -561 1020 -557
rect 986 -667 1020 -663
rect 986 -739 1020 -731
rect 986 -811 1020 -799
rect 986 -883 1020 -867
rect 986 -955 1020 -935
rect 986 -1027 1020 -1003
rect 986 -1099 1020 -1071
rect 986 -1171 1020 -1139
rect 986 -1241 1020 -1207
rect 986 -1309 1020 -1277
rect 986 -1377 1020 -1349
rect 986 -1445 1020 -1421
rect 986 -1513 1020 -1493
rect 986 -1581 1020 -1565
rect 986 -1649 1020 -1637
rect 986 -1717 1020 -1709
rect 986 -1785 1020 -1781
rect 986 -1891 1020 -1887
rect 986 -1963 1020 -1955
rect 986 -2035 1020 -2023
rect 986 -2107 1020 -2091
rect 986 -2179 1020 -2159
rect 986 -2251 1020 -2227
rect 986 -2323 1020 -2295
rect 986 -2395 1020 -2363
rect 986 -2465 1020 -2431
rect 986 -2533 1020 -2501
rect 986 -2601 1020 -2573
rect 986 -2669 1020 -2645
rect 986 -2737 1020 -2717
rect 986 -2805 1020 -2789
rect 986 -2873 1020 -2861
rect 986 -2941 1020 -2933
rect 986 -3009 1020 -3005
rect 986 -3115 1020 -3111
rect 986 -3187 1020 -3179
rect 986 -3259 1020 -3247
rect 986 -3331 1020 -3315
rect 986 -3403 1020 -3383
rect 986 -3475 1020 -3451
rect 986 -3547 1020 -3519
rect 986 -3619 1020 -3587
rect 986 -3689 1020 -3655
rect 986 -3757 1020 -3725
rect 986 -3825 1020 -3797
rect 986 -3893 1020 -3869
rect 986 -3961 1020 -3941
rect 986 -4029 1020 -4013
rect 986 -4097 1020 -4085
rect 986 -4165 1020 -4157
rect 986 -4233 1020 -4229
rect 986 -4339 1020 -4335
rect 986 -4411 1020 -4403
rect 986 -4483 1020 -4471
rect 986 -4555 1020 -4539
rect 986 -4627 1020 -4607
rect 986 -4699 1020 -4675
rect 986 -4771 1020 -4743
rect 986 -4843 1020 -4811
rect 986 -4913 1020 -4879
rect 986 -4981 1020 -4949
rect 986 -5049 1020 -5021
rect 986 -5117 1020 -5093
rect 986 -5185 1020 -5165
rect 986 -5253 1020 -5237
rect 986 -5321 1020 -5309
rect 986 -5389 1020 -5381
rect 986 -5457 1020 -5453
rect 986 -5563 1020 -5559
rect 986 -5635 1020 -5627
rect 986 -5707 1020 -5695
rect 986 -5779 1020 -5763
rect 986 -5851 1020 -5831
rect 986 -5923 1020 -5899
rect 986 -5995 1020 -5967
rect 986 -6067 1020 -6035
rect 986 -6137 1020 -6103
rect 986 -6205 1020 -6173
rect 986 -6273 1020 -6245
rect 986 -6341 1020 -6317
rect 986 -6409 1020 -6389
rect 986 -6477 1020 -6461
rect 986 -6545 1020 -6533
rect 986 -6613 1020 -6605
rect 986 -6681 1020 -6677
rect 986 -6787 1020 -6783
rect 986 -6859 1020 -6851
rect 986 -6931 1020 -6919
rect 986 -7003 1020 -6987
rect 986 -7075 1020 -7055
rect 986 -7147 1020 -7123
rect 986 -7219 1020 -7191
rect 986 -7291 1020 -7259
rect 986 -7361 1020 -7327
rect 986 -7429 1020 -7397
rect 986 -7497 1020 -7469
rect 986 -7565 1020 -7541
rect 986 -7633 1020 -7613
rect 986 -7701 1020 -7685
rect 986 -7769 1020 -7757
rect 986 -7837 1020 -7829
rect 986 -7905 1020 -7901
rect 986 -8011 1020 -8007
rect 986 -8083 1020 -8075
rect 986 -8155 1020 -8143
rect 986 -8227 1020 -8211
rect 986 -8299 1020 -8279
rect 986 -8371 1020 -8347
rect 986 -8443 1020 -8415
rect 986 -8515 1020 -8483
rect 986 -8585 1020 -8551
rect 986 -8653 1020 -8621
rect 986 -8721 1020 -8693
rect 986 -8789 1020 -8765
rect 986 -8857 1020 -8837
rect 986 -8925 1020 -8909
rect 986 -8993 1020 -8981
rect 986 -9061 1020 -9053
rect 986 -9129 1020 -9125
rect 986 -9235 1020 -9231
rect 986 -9307 1020 -9299
rect 986 -9379 1020 -9367
rect 986 -9451 1020 -9435
rect 986 -9523 1020 -9503
rect 986 -9604 1020 -9571
rect 1104 9571 1138 9604
rect 1104 9503 1138 9523
rect 1104 9435 1138 9451
rect 1104 9367 1138 9379
rect 1104 9299 1138 9307
rect 1104 9231 1138 9235
rect 1104 9125 1138 9129
rect 1104 9053 1138 9061
rect 1104 8981 1138 8993
rect 1104 8909 1138 8925
rect 1104 8837 1138 8857
rect 1104 8765 1138 8789
rect 1104 8693 1138 8721
rect 1104 8621 1138 8653
rect 1104 8551 1138 8585
rect 1104 8483 1138 8515
rect 1104 8415 1138 8443
rect 1104 8347 1138 8371
rect 1104 8279 1138 8299
rect 1104 8211 1138 8227
rect 1104 8143 1138 8155
rect 1104 8075 1138 8083
rect 1104 8007 1138 8011
rect 1104 7901 1138 7905
rect 1104 7829 1138 7837
rect 1104 7757 1138 7769
rect 1104 7685 1138 7701
rect 1104 7613 1138 7633
rect 1104 7541 1138 7565
rect 1104 7469 1138 7497
rect 1104 7397 1138 7429
rect 1104 7327 1138 7361
rect 1104 7259 1138 7291
rect 1104 7191 1138 7219
rect 1104 7123 1138 7147
rect 1104 7055 1138 7075
rect 1104 6987 1138 7003
rect 1104 6919 1138 6931
rect 1104 6851 1138 6859
rect 1104 6783 1138 6787
rect 1104 6677 1138 6681
rect 1104 6605 1138 6613
rect 1104 6533 1138 6545
rect 1104 6461 1138 6477
rect 1104 6389 1138 6409
rect 1104 6317 1138 6341
rect 1104 6245 1138 6273
rect 1104 6173 1138 6205
rect 1104 6103 1138 6137
rect 1104 6035 1138 6067
rect 1104 5967 1138 5995
rect 1104 5899 1138 5923
rect 1104 5831 1138 5851
rect 1104 5763 1138 5779
rect 1104 5695 1138 5707
rect 1104 5627 1138 5635
rect 1104 5559 1138 5563
rect 1104 5453 1138 5457
rect 1104 5381 1138 5389
rect 1104 5309 1138 5321
rect 1104 5237 1138 5253
rect 1104 5165 1138 5185
rect 1104 5093 1138 5117
rect 1104 5021 1138 5049
rect 1104 4949 1138 4981
rect 1104 4879 1138 4913
rect 1104 4811 1138 4843
rect 1104 4743 1138 4771
rect 1104 4675 1138 4699
rect 1104 4607 1138 4627
rect 1104 4539 1138 4555
rect 1104 4471 1138 4483
rect 1104 4403 1138 4411
rect 1104 4335 1138 4339
rect 1104 4229 1138 4233
rect 1104 4157 1138 4165
rect 1104 4085 1138 4097
rect 1104 4013 1138 4029
rect 1104 3941 1138 3961
rect 1104 3869 1138 3893
rect 1104 3797 1138 3825
rect 1104 3725 1138 3757
rect 1104 3655 1138 3689
rect 1104 3587 1138 3619
rect 1104 3519 1138 3547
rect 1104 3451 1138 3475
rect 1104 3383 1138 3403
rect 1104 3315 1138 3331
rect 1104 3247 1138 3259
rect 1104 3179 1138 3187
rect 1104 3111 1138 3115
rect 1104 3005 1138 3009
rect 1104 2933 1138 2941
rect 1104 2861 1138 2873
rect 1104 2789 1138 2805
rect 1104 2717 1138 2737
rect 1104 2645 1138 2669
rect 1104 2573 1138 2601
rect 1104 2501 1138 2533
rect 1104 2431 1138 2465
rect 1104 2363 1138 2395
rect 1104 2295 1138 2323
rect 1104 2227 1138 2251
rect 1104 2159 1138 2179
rect 1104 2091 1138 2107
rect 1104 2023 1138 2035
rect 1104 1955 1138 1963
rect 1104 1887 1138 1891
rect 1104 1781 1138 1785
rect 1104 1709 1138 1717
rect 1104 1637 1138 1649
rect 1104 1565 1138 1581
rect 1104 1493 1138 1513
rect 1104 1421 1138 1445
rect 1104 1349 1138 1377
rect 1104 1277 1138 1309
rect 1104 1207 1138 1241
rect 1104 1139 1138 1171
rect 1104 1071 1138 1099
rect 1104 1003 1138 1027
rect 1104 935 1138 955
rect 1104 867 1138 883
rect 1104 799 1138 811
rect 1104 731 1138 739
rect 1104 663 1138 667
rect 1104 557 1138 561
rect 1104 485 1138 493
rect 1104 413 1138 425
rect 1104 341 1138 357
rect 1104 269 1138 289
rect 1104 197 1138 221
rect 1104 125 1138 153
rect 1104 53 1138 85
rect 1104 -17 1138 17
rect 1104 -85 1138 -53
rect 1104 -153 1138 -125
rect 1104 -221 1138 -197
rect 1104 -289 1138 -269
rect 1104 -357 1138 -341
rect 1104 -425 1138 -413
rect 1104 -493 1138 -485
rect 1104 -561 1138 -557
rect 1104 -667 1138 -663
rect 1104 -739 1138 -731
rect 1104 -811 1138 -799
rect 1104 -883 1138 -867
rect 1104 -955 1138 -935
rect 1104 -1027 1138 -1003
rect 1104 -1099 1138 -1071
rect 1104 -1171 1138 -1139
rect 1104 -1241 1138 -1207
rect 1104 -1309 1138 -1277
rect 1104 -1377 1138 -1349
rect 1104 -1445 1138 -1421
rect 1104 -1513 1138 -1493
rect 1104 -1581 1138 -1565
rect 1104 -1649 1138 -1637
rect 1104 -1717 1138 -1709
rect 1104 -1785 1138 -1781
rect 1104 -1891 1138 -1887
rect 1104 -1963 1138 -1955
rect 1104 -2035 1138 -2023
rect 1104 -2107 1138 -2091
rect 1104 -2179 1138 -2159
rect 1104 -2251 1138 -2227
rect 1104 -2323 1138 -2295
rect 1104 -2395 1138 -2363
rect 1104 -2465 1138 -2431
rect 1104 -2533 1138 -2501
rect 1104 -2601 1138 -2573
rect 1104 -2669 1138 -2645
rect 1104 -2737 1138 -2717
rect 1104 -2805 1138 -2789
rect 1104 -2873 1138 -2861
rect 1104 -2941 1138 -2933
rect 1104 -3009 1138 -3005
rect 1104 -3115 1138 -3111
rect 1104 -3187 1138 -3179
rect 1104 -3259 1138 -3247
rect 1104 -3331 1138 -3315
rect 1104 -3403 1138 -3383
rect 1104 -3475 1138 -3451
rect 1104 -3547 1138 -3519
rect 1104 -3619 1138 -3587
rect 1104 -3689 1138 -3655
rect 1104 -3757 1138 -3725
rect 1104 -3825 1138 -3797
rect 1104 -3893 1138 -3869
rect 1104 -3961 1138 -3941
rect 1104 -4029 1138 -4013
rect 1104 -4097 1138 -4085
rect 1104 -4165 1138 -4157
rect 1104 -4233 1138 -4229
rect 1104 -4339 1138 -4335
rect 1104 -4411 1138 -4403
rect 1104 -4483 1138 -4471
rect 1104 -4555 1138 -4539
rect 1104 -4627 1138 -4607
rect 1104 -4699 1138 -4675
rect 1104 -4771 1138 -4743
rect 1104 -4843 1138 -4811
rect 1104 -4913 1138 -4879
rect 1104 -4981 1138 -4949
rect 1104 -5049 1138 -5021
rect 1104 -5117 1138 -5093
rect 1104 -5185 1138 -5165
rect 1104 -5253 1138 -5237
rect 1104 -5321 1138 -5309
rect 1104 -5389 1138 -5381
rect 1104 -5457 1138 -5453
rect 1104 -5563 1138 -5559
rect 1104 -5635 1138 -5627
rect 1104 -5707 1138 -5695
rect 1104 -5779 1138 -5763
rect 1104 -5851 1138 -5831
rect 1104 -5923 1138 -5899
rect 1104 -5995 1138 -5967
rect 1104 -6067 1138 -6035
rect 1104 -6137 1138 -6103
rect 1104 -6205 1138 -6173
rect 1104 -6273 1138 -6245
rect 1104 -6341 1138 -6317
rect 1104 -6409 1138 -6389
rect 1104 -6477 1138 -6461
rect 1104 -6545 1138 -6533
rect 1104 -6613 1138 -6605
rect 1104 -6681 1138 -6677
rect 1104 -6787 1138 -6783
rect 1104 -6859 1138 -6851
rect 1104 -6931 1138 -6919
rect 1104 -7003 1138 -6987
rect 1104 -7075 1138 -7055
rect 1104 -7147 1138 -7123
rect 1104 -7219 1138 -7191
rect 1104 -7291 1138 -7259
rect 1104 -7361 1138 -7327
rect 1104 -7429 1138 -7397
rect 1104 -7497 1138 -7469
rect 1104 -7565 1138 -7541
rect 1104 -7633 1138 -7613
rect 1104 -7701 1138 -7685
rect 1104 -7769 1138 -7757
rect 1104 -7837 1138 -7829
rect 1104 -7905 1138 -7901
rect 1104 -8011 1138 -8007
rect 1104 -8083 1138 -8075
rect 1104 -8155 1138 -8143
rect 1104 -8227 1138 -8211
rect 1104 -8299 1138 -8279
rect 1104 -8371 1138 -8347
rect 1104 -8443 1138 -8415
rect 1104 -8515 1138 -8483
rect 1104 -8585 1138 -8551
rect 1104 -8653 1138 -8621
rect 1104 -8721 1138 -8693
rect 1104 -8789 1138 -8765
rect 1104 -8857 1138 -8837
rect 1104 -8925 1138 -8909
rect 1104 -8993 1138 -8981
rect 1104 -9061 1138 -9053
rect 1104 -9129 1138 -9125
rect 1104 -9235 1138 -9231
rect 1104 -9307 1138 -9299
rect 1104 -9379 1138 -9367
rect 1104 -9451 1138 -9435
rect 1104 -9523 1138 -9503
rect 1104 -9604 1138 -9571
rect 1222 9571 1256 9604
rect 1222 9503 1256 9523
rect 1222 9435 1256 9451
rect 1222 9367 1256 9379
rect 1222 9299 1256 9307
rect 1222 9231 1256 9235
rect 1222 9125 1256 9129
rect 1222 9053 1256 9061
rect 1222 8981 1256 8993
rect 1222 8909 1256 8925
rect 1222 8837 1256 8857
rect 1222 8765 1256 8789
rect 1222 8693 1256 8721
rect 1222 8621 1256 8653
rect 1222 8551 1256 8585
rect 1222 8483 1256 8515
rect 1222 8415 1256 8443
rect 1222 8347 1256 8371
rect 1222 8279 1256 8299
rect 1222 8211 1256 8227
rect 1222 8143 1256 8155
rect 1222 8075 1256 8083
rect 1222 8007 1256 8011
rect 1222 7901 1256 7905
rect 1222 7829 1256 7837
rect 1222 7757 1256 7769
rect 1222 7685 1256 7701
rect 1222 7613 1256 7633
rect 1222 7541 1256 7565
rect 1222 7469 1256 7497
rect 1222 7397 1256 7429
rect 1222 7327 1256 7361
rect 1222 7259 1256 7291
rect 1222 7191 1256 7219
rect 1222 7123 1256 7147
rect 1222 7055 1256 7075
rect 1222 6987 1256 7003
rect 1222 6919 1256 6931
rect 1222 6851 1256 6859
rect 1222 6783 1256 6787
rect 1222 6677 1256 6681
rect 1222 6605 1256 6613
rect 1222 6533 1256 6545
rect 1222 6461 1256 6477
rect 1222 6389 1256 6409
rect 1222 6317 1256 6341
rect 1222 6245 1256 6273
rect 1222 6173 1256 6205
rect 1222 6103 1256 6137
rect 1222 6035 1256 6067
rect 1222 5967 1256 5995
rect 1222 5899 1256 5923
rect 1222 5831 1256 5851
rect 1222 5763 1256 5779
rect 1222 5695 1256 5707
rect 1222 5627 1256 5635
rect 1222 5559 1256 5563
rect 1222 5453 1256 5457
rect 1222 5381 1256 5389
rect 1222 5309 1256 5321
rect 1222 5237 1256 5253
rect 1222 5165 1256 5185
rect 1222 5093 1256 5117
rect 1222 5021 1256 5049
rect 1222 4949 1256 4981
rect 1222 4879 1256 4913
rect 1222 4811 1256 4843
rect 1222 4743 1256 4771
rect 1222 4675 1256 4699
rect 1222 4607 1256 4627
rect 1222 4539 1256 4555
rect 1222 4471 1256 4483
rect 1222 4403 1256 4411
rect 1222 4335 1256 4339
rect 1222 4229 1256 4233
rect 1222 4157 1256 4165
rect 1222 4085 1256 4097
rect 1222 4013 1256 4029
rect 1222 3941 1256 3961
rect 1222 3869 1256 3893
rect 1222 3797 1256 3825
rect 1222 3725 1256 3757
rect 1222 3655 1256 3689
rect 1222 3587 1256 3619
rect 1222 3519 1256 3547
rect 1222 3451 1256 3475
rect 1222 3383 1256 3403
rect 1222 3315 1256 3331
rect 1222 3247 1256 3259
rect 1222 3179 1256 3187
rect 1222 3111 1256 3115
rect 1222 3005 1256 3009
rect 1222 2933 1256 2941
rect 1222 2861 1256 2873
rect 1222 2789 1256 2805
rect 1222 2717 1256 2737
rect 1222 2645 1256 2669
rect 1222 2573 1256 2601
rect 1222 2501 1256 2533
rect 1222 2431 1256 2465
rect 1222 2363 1256 2395
rect 1222 2295 1256 2323
rect 1222 2227 1256 2251
rect 1222 2159 1256 2179
rect 1222 2091 1256 2107
rect 1222 2023 1256 2035
rect 1222 1955 1256 1963
rect 1222 1887 1256 1891
rect 1222 1781 1256 1785
rect 1222 1709 1256 1717
rect 1222 1637 1256 1649
rect 1222 1565 1256 1581
rect 1222 1493 1256 1513
rect 1222 1421 1256 1445
rect 1222 1349 1256 1377
rect 1222 1277 1256 1309
rect 1222 1207 1256 1241
rect 1222 1139 1256 1171
rect 1222 1071 1256 1099
rect 1222 1003 1256 1027
rect 1222 935 1256 955
rect 1222 867 1256 883
rect 1222 799 1256 811
rect 1222 731 1256 739
rect 1222 663 1256 667
rect 1222 557 1256 561
rect 1222 485 1256 493
rect 1222 413 1256 425
rect 1222 341 1256 357
rect 1222 269 1256 289
rect 1222 197 1256 221
rect 1222 125 1256 153
rect 1222 53 1256 85
rect 1222 -17 1256 17
rect 1222 -85 1256 -53
rect 1222 -153 1256 -125
rect 1222 -221 1256 -197
rect 1222 -289 1256 -269
rect 1222 -357 1256 -341
rect 1222 -425 1256 -413
rect 1222 -493 1256 -485
rect 1222 -561 1256 -557
rect 1222 -667 1256 -663
rect 1222 -739 1256 -731
rect 1222 -811 1256 -799
rect 1222 -883 1256 -867
rect 1222 -955 1256 -935
rect 1222 -1027 1256 -1003
rect 1222 -1099 1256 -1071
rect 1222 -1171 1256 -1139
rect 1222 -1241 1256 -1207
rect 1222 -1309 1256 -1277
rect 1222 -1377 1256 -1349
rect 1222 -1445 1256 -1421
rect 1222 -1513 1256 -1493
rect 1222 -1581 1256 -1565
rect 1222 -1649 1256 -1637
rect 1222 -1717 1256 -1709
rect 1222 -1785 1256 -1781
rect 1222 -1891 1256 -1887
rect 1222 -1963 1256 -1955
rect 1222 -2035 1256 -2023
rect 1222 -2107 1256 -2091
rect 1222 -2179 1256 -2159
rect 1222 -2251 1256 -2227
rect 1222 -2323 1256 -2295
rect 1222 -2395 1256 -2363
rect 1222 -2465 1256 -2431
rect 1222 -2533 1256 -2501
rect 1222 -2601 1256 -2573
rect 1222 -2669 1256 -2645
rect 1222 -2737 1256 -2717
rect 1222 -2805 1256 -2789
rect 1222 -2873 1256 -2861
rect 1222 -2941 1256 -2933
rect 1222 -3009 1256 -3005
rect 1222 -3115 1256 -3111
rect 1222 -3187 1256 -3179
rect 1222 -3259 1256 -3247
rect 1222 -3331 1256 -3315
rect 1222 -3403 1256 -3383
rect 1222 -3475 1256 -3451
rect 1222 -3547 1256 -3519
rect 1222 -3619 1256 -3587
rect 1222 -3689 1256 -3655
rect 1222 -3757 1256 -3725
rect 1222 -3825 1256 -3797
rect 1222 -3893 1256 -3869
rect 1222 -3961 1256 -3941
rect 1222 -4029 1256 -4013
rect 1222 -4097 1256 -4085
rect 1222 -4165 1256 -4157
rect 1222 -4233 1256 -4229
rect 1222 -4339 1256 -4335
rect 1222 -4411 1256 -4403
rect 1222 -4483 1256 -4471
rect 1222 -4555 1256 -4539
rect 1222 -4627 1256 -4607
rect 1222 -4699 1256 -4675
rect 1222 -4771 1256 -4743
rect 1222 -4843 1256 -4811
rect 1222 -4913 1256 -4879
rect 1222 -4981 1256 -4949
rect 1222 -5049 1256 -5021
rect 1222 -5117 1256 -5093
rect 1222 -5185 1256 -5165
rect 1222 -5253 1256 -5237
rect 1222 -5321 1256 -5309
rect 1222 -5389 1256 -5381
rect 1222 -5457 1256 -5453
rect 1222 -5563 1256 -5559
rect 1222 -5635 1256 -5627
rect 1222 -5707 1256 -5695
rect 1222 -5779 1256 -5763
rect 1222 -5851 1256 -5831
rect 1222 -5923 1256 -5899
rect 1222 -5995 1256 -5967
rect 1222 -6067 1256 -6035
rect 1222 -6137 1256 -6103
rect 1222 -6205 1256 -6173
rect 1222 -6273 1256 -6245
rect 1222 -6341 1256 -6317
rect 1222 -6409 1256 -6389
rect 1222 -6477 1256 -6461
rect 1222 -6545 1256 -6533
rect 1222 -6613 1256 -6605
rect 1222 -6681 1256 -6677
rect 1222 -6787 1256 -6783
rect 1222 -6859 1256 -6851
rect 1222 -6931 1256 -6919
rect 1222 -7003 1256 -6987
rect 1222 -7075 1256 -7055
rect 1222 -7147 1256 -7123
rect 1222 -7219 1256 -7191
rect 1222 -7291 1256 -7259
rect 1222 -7361 1256 -7327
rect 1222 -7429 1256 -7397
rect 1222 -7497 1256 -7469
rect 1222 -7565 1256 -7541
rect 1222 -7633 1256 -7613
rect 1222 -7701 1256 -7685
rect 1222 -7769 1256 -7757
rect 1222 -7837 1256 -7829
rect 1222 -7905 1256 -7901
rect 1222 -8011 1256 -8007
rect 1222 -8083 1256 -8075
rect 1222 -8155 1256 -8143
rect 1222 -8227 1256 -8211
rect 1222 -8299 1256 -8279
rect 1222 -8371 1256 -8347
rect 1222 -8443 1256 -8415
rect 1222 -8515 1256 -8483
rect 1222 -8585 1256 -8551
rect 1222 -8653 1256 -8621
rect 1222 -8721 1256 -8693
rect 1222 -8789 1256 -8765
rect 1222 -8857 1256 -8837
rect 1222 -8925 1256 -8909
rect 1222 -8993 1256 -8981
rect 1222 -9061 1256 -9053
rect 1222 -9129 1256 -9125
rect 1222 -9235 1256 -9231
rect 1222 -9307 1256 -9299
rect 1222 -9379 1256 -9367
rect 1222 -9451 1256 -9435
rect 1222 -9523 1256 -9503
rect 1222 -9604 1256 -9571
rect 1340 9571 1374 9604
rect 1340 9503 1374 9523
rect 1340 9435 1374 9451
rect 1340 9367 1374 9379
rect 1340 9299 1374 9307
rect 1340 9231 1374 9235
rect 1340 9125 1374 9129
rect 1340 9053 1374 9061
rect 1340 8981 1374 8993
rect 1340 8909 1374 8925
rect 1340 8837 1374 8857
rect 1340 8765 1374 8789
rect 1340 8693 1374 8721
rect 1340 8621 1374 8653
rect 1340 8551 1374 8585
rect 1340 8483 1374 8515
rect 1340 8415 1374 8443
rect 1340 8347 1374 8371
rect 1340 8279 1374 8299
rect 1340 8211 1374 8227
rect 1340 8143 1374 8155
rect 1340 8075 1374 8083
rect 1340 8007 1374 8011
rect 1340 7901 1374 7905
rect 1340 7829 1374 7837
rect 1340 7757 1374 7769
rect 1340 7685 1374 7701
rect 1340 7613 1374 7633
rect 1340 7541 1374 7565
rect 1340 7469 1374 7497
rect 1340 7397 1374 7429
rect 1340 7327 1374 7361
rect 1340 7259 1374 7291
rect 1340 7191 1374 7219
rect 1340 7123 1374 7147
rect 1340 7055 1374 7075
rect 1340 6987 1374 7003
rect 1340 6919 1374 6931
rect 1340 6851 1374 6859
rect 1340 6783 1374 6787
rect 1340 6677 1374 6681
rect 1340 6605 1374 6613
rect 1340 6533 1374 6545
rect 1340 6461 1374 6477
rect 1340 6389 1374 6409
rect 1340 6317 1374 6341
rect 1340 6245 1374 6273
rect 1340 6173 1374 6205
rect 1340 6103 1374 6137
rect 1340 6035 1374 6067
rect 1340 5967 1374 5995
rect 1340 5899 1374 5923
rect 1340 5831 1374 5851
rect 1340 5763 1374 5779
rect 1340 5695 1374 5707
rect 1340 5627 1374 5635
rect 1340 5559 1374 5563
rect 1340 5453 1374 5457
rect 1340 5381 1374 5389
rect 1340 5309 1374 5321
rect 1340 5237 1374 5253
rect 1340 5165 1374 5185
rect 1340 5093 1374 5117
rect 1340 5021 1374 5049
rect 1340 4949 1374 4981
rect 1340 4879 1374 4913
rect 1340 4811 1374 4843
rect 1340 4743 1374 4771
rect 1340 4675 1374 4699
rect 1340 4607 1374 4627
rect 1340 4539 1374 4555
rect 1340 4471 1374 4483
rect 1340 4403 1374 4411
rect 1340 4335 1374 4339
rect 1340 4229 1374 4233
rect 1340 4157 1374 4165
rect 1340 4085 1374 4097
rect 1340 4013 1374 4029
rect 1340 3941 1374 3961
rect 1340 3869 1374 3893
rect 1340 3797 1374 3825
rect 1340 3725 1374 3757
rect 1340 3655 1374 3689
rect 1340 3587 1374 3619
rect 1340 3519 1374 3547
rect 1340 3451 1374 3475
rect 1340 3383 1374 3403
rect 1340 3315 1374 3331
rect 1340 3247 1374 3259
rect 1340 3179 1374 3187
rect 1340 3111 1374 3115
rect 1340 3005 1374 3009
rect 1340 2933 1374 2941
rect 1340 2861 1374 2873
rect 1340 2789 1374 2805
rect 1340 2717 1374 2737
rect 1340 2645 1374 2669
rect 1340 2573 1374 2601
rect 1340 2501 1374 2533
rect 1340 2431 1374 2465
rect 1340 2363 1374 2395
rect 1340 2295 1374 2323
rect 1340 2227 1374 2251
rect 1340 2159 1374 2179
rect 1340 2091 1374 2107
rect 1340 2023 1374 2035
rect 1340 1955 1374 1963
rect 1340 1887 1374 1891
rect 1340 1781 1374 1785
rect 1340 1709 1374 1717
rect 1340 1637 1374 1649
rect 1340 1565 1374 1581
rect 1340 1493 1374 1513
rect 1340 1421 1374 1445
rect 1340 1349 1374 1377
rect 1340 1277 1374 1309
rect 1340 1207 1374 1241
rect 1340 1139 1374 1171
rect 1340 1071 1374 1099
rect 1340 1003 1374 1027
rect 1340 935 1374 955
rect 1340 867 1374 883
rect 1340 799 1374 811
rect 1340 731 1374 739
rect 1340 663 1374 667
rect 1340 557 1374 561
rect 1340 485 1374 493
rect 1340 413 1374 425
rect 1340 341 1374 357
rect 1340 269 1374 289
rect 1340 197 1374 221
rect 1340 125 1374 153
rect 1340 53 1374 85
rect 1340 -17 1374 17
rect 1340 -85 1374 -53
rect 1340 -153 1374 -125
rect 1340 -221 1374 -197
rect 1340 -289 1374 -269
rect 1340 -357 1374 -341
rect 1340 -425 1374 -413
rect 1340 -493 1374 -485
rect 1340 -561 1374 -557
rect 1340 -667 1374 -663
rect 1340 -739 1374 -731
rect 1340 -811 1374 -799
rect 1340 -883 1374 -867
rect 1340 -955 1374 -935
rect 1340 -1027 1374 -1003
rect 1340 -1099 1374 -1071
rect 1340 -1171 1374 -1139
rect 1340 -1241 1374 -1207
rect 1340 -1309 1374 -1277
rect 1340 -1377 1374 -1349
rect 1340 -1445 1374 -1421
rect 1340 -1513 1374 -1493
rect 1340 -1581 1374 -1565
rect 1340 -1649 1374 -1637
rect 1340 -1717 1374 -1709
rect 1340 -1785 1374 -1781
rect 1340 -1891 1374 -1887
rect 1340 -1963 1374 -1955
rect 1340 -2035 1374 -2023
rect 1340 -2107 1374 -2091
rect 1340 -2179 1374 -2159
rect 1340 -2251 1374 -2227
rect 1340 -2323 1374 -2295
rect 1340 -2395 1374 -2363
rect 1340 -2465 1374 -2431
rect 1340 -2533 1374 -2501
rect 1340 -2601 1374 -2573
rect 1340 -2669 1374 -2645
rect 1340 -2737 1374 -2717
rect 1340 -2805 1374 -2789
rect 1340 -2873 1374 -2861
rect 1340 -2941 1374 -2933
rect 1340 -3009 1374 -3005
rect 1340 -3115 1374 -3111
rect 1340 -3187 1374 -3179
rect 1340 -3259 1374 -3247
rect 1340 -3331 1374 -3315
rect 1340 -3403 1374 -3383
rect 1340 -3475 1374 -3451
rect 1340 -3547 1374 -3519
rect 1340 -3619 1374 -3587
rect 1340 -3689 1374 -3655
rect 1340 -3757 1374 -3725
rect 1340 -3825 1374 -3797
rect 1340 -3893 1374 -3869
rect 1340 -3961 1374 -3941
rect 1340 -4029 1374 -4013
rect 1340 -4097 1374 -4085
rect 1340 -4165 1374 -4157
rect 1340 -4233 1374 -4229
rect 1340 -4339 1374 -4335
rect 1340 -4411 1374 -4403
rect 1340 -4483 1374 -4471
rect 1340 -4555 1374 -4539
rect 1340 -4627 1374 -4607
rect 1340 -4699 1374 -4675
rect 1340 -4771 1374 -4743
rect 1340 -4843 1374 -4811
rect 1340 -4913 1374 -4879
rect 1340 -4981 1374 -4949
rect 1340 -5049 1374 -5021
rect 1340 -5117 1374 -5093
rect 1340 -5185 1374 -5165
rect 1340 -5253 1374 -5237
rect 1340 -5321 1374 -5309
rect 1340 -5389 1374 -5381
rect 1340 -5457 1374 -5453
rect 1340 -5563 1374 -5559
rect 1340 -5635 1374 -5627
rect 1340 -5707 1374 -5695
rect 1340 -5779 1374 -5763
rect 1340 -5851 1374 -5831
rect 1340 -5923 1374 -5899
rect 1340 -5995 1374 -5967
rect 1340 -6067 1374 -6035
rect 1340 -6137 1374 -6103
rect 1340 -6205 1374 -6173
rect 1340 -6273 1374 -6245
rect 1340 -6341 1374 -6317
rect 1340 -6409 1374 -6389
rect 1340 -6477 1374 -6461
rect 1340 -6545 1374 -6533
rect 1340 -6613 1374 -6605
rect 1340 -6681 1374 -6677
rect 1340 -6787 1374 -6783
rect 1340 -6859 1374 -6851
rect 1340 -6931 1374 -6919
rect 1340 -7003 1374 -6987
rect 1340 -7075 1374 -7055
rect 1340 -7147 1374 -7123
rect 1340 -7219 1374 -7191
rect 1340 -7291 1374 -7259
rect 1340 -7361 1374 -7327
rect 1340 -7429 1374 -7397
rect 1340 -7497 1374 -7469
rect 1340 -7565 1374 -7541
rect 1340 -7633 1374 -7613
rect 1340 -7701 1374 -7685
rect 1340 -7769 1374 -7757
rect 1340 -7837 1374 -7829
rect 1340 -7905 1374 -7901
rect 1340 -8011 1374 -8007
rect 1340 -8083 1374 -8075
rect 1340 -8155 1374 -8143
rect 1340 -8227 1374 -8211
rect 1340 -8299 1374 -8279
rect 1340 -8371 1374 -8347
rect 1340 -8443 1374 -8415
rect 1340 -8515 1374 -8483
rect 1340 -8585 1374 -8551
rect 1340 -8653 1374 -8621
rect 1340 -8721 1374 -8693
rect 1340 -8789 1374 -8765
rect 1340 -8857 1374 -8837
rect 1340 -8925 1374 -8909
rect 1340 -8993 1374 -8981
rect 1340 -9061 1374 -9053
rect 1340 -9129 1374 -9125
rect 1340 -9235 1374 -9231
rect 1340 -9307 1374 -9299
rect 1340 -9379 1374 -9367
rect 1340 -9451 1374 -9435
rect 1340 -9523 1374 -9503
rect 1340 -9604 1374 -9571
rect 1458 9571 1492 9604
rect 1458 9503 1492 9523
rect 1458 9435 1492 9451
rect 1458 9367 1492 9379
rect 1458 9299 1492 9307
rect 1458 9231 1492 9235
rect 1458 9125 1492 9129
rect 1458 9053 1492 9061
rect 1458 8981 1492 8993
rect 1458 8909 1492 8925
rect 1458 8837 1492 8857
rect 1458 8765 1492 8789
rect 1458 8693 1492 8721
rect 1458 8621 1492 8653
rect 1458 8551 1492 8585
rect 1458 8483 1492 8515
rect 1458 8415 1492 8443
rect 1458 8347 1492 8371
rect 1458 8279 1492 8299
rect 1458 8211 1492 8227
rect 1458 8143 1492 8155
rect 1458 8075 1492 8083
rect 1458 8007 1492 8011
rect 1458 7901 1492 7905
rect 1458 7829 1492 7837
rect 1458 7757 1492 7769
rect 1458 7685 1492 7701
rect 1458 7613 1492 7633
rect 1458 7541 1492 7565
rect 1458 7469 1492 7497
rect 1458 7397 1492 7429
rect 1458 7327 1492 7361
rect 1458 7259 1492 7291
rect 1458 7191 1492 7219
rect 1458 7123 1492 7147
rect 1458 7055 1492 7075
rect 1458 6987 1492 7003
rect 1458 6919 1492 6931
rect 1458 6851 1492 6859
rect 1458 6783 1492 6787
rect 1458 6677 1492 6681
rect 1458 6605 1492 6613
rect 1458 6533 1492 6545
rect 1458 6461 1492 6477
rect 1458 6389 1492 6409
rect 1458 6317 1492 6341
rect 1458 6245 1492 6273
rect 1458 6173 1492 6205
rect 1458 6103 1492 6137
rect 1458 6035 1492 6067
rect 1458 5967 1492 5995
rect 1458 5899 1492 5923
rect 1458 5831 1492 5851
rect 1458 5763 1492 5779
rect 1458 5695 1492 5707
rect 1458 5627 1492 5635
rect 1458 5559 1492 5563
rect 1458 5453 1492 5457
rect 1458 5381 1492 5389
rect 1458 5309 1492 5321
rect 1458 5237 1492 5253
rect 1458 5165 1492 5185
rect 1458 5093 1492 5117
rect 1458 5021 1492 5049
rect 1458 4949 1492 4981
rect 1458 4879 1492 4913
rect 1458 4811 1492 4843
rect 1458 4743 1492 4771
rect 1458 4675 1492 4699
rect 1458 4607 1492 4627
rect 1458 4539 1492 4555
rect 1458 4471 1492 4483
rect 1458 4403 1492 4411
rect 1458 4335 1492 4339
rect 1458 4229 1492 4233
rect 1458 4157 1492 4165
rect 1458 4085 1492 4097
rect 1458 4013 1492 4029
rect 1458 3941 1492 3961
rect 1458 3869 1492 3893
rect 1458 3797 1492 3825
rect 1458 3725 1492 3757
rect 1458 3655 1492 3689
rect 1458 3587 1492 3619
rect 1458 3519 1492 3547
rect 1458 3451 1492 3475
rect 1458 3383 1492 3403
rect 1458 3315 1492 3331
rect 1458 3247 1492 3259
rect 1458 3179 1492 3187
rect 1458 3111 1492 3115
rect 1458 3005 1492 3009
rect 1458 2933 1492 2941
rect 1458 2861 1492 2873
rect 1458 2789 1492 2805
rect 1458 2717 1492 2737
rect 1458 2645 1492 2669
rect 1458 2573 1492 2601
rect 1458 2501 1492 2533
rect 1458 2431 1492 2465
rect 1458 2363 1492 2395
rect 1458 2295 1492 2323
rect 1458 2227 1492 2251
rect 1458 2159 1492 2179
rect 1458 2091 1492 2107
rect 1458 2023 1492 2035
rect 1458 1955 1492 1963
rect 1458 1887 1492 1891
rect 1458 1781 1492 1785
rect 1458 1709 1492 1717
rect 1458 1637 1492 1649
rect 1458 1565 1492 1581
rect 1458 1493 1492 1513
rect 1458 1421 1492 1445
rect 1458 1349 1492 1377
rect 1458 1277 1492 1309
rect 1458 1207 1492 1241
rect 1458 1139 1492 1171
rect 1458 1071 1492 1099
rect 1458 1003 1492 1027
rect 1458 935 1492 955
rect 1458 867 1492 883
rect 1458 799 1492 811
rect 1458 731 1492 739
rect 1458 663 1492 667
rect 1458 557 1492 561
rect 1458 485 1492 493
rect 1458 413 1492 425
rect 1458 341 1492 357
rect 1458 269 1492 289
rect 1458 197 1492 221
rect 1458 125 1492 153
rect 1458 53 1492 85
rect 1458 -17 1492 17
rect 1458 -85 1492 -53
rect 1458 -153 1492 -125
rect 1458 -221 1492 -197
rect 1458 -289 1492 -269
rect 1458 -357 1492 -341
rect 1458 -425 1492 -413
rect 1458 -493 1492 -485
rect 1458 -561 1492 -557
rect 1458 -667 1492 -663
rect 1458 -739 1492 -731
rect 1458 -811 1492 -799
rect 1458 -883 1492 -867
rect 1458 -955 1492 -935
rect 1458 -1027 1492 -1003
rect 1458 -1099 1492 -1071
rect 1458 -1171 1492 -1139
rect 1458 -1241 1492 -1207
rect 1458 -1309 1492 -1277
rect 1458 -1377 1492 -1349
rect 1458 -1445 1492 -1421
rect 1458 -1513 1492 -1493
rect 1458 -1581 1492 -1565
rect 1458 -1649 1492 -1637
rect 1458 -1717 1492 -1709
rect 1458 -1785 1492 -1781
rect 1458 -1891 1492 -1887
rect 1458 -1963 1492 -1955
rect 1458 -2035 1492 -2023
rect 1458 -2107 1492 -2091
rect 1458 -2179 1492 -2159
rect 1458 -2251 1492 -2227
rect 1458 -2323 1492 -2295
rect 1458 -2395 1492 -2363
rect 1458 -2465 1492 -2431
rect 1458 -2533 1492 -2501
rect 1458 -2601 1492 -2573
rect 1458 -2669 1492 -2645
rect 1458 -2737 1492 -2717
rect 1458 -2805 1492 -2789
rect 1458 -2873 1492 -2861
rect 1458 -2941 1492 -2933
rect 1458 -3009 1492 -3005
rect 1458 -3115 1492 -3111
rect 1458 -3187 1492 -3179
rect 1458 -3259 1492 -3247
rect 1458 -3331 1492 -3315
rect 1458 -3403 1492 -3383
rect 1458 -3475 1492 -3451
rect 1458 -3547 1492 -3519
rect 1458 -3619 1492 -3587
rect 1458 -3689 1492 -3655
rect 1458 -3757 1492 -3725
rect 1458 -3825 1492 -3797
rect 1458 -3893 1492 -3869
rect 1458 -3961 1492 -3941
rect 1458 -4029 1492 -4013
rect 1458 -4097 1492 -4085
rect 1458 -4165 1492 -4157
rect 1458 -4233 1492 -4229
rect 1458 -4339 1492 -4335
rect 1458 -4411 1492 -4403
rect 1458 -4483 1492 -4471
rect 1458 -4555 1492 -4539
rect 1458 -4627 1492 -4607
rect 1458 -4699 1492 -4675
rect 1458 -4771 1492 -4743
rect 1458 -4843 1492 -4811
rect 1458 -4913 1492 -4879
rect 1458 -4981 1492 -4949
rect 1458 -5049 1492 -5021
rect 1458 -5117 1492 -5093
rect 1458 -5185 1492 -5165
rect 1458 -5253 1492 -5237
rect 1458 -5321 1492 -5309
rect 1458 -5389 1492 -5381
rect 1458 -5457 1492 -5453
rect 1458 -5563 1492 -5559
rect 1458 -5635 1492 -5627
rect 1458 -5707 1492 -5695
rect 1458 -5779 1492 -5763
rect 1458 -5851 1492 -5831
rect 1458 -5923 1492 -5899
rect 1458 -5995 1492 -5967
rect 1458 -6067 1492 -6035
rect 1458 -6137 1492 -6103
rect 1458 -6205 1492 -6173
rect 1458 -6273 1492 -6245
rect 1458 -6341 1492 -6317
rect 1458 -6409 1492 -6389
rect 1458 -6477 1492 -6461
rect 1458 -6545 1492 -6533
rect 1458 -6613 1492 -6605
rect 1458 -6681 1492 -6677
rect 1458 -6787 1492 -6783
rect 1458 -6859 1492 -6851
rect 1458 -6931 1492 -6919
rect 1458 -7003 1492 -6987
rect 1458 -7075 1492 -7055
rect 1458 -7147 1492 -7123
rect 1458 -7219 1492 -7191
rect 1458 -7291 1492 -7259
rect 1458 -7361 1492 -7327
rect 1458 -7429 1492 -7397
rect 1458 -7497 1492 -7469
rect 1458 -7565 1492 -7541
rect 1458 -7633 1492 -7613
rect 1458 -7701 1492 -7685
rect 1458 -7769 1492 -7757
rect 1458 -7837 1492 -7829
rect 1458 -7905 1492 -7901
rect 1458 -8011 1492 -8007
rect 1458 -8083 1492 -8075
rect 1458 -8155 1492 -8143
rect 1458 -8227 1492 -8211
rect 1458 -8299 1492 -8279
rect 1458 -8371 1492 -8347
rect 1458 -8443 1492 -8415
rect 1458 -8515 1492 -8483
rect 1458 -8585 1492 -8551
rect 1458 -8653 1492 -8621
rect 1458 -8721 1492 -8693
rect 1458 -8789 1492 -8765
rect 1458 -8857 1492 -8837
rect 1458 -8925 1492 -8909
rect 1458 -8993 1492 -8981
rect 1458 -9061 1492 -9053
rect 1458 -9129 1492 -9125
rect 1458 -9235 1492 -9231
rect 1458 -9307 1492 -9299
rect 1458 -9379 1492 -9367
rect 1458 -9451 1492 -9435
rect 1458 -9523 1492 -9503
rect 1458 -9604 1492 -9571
<< viali >>
rect -1492 9537 -1458 9557
rect -1492 9523 -1458 9537
rect -1492 9469 -1458 9485
rect -1492 9451 -1458 9469
rect -1492 9401 -1458 9413
rect -1492 9379 -1458 9401
rect -1492 9333 -1458 9341
rect -1492 9307 -1458 9333
rect -1492 9265 -1458 9269
rect -1492 9235 -1458 9265
rect -1492 9163 -1458 9197
rect -1492 9095 -1458 9125
rect -1492 9091 -1458 9095
rect -1492 9027 -1458 9053
rect -1492 9019 -1458 9027
rect -1492 8959 -1458 8981
rect -1492 8947 -1458 8959
rect -1492 8891 -1458 8909
rect -1492 8875 -1458 8891
rect -1492 8823 -1458 8837
rect -1492 8803 -1458 8823
rect -1492 8755 -1458 8765
rect -1492 8731 -1458 8755
rect -1492 8687 -1458 8693
rect -1492 8659 -1458 8687
rect -1492 8619 -1458 8621
rect -1492 8587 -1458 8619
rect -1492 8517 -1458 8549
rect -1492 8515 -1458 8517
rect -1492 8449 -1458 8477
rect -1492 8443 -1458 8449
rect -1492 8381 -1458 8405
rect -1492 8371 -1458 8381
rect -1492 8313 -1458 8333
rect -1492 8299 -1458 8313
rect -1492 8245 -1458 8261
rect -1492 8227 -1458 8245
rect -1492 8177 -1458 8189
rect -1492 8155 -1458 8177
rect -1492 8109 -1458 8117
rect -1492 8083 -1458 8109
rect -1492 8041 -1458 8045
rect -1492 8011 -1458 8041
rect -1492 7939 -1458 7973
rect -1492 7871 -1458 7901
rect -1492 7867 -1458 7871
rect -1492 7803 -1458 7829
rect -1492 7795 -1458 7803
rect -1492 7735 -1458 7757
rect -1492 7723 -1458 7735
rect -1492 7667 -1458 7685
rect -1492 7651 -1458 7667
rect -1492 7599 -1458 7613
rect -1492 7579 -1458 7599
rect -1492 7531 -1458 7541
rect -1492 7507 -1458 7531
rect -1492 7463 -1458 7469
rect -1492 7435 -1458 7463
rect -1492 7395 -1458 7397
rect -1492 7363 -1458 7395
rect -1492 7293 -1458 7325
rect -1492 7291 -1458 7293
rect -1492 7225 -1458 7253
rect -1492 7219 -1458 7225
rect -1492 7157 -1458 7181
rect -1492 7147 -1458 7157
rect -1492 7089 -1458 7109
rect -1492 7075 -1458 7089
rect -1492 7021 -1458 7037
rect -1492 7003 -1458 7021
rect -1492 6953 -1458 6965
rect -1492 6931 -1458 6953
rect -1492 6885 -1458 6893
rect -1492 6859 -1458 6885
rect -1492 6817 -1458 6821
rect -1492 6787 -1458 6817
rect -1492 6715 -1458 6749
rect -1492 6647 -1458 6677
rect -1492 6643 -1458 6647
rect -1492 6579 -1458 6605
rect -1492 6571 -1458 6579
rect -1492 6511 -1458 6533
rect -1492 6499 -1458 6511
rect -1492 6443 -1458 6461
rect -1492 6427 -1458 6443
rect -1492 6375 -1458 6389
rect -1492 6355 -1458 6375
rect -1492 6307 -1458 6317
rect -1492 6283 -1458 6307
rect -1492 6239 -1458 6245
rect -1492 6211 -1458 6239
rect -1492 6171 -1458 6173
rect -1492 6139 -1458 6171
rect -1492 6069 -1458 6101
rect -1492 6067 -1458 6069
rect -1492 6001 -1458 6029
rect -1492 5995 -1458 6001
rect -1492 5933 -1458 5957
rect -1492 5923 -1458 5933
rect -1492 5865 -1458 5885
rect -1492 5851 -1458 5865
rect -1492 5797 -1458 5813
rect -1492 5779 -1458 5797
rect -1492 5729 -1458 5741
rect -1492 5707 -1458 5729
rect -1492 5661 -1458 5669
rect -1492 5635 -1458 5661
rect -1492 5593 -1458 5597
rect -1492 5563 -1458 5593
rect -1492 5491 -1458 5525
rect -1492 5423 -1458 5453
rect -1492 5419 -1458 5423
rect -1492 5355 -1458 5381
rect -1492 5347 -1458 5355
rect -1492 5287 -1458 5309
rect -1492 5275 -1458 5287
rect -1492 5219 -1458 5237
rect -1492 5203 -1458 5219
rect -1492 5151 -1458 5165
rect -1492 5131 -1458 5151
rect -1492 5083 -1458 5093
rect -1492 5059 -1458 5083
rect -1492 5015 -1458 5021
rect -1492 4987 -1458 5015
rect -1492 4947 -1458 4949
rect -1492 4915 -1458 4947
rect -1492 4845 -1458 4877
rect -1492 4843 -1458 4845
rect -1492 4777 -1458 4805
rect -1492 4771 -1458 4777
rect -1492 4709 -1458 4733
rect -1492 4699 -1458 4709
rect -1492 4641 -1458 4661
rect -1492 4627 -1458 4641
rect -1492 4573 -1458 4589
rect -1492 4555 -1458 4573
rect -1492 4505 -1458 4517
rect -1492 4483 -1458 4505
rect -1492 4437 -1458 4445
rect -1492 4411 -1458 4437
rect -1492 4369 -1458 4373
rect -1492 4339 -1458 4369
rect -1492 4267 -1458 4301
rect -1492 4199 -1458 4229
rect -1492 4195 -1458 4199
rect -1492 4131 -1458 4157
rect -1492 4123 -1458 4131
rect -1492 4063 -1458 4085
rect -1492 4051 -1458 4063
rect -1492 3995 -1458 4013
rect -1492 3979 -1458 3995
rect -1492 3927 -1458 3941
rect -1492 3907 -1458 3927
rect -1492 3859 -1458 3869
rect -1492 3835 -1458 3859
rect -1492 3791 -1458 3797
rect -1492 3763 -1458 3791
rect -1492 3723 -1458 3725
rect -1492 3691 -1458 3723
rect -1492 3621 -1458 3653
rect -1492 3619 -1458 3621
rect -1492 3553 -1458 3581
rect -1492 3547 -1458 3553
rect -1492 3485 -1458 3509
rect -1492 3475 -1458 3485
rect -1492 3417 -1458 3437
rect -1492 3403 -1458 3417
rect -1492 3349 -1458 3365
rect -1492 3331 -1458 3349
rect -1492 3281 -1458 3293
rect -1492 3259 -1458 3281
rect -1492 3213 -1458 3221
rect -1492 3187 -1458 3213
rect -1492 3145 -1458 3149
rect -1492 3115 -1458 3145
rect -1492 3043 -1458 3077
rect -1492 2975 -1458 3005
rect -1492 2971 -1458 2975
rect -1492 2907 -1458 2933
rect -1492 2899 -1458 2907
rect -1492 2839 -1458 2861
rect -1492 2827 -1458 2839
rect -1492 2771 -1458 2789
rect -1492 2755 -1458 2771
rect -1492 2703 -1458 2717
rect -1492 2683 -1458 2703
rect -1492 2635 -1458 2645
rect -1492 2611 -1458 2635
rect -1492 2567 -1458 2573
rect -1492 2539 -1458 2567
rect -1492 2499 -1458 2501
rect -1492 2467 -1458 2499
rect -1492 2397 -1458 2429
rect -1492 2395 -1458 2397
rect -1492 2329 -1458 2357
rect -1492 2323 -1458 2329
rect -1492 2261 -1458 2285
rect -1492 2251 -1458 2261
rect -1492 2193 -1458 2213
rect -1492 2179 -1458 2193
rect -1492 2125 -1458 2141
rect -1492 2107 -1458 2125
rect -1492 2057 -1458 2069
rect -1492 2035 -1458 2057
rect -1492 1989 -1458 1997
rect -1492 1963 -1458 1989
rect -1492 1921 -1458 1925
rect -1492 1891 -1458 1921
rect -1492 1819 -1458 1853
rect -1492 1751 -1458 1781
rect -1492 1747 -1458 1751
rect -1492 1683 -1458 1709
rect -1492 1675 -1458 1683
rect -1492 1615 -1458 1637
rect -1492 1603 -1458 1615
rect -1492 1547 -1458 1565
rect -1492 1531 -1458 1547
rect -1492 1479 -1458 1493
rect -1492 1459 -1458 1479
rect -1492 1411 -1458 1421
rect -1492 1387 -1458 1411
rect -1492 1343 -1458 1349
rect -1492 1315 -1458 1343
rect -1492 1275 -1458 1277
rect -1492 1243 -1458 1275
rect -1492 1173 -1458 1205
rect -1492 1171 -1458 1173
rect -1492 1105 -1458 1133
rect -1492 1099 -1458 1105
rect -1492 1037 -1458 1061
rect -1492 1027 -1458 1037
rect -1492 969 -1458 989
rect -1492 955 -1458 969
rect -1492 901 -1458 917
rect -1492 883 -1458 901
rect -1492 833 -1458 845
rect -1492 811 -1458 833
rect -1492 765 -1458 773
rect -1492 739 -1458 765
rect -1492 697 -1458 701
rect -1492 667 -1458 697
rect -1492 595 -1458 629
rect -1492 527 -1458 557
rect -1492 523 -1458 527
rect -1492 459 -1458 485
rect -1492 451 -1458 459
rect -1492 391 -1458 413
rect -1492 379 -1458 391
rect -1492 323 -1458 341
rect -1492 307 -1458 323
rect -1492 255 -1458 269
rect -1492 235 -1458 255
rect -1492 187 -1458 197
rect -1492 163 -1458 187
rect -1492 119 -1458 125
rect -1492 91 -1458 119
rect -1492 51 -1458 53
rect -1492 19 -1458 51
rect -1492 -51 -1458 -19
rect -1492 -53 -1458 -51
rect -1492 -119 -1458 -91
rect -1492 -125 -1458 -119
rect -1492 -187 -1458 -163
rect -1492 -197 -1458 -187
rect -1492 -255 -1458 -235
rect -1492 -269 -1458 -255
rect -1492 -323 -1458 -307
rect -1492 -341 -1458 -323
rect -1492 -391 -1458 -379
rect -1492 -413 -1458 -391
rect -1492 -459 -1458 -451
rect -1492 -485 -1458 -459
rect -1492 -527 -1458 -523
rect -1492 -557 -1458 -527
rect -1492 -629 -1458 -595
rect -1492 -697 -1458 -667
rect -1492 -701 -1458 -697
rect -1492 -765 -1458 -739
rect -1492 -773 -1458 -765
rect -1492 -833 -1458 -811
rect -1492 -845 -1458 -833
rect -1492 -901 -1458 -883
rect -1492 -917 -1458 -901
rect -1492 -969 -1458 -955
rect -1492 -989 -1458 -969
rect -1492 -1037 -1458 -1027
rect -1492 -1061 -1458 -1037
rect -1492 -1105 -1458 -1099
rect -1492 -1133 -1458 -1105
rect -1492 -1173 -1458 -1171
rect -1492 -1205 -1458 -1173
rect -1492 -1275 -1458 -1243
rect -1492 -1277 -1458 -1275
rect -1492 -1343 -1458 -1315
rect -1492 -1349 -1458 -1343
rect -1492 -1411 -1458 -1387
rect -1492 -1421 -1458 -1411
rect -1492 -1479 -1458 -1459
rect -1492 -1493 -1458 -1479
rect -1492 -1547 -1458 -1531
rect -1492 -1565 -1458 -1547
rect -1492 -1615 -1458 -1603
rect -1492 -1637 -1458 -1615
rect -1492 -1683 -1458 -1675
rect -1492 -1709 -1458 -1683
rect -1492 -1751 -1458 -1747
rect -1492 -1781 -1458 -1751
rect -1492 -1853 -1458 -1819
rect -1492 -1921 -1458 -1891
rect -1492 -1925 -1458 -1921
rect -1492 -1989 -1458 -1963
rect -1492 -1997 -1458 -1989
rect -1492 -2057 -1458 -2035
rect -1492 -2069 -1458 -2057
rect -1492 -2125 -1458 -2107
rect -1492 -2141 -1458 -2125
rect -1492 -2193 -1458 -2179
rect -1492 -2213 -1458 -2193
rect -1492 -2261 -1458 -2251
rect -1492 -2285 -1458 -2261
rect -1492 -2329 -1458 -2323
rect -1492 -2357 -1458 -2329
rect -1492 -2397 -1458 -2395
rect -1492 -2429 -1458 -2397
rect -1492 -2499 -1458 -2467
rect -1492 -2501 -1458 -2499
rect -1492 -2567 -1458 -2539
rect -1492 -2573 -1458 -2567
rect -1492 -2635 -1458 -2611
rect -1492 -2645 -1458 -2635
rect -1492 -2703 -1458 -2683
rect -1492 -2717 -1458 -2703
rect -1492 -2771 -1458 -2755
rect -1492 -2789 -1458 -2771
rect -1492 -2839 -1458 -2827
rect -1492 -2861 -1458 -2839
rect -1492 -2907 -1458 -2899
rect -1492 -2933 -1458 -2907
rect -1492 -2975 -1458 -2971
rect -1492 -3005 -1458 -2975
rect -1492 -3077 -1458 -3043
rect -1492 -3145 -1458 -3115
rect -1492 -3149 -1458 -3145
rect -1492 -3213 -1458 -3187
rect -1492 -3221 -1458 -3213
rect -1492 -3281 -1458 -3259
rect -1492 -3293 -1458 -3281
rect -1492 -3349 -1458 -3331
rect -1492 -3365 -1458 -3349
rect -1492 -3417 -1458 -3403
rect -1492 -3437 -1458 -3417
rect -1492 -3485 -1458 -3475
rect -1492 -3509 -1458 -3485
rect -1492 -3553 -1458 -3547
rect -1492 -3581 -1458 -3553
rect -1492 -3621 -1458 -3619
rect -1492 -3653 -1458 -3621
rect -1492 -3723 -1458 -3691
rect -1492 -3725 -1458 -3723
rect -1492 -3791 -1458 -3763
rect -1492 -3797 -1458 -3791
rect -1492 -3859 -1458 -3835
rect -1492 -3869 -1458 -3859
rect -1492 -3927 -1458 -3907
rect -1492 -3941 -1458 -3927
rect -1492 -3995 -1458 -3979
rect -1492 -4013 -1458 -3995
rect -1492 -4063 -1458 -4051
rect -1492 -4085 -1458 -4063
rect -1492 -4131 -1458 -4123
rect -1492 -4157 -1458 -4131
rect -1492 -4199 -1458 -4195
rect -1492 -4229 -1458 -4199
rect -1492 -4301 -1458 -4267
rect -1492 -4369 -1458 -4339
rect -1492 -4373 -1458 -4369
rect -1492 -4437 -1458 -4411
rect -1492 -4445 -1458 -4437
rect -1492 -4505 -1458 -4483
rect -1492 -4517 -1458 -4505
rect -1492 -4573 -1458 -4555
rect -1492 -4589 -1458 -4573
rect -1492 -4641 -1458 -4627
rect -1492 -4661 -1458 -4641
rect -1492 -4709 -1458 -4699
rect -1492 -4733 -1458 -4709
rect -1492 -4777 -1458 -4771
rect -1492 -4805 -1458 -4777
rect -1492 -4845 -1458 -4843
rect -1492 -4877 -1458 -4845
rect -1492 -4947 -1458 -4915
rect -1492 -4949 -1458 -4947
rect -1492 -5015 -1458 -4987
rect -1492 -5021 -1458 -5015
rect -1492 -5083 -1458 -5059
rect -1492 -5093 -1458 -5083
rect -1492 -5151 -1458 -5131
rect -1492 -5165 -1458 -5151
rect -1492 -5219 -1458 -5203
rect -1492 -5237 -1458 -5219
rect -1492 -5287 -1458 -5275
rect -1492 -5309 -1458 -5287
rect -1492 -5355 -1458 -5347
rect -1492 -5381 -1458 -5355
rect -1492 -5423 -1458 -5419
rect -1492 -5453 -1458 -5423
rect -1492 -5525 -1458 -5491
rect -1492 -5593 -1458 -5563
rect -1492 -5597 -1458 -5593
rect -1492 -5661 -1458 -5635
rect -1492 -5669 -1458 -5661
rect -1492 -5729 -1458 -5707
rect -1492 -5741 -1458 -5729
rect -1492 -5797 -1458 -5779
rect -1492 -5813 -1458 -5797
rect -1492 -5865 -1458 -5851
rect -1492 -5885 -1458 -5865
rect -1492 -5933 -1458 -5923
rect -1492 -5957 -1458 -5933
rect -1492 -6001 -1458 -5995
rect -1492 -6029 -1458 -6001
rect -1492 -6069 -1458 -6067
rect -1492 -6101 -1458 -6069
rect -1492 -6171 -1458 -6139
rect -1492 -6173 -1458 -6171
rect -1492 -6239 -1458 -6211
rect -1492 -6245 -1458 -6239
rect -1492 -6307 -1458 -6283
rect -1492 -6317 -1458 -6307
rect -1492 -6375 -1458 -6355
rect -1492 -6389 -1458 -6375
rect -1492 -6443 -1458 -6427
rect -1492 -6461 -1458 -6443
rect -1492 -6511 -1458 -6499
rect -1492 -6533 -1458 -6511
rect -1492 -6579 -1458 -6571
rect -1492 -6605 -1458 -6579
rect -1492 -6647 -1458 -6643
rect -1492 -6677 -1458 -6647
rect -1492 -6749 -1458 -6715
rect -1492 -6817 -1458 -6787
rect -1492 -6821 -1458 -6817
rect -1492 -6885 -1458 -6859
rect -1492 -6893 -1458 -6885
rect -1492 -6953 -1458 -6931
rect -1492 -6965 -1458 -6953
rect -1492 -7021 -1458 -7003
rect -1492 -7037 -1458 -7021
rect -1492 -7089 -1458 -7075
rect -1492 -7109 -1458 -7089
rect -1492 -7157 -1458 -7147
rect -1492 -7181 -1458 -7157
rect -1492 -7225 -1458 -7219
rect -1492 -7253 -1458 -7225
rect -1492 -7293 -1458 -7291
rect -1492 -7325 -1458 -7293
rect -1492 -7395 -1458 -7363
rect -1492 -7397 -1458 -7395
rect -1492 -7463 -1458 -7435
rect -1492 -7469 -1458 -7463
rect -1492 -7531 -1458 -7507
rect -1492 -7541 -1458 -7531
rect -1492 -7599 -1458 -7579
rect -1492 -7613 -1458 -7599
rect -1492 -7667 -1458 -7651
rect -1492 -7685 -1458 -7667
rect -1492 -7735 -1458 -7723
rect -1492 -7757 -1458 -7735
rect -1492 -7803 -1458 -7795
rect -1492 -7829 -1458 -7803
rect -1492 -7871 -1458 -7867
rect -1492 -7901 -1458 -7871
rect -1492 -7973 -1458 -7939
rect -1492 -8041 -1458 -8011
rect -1492 -8045 -1458 -8041
rect -1492 -8109 -1458 -8083
rect -1492 -8117 -1458 -8109
rect -1492 -8177 -1458 -8155
rect -1492 -8189 -1458 -8177
rect -1492 -8245 -1458 -8227
rect -1492 -8261 -1458 -8245
rect -1492 -8313 -1458 -8299
rect -1492 -8333 -1458 -8313
rect -1492 -8381 -1458 -8371
rect -1492 -8405 -1458 -8381
rect -1492 -8449 -1458 -8443
rect -1492 -8477 -1458 -8449
rect -1492 -8517 -1458 -8515
rect -1492 -8549 -1458 -8517
rect -1492 -8619 -1458 -8587
rect -1492 -8621 -1458 -8619
rect -1492 -8687 -1458 -8659
rect -1492 -8693 -1458 -8687
rect -1492 -8755 -1458 -8731
rect -1492 -8765 -1458 -8755
rect -1492 -8823 -1458 -8803
rect -1492 -8837 -1458 -8823
rect -1492 -8891 -1458 -8875
rect -1492 -8909 -1458 -8891
rect -1492 -8959 -1458 -8947
rect -1492 -8981 -1458 -8959
rect -1492 -9027 -1458 -9019
rect -1492 -9053 -1458 -9027
rect -1492 -9095 -1458 -9091
rect -1492 -9125 -1458 -9095
rect -1492 -9197 -1458 -9163
rect -1492 -9265 -1458 -9235
rect -1492 -9269 -1458 -9265
rect -1492 -9333 -1458 -9307
rect -1492 -9341 -1458 -9333
rect -1492 -9401 -1458 -9379
rect -1492 -9413 -1458 -9401
rect -1492 -9469 -1458 -9451
rect -1492 -9485 -1458 -9469
rect -1492 -9537 -1458 -9523
rect -1492 -9557 -1458 -9537
rect -1374 9537 -1340 9557
rect -1374 9523 -1340 9537
rect -1374 9469 -1340 9485
rect -1374 9451 -1340 9469
rect -1374 9401 -1340 9413
rect -1374 9379 -1340 9401
rect -1374 9333 -1340 9341
rect -1374 9307 -1340 9333
rect -1374 9265 -1340 9269
rect -1374 9235 -1340 9265
rect -1374 9163 -1340 9197
rect -1374 9095 -1340 9125
rect -1374 9091 -1340 9095
rect -1374 9027 -1340 9053
rect -1374 9019 -1340 9027
rect -1374 8959 -1340 8981
rect -1374 8947 -1340 8959
rect -1374 8891 -1340 8909
rect -1374 8875 -1340 8891
rect -1374 8823 -1340 8837
rect -1374 8803 -1340 8823
rect -1374 8755 -1340 8765
rect -1374 8731 -1340 8755
rect -1374 8687 -1340 8693
rect -1374 8659 -1340 8687
rect -1374 8619 -1340 8621
rect -1374 8587 -1340 8619
rect -1374 8517 -1340 8549
rect -1374 8515 -1340 8517
rect -1374 8449 -1340 8477
rect -1374 8443 -1340 8449
rect -1374 8381 -1340 8405
rect -1374 8371 -1340 8381
rect -1374 8313 -1340 8333
rect -1374 8299 -1340 8313
rect -1374 8245 -1340 8261
rect -1374 8227 -1340 8245
rect -1374 8177 -1340 8189
rect -1374 8155 -1340 8177
rect -1374 8109 -1340 8117
rect -1374 8083 -1340 8109
rect -1374 8041 -1340 8045
rect -1374 8011 -1340 8041
rect -1374 7939 -1340 7973
rect -1374 7871 -1340 7901
rect -1374 7867 -1340 7871
rect -1374 7803 -1340 7829
rect -1374 7795 -1340 7803
rect -1374 7735 -1340 7757
rect -1374 7723 -1340 7735
rect -1374 7667 -1340 7685
rect -1374 7651 -1340 7667
rect -1374 7599 -1340 7613
rect -1374 7579 -1340 7599
rect -1374 7531 -1340 7541
rect -1374 7507 -1340 7531
rect -1374 7463 -1340 7469
rect -1374 7435 -1340 7463
rect -1374 7395 -1340 7397
rect -1374 7363 -1340 7395
rect -1374 7293 -1340 7325
rect -1374 7291 -1340 7293
rect -1374 7225 -1340 7253
rect -1374 7219 -1340 7225
rect -1374 7157 -1340 7181
rect -1374 7147 -1340 7157
rect -1374 7089 -1340 7109
rect -1374 7075 -1340 7089
rect -1374 7021 -1340 7037
rect -1374 7003 -1340 7021
rect -1374 6953 -1340 6965
rect -1374 6931 -1340 6953
rect -1374 6885 -1340 6893
rect -1374 6859 -1340 6885
rect -1374 6817 -1340 6821
rect -1374 6787 -1340 6817
rect -1374 6715 -1340 6749
rect -1374 6647 -1340 6677
rect -1374 6643 -1340 6647
rect -1374 6579 -1340 6605
rect -1374 6571 -1340 6579
rect -1374 6511 -1340 6533
rect -1374 6499 -1340 6511
rect -1374 6443 -1340 6461
rect -1374 6427 -1340 6443
rect -1374 6375 -1340 6389
rect -1374 6355 -1340 6375
rect -1374 6307 -1340 6317
rect -1374 6283 -1340 6307
rect -1374 6239 -1340 6245
rect -1374 6211 -1340 6239
rect -1374 6171 -1340 6173
rect -1374 6139 -1340 6171
rect -1374 6069 -1340 6101
rect -1374 6067 -1340 6069
rect -1374 6001 -1340 6029
rect -1374 5995 -1340 6001
rect -1374 5933 -1340 5957
rect -1374 5923 -1340 5933
rect -1374 5865 -1340 5885
rect -1374 5851 -1340 5865
rect -1374 5797 -1340 5813
rect -1374 5779 -1340 5797
rect -1374 5729 -1340 5741
rect -1374 5707 -1340 5729
rect -1374 5661 -1340 5669
rect -1374 5635 -1340 5661
rect -1374 5593 -1340 5597
rect -1374 5563 -1340 5593
rect -1374 5491 -1340 5525
rect -1374 5423 -1340 5453
rect -1374 5419 -1340 5423
rect -1374 5355 -1340 5381
rect -1374 5347 -1340 5355
rect -1374 5287 -1340 5309
rect -1374 5275 -1340 5287
rect -1374 5219 -1340 5237
rect -1374 5203 -1340 5219
rect -1374 5151 -1340 5165
rect -1374 5131 -1340 5151
rect -1374 5083 -1340 5093
rect -1374 5059 -1340 5083
rect -1374 5015 -1340 5021
rect -1374 4987 -1340 5015
rect -1374 4947 -1340 4949
rect -1374 4915 -1340 4947
rect -1374 4845 -1340 4877
rect -1374 4843 -1340 4845
rect -1374 4777 -1340 4805
rect -1374 4771 -1340 4777
rect -1374 4709 -1340 4733
rect -1374 4699 -1340 4709
rect -1374 4641 -1340 4661
rect -1374 4627 -1340 4641
rect -1374 4573 -1340 4589
rect -1374 4555 -1340 4573
rect -1374 4505 -1340 4517
rect -1374 4483 -1340 4505
rect -1374 4437 -1340 4445
rect -1374 4411 -1340 4437
rect -1374 4369 -1340 4373
rect -1374 4339 -1340 4369
rect -1374 4267 -1340 4301
rect -1374 4199 -1340 4229
rect -1374 4195 -1340 4199
rect -1374 4131 -1340 4157
rect -1374 4123 -1340 4131
rect -1374 4063 -1340 4085
rect -1374 4051 -1340 4063
rect -1374 3995 -1340 4013
rect -1374 3979 -1340 3995
rect -1374 3927 -1340 3941
rect -1374 3907 -1340 3927
rect -1374 3859 -1340 3869
rect -1374 3835 -1340 3859
rect -1374 3791 -1340 3797
rect -1374 3763 -1340 3791
rect -1374 3723 -1340 3725
rect -1374 3691 -1340 3723
rect -1374 3621 -1340 3653
rect -1374 3619 -1340 3621
rect -1374 3553 -1340 3581
rect -1374 3547 -1340 3553
rect -1374 3485 -1340 3509
rect -1374 3475 -1340 3485
rect -1374 3417 -1340 3437
rect -1374 3403 -1340 3417
rect -1374 3349 -1340 3365
rect -1374 3331 -1340 3349
rect -1374 3281 -1340 3293
rect -1374 3259 -1340 3281
rect -1374 3213 -1340 3221
rect -1374 3187 -1340 3213
rect -1374 3145 -1340 3149
rect -1374 3115 -1340 3145
rect -1374 3043 -1340 3077
rect -1374 2975 -1340 3005
rect -1374 2971 -1340 2975
rect -1374 2907 -1340 2933
rect -1374 2899 -1340 2907
rect -1374 2839 -1340 2861
rect -1374 2827 -1340 2839
rect -1374 2771 -1340 2789
rect -1374 2755 -1340 2771
rect -1374 2703 -1340 2717
rect -1374 2683 -1340 2703
rect -1374 2635 -1340 2645
rect -1374 2611 -1340 2635
rect -1374 2567 -1340 2573
rect -1374 2539 -1340 2567
rect -1374 2499 -1340 2501
rect -1374 2467 -1340 2499
rect -1374 2397 -1340 2429
rect -1374 2395 -1340 2397
rect -1374 2329 -1340 2357
rect -1374 2323 -1340 2329
rect -1374 2261 -1340 2285
rect -1374 2251 -1340 2261
rect -1374 2193 -1340 2213
rect -1374 2179 -1340 2193
rect -1374 2125 -1340 2141
rect -1374 2107 -1340 2125
rect -1374 2057 -1340 2069
rect -1374 2035 -1340 2057
rect -1374 1989 -1340 1997
rect -1374 1963 -1340 1989
rect -1374 1921 -1340 1925
rect -1374 1891 -1340 1921
rect -1374 1819 -1340 1853
rect -1374 1751 -1340 1781
rect -1374 1747 -1340 1751
rect -1374 1683 -1340 1709
rect -1374 1675 -1340 1683
rect -1374 1615 -1340 1637
rect -1374 1603 -1340 1615
rect -1374 1547 -1340 1565
rect -1374 1531 -1340 1547
rect -1374 1479 -1340 1493
rect -1374 1459 -1340 1479
rect -1374 1411 -1340 1421
rect -1374 1387 -1340 1411
rect -1374 1343 -1340 1349
rect -1374 1315 -1340 1343
rect -1374 1275 -1340 1277
rect -1374 1243 -1340 1275
rect -1374 1173 -1340 1205
rect -1374 1171 -1340 1173
rect -1374 1105 -1340 1133
rect -1374 1099 -1340 1105
rect -1374 1037 -1340 1061
rect -1374 1027 -1340 1037
rect -1374 969 -1340 989
rect -1374 955 -1340 969
rect -1374 901 -1340 917
rect -1374 883 -1340 901
rect -1374 833 -1340 845
rect -1374 811 -1340 833
rect -1374 765 -1340 773
rect -1374 739 -1340 765
rect -1374 697 -1340 701
rect -1374 667 -1340 697
rect -1374 595 -1340 629
rect -1374 527 -1340 557
rect -1374 523 -1340 527
rect -1374 459 -1340 485
rect -1374 451 -1340 459
rect -1374 391 -1340 413
rect -1374 379 -1340 391
rect -1374 323 -1340 341
rect -1374 307 -1340 323
rect -1374 255 -1340 269
rect -1374 235 -1340 255
rect -1374 187 -1340 197
rect -1374 163 -1340 187
rect -1374 119 -1340 125
rect -1374 91 -1340 119
rect -1374 51 -1340 53
rect -1374 19 -1340 51
rect -1374 -51 -1340 -19
rect -1374 -53 -1340 -51
rect -1374 -119 -1340 -91
rect -1374 -125 -1340 -119
rect -1374 -187 -1340 -163
rect -1374 -197 -1340 -187
rect -1374 -255 -1340 -235
rect -1374 -269 -1340 -255
rect -1374 -323 -1340 -307
rect -1374 -341 -1340 -323
rect -1374 -391 -1340 -379
rect -1374 -413 -1340 -391
rect -1374 -459 -1340 -451
rect -1374 -485 -1340 -459
rect -1374 -527 -1340 -523
rect -1374 -557 -1340 -527
rect -1374 -629 -1340 -595
rect -1374 -697 -1340 -667
rect -1374 -701 -1340 -697
rect -1374 -765 -1340 -739
rect -1374 -773 -1340 -765
rect -1374 -833 -1340 -811
rect -1374 -845 -1340 -833
rect -1374 -901 -1340 -883
rect -1374 -917 -1340 -901
rect -1374 -969 -1340 -955
rect -1374 -989 -1340 -969
rect -1374 -1037 -1340 -1027
rect -1374 -1061 -1340 -1037
rect -1374 -1105 -1340 -1099
rect -1374 -1133 -1340 -1105
rect -1374 -1173 -1340 -1171
rect -1374 -1205 -1340 -1173
rect -1374 -1275 -1340 -1243
rect -1374 -1277 -1340 -1275
rect -1374 -1343 -1340 -1315
rect -1374 -1349 -1340 -1343
rect -1374 -1411 -1340 -1387
rect -1374 -1421 -1340 -1411
rect -1374 -1479 -1340 -1459
rect -1374 -1493 -1340 -1479
rect -1374 -1547 -1340 -1531
rect -1374 -1565 -1340 -1547
rect -1374 -1615 -1340 -1603
rect -1374 -1637 -1340 -1615
rect -1374 -1683 -1340 -1675
rect -1374 -1709 -1340 -1683
rect -1374 -1751 -1340 -1747
rect -1374 -1781 -1340 -1751
rect -1374 -1853 -1340 -1819
rect -1374 -1921 -1340 -1891
rect -1374 -1925 -1340 -1921
rect -1374 -1989 -1340 -1963
rect -1374 -1997 -1340 -1989
rect -1374 -2057 -1340 -2035
rect -1374 -2069 -1340 -2057
rect -1374 -2125 -1340 -2107
rect -1374 -2141 -1340 -2125
rect -1374 -2193 -1340 -2179
rect -1374 -2213 -1340 -2193
rect -1374 -2261 -1340 -2251
rect -1374 -2285 -1340 -2261
rect -1374 -2329 -1340 -2323
rect -1374 -2357 -1340 -2329
rect -1374 -2397 -1340 -2395
rect -1374 -2429 -1340 -2397
rect -1374 -2499 -1340 -2467
rect -1374 -2501 -1340 -2499
rect -1374 -2567 -1340 -2539
rect -1374 -2573 -1340 -2567
rect -1374 -2635 -1340 -2611
rect -1374 -2645 -1340 -2635
rect -1374 -2703 -1340 -2683
rect -1374 -2717 -1340 -2703
rect -1374 -2771 -1340 -2755
rect -1374 -2789 -1340 -2771
rect -1374 -2839 -1340 -2827
rect -1374 -2861 -1340 -2839
rect -1374 -2907 -1340 -2899
rect -1374 -2933 -1340 -2907
rect -1374 -2975 -1340 -2971
rect -1374 -3005 -1340 -2975
rect -1374 -3077 -1340 -3043
rect -1374 -3145 -1340 -3115
rect -1374 -3149 -1340 -3145
rect -1374 -3213 -1340 -3187
rect -1374 -3221 -1340 -3213
rect -1374 -3281 -1340 -3259
rect -1374 -3293 -1340 -3281
rect -1374 -3349 -1340 -3331
rect -1374 -3365 -1340 -3349
rect -1374 -3417 -1340 -3403
rect -1374 -3437 -1340 -3417
rect -1374 -3485 -1340 -3475
rect -1374 -3509 -1340 -3485
rect -1374 -3553 -1340 -3547
rect -1374 -3581 -1340 -3553
rect -1374 -3621 -1340 -3619
rect -1374 -3653 -1340 -3621
rect -1374 -3723 -1340 -3691
rect -1374 -3725 -1340 -3723
rect -1374 -3791 -1340 -3763
rect -1374 -3797 -1340 -3791
rect -1374 -3859 -1340 -3835
rect -1374 -3869 -1340 -3859
rect -1374 -3927 -1340 -3907
rect -1374 -3941 -1340 -3927
rect -1374 -3995 -1340 -3979
rect -1374 -4013 -1340 -3995
rect -1374 -4063 -1340 -4051
rect -1374 -4085 -1340 -4063
rect -1374 -4131 -1340 -4123
rect -1374 -4157 -1340 -4131
rect -1374 -4199 -1340 -4195
rect -1374 -4229 -1340 -4199
rect -1374 -4301 -1340 -4267
rect -1374 -4369 -1340 -4339
rect -1374 -4373 -1340 -4369
rect -1374 -4437 -1340 -4411
rect -1374 -4445 -1340 -4437
rect -1374 -4505 -1340 -4483
rect -1374 -4517 -1340 -4505
rect -1374 -4573 -1340 -4555
rect -1374 -4589 -1340 -4573
rect -1374 -4641 -1340 -4627
rect -1374 -4661 -1340 -4641
rect -1374 -4709 -1340 -4699
rect -1374 -4733 -1340 -4709
rect -1374 -4777 -1340 -4771
rect -1374 -4805 -1340 -4777
rect -1374 -4845 -1340 -4843
rect -1374 -4877 -1340 -4845
rect -1374 -4947 -1340 -4915
rect -1374 -4949 -1340 -4947
rect -1374 -5015 -1340 -4987
rect -1374 -5021 -1340 -5015
rect -1374 -5083 -1340 -5059
rect -1374 -5093 -1340 -5083
rect -1374 -5151 -1340 -5131
rect -1374 -5165 -1340 -5151
rect -1374 -5219 -1340 -5203
rect -1374 -5237 -1340 -5219
rect -1374 -5287 -1340 -5275
rect -1374 -5309 -1340 -5287
rect -1374 -5355 -1340 -5347
rect -1374 -5381 -1340 -5355
rect -1374 -5423 -1340 -5419
rect -1374 -5453 -1340 -5423
rect -1374 -5525 -1340 -5491
rect -1374 -5593 -1340 -5563
rect -1374 -5597 -1340 -5593
rect -1374 -5661 -1340 -5635
rect -1374 -5669 -1340 -5661
rect -1374 -5729 -1340 -5707
rect -1374 -5741 -1340 -5729
rect -1374 -5797 -1340 -5779
rect -1374 -5813 -1340 -5797
rect -1374 -5865 -1340 -5851
rect -1374 -5885 -1340 -5865
rect -1374 -5933 -1340 -5923
rect -1374 -5957 -1340 -5933
rect -1374 -6001 -1340 -5995
rect -1374 -6029 -1340 -6001
rect -1374 -6069 -1340 -6067
rect -1374 -6101 -1340 -6069
rect -1374 -6171 -1340 -6139
rect -1374 -6173 -1340 -6171
rect -1374 -6239 -1340 -6211
rect -1374 -6245 -1340 -6239
rect -1374 -6307 -1340 -6283
rect -1374 -6317 -1340 -6307
rect -1374 -6375 -1340 -6355
rect -1374 -6389 -1340 -6375
rect -1374 -6443 -1340 -6427
rect -1374 -6461 -1340 -6443
rect -1374 -6511 -1340 -6499
rect -1374 -6533 -1340 -6511
rect -1374 -6579 -1340 -6571
rect -1374 -6605 -1340 -6579
rect -1374 -6647 -1340 -6643
rect -1374 -6677 -1340 -6647
rect -1374 -6749 -1340 -6715
rect -1374 -6817 -1340 -6787
rect -1374 -6821 -1340 -6817
rect -1374 -6885 -1340 -6859
rect -1374 -6893 -1340 -6885
rect -1374 -6953 -1340 -6931
rect -1374 -6965 -1340 -6953
rect -1374 -7021 -1340 -7003
rect -1374 -7037 -1340 -7021
rect -1374 -7089 -1340 -7075
rect -1374 -7109 -1340 -7089
rect -1374 -7157 -1340 -7147
rect -1374 -7181 -1340 -7157
rect -1374 -7225 -1340 -7219
rect -1374 -7253 -1340 -7225
rect -1374 -7293 -1340 -7291
rect -1374 -7325 -1340 -7293
rect -1374 -7395 -1340 -7363
rect -1374 -7397 -1340 -7395
rect -1374 -7463 -1340 -7435
rect -1374 -7469 -1340 -7463
rect -1374 -7531 -1340 -7507
rect -1374 -7541 -1340 -7531
rect -1374 -7599 -1340 -7579
rect -1374 -7613 -1340 -7599
rect -1374 -7667 -1340 -7651
rect -1374 -7685 -1340 -7667
rect -1374 -7735 -1340 -7723
rect -1374 -7757 -1340 -7735
rect -1374 -7803 -1340 -7795
rect -1374 -7829 -1340 -7803
rect -1374 -7871 -1340 -7867
rect -1374 -7901 -1340 -7871
rect -1374 -7973 -1340 -7939
rect -1374 -8041 -1340 -8011
rect -1374 -8045 -1340 -8041
rect -1374 -8109 -1340 -8083
rect -1374 -8117 -1340 -8109
rect -1374 -8177 -1340 -8155
rect -1374 -8189 -1340 -8177
rect -1374 -8245 -1340 -8227
rect -1374 -8261 -1340 -8245
rect -1374 -8313 -1340 -8299
rect -1374 -8333 -1340 -8313
rect -1374 -8381 -1340 -8371
rect -1374 -8405 -1340 -8381
rect -1374 -8449 -1340 -8443
rect -1374 -8477 -1340 -8449
rect -1374 -8517 -1340 -8515
rect -1374 -8549 -1340 -8517
rect -1374 -8619 -1340 -8587
rect -1374 -8621 -1340 -8619
rect -1374 -8687 -1340 -8659
rect -1374 -8693 -1340 -8687
rect -1374 -8755 -1340 -8731
rect -1374 -8765 -1340 -8755
rect -1374 -8823 -1340 -8803
rect -1374 -8837 -1340 -8823
rect -1374 -8891 -1340 -8875
rect -1374 -8909 -1340 -8891
rect -1374 -8959 -1340 -8947
rect -1374 -8981 -1340 -8959
rect -1374 -9027 -1340 -9019
rect -1374 -9053 -1340 -9027
rect -1374 -9095 -1340 -9091
rect -1374 -9125 -1340 -9095
rect -1374 -9197 -1340 -9163
rect -1374 -9265 -1340 -9235
rect -1374 -9269 -1340 -9265
rect -1374 -9333 -1340 -9307
rect -1374 -9341 -1340 -9333
rect -1374 -9401 -1340 -9379
rect -1374 -9413 -1340 -9401
rect -1374 -9469 -1340 -9451
rect -1374 -9485 -1340 -9469
rect -1374 -9537 -1340 -9523
rect -1374 -9557 -1340 -9537
rect -1256 9537 -1222 9557
rect -1256 9523 -1222 9537
rect -1256 9469 -1222 9485
rect -1256 9451 -1222 9469
rect -1256 9401 -1222 9413
rect -1256 9379 -1222 9401
rect -1256 9333 -1222 9341
rect -1256 9307 -1222 9333
rect -1256 9265 -1222 9269
rect -1256 9235 -1222 9265
rect -1256 9163 -1222 9197
rect -1256 9095 -1222 9125
rect -1256 9091 -1222 9095
rect -1256 9027 -1222 9053
rect -1256 9019 -1222 9027
rect -1256 8959 -1222 8981
rect -1256 8947 -1222 8959
rect -1256 8891 -1222 8909
rect -1256 8875 -1222 8891
rect -1256 8823 -1222 8837
rect -1256 8803 -1222 8823
rect -1256 8755 -1222 8765
rect -1256 8731 -1222 8755
rect -1256 8687 -1222 8693
rect -1256 8659 -1222 8687
rect -1256 8619 -1222 8621
rect -1256 8587 -1222 8619
rect -1256 8517 -1222 8549
rect -1256 8515 -1222 8517
rect -1256 8449 -1222 8477
rect -1256 8443 -1222 8449
rect -1256 8381 -1222 8405
rect -1256 8371 -1222 8381
rect -1256 8313 -1222 8333
rect -1256 8299 -1222 8313
rect -1256 8245 -1222 8261
rect -1256 8227 -1222 8245
rect -1256 8177 -1222 8189
rect -1256 8155 -1222 8177
rect -1256 8109 -1222 8117
rect -1256 8083 -1222 8109
rect -1256 8041 -1222 8045
rect -1256 8011 -1222 8041
rect -1256 7939 -1222 7973
rect -1256 7871 -1222 7901
rect -1256 7867 -1222 7871
rect -1256 7803 -1222 7829
rect -1256 7795 -1222 7803
rect -1256 7735 -1222 7757
rect -1256 7723 -1222 7735
rect -1256 7667 -1222 7685
rect -1256 7651 -1222 7667
rect -1256 7599 -1222 7613
rect -1256 7579 -1222 7599
rect -1256 7531 -1222 7541
rect -1256 7507 -1222 7531
rect -1256 7463 -1222 7469
rect -1256 7435 -1222 7463
rect -1256 7395 -1222 7397
rect -1256 7363 -1222 7395
rect -1256 7293 -1222 7325
rect -1256 7291 -1222 7293
rect -1256 7225 -1222 7253
rect -1256 7219 -1222 7225
rect -1256 7157 -1222 7181
rect -1256 7147 -1222 7157
rect -1256 7089 -1222 7109
rect -1256 7075 -1222 7089
rect -1256 7021 -1222 7037
rect -1256 7003 -1222 7021
rect -1256 6953 -1222 6965
rect -1256 6931 -1222 6953
rect -1256 6885 -1222 6893
rect -1256 6859 -1222 6885
rect -1256 6817 -1222 6821
rect -1256 6787 -1222 6817
rect -1256 6715 -1222 6749
rect -1256 6647 -1222 6677
rect -1256 6643 -1222 6647
rect -1256 6579 -1222 6605
rect -1256 6571 -1222 6579
rect -1256 6511 -1222 6533
rect -1256 6499 -1222 6511
rect -1256 6443 -1222 6461
rect -1256 6427 -1222 6443
rect -1256 6375 -1222 6389
rect -1256 6355 -1222 6375
rect -1256 6307 -1222 6317
rect -1256 6283 -1222 6307
rect -1256 6239 -1222 6245
rect -1256 6211 -1222 6239
rect -1256 6171 -1222 6173
rect -1256 6139 -1222 6171
rect -1256 6069 -1222 6101
rect -1256 6067 -1222 6069
rect -1256 6001 -1222 6029
rect -1256 5995 -1222 6001
rect -1256 5933 -1222 5957
rect -1256 5923 -1222 5933
rect -1256 5865 -1222 5885
rect -1256 5851 -1222 5865
rect -1256 5797 -1222 5813
rect -1256 5779 -1222 5797
rect -1256 5729 -1222 5741
rect -1256 5707 -1222 5729
rect -1256 5661 -1222 5669
rect -1256 5635 -1222 5661
rect -1256 5593 -1222 5597
rect -1256 5563 -1222 5593
rect -1256 5491 -1222 5525
rect -1256 5423 -1222 5453
rect -1256 5419 -1222 5423
rect -1256 5355 -1222 5381
rect -1256 5347 -1222 5355
rect -1256 5287 -1222 5309
rect -1256 5275 -1222 5287
rect -1256 5219 -1222 5237
rect -1256 5203 -1222 5219
rect -1256 5151 -1222 5165
rect -1256 5131 -1222 5151
rect -1256 5083 -1222 5093
rect -1256 5059 -1222 5083
rect -1256 5015 -1222 5021
rect -1256 4987 -1222 5015
rect -1256 4947 -1222 4949
rect -1256 4915 -1222 4947
rect -1256 4845 -1222 4877
rect -1256 4843 -1222 4845
rect -1256 4777 -1222 4805
rect -1256 4771 -1222 4777
rect -1256 4709 -1222 4733
rect -1256 4699 -1222 4709
rect -1256 4641 -1222 4661
rect -1256 4627 -1222 4641
rect -1256 4573 -1222 4589
rect -1256 4555 -1222 4573
rect -1256 4505 -1222 4517
rect -1256 4483 -1222 4505
rect -1256 4437 -1222 4445
rect -1256 4411 -1222 4437
rect -1256 4369 -1222 4373
rect -1256 4339 -1222 4369
rect -1256 4267 -1222 4301
rect -1256 4199 -1222 4229
rect -1256 4195 -1222 4199
rect -1256 4131 -1222 4157
rect -1256 4123 -1222 4131
rect -1256 4063 -1222 4085
rect -1256 4051 -1222 4063
rect -1256 3995 -1222 4013
rect -1256 3979 -1222 3995
rect -1256 3927 -1222 3941
rect -1256 3907 -1222 3927
rect -1256 3859 -1222 3869
rect -1256 3835 -1222 3859
rect -1256 3791 -1222 3797
rect -1256 3763 -1222 3791
rect -1256 3723 -1222 3725
rect -1256 3691 -1222 3723
rect -1256 3621 -1222 3653
rect -1256 3619 -1222 3621
rect -1256 3553 -1222 3581
rect -1256 3547 -1222 3553
rect -1256 3485 -1222 3509
rect -1256 3475 -1222 3485
rect -1256 3417 -1222 3437
rect -1256 3403 -1222 3417
rect -1256 3349 -1222 3365
rect -1256 3331 -1222 3349
rect -1256 3281 -1222 3293
rect -1256 3259 -1222 3281
rect -1256 3213 -1222 3221
rect -1256 3187 -1222 3213
rect -1256 3145 -1222 3149
rect -1256 3115 -1222 3145
rect -1256 3043 -1222 3077
rect -1256 2975 -1222 3005
rect -1256 2971 -1222 2975
rect -1256 2907 -1222 2933
rect -1256 2899 -1222 2907
rect -1256 2839 -1222 2861
rect -1256 2827 -1222 2839
rect -1256 2771 -1222 2789
rect -1256 2755 -1222 2771
rect -1256 2703 -1222 2717
rect -1256 2683 -1222 2703
rect -1256 2635 -1222 2645
rect -1256 2611 -1222 2635
rect -1256 2567 -1222 2573
rect -1256 2539 -1222 2567
rect -1256 2499 -1222 2501
rect -1256 2467 -1222 2499
rect -1256 2397 -1222 2429
rect -1256 2395 -1222 2397
rect -1256 2329 -1222 2357
rect -1256 2323 -1222 2329
rect -1256 2261 -1222 2285
rect -1256 2251 -1222 2261
rect -1256 2193 -1222 2213
rect -1256 2179 -1222 2193
rect -1256 2125 -1222 2141
rect -1256 2107 -1222 2125
rect -1256 2057 -1222 2069
rect -1256 2035 -1222 2057
rect -1256 1989 -1222 1997
rect -1256 1963 -1222 1989
rect -1256 1921 -1222 1925
rect -1256 1891 -1222 1921
rect -1256 1819 -1222 1853
rect -1256 1751 -1222 1781
rect -1256 1747 -1222 1751
rect -1256 1683 -1222 1709
rect -1256 1675 -1222 1683
rect -1256 1615 -1222 1637
rect -1256 1603 -1222 1615
rect -1256 1547 -1222 1565
rect -1256 1531 -1222 1547
rect -1256 1479 -1222 1493
rect -1256 1459 -1222 1479
rect -1256 1411 -1222 1421
rect -1256 1387 -1222 1411
rect -1256 1343 -1222 1349
rect -1256 1315 -1222 1343
rect -1256 1275 -1222 1277
rect -1256 1243 -1222 1275
rect -1256 1173 -1222 1205
rect -1256 1171 -1222 1173
rect -1256 1105 -1222 1133
rect -1256 1099 -1222 1105
rect -1256 1037 -1222 1061
rect -1256 1027 -1222 1037
rect -1256 969 -1222 989
rect -1256 955 -1222 969
rect -1256 901 -1222 917
rect -1256 883 -1222 901
rect -1256 833 -1222 845
rect -1256 811 -1222 833
rect -1256 765 -1222 773
rect -1256 739 -1222 765
rect -1256 697 -1222 701
rect -1256 667 -1222 697
rect -1256 595 -1222 629
rect -1256 527 -1222 557
rect -1256 523 -1222 527
rect -1256 459 -1222 485
rect -1256 451 -1222 459
rect -1256 391 -1222 413
rect -1256 379 -1222 391
rect -1256 323 -1222 341
rect -1256 307 -1222 323
rect -1256 255 -1222 269
rect -1256 235 -1222 255
rect -1256 187 -1222 197
rect -1256 163 -1222 187
rect -1256 119 -1222 125
rect -1256 91 -1222 119
rect -1256 51 -1222 53
rect -1256 19 -1222 51
rect -1256 -51 -1222 -19
rect -1256 -53 -1222 -51
rect -1256 -119 -1222 -91
rect -1256 -125 -1222 -119
rect -1256 -187 -1222 -163
rect -1256 -197 -1222 -187
rect -1256 -255 -1222 -235
rect -1256 -269 -1222 -255
rect -1256 -323 -1222 -307
rect -1256 -341 -1222 -323
rect -1256 -391 -1222 -379
rect -1256 -413 -1222 -391
rect -1256 -459 -1222 -451
rect -1256 -485 -1222 -459
rect -1256 -527 -1222 -523
rect -1256 -557 -1222 -527
rect -1256 -629 -1222 -595
rect -1256 -697 -1222 -667
rect -1256 -701 -1222 -697
rect -1256 -765 -1222 -739
rect -1256 -773 -1222 -765
rect -1256 -833 -1222 -811
rect -1256 -845 -1222 -833
rect -1256 -901 -1222 -883
rect -1256 -917 -1222 -901
rect -1256 -969 -1222 -955
rect -1256 -989 -1222 -969
rect -1256 -1037 -1222 -1027
rect -1256 -1061 -1222 -1037
rect -1256 -1105 -1222 -1099
rect -1256 -1133 -1222 -1105
rect -1256 -1173 -1222 -1171
rect -1256 -1205 -1222 -1173
rect -1256 -1275 -1222 -1243
rect -1256 -1277 -1222 -1275
rect -1256 -1343 -1222 -1315
rect -1256 -1349 -1222 -1343
rect -1256 -1411 -1222 -1387
rect -1256 -1421 -1222 -1411
rect -1256 -1479 -1222 -1459
rect -1256 -1493 -1222 -1479
rect -1256 -1547 -1222 -1531
rect -1256 -1565 -1222 -1547
rect -1256 -1615 -1222 -1603
rect -1256 -1637 -1222 -1615
rect -1256 -1683 -1222 -1675
rect -1256 -1709 -1222 -1683
rect -1256 -1751 -1222 -1747
rect -1256 -1781 -1222 -1751
rect -1256 -1853 -1222 -1819
rect -1256 -1921 -1222 -1891
rect -1256 -1925 -1222 -1921
rect -1256 -1989 -1222 -1963
rect -1256 -1997 -1222 -1989
rect -1256 -2057 -1222 -2035
rect -1256 -2069 -1222 -2057
rect -1256 -2125 -1222 -2107
rect -1256 -2141 -1222 -2125
rect -1256 -2193 -1222 -2179
rect -1256 -2213 -1222 -2193
rect -1256 -2261 -1222 -2251
rect -1256 -2285 -1222 -2261
rect -1256 -2329 -1222 -2323
rect -1256 -2357 -1222 -2329
rect -1256 -2397 -1222 -2395
rect -1256 -2429 -1222 -2397
rect -1256 -2499 -1222 -2467
rect -1256 -2501 -1222 -2499
rect -1256 -2567 -1222 -2539
rect -1256 -2573 -1222 -2567
rect -1256 -2635 -1222 -2611
rect -1256 -2645 -1222 -2635
rect -1256 -2703 -1222 -2683
rect -1256 -2717 -1222 -2703
rect -1256 -2771 -1222 -2755
rect -1256 -2789 -1222 -2771
rect -1256 -2839 -1222 -2827
rect -1256 -2861 -1222 -2839
rect -1256 -2907 -1222 -2899
rect -1256 -2933 -1222 -2907
rect -1256 -2975 -1222 -2971
rect -1256 -3005 -1222 -2975
rect -1256 -3077 -1222 -3043
rect -1256 -3145 -1222 -3115
rect -1256 -3149 -1222 -3145
rect -1256 -3213 -1222 -3187
rect -1256 -3221 -1222 -3213
rect -1256 -3281 -1222 -3259
rect -1256 -3293 -1222 -3281
rect -1256 -3349 -1222 -3331
rect -1256 -3365 -1222 -3349
rect -1256 -3417 -1222 -3403
rect -1256 -3437 -1222 -3417
rect -1256 -3485 -1222 -3475
rect -1256 -3509 -1222 -3485
rect -1256 -3553 -1222 -3547
rect -1256 -3581 -1222 -3553
rect -1256 -3621 -1222 -3619
rect -1256 -3653 -1222 -3621
rect -1256 -3723 -1222 -3691
rect -1256 -3725 -1222 -3723
rect -1256 -3791 -1222 -3763
rect -1256 -3797 -1222 -3791
rect -1256 -3859 -1222 -3835
rect -1256 -3869 -1222 -3859
rect -1256 -3927 -1222 -3907
rect -1256 -3941 -1222 -3927
rect -1256 -3995 -1222 -3979
rect -1256 -4013 -1222 -3995
rect -1256 -4063 -1222 -4051
rect -1256 -4085 -1222 -4063
rect -1256 -4131 -1222 -4123
rect -1256 -4157 -1222 -4131
rect -1256 -4199 -1222 -4195
rect -1256 -4229 -1222 -4199
rect -1256 -4301 -1222 -4267
rect -1256 -4369 -1222 -4339
rect -1256 -4373 -1222 -4369
rect -1256 -4437 -1222 -4411
rect -1256 -4445 -1222 -4437
rect -1256 -4505 -1222 -4483
rect -1256 -4517 -1222 -4505
rect -1256 -4573 -1222 -4555
rect -1256 -4589 -1222 -4573
rect -1256 -4641 -1222 -4627
rect -1256 -4661 -1222 -4641
rect -1256 -4709 -1222 -4699
rect -1256 -4733 -1222 -4709
rect -1256 -4777 -1222 -4771
rect -1256 -4805 -1222 -4777
rect -1256 -4845 -1222 -4843
rect -1256 -4877 -1222 -4845
rect -1256 -4947 -1222 -4915
rect -1256 -4949 -1222 -4947
rect -1256 -5015 -1222 -4987
rect -1256 -5021 -1222 -5015
rect -1256 -5083 -1222 -5059
rect -1256 -5093 -1222 -5083
rect -1256 -5151 -1222 -5131
rect -1256 -5165 -1222 -5151
rect -1256 -5219 -1222 -5203
rect -1256 -5237 -1222 -5219
rect -1256 -5287 -1222 -5275
rect -1256 -5309 -1222 -5287
rect -1256 -5355 -1222 -5347
rect -1256 -5381 -1222 -5355
rect -1256 -5423 -1222 -5419
rect -1256 -5453 -1222 -5423
rect -1256 -5525 -1222 -5491
rect -1256 -5593 -1222 -5563
rect -1256 -5597 -1222 -5593
rect -1256 -5661 -1222 -5635
rect -1256 -5669 -1222 -5661
rect -1256 -5729 -1222 -5707
rect -1256 -5741 -1222 -5729
rect -1256 -5797 -1222 -5779
rect -1256 -5813 -1222 -5797
rect -1256 -5865 -1222 -5851
rect -1256 -5885 -1222 -5865
rect -1256 -5933 -1222 -5923
rect -1256 -5957 -1222 -5933
rect -1256 -6001 -1222 -5995
rect -1256 -6029 -1222 -6001
rect -1256 -6069 -1222 -6067
rect -1256 -6101 -1222 -6069
rect -1256 -6171 -1222 -6139
rect -1256 -6173 -1222 -6171
rect -1256 -6239 -1222 -6211
rect -1256 -6245 -1222 -6239
rect -1256 -6307 -1222 -6283
rect -1256 -6317 -1222 -6307
rect -1256 -6375 -1222 -6355
rect -1256 -6389 -1222 -6375
rect -1256 -6443 -1222 -6427
rect -1256 -6461 -1222 -6443
rect -1256 -6511 -1222 -6499
rect -1256 -6533 -1222 -6511
rect -1256 -6579 -1222 -6571
rect -1256 -6605 -1222 -6579
rect -1256 -6647 -1222 -6643
rect -1256 -6677 -1222 -6647
rect -1256 -6749 -1222 -6715
rect -1256 -6817 -1222 -6787
rect -1256 -6821 -1222 -6817
rect -1256 -6885 -1222 -6859
rect -1256 -6893 -1222 -6885
rect -1256 -6953 -1222 -6931
rect -1256 -6965 -1222 -6953
rect -1256 -7021 -1222 -7003
rect -1256 -7037 -1222 -7021
rect -1256 -7089 -1222 -7075
rect -1256 -7109 -1222 -7089
rect -1256 -7157 -1222 -7147
rect -1256 -7181 -1222 -7157
rect -1256 -7225 -1222 -7219
rect -1256 -7253 -1222 -7225
rect -1256 -7293 -1222 -7291
rect -1256 -7325 -1222 -7293
rect -1256 -7395 -1222 -7363
rect -1256 -7397 -1222 -7395
rect -1256 -7463 -1222 -7435
rect -1256 -7469 -1222 -7463
rect -1256 -7531 -1222 -7507
rect -1256 -7541 -1222 -7531
rect -1256 -7599 -1222 -7579
rect -1256 -7613 -1222 -7599
rect -1256 -7667 -1222 -7651
rect -1256 -7685 -1222 -7667
rect -1256 -7735 -1222 -7723
rect -1256 -7757 -1222 -7735
rect -1256 -7803 -1222 -7795
rect -1256 -7829 -1222 -7803
rect -1256 -7871 -1222 -7867
rect -1256 -7901 -1222 -7871
rect -1256 -7973 -1222 -7939
rect -1256 -8041 -1222 -8011
rect -1256 -8045 -1222 -8041
rect -1256 -8109 -1222 -8083
rect -1256 -8117 -1222 -8109
rect -1256 -8177 -1222 -8155
rect -1256 -8189 -1222 -8177
rect -1256 -8245 -1222 -8227
rect -1256 -8261 -1222 -8245
rect -1256 -8313 -1222 -8299
rect -1256 -8333 -1222 -8313
rect -1256 -8381 -1222 -8371
rect -1256 -8405 -1222 -8381
rect -1256 -8449 -1222 -8443
rect -1256 -8477 -1222 -8449
rect -1256 -8517 -1222 -8515
rect -1256 -8549 -1222 -8517
rect -1256 -8619 -1222 -8587
rect -1256 -8621 -1222 -8619
rect -1256 -8687 -1222 -8659
rect -1256 -8693 -1222 -8687
rect -1256 -8755 -1222 -8731
rect -1256 -8765 -1222 -8755
rect -1256 -8823 -1222 -8803
rect -1256 -8837 -1222 -8823
rect -1256 -8891 -1222 -8875
rect -1256 -8909 -1222 -8891
rect -1256 -8959 -1222 -8947
rect -1256 -8981 -1222 -8959
rect -1256 -9027 -1222 -9019
rect -1256 -9053 -1222 -9027
rect -1256 -9095 -1222 -9091
rect -1256 -9125 -1222 -9095
rect -1256 -9197 -1222 -9163
rect -1256 -9265 -1222 -9235
rect -1256 -9269 -1222 -9265
rect -1256 -9333 -1222 -9307
rect -1256 -9341 -1222 -9333
rect -1256 -9401 -1222 -9379
rect -1256 -9413 -1222 -9401
rect -1256 -9469 -1222 -9451
rect -1256 -9485 -1222 -9469
rect -1256 -9537 -1222 -9523
rect -1256 -9557 -1222 -9537
rect -1138 9537 -1104 9557
rect -1138 9523 -1104 9537
rect -1138 9469 -1104 9485
rect -1138 9451 -1104 9469
rect -1138 9401 -1104 9413
rect -1138 9379 -1104 9401
rect -1138 9333 -1104 9341
rect -1138 9307 -1104 9333
rect -1138 9265 -1104 9269
rect -1138 9235 -1104 9265
rect -1138 9163 -1104 9197
rect -1138 9095 -1104 9125
rect -1138 9091 -1104 9095
rect -1138 9027 -1104 9053
rect -1138 9019 -1104 9027
rect -1138 8959 -1104 8981
rect -1138 8947 -1104 8959
rect -1138 8891 -1104 8909
rect -1138 8875 -1104 8891
rect -1138 8823 -1104 8837
rect -1138 8803 -1104 8823
rect -1138 8755 -1104 8765
rect -1138 8731 -1104 8755
rect -1138 8687 -1104 8693
rect -1138 8659 -1104 8687
rect -1138 8619 -1104 8621
rect -1138 8587 -1104 8619
rect -1138 8517 -1104 8549
rect -1138 8515 -1104 8517
rect -1138 8449 -1104 8477
rect -1138 8443 -1104 8449
rect -1138 8381 -1104 8405
rect -1138 8371 -1104 8381
rect -1138 8313 -1104 8333
rect -1138 8299 -1104 8313
rect -1138 8245 -1104 8261
rect -1138 8227 -1104 8245
rect -1138 8177 -1104 8189
rect -1138 8155 -1104 8177
rect -1138 8109 -1104 8117
rect -1138 8083 -1104 8109
rect -1138 8041 -1104 8045
rect -1138 8011 -1104 8041
rect -1138 7939 -1104 7973
rect -1138 7871 -1104 7901
rect -1138 7867 -1104 7871
rect -1138 7803 -1104 7829
rect -1138 7795 -1104 7803
rect -1138 7735 -1104 7757
rect -1138 7723 -1104 7735
rect -1138 7667 -1104 7685
rect -1138 7651 -1104 7667
rect -1138 7599 -1104 7613
rect -1138 7579 -1104 7599
rect -1138 7531 -1104 7541
rect -1138 7507 -1104 7531
rect -1138 7463 -1104 7469
rect -1138 7435 -1104 7463
rect -1138 7395 -1104 7397
rect -1138 7363 -1104 7395
rect -1138 7293 -1104 7325
rect -1138 7291 -1104 7293
rect -1138 7225 -1104 7253
rect -1138 7219 -1104 7225
rect -1138 7157 -1104 7181
rect -1138 7147 -1104 7157
rect -1138 7089 -1104 7109
rect -1138 7075 -1104 7089
rect -1138 7021 -1104 7037
rect -1138 7003 -1104 7021
rect -1138 6953 -1104 6965
rect -1138 6931 -1104 6953
rect -1138 6885 -1104 6893
rect -1138 6859 -1104 6885
rect -1138 6817 -1104 6821
rect -1138 6787 -1104 6817
rect -1138 6715 -1104 6749
rect -1138 6647 -1104 6677
rect -1138 6643 -1104 6647
rect -1138 6579 -1104 6605
rect -1138 6571 -1104 6579
rect -1138 6511 -1104 6533
rect -1138 6499 -1104 6511
rect -1138 6443 -1104 6461
rect -1138 6427 -1104 6443
rect -1138 6375 -1104 6389
rect -1138 6355 -1104 6375
rect -1138 6307 -1104 6317
rect -1138 6283 -1104 6307
rect -1138 6239 -1104 6245
rect -1138 6211 -1104 6239
rect -1138 6171 -1104 6173
rect -1138 6139 -1104 6171
rect -1138 6069 -1104 6101
rect -1138 6067 -1104 6069
rect -1138 6001 -1104 6029
rect -1138 5995 -1104 6001
rect -1138 5933 -1104 5957
rect -1138 5923 -1104 5933
rect -1138 5865 -1104 5885
rect -1138 5851 -1104 5865
rect -1138 5797 -1104 5813
rect -1138 5779 -1104 5797
rect -1138 5729 -1104 5741
rect -1138 5707 -1104 5729
rect -1138 5661 -1104 5669
rect -1138 5635 -1104 5661
rect -1138 5593 -1104 5597
rect -1138 5563 -1104 5593
rect -1138 5491 -1104 5525
rect -1138 5423 -1104 5453
rect -1138 5419 -1104 5423
rect -1138 5355 -1104 5381
rect -1138 5347 -1104 5355
rect -1138 5287 -1104 5309
rect -1138 5275 -1104 5287
rect -1138 5219 -1104 5237
rect -1138 5203 -1104 5219
rect -1138 5151 -1104 5165
rect -1138 5131 -1104 5151
rect -1138 5083 -1104 5093
rect -1138 5059 -1104 5083
rect -1138 5015 -1104 5021
rect -1138 4987 -1104 5015
rect -1138 4947 -1104 4949
rect -1138 4915 -1104 4947
rect -1138 4845 -1104 4877
rect -1138 4843 -1104 4845
rect -1138 4777 -1104 4805
rect -1138 4771 -1104 4777
rect -1138 4709 -1104 4733
rect -1138 4699 -1104 4709
rect -1138 4641 -1104 4661
rect -1138 4627 -1104 4641
rect -1138 4573 -1104 4589
rect -1138 4555 -1104 4573
rect -1138 4505 -1104 4517
rect -1138 4483 -1104 4505
rect -1138 4437 -1104 4445
rect -1138 4411 -1104 4437
rect -1138 4369 -1104 4373
rect -1138 4339 -1104 4369
rect -1138 4267 -1104 4301
rect -1138 4199 -1104 4229
rect -1138 4195 -1104 4199
rect -1138 4131 -1104 4157
rect -1138 4123 -1104 4131
rect -1138 4063 -1104 4085
rect -1138 4051 -1104 4063
rect -1138 3995 -1104 4013
rect -1138 3979 -1104 3995
rect -1138 3927 -1104 3941
rect -1138 3907 -1104 3927
rect -1138 3859 -1104 3869
rect -1138 3835 -1104 3859
rect -1138 3791 -1104 3797
rect -1138 3763 -1104 3791
rect -1138 3723 -1104 3725
rect -1138 3691 -1104 3723
rect -1138 3621 -1104 3653
rect -1138 3619 -1104 3621
rect -1138 3553 -1104 3581
rect -1138 3547 -1104 3553
rect -1138 3485 -1104 3509
rect -1138 3475 -1104 3485
rect -1138 3417 -1104 3437
rect -1138 3403 -1104 3417
rect -1138 3349 -1104 3365
rect -1138 3331 -1104 3349
rect -1138 3281 -1104 3293
rect -1138 3259 -1104 3281
rect -1138 3213 -1104 3221
rect -1138 3187 -1104 3213
rect -1138 3145 -1104 3149
rect -1138 3115 -1104 3145
rect -1138 3043 -1104 3077
rect -1138 2975 -1104 3005
rect -1138 2971 -1104 2975
rect -1138 2907 -1104 2933
rect -1138 2899 -1104 2907
rect -1138 2839 -1104 2861
rect -1138 2827 -1104 2839
rect -1138 2771 -1104 2789
rect -1138 2755 -1104 2771
rect -1138 2703 -1104 2717
rect -1138 2683 -1104 2703
rect -1138 2635 -1104 2645
rect -1138 2611 -1104 2635
rect -1138 2567 -1104 2573
rect -1138 2539 -1104 2567
rect -1138 2499 -1104 2501
rect -1138 2467 -1104 2499
rect -1138 2397 -1104 2429
rect -1138 2395 -1104 2397
rect -1138 2329 -1104 2357
rect -1138 2323 -1104 2329
rect -1138 2261 -1104 2285
rect -1138 2251 -1104 2261
rect -1138 2193 -1104 2213
rect -1138 2179 -1104 2193
rect -1138 2125 -1104 2141
rect -1138 2107 -1104 2125
rect -1138 2057 -1104 2069
rect -1138 2035 -1104 2057
rect -1138 1989 -1104 1997
rect -1138 1963 -1104 1989
rect -1138 1921 -1104 1925
rect -1138 1891 -1104 1921
rect -1138 1819 -1104 1853
rect -1138 1751 -1104 1781
rect -1138 1747 -1104 1751
rect -1138 1683 -1104 1709
rect -1138 1675 -1104 1683
rect -1138 1615 -1104 1637
rect -1138 1603 -1104 1615
rect -1138 1547 -1104 1565
rect -1138 1531 -1104 1547
rect -1138 1479 -1104 1493
rect -1138 1459 -1104 1479
rect -1138 1411 -1104 1421
rect -1138 1387 -1104 1411
rect -1138 1343 -1104 1349
rect -1138 1315 -1104 1343
rect -1138 1275 -1104 1277
rect -1138 1243 -1104 1275
rect -1138 1173 -1104 1205
rect -1138 1171 -1104 1173
rect -1138 1105 -1104 1133
rect -1138 1099 -1104 1105
rect -1138 1037 -1104 1061
rect -1138 1027 -1104 1037
rect -1138 969 -1104 989
rect -1138 955 -1104 969
rect -1138 901 -1104 917
rect -1138 883 -1104 901
rect -1138 833 -1104 845
rect -1138 811 -1104 833
rect -1138 765 -1104 773
rect -1138 739 -1104 765
rect -1138 697 -1104 701
rect -1138 667 -1104 697
rect -1138 595 -1104 629
rect -1138 527 -1104 557
rect -1138 523 -1104 527
rect -1138 459 -1104 485
rect -1138 451 -1104 459
rect -1138 391 -1104 413
rect -1138 379 -1104 391
rect -1138 323 -1104 341
rect -1138 307 -1104 323
rect -1138 255 -1104 269
rect -1138 235 -1104 255
rect -1138 187 -1104 197
rect -1138 163 -1104 187
rect -1138 119 -1104 125
rect -1138 91 -1104 119
rect -1138 51 -1104 53
rect -1138 19 -1104 51
rect -1138 -51 -1104 -19
rect -1138 -53 -1104 -51
rect -1138 -119 -1104 -91
rect -1138 -125 -1104 -119
rect -1138 -187 -1104 -163
rect -1138 -197 -1104 -187
rect -1138 -255 -1104 -235
rect -1138 -269 -1104 -255
rect -1138 -323 -1104 -307
rect -1138 -341 -1104 -323
rect -1138 -391 -1104 -379
rect -1138 -413 -1104 -391
rect -1138 -459 -1104 -451
rect -1138 -485 -1104 -459
rect -1138 -527 -1104 -523
rect -1138 -557 -1104 -527
rect -1138 -629 -1104 -595
rect -1138 -697 -1104 -667
rect -1138 -701 -1104 -697
rect -1138 -765 -1104 -739
rect -1138 -773 -1104 -765
rect -1138 -833 -1104 -811
rect -1138 -845 -1104 -833
rect -1138 -901 -1104 -883
rect -1138 -917 -1104 -901
rect -1138 -969 -1104 -955
rect -1138 -989 -1104 -969
rect -1138 -1037 -1104 -1027
rect -1138 -1061 -1104 -1037
rect -1138 -1105 -1104 -1099
rect -1138 -1133 -1104 -1105
rect -1138 -1173 -1104 -1171
rect -1138 -1205 -1104 -1173
rect -1138 -1275 -1104 -1243
rect -1138 -1277 -1104 -1275
rect -1138 -1343 -1104 -1315
rect -1138 -1349 -1104 -1343
rect -1138 -1411 -1104 -1387
rect -1138 -1421 -1104 -1411
rect -1138 -1479 -1104 -1459
rect -1138 -1493 -1104 -1479
rect -1138 -1547 -1104 -1531
rect -1138 -1565 -1104 -1547
rect -1138 -1615 -1104 -1603
rect -1138 -1637 -1104 -1615
rect -1138 -1683 -1104 -1675
rect -1138 -1709 -1104 -1683
rect -1138 -1751 -1104 -1747
rect -1138 -1781 -1104 -1751
rect -1138 -1853 -1104 -1819
rect -1138 -1921 -1104 -1891
rect -1138 -1925 -1104 -1921
rect -1138 -1989 -1104 -1963
rect -1138 -1997 -1104 -1989
rect -1138 -2057 -1104 -2035
rect -1138 -2069 -1104 -2057
rect -1138 -2125 -1104 -2107
rect -1138 -2141 -1104 -2125
rect -1138 -2193 -1104 -2179
rect -1138 -2213 -1104 -2193
rect -1138 -2261 -1104 -2251
rect -1138 -2285 -1104 -2261
rect -1138 -2329 -1104 -2323
rect -1138 -2357 -1104 -2329
rect -1138 -2397 -1104 -2395
rect -1138 -2429 -1104 -2397
rect -1138 -2499 -1104 -2467
rect -1138 -2501 -1104 -2499
rect -1138 -2567 -1104 -2539
rect -1138 -2573 -1104 -2567
rect -1138 -2635 -1104 -2611
rect -1138 -2645 -1104 -2635
rect -1138 -2703 -1104 -2683
rect -1138 -2717 -1104 -2703
rect -1138 -2771 -1104 -2755
rect -1138 -2789 -1104 -2771
rect -1138 -2839 -1104 -2827
rect -1138 -2861 -1104 -2839
rect -1138 -2907 -1104 -2899
rect -1138 -2933 -1104 -2907
rect -1138 -2975 -1104 -2971
rect -1138 -3005 -1104 -2975
rect -1138 -3077 -1104 -3043
rect -1138 -3145 -1104 -3115
rect -1138 -3149 -1104 -3145
rect -1138 -3213 -1104 -3187
rect -1138 -3221 -1104 -3213
rect -1138 -3281 -1104 -3259
rect -1138 -3293 -1104 -3281
rect -1138 -3349 -1104 -3331
rect -1138 -3365 -1104 -3349
rect -1138 -3417 -1104 -3403
rect -1138 -3437 -1104 -3417
rect -1138 -3485 -1104 -3475
rect -1138 -3509 -1104 -3485
rect -1138 -3553 -1104 -3547
rect -1138 -3581 -1104 -3553
rect -1138 -3621 -1104 -3619
rect -1138 -3653 -1104 -3621
rect -1138 -3723 -1104 -3691
rect -1138 -3725 -1104 -3723
rect -1138 -3791 -1104 -3763
rect -1138 -3797 -1104 -3791
rect -1138 -3859 -1104 -3835
rect -1138 -3869 -1104 -3859
rect -1138 -3927 -1104 -3907
rect -1138 -3941 -1104 -3927
rect -1138 -3995 -1104 -3979
rect -1138 -4013 -1104 -3995
rect -1138 -4063 -1104 -4051
rect -1138 -4085 -1104 -4063
rect -1138 -4131 -1104 -4123
rect -1138 -4157 -1104 -4131
rect -1138 -4199 -1104 -4195
rect -1138 -4229 -1104 -4199
rect -1138 -4301 -1104 -4267
rect -1138 -4369 -1104 -4339
rect -1138 -4373 -1104 -4369
rect -1138 -4437 -1104 -4411
rect -1138 -4445 -1104 -4437
rect -1138 -4505 -1104 -4483
rect -1138 -4517 -1104 -4505
rect -1138 -4573 -1104 -4555
rect -1138 -4589 -1104 -4573
rect -1138 -4641 -1104 -4627
rect -1138 -4661 -1104 -4641
rect -1138 -4709 -1104 -4699
rect -1138 -4733 -1104 -4709
rect -1138 -4777 -1104 -4771
rect -1138 -4805 -1104 -4777
rect -1138 -4845 -1104 -4843
rect -1138 -4877 -1104 -4845
rect -1138 -4947 -1104 -4915
rect -1138 -4949 -1104 -4947
rect -1138 -5015 -1104 -4987
rect -1138 -5021 -1104 -5015
rect -1138 -5083 -1104 -5059
rect -1138 -5093 -1104 -5083
rect -1138 -5151 -1104 -5131
rect -1138 -5165 -1104 -5151
rect -1138 -5219 -1104 -5203
rect -1138 -5237 -1104 -5219
rect -1138 -5287 -1104 -5275
rect -1138 -5309 -1104 -5287
rect -1138 -5355 -1104 -5347
rect -1138 -5381 -1104 -5355
rect -1138 -5423 -1104 -5419
rect -1138 -5453 -1104 -5423
rect -1138 -5525 -1104 -5491
rect -1138 -5593 -1104 -5563
rect -1138 -5597 -1104 -5593
rect -1138 -5661 -1104 -5635
rect -1138 -5669 -1104 -5661
rect -1138 -5729 -1104 -5707
rect -1138 -5741 -1104 -5729
rect -1138 -5797 -1104 -5779
rect -1138 -5813 -1104 -5797
rect -1138 -5865 -1104 -5851
rect -1138 -5885 -1104 -5865
rect -1138 -5933 -1104 -5923
rect -1138 -5957 -1104 -5933
rect -1138 -6001 -1104 -5995
rect -1138 -6029 -1104 -6001
rect -1138 -6069 -1104 -6067
rect -1138 -6101 -1104 -6069
rect -1138 -6171 -1104 -6139
rect -1138 -6173 -1104 -6171
rect -1138 -6239 -1104 -6211
rect -1138 -6245 -1104 -6239
rect -1138 -6307 -1104 -6283
rect -1138 -6317 -1104 -6307
rect -1138 -6375 -1104 -6355
rect -1138 -6389 -1104 -6375
rect -1138 -6443 -1104 -6427
rect -1138 -6461 -1104 -6443
rect -1138 -6511 -1104 -6499
rect -1138 -6533 -1104 -6511
rect -1138 -6579 -1104 -6571
rect -1138 -6605 -1104 -6579
rect -1138 -6647 -1104 -6643
rect -1138 -6677 -1104 -6647
rect -1138 -6749 -1104 -6715
rect -1138 -6817 -1104 -6787
rect -1138 -6821 -1104 -6817
rect -1138 -6885 -1104 -6859
rect -1138 -6893 -1104 -6885
rect -1138 -6953 -1104 -6931
rect -1138 -6965 -1104 -6953
rect -1138 -7021 -1104 -7003
rect -1138 -7037 -1104 -7021
rect -1138 -7089 -1104 -7075
rect -1138 -7109 -1104 -7089
rect -1138 -7157 -1104 -7147
rect -1138 -7181 -1104 -7157
rect -1138 -7225 -1104 -7219
rect -1138 -7253 -1104 -7225
rect -1138 -7293 -1104 -7291
rect -1138 -7325 -1104 -7293
rect -1138 -7395 -1104 -7363
rect -1138 -7397 -1104 -7395
rect -1138 -7463 -1104 -7435
rect -1138 -7469 -1104 -7463
rect -1138 -7531 -1104 -7507
rect -1138 -7541 -1104 -7531
rect -1138 -7599 -1104 -7579
rect -1138 -7613 -1104 -7599
rect -1138 -7667 -1104 -7651
rect -1138 -7685 -1104 -7667
rect -1138 -7735 -1104 -7723
rect -1138 -7757 -1104 -7735
rect -1138 -7803 -1104 -7795
rect -1138 -7829 -1104 -7803
rect -1138 -7871 -1104 -7867
rect -1138 -7901 -1104 -7871
rect -1138 -7973 -1104 -7939
rect -1138 -8041 -1104 -8011
rect -1138 -8045 -1104 -8041
rect -1138 -8109 -1104 -8083
rect -1138 -8117 -1104 -8109
rect -1138 -8177 -1104 -8155
rect -1138 -8189 -1104 -8177
rect -1138 -8245 -1104 -8227
rect -1138 -8261 -1104 -8245
rect -1138 -8313 -1104 -8299
rect -1138 -8333 -1104 -8313
rect -1138 -8381 -1104 -8371
rect -1138 -8405 -1104 -8381
rect -1138 -8449 -1104 -8443
rect -1138 -8477 -1104 -8449
rect -1138 -8517 -1104 -8515
rect -1138 -8549 -1104 -8517
rect -1138 -8619 -1104 -8587
rect -1138 -8621 -1104 -8619
rect -1138 -8687 -1104 -8659
rect -1138 -8693 -1104 -8687
rect -1138 -8755 -1104 -8731
rect -1138 -8765 -1104 -8755
rect -1138 -8823 -1104 -8803
rect -1138 -8837 -1104 -8823
rect -1138 -8891 -1104 -8875
rect -1138 -8909 -1104 -8891
rect -1138 -8959 -1104 -8947
rect -1138 -8981 -1104 -8959
rect -1138 -9027 -1104 -9019
rect -1138 -9053 -1104 -9027
rect -1138 -9095 -1104 -9091
rect -1138 -9125 -1104 -9095
rect -1138 -9197 -1104 -9163
rect -1138 -9265 -1104 -9235
rect -1138 -9269 -1104 -9265
rect -1138 -9333 -1104 -9307
rect -1138 -9341 -1104 -9333
rect -1138 -9401 -1104 -9379
rect -1138 -9413 -1104 -9401
rect -1138 -9469 -1104 -9451
rect -1138 -9485 -1104 -9469
rect -1138 -9537 -1104 -9523
rect -1138 -9557 -1104 -9537
rect -1020 9537 -986 9557
rect -1020 9523 -986 9537
rect -1020 9469 -986 9485
rect -1020 9451 -986 9469
rect -1020 9401 -986 9413
rect -1020 9379 -986 9401
rect -1020 9333 -986 9341
rect -1020 9307 -986 9333
rect -1020 9265 -986 9269
rect -1020 9235 -986 9265
rect -1020 9163 -986 9197
rect -1020 9095 -986 9125
rect -1020 9091 -986 9095
rect -1020 9027 -986 9053
rect -1020 9019 -986 9027
rect -1020 8959 -986 8981
rect -1020 8947 -986 8959
rect -1020 8891 -986 8909
rect -1020 8875 -986 8891
rect -1020 8823 -986 8837
rect -1020 8803 -986 8823
rect -1020 8755 -986 8765
rect -1020 8731 -986 8755
rect -1020 8687 -986 8693
rect -1020 8659 -986 8687
rect -1020 8619 -986 8621
rect -1020 8587 -986 8619
rect -1020 8517 -986 8549
rect -1020 8515 -986 8517
rect -1020 8449 -986 8477
rect -1020 8443 -986 8449
rect -1020 8381 -986 8405
rect -1020 8371 -986 8381
rect -1020 8313 -986 8333
rect -1020 8299 -986 8313
rect -1020 8245 -986 8261
rect -1020 8227 -986 8245
rect -1020 8177 -986 8189
rect -1020 8155 -986 8177
rect -1020 8109 -986 8117
rect -1020 8083 -986 8109
rect -1020 8041 -986 8045
rect -1020 8011 -986 8041
rect -1020 7939 -986 7973
rect -1020 7871 -986 7901
rect -1020 7867 -986 7871
rect -1020 7803 -986 7829
rect -1020 7795 -986 7803
rect -1020 7735 -986 7757
rect -1020 7723 -986 7735
rect -1020 7667 -986 7685
rect -1020 7651 -986 7667
rect -1020 7599 -986 7613
rect -1020 7579 -986 7599
rect -1020 7531 -986 7541
rect -1020 7507 -986 7531
rect -1020 7463 -986 7469
rect -1020 7435 -986 7463
rect -1020 7395 -986 7397
rect -1020 7363 -986 7395
rect -1020 7293 -986 7325
rect -1020 7291 -986 7293
rect -1020 7225 -986 7253
rect -1020 7219 -986 7225
rect -1020 7157 -986 7181
rect -1020 7147 -986 7157
rect -1020 7089 -986 7109
rect -1020 7075 -986 7089
rect -1020 7021 -986 7037
rect -1020 7003 -986 7021
rect -1020 6953 -986 6965
rect -1020 6931 -986 6953
rect -1020 6885 -986 6893
rect -1020 6859 -986 6885
rect -1020 6817 -986 6821
rect -1020 6787 -986 6817
rect -1020 6715 -986 6749
rect -1020 6647 -986 6677
rect -1020 6643 -986 6647
rect -1020 6579 -986 6605
rect -1020 6571 -986 6579
rect -1020 6511 -986 6533
rect -1020 6499 -986 6511
rect -1020 6443 -986 6461
rect -1020 6427 -986 6443
rect -1020 6375 -986 6389
rect -1020 6355 -986 6375
rect -1020 6307 -986 6317
rect -1020 6283 -986 6307
rect -1020 6239 -986 6245
rect -1020 6211 -986 6239
rect -1020 6171 -986 6173
rect -1020 6139 -986 6171
rect -1020 6069 -986 6101
rect -1020 6067 -986 6069
rect -1020 6001 -986 6029
rect -1020 5995 -986 6001
rect -1020 5933 -986 5957
rect -1020 5923 -986 5933
rect -1020 5865 -986 5885
rect -1020 5851 -986 5865
rect -1020 5797 -986 5813
rect -1020 5779 -986 5797
rect -1020 5729 -986 5741
rect -1020 5707 -986 5729
rect -1020 5661 -986 5669
rect -1020 5635 -986 5661
rect -1020 5593 -986 5597
rect -1020 5563 -986 5593
rect -1020 5491 -986 5525
rect -1020 5423 -986 5453
rect -1020 5419 -986 5423
rect -1020 5355 -986 5381
rect -1020 5347 -986 5355
rect -1020 5287 -986 5309
rect -1020 5275 -986 5287
rect -1020 5219 -986 5237
rect -1020 5203 -986 5219
rect -1020 5151 -986 5165
rect -1020 5131 -986 5151
rect -1020 5083 -986 5093
rect -1020 5059 -986 5083
rect -1020 5015 -986 5021
rect -1020 4987 -986 5015
rect -1020 4947 -986 4949
rect -1020 4915 -986 4947
rect -1020 4845 -986 4877
rect -1020 4843 -986 4845
rect -1020 4777 -986 4805
rect -1020 4771 -986 4777
rect -1020 4709 -986 4733
rect -1020 4699 -986 4709
rect -1020 4641 -986 4661
rect -1020 4627 -986 4641
rect -1020 4573 -986 4589
rect -1020 4555 -986 4573
rect -1020 4505 -986 4517
rect -1020 4483 -986 4505
rect -1020 4437 -986 4445
rect -1020 4411 -986 4437
rect -1020 4369 -986 4373
rect -1020 4339 -986 4369
rect -1020 4267 -986 4301
rect -1020 4199 -986 4229
rect -1020 4195 -986 4199
rect -1020 4131 -986 4157
rect -1020 4123 -986 4131
rect -1020 4063 -986 4085
rect -1020 4051 -986 4063
rect -1020 3995 -986 4013
rect -1020 3979 -986 3995
rect -1020 3927 -986 3941
rect -1020 3907 -986 3927
rect -1020 3859 -986 3869
rect -1020 3835 -986 3859
rect -1020 3791 -986 3797
rect -1020 3763 -986 3791
rect -1020 3723 -986 3725
rect -1020 3691 -986 3723
rect -1020 3621 -986 3653
rect -1020 3619 -986 3621
rect -1020 3553 -986 3581
rect -1020 3547 -986 3553
rect -1020 3485 -986 3509
rect -1020 3475 -986 3485
rect -1020 3417 -986 3437
rect -1020 3403 -986 3417
rect -1020 3349 -986 3365
rect -1020 3331 -986 3349
rect -1020 3281 -986 3293
rect -1020 3259 -986 3281
rect -1020 3213 -986 3221
rect -1020 3187 -986 3213
rect -1020 3145 -986 3149
rect -1020 3115 -986 3145
rect -1020 3043 -986 3077
rect -1020 2975 -986 3005
rect -1020 2971 -986 2975
rect -1020 2907 -986 2933
rect -1020 2899 -986 2907
rect -1020 2839 -986 2861
rect -1020 2827 -986 2839
rect -1020 2771 -986 2789
rect -1020 2755 -986 2771
rect -1020 2703 -986 2717
rect -1020 2683 -986 2703
rect -1020 2635 -986 2645
rect -1020 2611 -986 2635
rect -1020 2567 -986 2573
rect -1020 2539 -986 2567
rect -1020 2499 -986 2501
rect -1020 2467 -986 2499
rect -1020 2397 -986 2429
rect -1020 2395 -986 2397
rect -1020 2329 -986 2357
rect -1020 2323 -986 2329
rect -1020 2261 -986 2285
rect -1020 2251 -986 2261
rect -1020 2193 -986 2213
rect -1020 2179 -986 2193
rect -1020 2125 -986 2141
rect -1020 2107 -986 2125
rect -1020 2057 -986 2069
rect -1020 2035 -986 2057
rect -1020 1989 -986 1997
rect -1020 1963 -986 1989
rect -1020 1921 -986 1925
rect -1020 1891 -986 1921
rect -1020 1819 -986 1853
rect -1020 1751 -986 1781
rect -1020 1747 -986 1751
rect -1020 1683 -986 1709
rect -1020 1675 -986 1683
rect -1020 1615 -986 1637
rect -1020 1603 -986 1615
rect -1020 1547 -986 1565
rect -1020 1531 -986 1547
rect -1020 1479 -986 1493
rect -1020 1459 -986 1479
rect -1020 1411 -986 1421
rect -1020 1387 -986 1411
rect -1020 1343 -986 1349
rect -1020 1315 -986 1343
rect -1020 1275 -986 1277
rect -1020 1243 -986 1275
rect -1020 1173 -986 1205
rect -1020 1171 -986 1173
rect -1020 1105 -986 1133
rect -1020 1099 -986 1105
rect -1020 1037 -986 1061
rect -1020 1027 -986 1037
rect -1020 969 -986 989
rect -1020 955 -986 969
rect -1020 901 -986 917
rect -1020 883 -986 901
rect -1020 833 -986 845
rect -1020 811 -986 833
rect -1020 765 -986 773
rect -1020 739 -986 765
rect -1020 697 -986 701
rect -1020 667 -986 697
rect -1020 595 -986 629
rect -1020 527 -986 557
rect -1020 523 -986 527
rect -1020 459 -986 485
rect -1020 451 -986 459
rect -1020 391 -986 413
rect -1020 379 -986 391
rect -1020 323 -986 341
rect -1020 307 -986 323
rect -1020 255 -986 269
rect -1020 235 -986 255
rect -1020 187 -986 197
rect -1020 163 -986 187
rect -1020 119 -986 125
rect -1020 91 -986 119
rect -1020 51 -986 53
rect -1020 19 -986 51
rect -1020 -51 -986 -19
rect -1020 -53 -986 -51
rect -1020 -119 -986 -91
rect -1020 -125 -986 -119
rect -1020 -187 -986 -163
rect -1020 -197 -986 -187
rect -1020 -255 -986 -235
rect -1020 -269 -986 -255
rect -1020 -323 -986 -307
rect -1020 -341 -986 -323
rect -1020 -391 -986 -379
rect -1020 -413 -986 -391
rect -1020 -459 -986 -451
rect -1020 -485 -986 -459
rect -1020 -527 -986 -523
rect -1020 -557 -986 -527
rect -1020 -629 -986 -595
rect -1020 -697 -986 -667
rect -1020 -701 -986 -697
rect -1020 -765 -986 -739
rect -1020 -773 -986 -765
rect -1020 -833 -986 -811
rect -1020 -845 -986 -833
rect -1020 -901 -986 -883
rect -1020 -917 -986 -901
rect -1020 -969 -986 -955
rect -1020 -989 -986 -969
rect -1020 -1037 -986 -1027
rect -1020 -1061 -986 -1037
rect -1020 -1105 -986 -1099
rect -1020 -1133 -986 -1105
rect -1020 -1173 -986 -1171
rect -1020 -1205 -986 -1173
rect -1020 -1275 -986 -1243
rect -1020 -1277 -986 -1275
rect -1020 -1343 -986 -1315
rect -1020 -1349 -986 -1343
rect -1020 -1411 -986 -1387
rect -1020 -1421 -986 -1411
rect -1020 -1479 -986 -1459
rect -1020 -1493 -986 -1479
rect -1020 -1547 -986 -1531
rect -1020 -1565 -986 -1547
rect -1020 -1615 -986 -1603
rect -1020 -1637 -986 -1615
rect -1020 -1683 -986 -1675
rect -1020 -1709 -986 -1683
rect -1020 -1751 -986 -1747
rect -1020 -1781 -986 -1751
rect -1020 -1853 -986 -1819
rect -1020 -1921 -986 -1891
rect -1020 -1925 -986 -1921
rect -1020 -1989 -986 -1963
rect -1020 -1997 -986 -1989
rect -1020 -2057 -986 -2035
rect -1020 -2069 -986 -2057
rect -1020 -2125 -986 -2107
rect -1020 -2141 -986 -2125
rect -1020 -2193 -986 -2179
rect -1020 -2213 -986 -2193
rect -1020 -2261 -986 -2251
rect -1020 -2285 -986 -2261
rect -1020 -2329 -986 -2323
rect -1020 -2357 -986 -2329
rect -1020 -2397 -986 -2395
rect -1020 -2429 -986 -2397
rect -1020 -2499 -986 -2467
rect -1020 -2501 -986 -2499
rect -1020 -2567 -986 -2539
rect -1020 -2573 -986 -2567
rect -1020 -2635 -986 -2611
rect -1020 -2645 -986 -2635
rect -1020 -2703 -986 -2683
rect -1020 -2717 -986 -2703
rect -1020 -2771 -986 -2755
rect -1020 -2789 -986 -2771
rect -1020 -2839 -986 -2827
rect -1020 -2861 -986 -2839
rect -1020 -2907 -986 -2899
rect -1020 -2933 -986 -2907
rect -1020 -2975 -986 -2971
rect -1020 -3005 -986 -2975
rect -1020 -3077 -986 -3043
rect -1020 -3145 -986 -3115
rect -1020 -3149 -986 -3145
rect -1020 -3213 -986 -3187
rect -1020 -3221 -986 -3213
rect -1020 -3281 -986 -3259
rect -1020 -3293 -986 -3281
rect -1020 -3349 -986 -3331
rect -1020 -3365 -986 -3349
rect -1020 -3417 -986 -3403
rect -1020 -3437 -986 -3417
rect -1020 -3485 -986 -3475
rect -1020 -3509 -986 -3485
rect -1020 -3553 -986 -3547
rect -1020 -3581 -986 -3553
rect -1020 -3621 -986 -3619
rect -1020 -3653 -986 -3621
rect -1020 -3723 -986 -3691
rect -1020 -3725 -986 -3723
rect -1020 -3791 -986 -3763
rect -1020 -3797 -986 -3791
rect -1020 -3859 -986 -3835
rect -1020 -3869 -986 -3859
rect -1020 -3927 -986 -3907
rect -1020 -3941 -986 -3927
rect -1020 -3995 -986 -3979
rect -1020 -4013 -986 -3995
rect -1020 -4063 -986 -4051
rect -1020 -4085 -986 -4063
rect -1020 -4131 -986 -4123
rect -1020 -4157 -986 -4131
rect -1020 -4199 -986 -4195
rect -1020 -4229 -986 -4199
rect -1020 -4301 -986 -4267
rect -1020 -4369 -986 -4339
rect -1020 -4373 -986 -4369
rect -1020 -4437 -986 -4411
rect -1020 -4445 -986 -4437
rect -1020 -4505 -986 -4483
rect -1020 -4517 -986 -4505
rect -1020 -4573 -986 -4555
rect -1020 -4589 -986 -4573
rect -1020 -4641 -986 -4627
rect -1020 -4661 -986 -4641
rect -1020 -4709 -986 -4699
rect -1020 -4733 -986 -4709
rect -1020 -4777 -986 -4771
rect -1020 -4805 -986 -4777
rect -1020 -4845 -986 -4843
rect -1020 -4877 -986 -4845
rect -1020 -4947 -986 -4915
rect -1020 -4949 -986 -4947
rect -1020 -5015 -986 -4987
rect -1020 -5021 -986 -5015
rect -1020 -5083 -986 -5059
rect -1020 -5093 -986 -5083
rect -1020 -5151 -986 -5131
rect -1020 -5165 -986 -5151
rect -1020 -5219 -986 -5203
rect -1020 -5237 -986 -5219
rect -1020 -5287 -986 -5275
rect -1020 -5309 -986 -5287
rect -1020 -5355 -986 -5347
rect -1020 -5381 -986 -5355
rect -1020 -5423 -986 -5419
rect -1020 -5453 -986 -5423
rect -1020 -5525 -986 -5491
rect -1020 -5593 -986 -5563
rect -1020 -5597 -986 -5593
rect -1020 -5661 -986 -5635
rect -1020 -5669 -986 -5661
rect -1020 -5729 -986 -5707
rect -1020 -5741 -986 -5729
rect -1020 -5797 -986 -5779
rect -1020 -5813 -986 -5797
rect -1020 -5865 -986 -5851
rect -1020 -5885 -986 -5865
rect -1020 -5933 -986 -5923
rect -1020 -5957 -986 -5933
rect -1020 -6001 -986 -5995
rect -1020 -6029 -986 -6001
rect -1020 -6069 -986 -6067
rect -1020 -6101 -986 -6069
rect -1020 -6171 -986 -6139
rect -1020 -6173 -986 -6171
rect -1020 -6239 -986 -6211
rect -1020 -6245 -986 -6239
rect -1020 -6307 -986 -6283
rect -1020 -6317 -986 -6307
rect -1020 -6375 -986 -6355
rect -1020 -6389 -986 -6375
rect -1020 -6443 -986 -6427
rect -1020 -6461 -986 -6443
rect -1020 -6511 -986 -6499
rect -1020 -6533 -986 -6511
rect -1020 -6579 -986 -6571
rect -1020 -6605 -986 -6579
rect -1020 -6647 -986 -6643
rect -1020 -6677 -986 -6647
rect -1020 -6749 -986 -6715
rect -1020 -6817 -986 -6787
rect -1020 -6821 -986 -6817
rect -1020 -6885 -986 -6859
rect -1020 -6893 -986 -6885
rect -1020 -6953 -986 -6931
rect -1020 -6965 -986 -6953
rect -1020 -7021 -986 -7003
rect -1020 -7037 -986 -7021
rect -1020 -7089 -986 -7075
rect -1020 -7109 -986 -7089
rect -1020 -7157 -986 -7147
rect -1020 -7181 -986 -7157
rect -1020 -7225 -986 -7219
rect -1020 -7253 -986 -7225
rect -1020 -7293 -986 -7291
rect -1020 -7325 -986 -7293
rect -1020 -7395 -986 -7363
rect -1020 -7397 -986 -7395
rect -1020 -7463 -986 -7435
rect -1020 -7469 -986 -7463
rect -1020 -7531 -986 -7507
rect -1020 -7541 -986 -7531
rect -1020 -7599 -986 -7579
rect -1020 -7613 -986 -7599
rect -1020 -7667 -986 -7651
rect -1020 -7685 -986 -7667
rect -1020 -7735 -986 -7723
rect -1020 -7757 -986 -7735
rect -1020 -7803 -986 -7795
rect -1020 -7829 -986 -7803
rect -1020 -7871 -986 -7867
rect -1020 -7901 -986 -7871
rect -1020 -7973 -986 -7939
rect -1020 -8041 -986 -8011
rect -1020 -8045 -986 -8041
rect -1020 -8109 -986 -8083
rect -1020 -8117 -986 -8109
rect -1020 -8177 -986 -8155
rect -1020 -8189 -986 -8177
rect -1020 -8245 -986 -8227
rect -1020 -8261 -986 -8245
rect -1020 -8313 -986 -8299
rect -1020 -8333 -986 -8313
rect -1020 -8381 -986 -8371
rect -1020 -8405 -986 -8381
rect -1020 -8449 -986 -8443
rect -1020 -8477 -986 -8449
rect -1020 -8517 -986 -8515
rect -1020 -8549 -986 -8517
rect -1020 -8619 -986 -8587
rect -1020 -8621 -986 -8619
rect -1020 -8687 -986 -8659
rect -1020 -8693 -986 -8687
rect -1020 -8755 -986 -8731
rect -1020 -8765 -986 -8755
rect -1020 -8823 -986 -8803
rect -1020 -8837 -986 -8823
rect -1020 -8891 -986 -8875
rect -1020 -8909 -986 -8891
rect -1020 -8959 -986 -8947
rect -1020 -8981 -986 -8959
rect -1020 -9027 -986 -9019
rect -1020 -9053 -986 -9027
rect -1020 -9095 -986 -9091
rect -1020 -9125 -986 -9095
rect -1020 -9197 -986 -9163
rect -1020 -9265 -986 -9235
rect -1020 -9269 -986 -9265
rect -1020 -9333 -986 -9307
rect -1020 -9341 -986 -9333
rect -1020 -9401 -986 -9379
rect -1020 -9413 -986 -9401
rect -1020 -9469 -986 -9451
rect -1020 -9485 -986 -9469
rect -1020 -9537 -986 -9523
rect -1020 -9557 -986 -9537
rect -902 9537 -868 9557
rect -902 9523 -868 9537
rect -902 9469 -868 9485
rect -902 9451 -868 9469
rect -902 9401 -868 9413
rect -902 9379 -868 9401
rect -902 9333 -868 9341
rect -902 9307 -868 9333
rect -902 9265 -868 9269
rect -902 9235 -868 9265
rect -902 9163 -868 9197
rect -902 9095 -868 9125
rect -902 9091 -868 9095
rect -902 9027 -868 9053
rect -902 9019 -868 9027
rect -902 8959 -868 8981
rect -902 8947 -868 8959
rect -902 8891 -868 8909
rect -902 8875 -868 8891
rect -902 8823 -868 8837
rect -902 8803 -868 8823
rect -902 8755 -868 8765
rect -902 8731 -868 8755
rect -902 8687 -868 8693
rect -902 8659 -868 8687
rect -902 8619 -868 8621
rect -902 8587 -868 8619
rect -902 8517 -868 8549
rect -902 8515 -868 8517
rect -902 8449 -868 8477
rect -902 8443 -868 8449
rect -902 8381 -868 8405
rect -902 8371 -868 8381
rect -902 8313 -868 8333
rect -902 8299 -868 8313
rect -902 8245 -868 8261
rect -902 8227 -868 8245
rect -902 8177 -868 8189
rect -902 8155 -868 8177
rect -902 8109 -868 8117
rect -902 8083 -868 8109
rect -902 8041 -868 8045
rect -902 8011 -868 8041
rect -902 7939 -868 7973
rect -902 7871 -868 7901
rect -902 7867 -868 7871
rect -902 7803 -868 7829
rect -902 7795 -868 7803
rect -902 7735 -868 7757
rect -902 7723 -868 7735
rect -902 7667 -868 7685
rect -902 7651 -868 7667
rect -902 7599 -868 7613
rect -902 7579 -868 7599
rect -902 7531 -868 7541
rect -902 7507 -868 7531
rect -902 7463 -868 7469
rect -902 7435 -868 7463
rect -902 7395 -868 7397
rect -902 7363 -868 7395
rect -902 7293 -868 7325
rect -902 7291 -868 7293
rect -902 7225 -868 7253
rect -902 7219 -868 7225
rect -902 7157 -868 7181
rect -902 7147 -868 7157
rect -902 7089 -868 7109
rect -902 7075 -868 7089
rect -902 7021 -868 7037
rect -902 7003 -868 7021
rect -902 6953 -868 6965
rect -902 6931 -868 6953
rect -902 6885 -868 6893
rect -902 6859 -868 6885
rect -902 6817 -868 6821
rect -902 6787 -868 6817
rect -902 6715 -868 6749
rect -902 6647 -868 6677
rect -902 6643 -868 6647
rect -902 6579 -868 6605
rect -902 6571 -868 6579
rect -902 6511 -868 6533
rect -902 6499 -868 6511
rect -902 6443 -868 6461
rect -902 6427 -868 6443
rect -902 6375 -868 6389
rect -902 6355 -868 6375
rect -902 6307 -868 6317
rect -902 6283 -868 6307
rect -902 6239 -868 6245
rect -902 6211 -868 6239
rect -902 6171 -868 6173
rect -902 6139 -868 6171
rect -902 6069 -868 6101
rect -902 6067 -868 6069
rect -902 6001 -868 6029
rect -902 5995 -868 6001
rect -902 5933 -868 5957
rect -902 5923 -868 5933
rect -902 5865 -868 5885
rect -902 5851 -868 5865
rect -902 5797 -868 5813
rect -902 5779 -868 5797
rect -902 5729 -868 5741
rect -902 5707 -868 5729
rect -902 5661 -868 5669
rect -902 5635 -868 5661
rect -902 5593 -868 5597
rect -902 5563 -868 5593
rect -902 5491 -868 5525
rect -902 5423 -868 5453
rect -902 5419 -868 5423
rect -902 5355 -868 5381
rect -902 5347 -868 5355
rect -902 5287 -868 5309
rect -902 5275 -868 5287
rect -902 5219 -868 5237
rect -902 5203 -868 5219
rect -902 5151 -868 5165
rect -902 5131 -868 5151
rect -902 5083 -868 5093
rect -902 5059 -868 5083
rect -902 5015 -868 5021
rect -902 4987 -868 5015
rect -902 4947 -868 4949
rect -902 4915 -868 4947
rect -902 4845 -868 4877
rect -902 4843 -868 4845
rect -902 4777 -868 4805
rect -902 4771 -868 4777
rect -902 4709 -868 4733
rect -902 4699 -868 4709
rect -902 4641 -868 4661
rect -902 4627 -868 4641
rect -902 4573 -868 4589
rect -902 4555 -868 4573
rect -902 4505 -868 4517
rect -902 4483 -868 4505
rect -902 4437 -868 4445
rect -902 4411 -868 4437
rect -902 4369 -868 4373
rect -902 4339 -868 4369
rect -902 4267 -868 4301
rect -902 4199 -868 4229
rect -902 4195 -868 4199
rect -902 4131 -868 4157
rect -902 4123 -868 4131
rect -902 4063 -868 4085
rect -902 4051 -868 4063
rect -902 3995 -868 4013
rect -902 3979 -868 3995
rect -902 3927 -868 3941
rect -902 3907 -868 3927
rect -902 3859 -868 3869
rect -902 3835 -868 3859
rect -902 3791 -868 3797
rect -902 3763 -868 3791
rect -902 3723 -868 3725
rect -902 3691 -868 3723
rect -902 3621 -868 3653
rect -902 3619 -868 3621
rect -902 3553 -868 3581
rect -902 3547 -868 3553
rect -902 3485 -868 3509
rect -902 3475 -868 3485
rect -902 3417 -868 3437
rect -902 3403 -868 3417
rect -902 3349 -868 3365
rect -902 3331 -868 3349
rect -902 3281 -868 3293
rect -902 3259 -868 3281
rect -902 3213 -868 3221
rect -902 3187 -868 3213
rect -902 3145 -868 3149
rect -902 3115 -868 3145
rect -902 3043 -868 3077
rect -902 2975 -868 3005
rect -902 2971 -868 2975
rect -902 2907 -868 2933
rect -902 2899 -868 2907
rect -902 2839 -868 2861
rect -902 2827 -868 2839
rect -902 2771 -868 2789
rect -902 2755 -868 2771
rect -902 2703 -868 2717
rect -902 2683 -868 2703
rect -902 2635 -868 2645
rect -902 2611 -868 2635
rect -902 2567 -868 2573
rect -902 2539 -868 2567
rect -902 2499 -868 2501
rect -902 2467 -868 2499
rect -902 2397 -868 2429
rect -902 2395 -868 2397
rect -902 2329 -868 2357
rect -902 2323 -868 2329
rect -902 2261 -868 2285
rect -902 2251 -868 2261
rect -902 2193 -868 2213
rect -902 2179 -868 2193
rect -902 2125 -868 2141
rect -902 2107 -868 2125
rect -902 2057 -868 2069
rect -902 2035 -868 2057
rect -902 1989 -868 1997
rect -902 1963 -868 1989
rect -902 1921 -868 1925
rect -902 1891 -868 1921
rect -902 1819 -868 1853
rect -902 1751 -868 1781
rect -902 1747 -868 1751
rect -902 1683 -868 1709
rect -902 1675 -868 1683
rect -902 1615 -868 1637
rect -902 1603 -868 1615
rect -902 1547 -868 1565
rect -902 1531 -868 1547
rect -902 1479 -868 1493
rect -902 1459 -868 1479
rect -902 1411 -868 1421
rect -902 1387 -868 1411
rect -902 1343 -868 1349
rect -902 1315 -868 1343
rect -902 1275 -868 1277
rect -902 1243 -868 1275
rect -902 1173 -868 1205
rect -902 1171 -868 1173
rect -902 1105 -868 1133
rect -902 1099 -868 1105
rect -902 1037 -868 1061
rect -902 1027 -868 1037
rect -902 969 -868 989
rect -902 955 -868 969
rect -902 901 -868 917
rect -902 883 -868 901
rect -902 833 -868 845
rect -902 811 -868 833
rect -902 765 -868 773
rect -902 739 -868 765
rect -902 697 -868 701
rect -902 667 -868 697
rect -902 595 -868 629
rect -902 527 -868 557
rect -902 523 -868 527
rect -902 459 -868 485
rect -902 451 -868 459
rect -902 391 -868 413
rect -902 379 -868 391
rect -902 323 -868 341
rect -902 307 -868 323
rect -902 255 -868 269
rect -902 235 -868 255
rect -902 187 -868 197
rect -902 163 -868 187
rect -902 119 -868 125
rect -902 91 -868 119
rect -902 51 -868 53
rect -902 19 -868 51
rect -902 -51 -868 -19
rect -902 -53 -868 -51
rect -902 -119 -868 -91
rect -902 -125 -868 -119
rect -902 -187 -868 -163
rect -902 -197 -868 -187
rect -902 -255 -868 -235
rect -902 -269 -868 -255
rect -902 -323 -868 -307
rect -902 -341 -868 -323
rect -902 -391 -868 -379
rect -902 -413 -868 -391
rect -902 -459 -868 -451
rect -902 -485 -868 -459
rect -902 -527 -868 -523
rect -902 -557 -868 -527
rect -902 -629 -868 -595
rect -902 -697 -868 -667
rect -902 -701 -868 -697
rect -902 -765 -868 -739
rect -902 -773 -868 -765
rect -902 -833 -868 -811
rect -902 -845 -868 -833
rect -902 -901 -868 -883
rect -902 -917 -868 -901
rect -902 -969 -868 -955
rect -902 -989 -868 -969
rect -902 -1037 -868 -1027
rect -902 -1061 -868 -1037
rect -902 -1105 -868 -1099
rect -902 -1133 -868 -1105
rect -902 -1173 -868 -1171
rect -902 -1205 -868 -1173
rect -902 -1275 -868 -1243
rect -902 -1277 -868 -1275
rect -902 -1343 -868 -1315
rect -902 -1349 -868 -1343
rect -902 -1411 -868 -1387
rect -902 -1421 -868 -1411
rect -902 -1479 -868 -1459
rect -902 -1493 -868 -1479
rect -902 -1547 -868 -1531
rect -902 -1565 -868 -1547
rect -902 -1615 -868 -1603
rect -902 -1637 -868 -1615
rect -902 -1683 -868 -1675
rect -902 -1709 -868 -1683
rect -902 -1751 -868 -1747
rect -902 -1781 -868 -1751
rect -902 -1853 -868 -1819
rect -902 -1921 -868 -1891
rect -902 -1925 -868 -1921
rect -902 -1989 -868 -1963
rect -902 -1997 -868 -1989
rect -902 -2057 -868 -2035
rect -902 -2069 -868 -2057
rect -902 -2125 -868 -2107
rect -902 -2141 -868 -2125
rect -902 -2193 -868 -2179
rect -902 -2213 -868 -2193
rect -902 -2261 -868 -2251
rect -902 -2285 -868 -2261
rect -902 -2329 -868 -2323
rect -902 -2357 -868 -2329
rect -902 -2397 -868 -2395
rect -902 -2429 -868 -2397
rect -902 -2499 -868 -2467
rect -902 -2501 -868 -2499
rect -902 -2567 -868 -2539
rect -902 -2573 -868 -2567
rect -902 -2635 -868 -2611
rect -902 -2645 -868 -2635
rect -902 -2703 -868 -2683
rect -902 -2717 -868 -2703
rect -902 -2771 -868 -2755
rect -902 -2789 -868 -2771
rect -902 -2839 -868 -2827
rect -902 -2861 -868 -2839
rect -902 -2907 -868 -2899
rect -902 -2933 -868 -2907
rect -902 -2975 -868 -2971
rect -902 -3005 -868 -2975
rect -902 -3077 -868 -3043
rect -902 -3145 -868 -3115
rect -902 -3149 -868 -3145
rect -902 -3213 -868 -3187
rect -902 -3221 -868 -3213
rect -902 -3281 -868 -3259
rect -902 -3293 -868 -3281
rect -902 -3349 -868 -3331
rect -902 -3365 -868 -3349
rect -902 -3417 -868 -3403
rect -902 -3437 -868 -3417
rect -902 -3485 -868 -3475
rect -902 -3509 -868 -3485
rect -902 -3553 -868 -3547
rect -902 -3581 -868 -3553
rect -902 -3621 -868 -3619
rect -902 -3653 -868 -3621
rect -902 -3723 -868 -3691
rect -902 -3725 -868 -3723
rect -902 -3791 -868 -3763
rect -902 -3797 -868 -3791
rect -902 -3859 -868 -3835
rect -902 -3869 -868 -3859
rect -902 -3927 -868 -3907
rect -902 -3941 -868 -3927
rect -902 -3995 -868 -3979
rect -902 -4013 -868 -3995
rect -902 -4063 -868 -4051
rect -902 -4085 -868 -4063
rect -902 -4131 -868 -4123
rect -902 -4157 -868 -4131
rect -902 -4199 -868 -4195
rect -902 -4229 -868 -4199
rect -902 -4301 -868 -4267
rect -902 -4369 -868 -4339
rect -902 -4373 -868 -4369
rect -902 -4437 -868 -4411
rect -902 -4445 -868 -4437
rect -902 -4505 -868 -4483
rect -902 -4517 -868 -4505
rect -902 -4573 -868 -4555
rect -902 -4589 -868 -4573
rect -902 -4641 -868 -4627
rect -902 -4661 -868 -4641
rect -902 -4709 -868 -4699
rect -902 -4733 -868 -4709
rect -902 -4777 -868 -4771
rect -902 -4805 -868 -4777
rect -902 -4845 -868 -4843
rect -902 -4877 -868 -4845
rect -902 -4947 -868 -4915
rect -902 -4949 -868 -4947
rect -902 -5015 -868 -4987
rect -902 -5021 -868 -5015
rect -902 -5083 -868 -5059
rect -902 -5093 -868 -5083
rect -902 -5151 -868 -5131
rect -902 -5165 -868 -5151
rect -902 -5219 -868 -5203
rect -902 -5237 -868 -5219
rect -902 -5287 -868 -5275
rect -902 -5309 -868 -5287
rect -902 -5355 -868 -5347
rect -902 -5381 -868 -5355
rect -902 -5423 -868 -5419
rect -902 -5453 -868 -5423
rect -902 -5525 -868 -5491
rect -902 -5593 -868 -5563
rect -902 -5597 -868 -5593
rect -902 -5661 -868 -5635
rect -902 -5669 -868 -5661
rect -902 -5729 -868 -5707
rect -902 -5741 -868 -5729
rect -902 -5797 -868 -5779
rect -902 -5813 -868 -5797
rect -902 -5865 -868 -5851
rect -902 -5885 -868 -5865
rect -902 -5933 -868 -5923
rect -902 -5957 -868 -5933
rect -902 -6001 -868 -5995
rect -902 -6029 -868 -6001
rect -902 -6069 -868 -6067
rect -902 -6101 -868 -6069
rect -902 -6171 -868 -6139
rect -902 -6173 -868 -6171
rect -902 -6239 -868 -6211
rect -902 -6245 -868 -6239
rect -902 -6307 -868 -6283
rect -902 -6317 -868 -6307
rect -902 -6375 -868 -6355
rect -902 -6389 -868 -6375
rect -902 -6443 -868 -6427
rect -902 -6461 -868 -6443
rect -902 -6511 -868 -6499
rect -902 -6533 -868 -6511
rect -902 -6579 -868 -6571
rect -902 -6605 -868 -6579
rect -902 -6647 -868 -6643
rect -902 -6677 -868 -6647
rect -902 -6749 -868 -6715
rect -902 -6817 -868 -6787
rect -902 -6821 -868 -6817
rect -902 -6885 -868 -6859
rect -902 -6893 -868 -6885
rect -902 -6953 -868 -6931
rect -902 -6965 -868 -6953
rect -902 -7021 -868 -7003
rect -902 -7037 -868 -7021
rect -902 -7089 -868 -7075
rect -902 -7109 -868 -7089
rect -902 -7157 -868 -7147
rect -902 -7181 -868 -7157
rect -902 -7225 -868 -7219
rect -902 -7253 -868 -7225
rect -902 -7293 -868 -7291
rect -902 -7325 -868 -7293
rect -902 -7395 -868 -7363
rect -902 -7397 -868 -7395
rect -902 -7463 -868 -7435
rect -902 -7469 -868 -7463
rect -902 -7531 -868 -7507
rect -902 -7541 -868 -7531
rect -902 -7599 -868 -7579
rect -902 -7613 -868 -7599
rect -902 -7667 -868 -7651
rect -902 -7685 -868 -7667
rect -902 -7735 -868 -7723
rect -902 -7757 -868 -7735
rect -902 -7803 -868 -7795
rect -902 -7829 -868 -7803
rect -902 -7871 -868 -7867
rect -902 -7901 -868 -7871
rect -902 -7973 -868 -7939
rect -902 -8041 -868 -8011
rect -902 -8045 -868 -8041
rect -902 -8109 -868 -8083
rect -902 -8117 -868 -8109
rect -902 -8177 -868 -8155
rect -902 -8189 -868 -8177
rect -902 -8245 -868 -8227
rect -902 -8261 -868 -8245
rect -902 -8313 -868 -8299
rect -902 -8333 -868 -8313
rect -902 -8381 -868 -8371
rect -902 -8405 -868 -8381
rect -902 -8449 -868 -8443
rect -902 -8477 -868 -8449
rect -902 -8517 -868 -8515
rect -902 -8549 -868 -8517
rect -902 -8619 -868 -8587
rect -902 -8621 -868 -8619
rect -902 -8687 -868 -8659
rect -902 -8693 -868 -8687
rect -902 -8755 -868 -8731
rect -902 -8765 -868 -8755
rect -902 -8823 -868 -8803
rect -902 -8837 -868 -8823
rect -902 -8891 -868 -8875
rect -902 -8909 -868 -8891
rect -902 -8959 -868 -8947
rect -902 -8981 -868 -8959
rect -902 -9027 -868 -9019
rect -902 -9053 -868 -9027
rect -902 -9095 -868 -9091
rect -902 -9125 -868 -9095
rect -902 -9197 -868 -9163
rect -902 -9265 -868 -9235
rect -902 -9269 -868 -9265
rect -902 -9333 -868 -9307
rect -902 -9341 -868 -9333
rect -902 -9401 -868 -9379
rect -902 -9413 -868 -9401
rect -902 -9469 -868 -9451
rect -902 -9485 -868 -9469
rect -902 -9537 -868 -9523
rect -902 -9557 -868 -9537
rect -784 9537 -750 9557
rect -784 9523 -750 9537
rect -784 9469 -750 9485
rect -784 9451 -750 9469
rect -784 9401 -750 9413
rect -784 9379 -750 9401
rect -784 9333 -750 9341
rect -784 9307 -750 9333
rect -784 9265 -750 9269
rect -784 9235 -750 9265
rect -784 9163 -750 9197
rect -784 9095 -750 9125
rect -784 9091 -750 9095
rect -784 9027 -750 9053
rect -784 9019 -750 9027
rect -784 8959 -750 8981
rect -784 8947 -750 8959
rect -784 8891 -750 8909
rect -784 8875 -750 8891
rect -784 8823 -750 8837
rect -784 8803 -750 8823
rect -784 8755 -750 8765
rect -784 8731 -750 8755
rect -784 8687 -750 8693
rect -784 8659 -750 8687
rect -784 8619 -750 8621
rect -784 8587 -750 8619
rect -784 8517 -750 8549
rect -784 8515 -750 8517
rect -784 8449 -750 8477
rect -784 8443 -750 8449
rect -784 8381 -750 8405
rect -784 8371 -750 8381
rect -784 8313 -750 8333
rect -784 8299 -750 8313
rect -784 8245 -750 8261
rect -784 8227 -750 8245
rect -784 8177 -750 8189
rect -784 8155 -750 8177
rect -784 8109 -750 8117
rect -784 8083 -750 8109
rect -784 8041 -750 8045
rect -784 8011 -750 8041
rect -784 7939 -750 7973
rect -784 7871 -750 7901
rect -784 7867 -750 7871
rect -784 7803 -750 7829
rect -784 7795 -750 7803
rect -784 7735 -750 7757
rect -784 7723 -750 7735
rect -784 7667 -750 7685
rect -784 7651 -750 7667
rect -784 7599 -750 7613
rect -784 7579 -750 7599
rect -784 7531 -750 7541
rect -784 7507 -750 7531
rect -784 7463 -750 7469
rect -784 7435 -750 7463
rect -784 7395 -750 7397
rect -784 7363 -750 7395
rect -784 7293 -750 7325
rect -784 7291 -750 7293
rect -784 7225 -750 7253
rect -784 7219 -750 7225
rect -784 7157 -750 7181
rect -784 7147 -750 7157
rect -784 7089 -750 7109
rect -784 7075 -750 7089
rect -784 7021 -750 7037
rect -784 7003 -750 7021
rect -784 6953 -750 6965
rect -784 6931 -750 6953
rect -784 6885 -750 6893
rect -784 6859 -750 6885
rect -784 6817 -750 6821
rect -784 6787 -750 6817
rect -784 6715 -750 6749
rect -784 6647 -750 6677
rect -784 6643 -750 6647
rect -784 6579 -750 6605
rect -784 6571 -750 6579
rect -784 6511 -750 6533
rect -784 6499 -750 6511
rect -784 6443 -750 6461
rect -784 6427 -750 6443
rect -784 6375 -750 6389
rect -784 6355 -750 6375
rect -784 6307 -750 6317
rect -784 6283 -750 6307
rect -784 6239 -750 6245
rect -784 6211 -750 6239
rect -784 6171 -750 6173
rect -784 6139 -750 6171
rect -784 6069 -750 6101
rect -784 6067 -750 6069
rect -784 6001 -750 6029
rect -784 5995 -750 6001
rect -784 5933 -750 5957
rect -784 5923 -750 5933
rect -784 5865 -750 5885
rect -784 5851 -750 5865
rect -784 5797 -750 5813
rect -784 5779 -750 5797
rect -784 5729 -750 5741
rect -784 5707 -750 5729
rect -784 5661 -750 5669
rect -784 5635 -750 5661
rect -784 5593 -750 5597
rect -784 5563 -750 5593
rect -784 5491 -750 5525
rect -784 5423 -750 5453
rect -784 5419 -750 5423
rect -784 5355 -750 5381
rect -784 5347 -750 5355
rect -784 5287 -750 5309
rect -784 5275 -750 5287
rect -784 5219 -750 5237
rect -784 5203 -750 5219
rect -784 5151 -750 5165
rect -784 5131 -750 5151
rect -784 5083 -750 5093
rect -784 5059 -750 5083
rect -784 5015 -750 5021
rect -784 4987 -750 5015
rect -784 4947 -750 4949
rect -784 4915 -750 4947
rect -784 4845 -750 4877
rect -784 4843 -750 4845
rect -784 4777 -750 4805
rect -784 4771 -750 4777
rect -784 4709 -750 4733
rect -784 4699 -750 4709
rect -784 4641 -750 4661
rect -784 4627 -750 4641
rect -784 4573 -750 4589
rect -784 4555 -750 4573
rect -784 4505 -750 4517
rect -784 4483 -750 4505
rect -784 4437 -750 4445
rect -784 4411 -750 4437
rect -784 4369 -750 4373
rect -784 4339 -750 4369
rect -784 4267 -750 4301
rect -784 4199 -750 4229
rect -784 4195 -750 4199
rect -784 4131 -750 4157
rect -784 4123 -750 4131
rect -784 4063 -750 4085
rect -784 4051 -750 4063
rect -784 3995 -750 4013
rect -784 3979 -750 3995
rect -784 3927 -750 3941
rect -784 3907 -750 3927
rect -784 3859 -750 3869
rect -784 3835 -750 3859
rect -784 3791 -750 3797
rect -784 3763 -750 3791
rect -784 3723 -750 3725
rect -784 3691 -750 3723
rect -784 3621 -750 3653
rect -784 3619 -750 3621
rect -784 3553 -750 3581
rect -784 3547 -750 3553
rect -784 3485 -750 3509
rect -784 3475 -750 3485
rect -784 3417 -750 3437
rect -784 3403 -750 3417
rect -784 3349 -750 3365
rect -784 3331 -750 3349
rect -784 3281 -750 3293
rect -784 3259 -750 3281
rect -784 3213 -750 3221
rect -784 3187 -750 3213
rect -784 3145 -750 3149
rect -784 3115 -750 3145
rect -784 3043 -750 3077
rect -784 2975 -750 3005
rect -784 2971 -750 2975
rect -784 2907 -750 2933
rect -784 2899 -750 2907
rect -784 2839 -750 2861
rect -784 2827 -750 2839
rect -784 2771 -750 2789
rect -784 2755 -750 2771
rect -784 2703 -750 2717
rect -784 2683 -750 2703
rect -784 2635 -750 2645
rect -784 2611 -750 2635
rect -784 2567 -750 2573
rect -784 2539 -750 2567
rect -784 2499 -750 2501
rect -784 2467 -750 2499
rect -784 2397 -750 2429
rect -784 2395 -750 2397
rect -784 2329 -750 2357
rect -784 2323 -750 2329
rect -784 2261 -750 2285
rect -784 2251 -750 2261
rect -784 2193 -750 2213
rect -784 2179 -750 2193
rect -784 2125 -750 2141
rect -784 2107 -750 2125
rect -784 2057 -750 2069
rect -784 2035 -750 2057
rect -784 1989 -750 1997
rect -784 1963 -750 1989
rect -784 1921 -750 1925
rect -784 1891 -750 1921
rect -784 1819 -750 1853
rect -784 1751 -750 1781
rect -784 1747 -750 1751
rect -784 1683 -750 1709
rect -784 1675 -750 1683
rect -784 1615 -750 1637
rect -784 1603 -750 1615
rect -784 1547 -750 1565
rect -784 1531 -750 1547
rect -784 1479 -750 1493
rect -784 1459 -750 1479
rect -784 1411 -750 1421
rect -784 1387 -750 1411
rect -784 1343 -750 1349
rect -784 1315 -750 1343
rect -784 1275 -750 1277
rect -784 1243 -750 1275
rect -784 1173 -750 1205
rect -784 1171 -750 1173
rect -784 1105 -750 1133
rect -784 1099 -750 1105
rect -784 1037 -750 1061
rect -784 1027 -750 1037
rect -784 969 -750 989
rect -784 955 -750 969
rect -784 901 -750 917
rect -784 883 -750 901
rect -784 833 -750 845
rect -784 811 -750 833
rect -784 765 -750 773
rect -784 739 -750 765
rect -784 697 -750 701
rect -784 667 -750 697
rect -784 595 -750 629
rect -784 527 -750 557
rect -784 523 -750 527
rect -784 459 -750 485
rect -784 451 -750 459
rect -784 391 -750 413
rect -784 379 -750 391
rect -784 323 -750 341
rect -784 307 -750 323
rect -784 255 -750 269
rect -784 235 -750 255
rect -784 187 -750 197
rect -784 163 -750 187
rect -784 119 -750 125
rect -784 91 -750 119
rect -784 51 -750 53
rect -784 19 -750 51
rect -784 -51 -750 -19
rect -784 -53 -750 -51
rect -784 -119 -750 -91
rect -784 -125 -750 -119
rect -784 -187 -750 -163
rect -784 -197 -750 -187
rect -784 -255 -750 -235
rect -784 -269 -750 -255
rect -784 -323 -750 -307
rect -784 -341 -750 -323
rect -784 -391 -750 -379
rect -784 -413 -750 -391
rect -784 -459 -750 -451
rect -784 -485 -750 -459
rect -784 -527 -750 -523
rect -784 -557 -750 -527
rect -784 -629 -750 -595
rect -784 -697 -750 -667
rect -784 -701 -750 -697
rect -784 -765 -750 -739
rect -784 -773 -750 -765
rect -784 -833 -750 -811
rect -784 -845 -750 -833
rect -784 -901 -750 -883
rect -784 -917 -750 -901
rect -784 -969 -750 -955
rect -784 -989 -750 -969
rect -784 -1037 -750 -1027
rect -784 -1061 -750 -1037
rect -784 -1105 -750 -1099
rect -784 -1133 -750 -1105
rect -784 -1173 -750 -1171
rect -784 -1205 -750 -1173
rect -784 -1275 -750 -1243
rect -784 -1277 -750 -1275
rect -784 -1343 -750 -1315
rect -784 -1349 -750 -1343
rect -784 -1411 -750 -1387
rect -784 -1421 -750 -1411
rect -784 -1479 -750 -1459
rect -784 -1493 -750 -1479
rect -784 -1547 -750 -1531
rect -784 -1565 -750 -1547
rect -784 -1615 -750 -1603
rect -784 -1637 -750 -1615
rect -784 -1683 -750 -1675
rect -784 -1709 -750 -1683
rect -784 -1751 -750 -1747
rect -784 -1781 -750 -1751
rect -784 -1853 -750 -1819
rect -784 -1921 -750 -1891
rect -784 -1925 -750 -1921
rect -784 -1989 -750 -1963
rect -784 -1997 -750 -1989
rect -784 -2057 -750 -2035
rect -784 -2069 -750 -2057
rect -784 -2125 -750 -2107
rect -784 -2141 -750 -2125
rect -784 -2193 -750 -2179
rect -784 -2213 -750 -2193
rect -784 -2261 -750 -2251
rect -784 -2285 -750 -2261
rect -784 -2329 -750 -2323
rect -784 -2357 -750 -2329
rect -784 -2397 -750 -2395
rect -784 -2429 -750 -2397
rect -784 -2499 -750 -2467
rect -784 -2501 -750 -2499
rect -784 -2567 -750 -2539
rect -784 -2573 -750 -2567
rect -784 -2635 -750 -2611
rect -784 -2645 -750 -2635
rect -784 -2703 -750 -2683
rect -784 -2717 -750 -2703
rect -784 -2771 -750 -2755
rect -784 -2789 -750 -2771
rect -784 -2839 -750 -2827
rect -784 -2861 -750 -2839
rect -784 -2907 -750 -2899
rect -784 -2933 -750 -2907
rect -784 -2975 -750 -2971
rect -784 -3005 -750 -2975
rect -784 -3077 -750 -3043
rect -784 -3145 -750 -3115
rect -784 -3149 -750 -3145
rect -784 -3213 -750 -3187
rect -784 -3221 -750 -3213
rect -784 -3281 -750 -3259
rect -784 -3293 -750 -3281
rect -784 -3349 -750 -3331
rect -784 -3365 -750 -3349
rect -784 -3417 -750 -3403
rect -784 -3437 -750 -3417
rect -784 -3485 -750 -3475
rect -784 -3509 -750 -3485
rect -784 -3553 -750 -3547
rect -784 -3581 -750 -3553
rect -784 -3621 -750 -3619
rect -784 -3653 -750 -3621
rect -784 -3723 -750 -3691
rect -784 -3725 -750 -3723
rect -784 -3791 -750 -3763
rect -784 -3797 -750 -3791
rect -784 -3859 -750 -3835
rect -784 -3869 -750 -3859
rect -784 -3927 -750 -3907
rect -784 -3941 -750 -3927
rect -784 -3995 -750 -3979
rect -784 -4013 -750 -3995
rect -784 -4063 -750 -4051
rect -784 -4085 -750 -4063
rect -784 -4131 -750 -4123
rect -784 -4157 -750 -4131
rect -784 -4199 -750 -4195
rect -784 -4229 -750 -4199
rect -784 -4301 -750 -4267
rect -784 -4369 -750 -4339
rect -784 -4373 -750 -4369
rect -784 -4437 -750 -4411
rect -784 -4445 -750 -4437
rect -784 -4505 -750 -4483
rect -784 -4517 -750 -4505
rect -784 -4573 -750 -4555
rect -784 -4589 -750 -4573
rect -784 -4641 -750 -4627
rect -784 -4661 -750 -4641
rect -784 -4709 -750 -4699
rect -784 -4733 -750 -4709
rect -784 -4777 -750 -4771
rect -784 -4805 -750 -4777
rect -784 -4845 -750 -4843
rect -784 -4877 -750 -4845
rect -784 -4947 -750 -4915
rect -784 -4949 -750 -4947
rect -784 -5015 -750 -4987
rect -784 -5021 -750 -5015
rect -784 -5083 -750 -5059
rect -784 -5093 -750 -5083
rect -784 -5151 -750 -5131
rect -784 -5165 -750 -5151
rect -784 -5219 -750 -5203
rect -784 -5237 -750 -5219
rect -784 -5287 -750 -5275
rect -784 -5309 -750 -5287
rect -784 -5355 -750 -5347
rect -784 -5381 -750 -5355
rect -784 -5423 -750 -5419
rect -784 -5453 -750 -5423
rect -784 -5525 -750 -5491
rect -784 -5593 -750 -5563
rect -784 -5597 -750 -5593
rect -784 -5661 -750 -5635
rect -784 -5669 -750 -5661
rect -784 -5729 -750 -5707
rect -784 -5741 -750 -5729
rect -784 -5797 -750 -5779
rect -784 -5813 -750 -5797
rect -784 -5865 -750 -5851
rect -784 -5885 -750 -5865
rect -784 -5933 -750 -5923
rect -784 -5957 -750 -5933
rect -784 -6001 -750 -5995
rect -784 -6029 -750 -6001
rect -784 -6069 -750 -6067
rect -784 -6101 -750 -6069
rect -784 -6171 -750 -6139
rect -784 -6173 -750 -6171
rect -784 -6239 -750 -6211
rect -784 -6245 -750 -6239
rect -784 -6307 -750 -6283
rect -784 -6317 -750 -6307
rect -784 -6375 -750 -6355
rect -784 -6389 -750 -6375
rect -784 -6443 -750 -6427
rect -784 -6461 -750 -6443
rect -784 -6511 -750 -6499
rect -784 -6533 -750 -6511
rect -784 -6579 -750 -6571
rect -784 -6605 -750 -6579
rect -784 -6647 -750 -6643
rect -784 -6677 -750 -6647
rect -784 -6749 -750 -6715
rect -784 -6817 -750 -6787
rect -784 -6821 -750 -6817
rect -784 -6885 -750 -6859
rect -784 -6893 -750 -6885
rect -784 -6953 -750 -6931
rect -784 -6965 -750 -6953
rect -784 -7021 -750 -7003
rect -784 -7037 -750 -7021
rect -784 -7089 -750 -7075
rect -784 -7109 -750 -7089
rect -784 -7157 -750 -7147
rect -784 -7181 -750 -7157
rect -784 -7225 -750 -7219
rect -784 -7253 -750 -7225
rect -784 -7293 -750 -7291
rect -784 -7325 -750 -7293
rect -784 -7395 -750 -7363
rect -784 -7397 -750 -7395
rect -784 -7463 -750 -7435
rect -784 -7469 -750 -7463
rect -784 -7531 -750 -7507
rect -784 -7541 -750 -7531
rect -784 -7599 -750 -7579
rect -784 -7613 -750 -7599
rect -784 -7667 -750 -7651
rect -784 -7685 -750 -7667
rect -784 -7735 -750 -7723
rect -784 -7757 -750 -7735
rect -784 -7803 -750 -7795
rect -784 -7829 -750 -7803
rect -784 -7871 -750 -7867
rect -784 -7901 -750 -7871
rect -784 -7973 -750 -7939
rect -784 -8041 -750 -8011
rect -784 -8045 -750 -8041
rect -784 -8109 -750 -8083
rect -784 -8117 -750 -8109
rect -784 -8177 -750 -8155
rect -784 -8189 -750 -8177
rect -784 -8245 -750 -8227
rect -784 -8261 -750 -8245
rect -784 -8313 -750 -8299
rect -784 -8333 -750 -8313
rect -784 -8381 -750 -8371
rect -784 -8405 -750 -8381
rect -784 -8449 -750 -8443
rect -784 -8477 -750 -8449
rect -784 -8517 -750 -8515
rect -784 -8549 -750 -8517
rect -784 -8619 -750 -8587
rect -784 -8621 -750 -8619
rect -784 -8687 -750 -8659
rect -784 -8693 -750 -8687
rect -784 -8755 -750 -8731
rect -784 -8765 -750 -8755
rect -784 -8823 -750 -8803
rect -784 -8837 -750 -8823
rect -784 -8891 -750 -8875
rect -784 -8909 -750 -8891
rect -784 -8959 -750 -8947
rect -784 -8981 -750 -8959
rect -784 -9027 -750 -9019
rect -784 -9053 -750 -9027
rect -784 -9095 -750 -9091
rect -784 -9125 -750 -9095
rect -784 -9197 -750 -9163
rect -784 -9265 -750 -9235
rect -784 -9269 -750 -9265
rect -784 -9333 -750 -9307
rect -784 -9341 -750 -9333
rect -784 -9401 -750 -9379
rect -784 -9413 -750 -9401
rect -784 -9469 -750 -9451
rect -784 -9485 -750 -9469
rect -784 -9537 -750 -9523
rect -784 -9557 -750 -9537
rect -666 9537 -632 9557
rect -666 9523 -632 9537
rect -666 9469 -632 9485
rect -666 9451 -632 9469
rect -666 9401 -632 9413
rect -666 9379 -632 9401
rect -666 9333 -632 9341
rect -666 9307 -632 9333
rect -666 9265 -632 9269
rect -666 9235 -632 9265
rect -666 9163 -632 9197
rect -666 9095 -632 9125
rect -666 9091 -632 9095
rect -666 9027 -632 9053
rect -666 9019 -632 9027
rect -666 8959 -632 8981
rect -666 8947 -632 8959
rect -666 8891 -632 8909
rect -666 8875 -632 8891
rect -666 8823 -632 8837
rect -666 8803 -632 8823
rect -666 8755 -632 8765
rect -666 8731 -632 8755
rect -666 8687 -632 8693
rect -666 8659 -632 8687
rect -666 8619 -632 8621
rect -666 8587 -632 8619
rect -666 8517 -632 8549
rect -666 8515 -632 8517
rect -666 8449 -632 8477
rect -666 8443 -632 8449
rect -666 8381 -632 8405
rect -666 8371 -632 8381
rect -666 8313 -632 8333
rect -666 8299 -632 8313
rect -666 8245 -632 8261
rect -666 8227 -632 8245
rect -666 8177 -632 8189
rect -666 8155 -632 8177
rect -666 8109 -632 8117
rect -666 8083 -632 8109
rect -666 8041 -632 8045
rect -666 8011 -632 8041
rect -666 7939 -632 7973
rect -666 7871 -632 7901
rect -666 7867 -632 7871
rect -666 7803 -632 7829
rect -666 7795 -632 7803
rect -666 7735 -632 7757
rect -666 7723 -632 7735
rect -666 7667 -632 7685
rect -666 7651 -632 7667
rect -666 7599 -632 7613
rect -666 7579 -632 7599
rect -666 7531 -632 7541
rect -666 7507 -632 7531
rect -666 7463 -632 7469
rect -666 7435 -632 7463
rect -666 7395 -632 7397
rect -666 7363 -632 7395
rect -666 7293 -632 7325
rect -666 7291 -632 7293
rect -666 7225 -632 7253
rect -666 7219 -632 7225
rect -666 7157 -632 7181
rect -666 7147 -632 7157
rect -666 7089 -632 7109
rect -666 7075 -632 7089
rect -666 7021 -632 7037
rect -666 7003 -632 7021
rect -666 6953 -632 6965
rect -666 6931 -632 6953
rect -666 6885 -632 6893
rect -666 6859 -632 6885
rect -666 6817 -632 6821
rect -666 6787 -632 6817
rect -666 6715 -632 6749
rect -666 6647 -632 6677
rect -666 6643 -632 6647
rect -666 6579 -632 6605
rect -666 6571 -632 6579
rect -666 6511 -632 6533
rect -666 6499 -632 6511
rect -666 6443 -632 6461
rect -666 6427 -632 6443
rect -666 6375 -632 6389
rect -666 6355 -632 6375
rect -666 6307 -632 6317
rect -666 6283 -632 6307
rect -666 6239 -632 6245
rect -666 6211 -632 6239
rect -666 6171 -632 6173
rect -666 6139 -632 6171
rect -666 6069 -632 6101
rect -666 6067 -632 6069
rect -666 6001 -632 6029
rect -666 5995 -632 6001
rect -666 5933 -632 5957
rect -666 5923 -632 5933
rect -666 5865 -632 5885
rect -666 5851 -632 5865
rect -666 5797 -632 5813
rect -666 5779 -632 5797
rect -666 5729 -632 5741
rect -666 5707 -632 5729
rect -666 5661 -632 5669
rect -666 5635 -632 5661
rect -666 5593 -632 5597
rect -666 5563 -632 5593
rect -666 5491 -632 5525
rect -666 5423 -632 5453
rect -666 5419 -632 5423
rect -666 5355 -632 5381
rect -666 5347 -632 5355
rect -666 5287 -632 5309
rect -666 5275 -632 5287
rect -666 5219 -632 5237
rect -666 5203 -632 5219
rect -666 5151 -632 5165
rect -666 5131 -632 5151
rect -666 5083 -632 5093
rect -666 5059 -632 5083
rect -666 5015 -632 5021
rect -666 4987 -632 5015
rect -666 4947 -632 4949
rect -666 4915 -632 4947
rect -666 4845 -632 4877
rect -666 4843 -632 4845
rect -666 4777 -632 4805
rect -666 4771 -632 4777
rect -666 4709 -632 4733
rect -666 4699 -632 4709
rect -666 4641 -632 4661
rect -666 4627 -632 4641
rect -666 4573 -632 4589
rect -666 4555 -632 4573
rect -666 4505 -632 4517
rect -666 4483 -632 4505
rect -666 4437 -632 4445
rect -666 4411 -632 4437
rect -666 4369 -632 4373
rect -666 4339 -632 4369
rect -666 4267 -632 4301
rect -666 4199 -632 4229
rect -666 4195 -632 4199
rect -666 4131 -632 4157
rect -666 4123 -632 4131
rect -666 4063 -632 4085
rect -666 4051 -632 4063
rect -666 3995 -632 4013
rect -666 3979 -632 3995
rect -666 3927 -632 3941
rect -666 3907 -632 3927
rect -666 3859 -632 3869
rect -666 3835 -632 3859
rect -666 3791 -632 3797
rect -666 3763 -632 3791
rect -666 3723 -632 3725
rect -666 3691 -632 3723
rect -666 3621 -632 3653
rect -666 3619 -632 3621
rect -666 3553 -632 3581
rect -666 3547 -632 3553
rect -666 3485 -632 3509
rect -666 3475 -632 3485
rect -666 3417 -632 3437
rect -666 3403 -632 3417
rect -666 3349 -632 3365
rect -666 3331 -632 3349
rect -666 3281 -632 3293
rect -666 3259 -632 3281
rect -666 3213 -632 3221
rect -666 3187 -632 3213
rect -666 3145 -632 3149
rect -666 3115 -632 3145
rect -666 3043 -632 3077
rect -666 2975 -632 3005
rect -666 2971 -632 2975
rect -666 2907 -632 2933
rect -666 2899 -632 2907
rect -666 2839 -632 2861
rect -666 2827 -632 2839
rect -666 2771 -632 2789
rect -666 2755 -632 2771
rect -666 2703 -632 2717
rect -666 2683 -632 2703
rect -666 2635 -632 2645
rect -666 2611 -632 2635
rect -666 2567 -632 2573
rect -666 2539 -632 2567
rect -666 2499 -632 2501
rect -666 2467 -632 2499
rect -666 2397 -632 2429
rect -666 2395 -632 2397
rect -666 2329 -632 2357
rect -666 2323 -632 2329
rect -666 2261 -632 2285
rect -666 2251 -632 2261
rect -666 2193 -632 2213
rect -666 2179 -632 2193
rect -666 2125 -632 2141
rect -666 2107 -632 2125
rect -666 2057 -632 2069
rect -666 2035 -632 2057
rect -666 1989 -632 1997
rect -666 1963 -632 1989
rect -666 1921 -632 1925
rect -666 1891 -632 1921
rect -666 1819 -632 1853
rect -666 1751 -632 1781
rect -666 1747 -632 1751
rect -666 1683 -632 1709
rect -666 1675 -632 1683
rect -666 1615 -632 1637
rect -666 1603 -632 1615
rect -666 1547 -632 1565
rect -666 1531 -632 1547
rect -666 1479 -632 1493
rect -666 1459 -632 1479
rect -666 1411 -632 1421
rect -666 1387 -632 1411
rect -666 1343 -632 1349
rect -666 1315 -632 1343
rect -666 1275 -632 1277
rect -666 1243 -632 1275
rect -666 1173 -632 1205
rect -666 1171 -632 1173
rect -666 1105 -632 1133
rect -666 1099 -632 1105
rect -666 1037 -632 1061
rect -666 1027 -632 1037
rect -666 969 -632 989
rect -666 955 -632 969
rect -666 901 -632 917
rect -666 883 -632 901
rect -666 833 -632 845
rect -666 811 -632 833
rect -666 765 -632 773
rect -666 739 -632 765
rect -666 697 -632 701
rect -666 667 -632 697
rect -666 595 -632 629
rect -666 527 -632 557
rect -666 523 -632 527
rect -666 459 -632 485
rect -666 451 -632 459
rect -666 391 -632 413
rect -666 379 -632 391
rect -666 323 -632 341
rect -666 307 -632 323
rect -666 255 -632 269
rect -666 235 -632 255
rect -666 187 -632 197
rect -666 163 -632 187
rect -666 119 -632 125
rect -666 91 -632 119
rect -666 51 -632 53
rect -666 19 -632 51
rect -666 -51 -632 -19
rect -666 -53 -632 -51
rect -666 -119 -632 -91
rect -666 -125 -632 -119
rect -666 -187 -632 -163
rect -666 -197 -632 -187
rect -666 -255 -632 -235
rect -666 -269 -632 -255
rect -666 -323 -632 -307
rect -666 -341 -632 -323
rect -666 -391 -632 -379
rect -666 -413 -632 -391
rect -666 -459 -632 -451
rect -666 -485 -632 -459
rect -666 -527 -632 -523
rect -666 -557 -632 -527
rect -666 -629 -632 -595
rect -666 -697 -632 -667
rect -666 -701 -632 -697
rect -666 -765 -632 -739
rect -666 -773 -632 -765
rect -666 -833 -632 -811
rect -666 -845 -632 -833
rect -666 -901 -632 -883
rect -666 -917 -632 -901
rect -666 -969 -632 -955
rect -666 -989 -632 -969
rect -666 -1037 -632 -1027
rect -666 -1061 -632 -1037
rect -666 -1105 -632 -1099
rect -666 -1133 -632 -1105
rect -666 -1173 -632 -1171
rect -666 -1205 -632 -1173
rect -666 -1275 -632 -1243
rect -666 -1277 -632 -1275
rect -666 -1343 -632 -1315
rect -666 -1349 -632 -1343
rect -666 -1411 -632 -1387
rect -666 -1421 -632 -1411
rect -666 -1479 -632 -1459
rect -666 -1493 -632 -1479
rect -666 -1547 -632 -1531
rect -666 -1565 -632 -1547
rect -666 -1615 -632 -1603
rect -666 -1637 -632 -1615
rect -666 -1683 -632 -1675
rect -666 -1709 -632 -1683
rect -666 -1751 -632 -1747
rect -666 -1781 -632 -1751
rect -666 -1853 -632 -1819
rect -666 -1921 -632 -1891
rect -666 -1925 -632 -1921
rect -666 -1989 -632 -1963
rect -666 -1997 -632 -1989
rect -666 -2057 -632 -2035
rect -666 -2069 -632 -2057
rect -666 -2125 -632 -2107
rect -666 -2141 -632 -2125
rect -666 -2193 -632 -2179
rect -666 -2213 -632 -2193
rect -666 -2261 -632 -2251
rect -666 -2285 -632 -2261
rect -666 -2329 -632 -2323
rect -666 -2357 -632 -2329
rect -666 -2397 -632 -2395
rect -666 -2429 -632 -2397
rect -666 -2499 -632 -2467
rect -666 -2501 -632 -2499
rect -666 -2567 -632 -2539
rect -666 -2573 -632 -2567
rect -666 -2635 -632 -2611
rect -666 -2645 -632 -2635
rect -666 -2703 -632 -2683
rect -666 -2717 -632 -2703
rect -666 -2771 -632 -2755
rect -666 -2789 -632 -2771
rect -666 -2839 -632 -2827
rect -666 -2861 -632 -2839
rect -666 -2907 -632 -2899
rect -666 -2933 -632 -2907
rect -666 -2975 -632 -2971
rect -666 -3005 -632 -2975
rect -666 -3077 -632 -3043
rect -666 -3145 -632 -3115
rect -666 -3149 -632 -3145
rect -666 -3213 -632 -3187
rect -666 -3221 -632 -3213
rect -666 -3281 -632 -3259
rect -666 -3293 -632 -3281
rect -666 -3349 -632 -3331
rect -666 -3365 -632 -3349
rect -666 -3417 -632 -3403
rect -666 -3437 -632 -3417
rect -666 -3485 -632 -3475
rect -666 -3509 -632 -3485
rect -666 -3553 -632 -3547
rect -666 -3581 -632 -3553
rect -666 -3621 -632 -3619
rect -666 -3653 -632 -3621
rect -666 -3723 -632 -3691
rect -666 -3725 -632 -3723
rect -666 -3791 -632 -3763
rect -666 -3797 -632 -3791
rect -666 -3859 -632 -3835
rect -666 -3869 -632 -3859
rect -666 -3927 -632 -3907
rect -666 -3941 -632 -3927
rect -666 -3995 -632 -3979
rect -666 -4013 -632 -3995
rect -666 -4063 -632 -4051
rect -666 -4085 -632 -4063
rect -666 -4131 -632 -4123
rect -666 -4157 -632 -4131
rect -666 -4199 -632 -4195
rect -666 -4229 -632 -4199
rect -666 -4301 -632 -4267
rect -666 -4369 -632 -4339
rect -666 -4373 -632 -4369
rect -666 -4437 -632 -4411
rect -666 -4445 -632 -4437
rect -666 -4505 -632 -4483
rect -666 -4517 -632 -4505
rect -666 -4573 -632 -4555
rect -666 -4589 -632 -4573
rect -666 -4641 -632 -4627
rect -666 -4661 -632 -4641
rect -666 -4709 -632 -4699
rect -666 -4733 -632 -4709
rect -666 -4777 -632 -4771
rect -666 -4805 -632 -4777
rect -666 -4845 -632 -4843
rect -666 -4877 -632 -4845
rect -666 -4947 -632 -4915
rect -666 -4949 -632 -4947
rect -666 -5015 -632 -4987
rect -666 -5021 -632 -5015
rect -666 -5083 -632 -5059
rect -666 -5093 -632 -5083
rect -666 -5151 -632 -5131
rect -666 -5165 -632 -5151
rect -666 -5219 -632 -5203
rect -666 -5237 -632 -5219
rect -666 -5287 -632 -5275
rect -666 -5309 -632 -5287
rect -666 -5355 -632 -5347
rect -666 -5381 -632 -5355
rect -666 -5423 -632 -5419
rect -666 -5453 -632 -5423
rect -666 -5525 -632 -5491
rect -666 -5593 -632 -5563
rect -666 -5597 -632 -5593
rect -666 -5661 -632 -5635
rect -666 -5669 -632 -5661
rect -666 -5729 -632 -5707
rect -666 -5741 -632 -5729
rect -666 -5797 -632 -5779
rect -666 -5813 -632 -5797
rect -666 -5865 -632 -5851
rect -666 -5885 -632 -5865
rect -666 -5933 -632 -5923
rect -666 -5957 -632 -5933
rect -666 -6001 -632 -5995
rect -666 -6029 -632 -6001
rect -666 -6069 -632 -6067
rect -666 -6101 -632 -6069
rect -666 -6171 -632 -6139
rect -666 -6173 -632 -6171
rect -666 -6239 -632 -6211
rect -666 -6245 -632 -6239
rect -666 -6307 -632 -6283
rect -666 -6317 -632 -6307
rect -666 -6375 -632 -6355
rect -666 -6389 -632 -6375
rect -666 -6443 -632 -6427
rect -666 -6461 -632 -6443
rect -666 -6511 -632 -6499
rect -666 -6533 -632 -6511
rect -666 -6579 -632 -6571
rect -666 -6605 -632 -6579
rect -666 -6647 -632 -6643
rect -666 -6677 -632 -6647
rect -666 -6749 -632 -6715
rect -666 -6817 -632 -6787
rect -666 -6821 -632 -6817
rect -666 -6885 -632 -6859
rect -666 -6893 -632 -6885
rect -666 -6953 -632 -6931
rect -666 -6965 -632 -6953
rect -666 -7021 -632 -7003
rect -666 -7037 -632 -7021
rect -666 -7089 -632 -7075
rect -666 -7109 -632 -7089
rect -666 -7157 -632 -7147
rect -666 -7181 -632 -7157
rect -666 -7225 -632 -7219
rect -666 -7253 -632 -7225
rect -666 -7293 -632 -7291
rect -666 -7325 -632 -7293
rect -666 -7395 -632 -7363
rect -666 -7397 -632 -7395
rect -666 -7463 -632 -7435
rect -666 -7469 -632 -7463
rect -666 -7531 -632 -7507
rect -666 -7541 -632 -7531
rect -666 -7599 -632 -7579
rect -666 -7613 -632 -7599
rect -666 -7667 -632 -7651
rect -666 -7685 -632 -7667
rect -666 -7735 -632 -7723
rect -666 -7757 -632 -7735
rect -666 -7803 -632 -7795
rect -666 -7829 -632 -7803
rect -666 -7871 -632 -7867
rect -666 -7901 -632 -7871
rect -666 -7973 -632 -7939
rect -666 -8041 -632 -8011
rect -666 -8045 -632 -8041
rect -666 -8109 -632 -8083
rect -666 -8117 -632 -8109
rect -666 -8177 -632 -8155
rect -666 -8189 -632 -8177
rect -666 -8245 -632 -8227
rect -666 -8261 -632 -8245
rect -666 -8313 -632 -8299
rect -666 -8333 -632 -8313
rect -666 -8381 -632 -8371
rect -666 -8405 -632 -8381
rect -666 -8449 -632 -8443
rect -666 -8477 -632 -8449
rect -666 -8517 -632 -8515
rect -666 -8549 -632 -8517
rect -666 -8619 -632 -8587
rect -666 -8621 -632 -8619
rect -666 -8687 -632 -8659
rect -666 -8693 -632 -8687
rect -666 -8755 -632 -8731
rect -666 -8765 -632 -8755
rect -666 -8823 -632 -8803
rect -666 -8837 -632 -8823
rect -666 -8891 -632 -8875
rect -666 -8909 -632 -8891
rect -666 -8959 -632 -8947
rect -666 -8981 -632 -8959
rect -666 -9027 -632 -9019
rect -666 -9053 -632 -9027
rect -666 -9095 -632 -9091
rect -666 -9125 -632 -9095
rect -666 -9197 -632 -9163
rect -666 -9265 -632 -9235
rect -666 -9269 -632 -9265
rect -666 -9333 -632 -9307
rect -666 -9341 -632 -9333
rect -666 -9401 -632 -9379
rect -666 -9413 -632 -9401
rect -666 -9469 -632 -9451
rect -666 -9485 -632 -9469
rect -666 -9537 -632 -9523
rect -666 -9557 -632 -9537
rect -548 9537 -514 9557
rect -548 9523 -514 9537
rect -548 9469 -514 9485
rect -548 9451 -514 9469
rect -548 9401 -514 9413
rect -548 9379 -514 9401
rect -548 9333 -514 9341
rect -548 9307 -514 9333
rect -548 9265 -514 9269
rect -548 9235 -514 9265
rect -548 9163 -514 9197
rect -548 9095 -514 9125
rect -548 9091 -514 9095
rect -548 9027 -514 9053
rect -548 9019 -514 9027
rect -548 8959 -514 8981
rect -548 8947 -514 8959
rect -548 8891 -514 8909
rect -548 8875 -514 8891
rect -548 8823 -514 8837
rect -548 8803 -514 8823
rect -548 8755 -514 8765
rect -548 8731 -514 8755
rect -548 8687 -514 8693
rect -548 8659 -514 8687
rect -548 8619 -514 8621
rect -548 8587 -514 8619
rect -548 8517 -514 8549
rect -548 8515 -514 8517
rect -548 8449 -514 8477
rect -548 8443 -514 8449
rect -548 8381 -514 8405
rect -548 8371 -514 8381
rect -548 8313 -514 8333
rect -548 8299 -514 8313
rect -548 8245 -514 8261
rect -548 8227 -514 8245
rect -548 8177 -514 8189
rect -548 8155 -514 8177
rect -548 8109 -514 8117
rect -548 8083 -514 8109
rect -548 8041 -514 8045
rect -548 8011 -514 8041
rect -548 7939 -514 7973
rect -548 7871 -514 7901
rect -548 7867 -514 7871
rect -548 7803 -514 7829
rect -548 7795 -514 7803
rect -548 7735 -514 7757
rect -548 7723 -514 7735
rect -548 7667 -514 7685
rect -548 7651 -514 7667
rect -548 7599 -514 7613
rect -548 7579 -514 7599
rect -548 7531 -514 7541
rect -548 7507 -514 7531
rect -548 7463 -514 7469
rect -548 7435 -514 7463
rect -548 7395 -514 7397
rect -548 7363 -514 7395
rect -548 7293 -514 7325
rect -548 7291 -514 7293
rect -548 7225 -514 7253
rect -548 7219 -514 7225
rect -548 7157 -514 7181
rect -548 7147 -514 7157
rect -548 7089 -514 7109
rect -548 7075 -514 7089
rect -548 7021 -514 7037
rect -548 7003 -514 7021
rect -548 6953 -514 6965
rect -548 6931 -514 6953
rect -548 6885 -514 6893
rect -548 6859 -514 6885
rect -548 6817 -514 6821
rect -548 6787 -514 6817
rect -548 6715 -514 6749
rect -548 6647 -514 6677
rect -548 6643 -514 6647
rect -548 6579 -514 6605
rect -548 6571 -514 6579
rect -548 6511 -514 6533
rect -548 6499 -514 6511
rect -548 6443 -514 6461
rect -548 6427 -514 6443
rect -548 6375 -514 6389
rect -548 6355 -514 6375
rect -548 6307 -514 6317
rect -548 6283 -514 6307
rect -548 6239 -514 6245
rect -548 6211 -514 6239
rect -548 6171 -514 6173
rect -548 6139 -514 6171
rect -548 6069 -514 6101
rect -548 6067 -514 6069
rect -548 6001 -514 6029
rect -548 5995 -514 6001
rect -548 5933 -514 5957
rect -548 5923 -514 5933
rect -548 5865 -514 5885
rect -548 5851 -514 5865
rect -548 5797 -514 5813
rect -548 5779 -514 5797
rect -548 5729 -514 5741
rect -548 5707 -514 5729
rect -548 5661 -514 5669
rect -548 5635 -514 5661
rect -548 5593 -514 5597
rect -548 5563 -514 5593
rect -548 5491 -514 5525
rect -548 5423 -514 5453
rect -548 5419 -514 5423
rect -548 5355 -514 5381
rect -548 5347 -514 5355
rect -548 5287 -514 5309
rect -548 5275 -514 5287
rect -548 5219 -514 5237
rect -548 5203 -514 5219
rect -548 5151 -514 5165
rect -548 5131 -514 5151
rect -548 5083 -514 5093
rect -548 5059 -514 5083
rect -548 5015 -514 5021
rect -548 4987 -514 5015
rect -548 4947 -514 4949
rect -548 4915 -514 4947
rect -548 4845 -514 4877
rect -548 4843 -514 4845
rect -548 4777 -514 4805
rect -548 4771 -514 4777
rect -548 4709 -514 4733
rect -548 4699 -514 4709
rect -548 4641 -514 4661
rect -548 4627 -514 4641
rect -548 4573 -514 4589
rect -548 4555 -514 4573
rect -548 4505 -514 4517
rect -548 4483 -514 4505
rect -548 4437 -514 4445
rect -548 4411 -514 4437
rect -548 4369 -514 4373
rect -548 4339 -514 4369
rect -548 4267 -514 4301
rect -548 4199 -514 4229
rect -548 4195 -514 4199
rect -548 4131 -514 4157
rect -548 4123 -514 4131
rect -548 4063 -514 4085
rect -548 4051 -514 4063
rect -548 3995 -514 4013
rect -548 3979 -514 3995
rect -548 3927 -514 3941
rect -548 3907 -514 3927
rect -548 3859 -514 3869
rect -548 3835 -514 3859
rect -548 3791 -514 3797
rect -548 3763 -514 3791
rect -548 3723 -514 3725
rect -548 3691 -514 3723
rect -548 3621 -514 3653
rect -548 3619 -514 3621
rect -548 3553 -514 3581
rect -548 3547 -514 3553
rect -548 3485 -514 3509
rect -548 3475 -514 3485
rect -548 3417 -514 3437
rect -548 3403 -514 3417
rect -548 3349 -514 3365
rect -548 3331 -514 3349
rect -548 3281 -514 3293
rect -548 3259 -514 3281
rect -548 3213 -514 3221
rect -548 3187 -514 3213
rect -548 3145 -514 3149
rect -548 3115 -514 3145
rect -548 3043 -514 3077
rect -548 2975 -514 3005
rect -548 2971 -514 2975
rect -548 2907 -514 2933
rect -548 2899 -514 2907
rect -548 2839 -514 2861
rect -548 2827 -514 2839
rect -548 2771 -514 2789
rect -548 2755 -514 2771
rect -548 2703 -514 2717
rect -548 2683 -514 2703
rect -548 2635 -514 2645
rect -548 2611 -514 2635
rect -548 2567 -514 2573
rect -548 2539 -514 2567
rect -548 2499 -514 2501
rect -548 2467 -514 2499
rect -548 2397 -514 2429
rect -548 2395 -514 2397
rect -548 2329 -514 2357
rect -548 2323 -514 2329
rect -548 2261 -514 2285
rect -548 2251 -514 2261
rect -548 2193 -514 2213
rect -548 2179 -514 2193
rect -548 2125 -514 2141
rect -548 2107 -514 2125
rect -548 2057 -514 2069
rect -548 2035 -514 2057
rect -548 1989 -514 1997
rect -548 1963 -514 1989
rect -548 1921 -514 1925
rect -548 1891 -514 1921
rect -548 1819 -514 1853
rect -548 1751 -514 1781
rect -548 1747 -514 1751
rect -548 1683 -514 1709
rect -548 1675 -514 1683
rect -548 1615 -514 1637
rect -548 1603 -514 1615
rect -548 1547 -514 1565
rect -548 1531 -514 1547
rect -548 1479 -514 1493
rect -548 1459 -514 1479
rect -548 1411 -514 1421
rect -548 1387 -514 1411
rect -548 1343 -514 1349
rect -548 1315 -514 1343
rect -548 1275 -514 1277
rect -548 1243 -514 1275
rect -548 1173 -514 1205
rect -548 1171 -514 1173
rect -548 1105 -514 1133
rect -548 1099 -514 1105
rect -548 1037 -514 1061
rect -548 1027 -514 1037
rect -548 969 -514 989
rect -548 955 -514 969
rect -548 901 -514 917
rect -548 883 -514 901
rect -548 833 -514 845
rect -548 811 -514 833
rect -548 765 -514 773
rect -548 739 -514 765
rect -548 697 -514 701
rect -548 667 -514 697
rect -548 595 -514 629
rect -548 527 -514 557
rect -548 523 -514 527
rect -548 459 -514 485
rect -548 451 -514 459
rect -548 391 -514 413
rect -548 379 -514 391
rect -548 323 -514 341
rect -548 307 -514 323
rect -548 255 -514 269
rect -548 235 -514 255
rect -548 187 -514 197
rect -548 163 -514 187
rect -548 119 -514 125
rect -548 91 -514 119
rect -548 51 -514 53
rect -548 19 -514 51
rect -548 -51 -514 -19
rect -548 -53 -514 -51
rect -548 -119 -514 -91
rect -548 -125 -514 -119
rect -548 -187 -514 -163
rect -548 -197 -514 -187
rect -548 -255 -514 -235
rect -548 -269 -514 -255
rect -548 -323 -514 -307
rect -548 -341 -514 -323
rect -548 -391 -514 -379
rect -548 -413 -514 -391
rect -548 -459 -514 -451
rect -548 -485 -514 -459
rect -548 -527 -514 -523
rect -548 -557 -514 -527
rect -548 -629 -514 -595
rect -548 -697 -514 -667
rect -548 -701 -514 -697
rect -548 -765 -514 -739
rect -548 -773 -514 -765
rect -548 -833 -514 -811
rect -548 -845 -514 -833
rect -548 -901 -514 -883
rect -548 -917 -514 -901
rect -548 -969 -514 -955
rect -548 -989 -514 -969
rect -548 -1037 -514 -1027
rect -548 -1061 -514 -1037
rect -548 -1105 -514 -1099
rect -548 -1133 -514 -1105
rect -548 -1173 -514 -1171
rect -548 -1205 -514 -1173
rect -548 -1275 -514 -1243
rect -548 -1277 -514 -1275
rect -548 -1343 -514 -1315
rect -548 -1349 -514 -1343
rect -548 -1411 -514 -1387
rect -548 -1421 -514 -1411
rect -548 -1479 -514 -1459
rect -548 -1493 -514 -1479
rect -548 -1547 -514 -1531
rect -548 -1565 -514 -1547
rect -548 -1615 -514 -1603
rect -548 -1637 -514 -1615
rect -548 -1683 -514 -1675
rect -548 -1709 -514 -1683
rect -548 -1751 -514 -1747
rect -548 -1781 -514 -1751
rect -548 -1853 -514 -1819
rect -548 -1921 -514 -1891
rect -548 -1925 -514 -1921
rect -548 -1989 -514 -1963
rect -548 -1997 -514 -1989
rect -548 -2057 -514 -2035
rect -548 -2069 -514 -2057
rect -548 -2125 -514 -2107
rect -548 -2141 -514 -2125
rect -548 -2193 -514 -2179
rect -548 -2213 -514 -2193
rect -548 -2261 -514 -2251
rect -548 -2285 -514 -2261
rect -548 -2329 -514 -2323
rect -548 -2357 -514 -2329
rect -548 -2397 -514 -2395
rect -548 -2429 -514 -2397
rect -548 -2499 -514 -2467
rect -548 -2501 -514 -2499
rect -548 -2567 -514 -2539
rect -548 -2573 -514 -2567
rect -548 -2635 -514 -2611
rect -548 -2645 -514 -2635
rect -548 -2703 -514 -2683
rect -548 -2717 -514 -2703
rect -548 -2771 -514 -2755
rect -548 -2789 -514 -2771
rect -548 -2839 -514 -2827
rect -548 -2861 -514 -2839
rect -548 -2907 -514 -2899
rect -548 -2933 -514 -2907
rect -548 -2975 -514 -2971
rect -548 -3005 -514 -2975
rect -548 -3077 -514 -3043
rect -548 -3145 -514 -3115
rect -548 -3149 -514 -3145
rect -548 -3213 -514 -3187
rect -548 -3221 -514 -3213
rect -548 -3281 -514 -3259
rect -548 -3293 -514 -3281
rect -548 -3349 -514 -3331
rect -548 -3365 -514 -3349
rect -548 -3417 -514 -3403
rect -548 -3437 -514 -3417
rect -548 -3485 -514 -3475
rect -548 -3509 -514 -3485
rect -548 -3553 -514 -3547
rect -548 -3581 -514 -3553
rect -548 -3621 -514 -3619
rect -548 -3653 -514 -3621
rect -548 -3723 -514 -3691
rect -548 -3725 -514 -3723
rect -548 -3791 -514 -3763
rect -548 -3797 -514 -3791
rect -548 -3859 -514 -3835
rect -548 -3869 -514 -3859
rect -548 -3927 -514 -3907
rect -548 -3941 -514 -3927
rect -548 -3995 -514 -3979
rect -548 -4013 -514 -3995
rect -548 -4063 -514 -4051
rect -548 -4085 -514 -4063
rect -548 -4131 -514 -4123
rect -548 -4157 -514 -4131
rect -548 -4199 -514 -4195
rect -548 -4229 -514 -4199
rect -548 -4301 -514 -4267
rect -548 -4369 -514 -4339
rect -548 -4373 -514 -4369
rect -548 -4437 -514 -4411
rect -548 -4445 -514 -4437
rect -548 -4505 -514 -4483
rect -548 -4517 -514 -4505
rect -548 -4573 -514 -4555
rect -548 -4589 -514 -4573
rect -548 -4641 -514 -4627
rect -548 -4661 -514 -4641
rect -548 -4709 -514 -4699
rect -548 -4733 -514 -4709
rect -548 -4777 -514 -4771
rect -548 -4805 -514 -4777
rect -548 -4845 -514 -4843
rect -548 -4877 -514 -4845
rect -548 -4947 -514 -4915
rect -548 -4949 -514 -4947
rect -548 -5015 -514 -4987
rect -548 -5021 -514 -5015
rect -548 -5083 -514 -5059
rect -548 -5093 -514 -5083
rect -548 -5151 -514 -5131
rect -548 -5165 -514 -5151
rect -548 -5219 -514 -5203
rect -548 -5237 -514 -5219
rect -548 -5287 -514 -5275
rect -548 -5309 -514 -5287
rect -548 -5355 -514 -5347
rect -548 -5381 -514 -5355
rect -548 -5423 -514 -5419
rect -548 -5453 -514 -5423
rect -548 -5525 -514 -5491
rect -548 -5593 -514 -5563
rect -548 -5597 -514 -5593
rect -548 -5661 -514 -5635
rect -548 -5669 -514 -5661
rect -548 -5729 -514 -5707
rect -548 -5741 -514 -5729
rect -548 -5797 -514 -5779
rect -548 -5813 -514 -5797
rect -548 -5865 -514 -5851
rect -548 -5885 -514 -5865
rect -548 -5933 -514 -5923
rect -548 -5957 -514 -5933
rect -548 -6001 -514 -5995
rect -548 -6029 -514 -6001
rect -548 -6069 -514 -6067
rect -548 -6101 -514 -6069
rect -548 -6171 -514 -6139
rect -548 -6173 -514 -6171
rect -548 -6239 -514 -6211
rect -548 -6245 -514 -6239
rect -548 -6307 -514 -6283
rect -548 -6317 -514 -6307
rect -548 -6375 -514 -6355
rect -548 -6389 -514 -6375
rect -548 -6443 -514 -6427
rect -548 -6461 -514 -6443
rect -548 -6511 -514 -6499
rect -548 -6533 -514 -6511
rect -548 -6579 -514 -6571
rect -548 -6605 -514 -6579
rect -548 -6647 -514 -6643
rect -548 -6677 -514 -6647
rect -548 -6749 -514 -6715
rect -548 -6817 -514 -6787
rect -548 -6821 -514 -6817
rect -548 -6885 -514 -6859
rect -548 -6893 -514 -6885
rect -548 -6953 -514 -6931
rect -548 -6965 -514 -6953
rect -548 -7021 -514 -7003
rect -548 -7037 -514 -7021
rect -548 -7089 -514 -7075
rect -548 -7109 -514 -7089
rect -548 -7157 -514 -7147
rect -548 -7181 -514 -7157
rect -548 -7225 -514 -7219
rect -548 -7253 -514 -7225
rect -548 -7293 -514 -7291
rect -548 -7325 -514 -7293
rect -548 -7395 -514 -7363
rect -548 -7397 -514 -7395
rect -548 -7463 -514 -7435
rect -548 -7469 -514 -7463
rect -548 -7531 -514 -7507
rect -548 -7541 -514 -7531
rect -548 -7599 -514 -7579
rect -548 -7613 -514 -7599
rect -548 -7667 -514 -7651
rect -548 -7685 -514 -7667
rect -548 -7735 -514 -7723
rect -548 -7757 -514 -7735
rect -548 -7803 -514 -7795
rect -548 -7829 -514 -7803
rect -548 -7871 -514 -7867
rect -548 -7901 -514 -7871
rect -548 -7973 -514 -7939
rect -548 -8041 -514 -8011
rect -548 -8045 -514 -8041
rect -548 -8109 -514 -8083
rect -548 -8117 -514 -8109
rect -548 -8177 -514 -8155
rect -548 -8189 -514 -8177
rect -548 -8245 -514 -8227
rect -548 -8261 -514 -8245
rect -548 -8313 -514 -8299
rect -548 -8333 -514 -8313
rect -548 -8381 -514 -8371
rect -548 -8405 -514 -8381
rect -548 -8449 -514 -8443
rect -548 -8477 -514 -8449
rect -548 -8517 -514 -8515
rect -548 -8549 -514 -8517
rect -548 -8619 -514 -8587
rect -548 -8621 -514 -8619
rect -548 -8687 -514 -8659
rect -548 -8693 -514 -8687
rect -548 -8755 -514 -8731
rect -548 -8765 -514 -8755
rect -548 -8823 -514 -8803
rect -548 -8837 -514 -8823
rect -548 -8891 -514 -8875
rect -548 -8909 -514 -8891
rect -548 -8959 -514 -8947
rect -548 -8981 -514 -8959
rect -548 -9027 -514 -9019
rect -548 -9053 -514 -9027
rect -548 -9095 -514 -9091
rect -548 -9125 -514 -9095
rect -548 -9197 -514 -9163
rect -548 -9265 -514 -9235
rect -548 -9269 -514 -9265
rect -548 -9333 -514 -9307
rect -548 -9341 -514 -9333
rect -548 -9401 -514 -9379
rect -548 -9413 -514 -9401
rect -548 -9469 -514 -9451
rect -548 -9485 -514 -9469
rect -548 -9537 -514 -9523
rect -548 -9557 -514 -9537
rect -430 9537 -396 9557
rect -430 9523 -396 9537
rect -430 9469 -396 9485
rect -430 9451 -396 9469
rect -430 9401 -396 9413
rect -430 9379 -396 9401
rect -430 9333 -396 9341
rect -430 9307 -396 9333
rect -430 9265 -396 9269
rect -430 9235 -396 9265
rect -430 9163 -396 9197
rect -430 9095 -396 9125
rect -430 9091 -396 9095
rect -430 9027 -396 9053
rect -430 9019 -396 9027
rect -430 8959 -396 8981
rect -430 8947 -396 8959
rect -430 8891 -396 8909
rect -430 8875 -396 8891
rect -430 8823 -396 8837
rect -430 8803 -396 8823
rect -430 8755 -396 8765
rect -430 8731 -396 8755
rect -430 8687 -396 8693
rect -430 8659 -396 8687
rect -430 8619 -396 8621
rect -430 8587 -396 8619
rect -430 8517 -396 8549
rect -430 8515 -396 8517
rect -430 8449 -396 8477
rect -430 8443 -396 8449
rect -430 8381 -396 8405
rect -430 8371 -396 8381
rect -430 8313 -396 8333
rect -430 8299 -396 8313
rect -430 8245 -396 8261
rect -430 8227 -396 8245
rect -430 8177 -396 8189
rect -430 8155 -396 8177
rect -430 8109 -396 8117
rect -430 8083 -396 8109
rect -430 8041 -396 8045
rect -430 8011 -396 8041
rect -430 7939 -396 7973
rect -430 7871 -396 7901
rect -430 7867 -396 7871
rect -430 7803 -396 7829
rect -430 7795 -396 7803
rect -430 7735 -396 7757
rect -430 7723 -396 7735
rect -430 7667 -396 7685
rect -430 7651 -396 7667
rect -430 7599 -396 7613
rect -430 7579 -396 7599
rect -430 7531 -396 7541
rect -430 7507 -396 7531
rect -430 7463 -396 7469
rect -430 7435 -396 7463
rect -430 7395 -396 7397
rect -430 7363 -396 7395
rect -430 7293 -396 7325
rect -430 7291 -396 7293
rect -430 7225 -396 7253
rect -430 7219 -396 7225
rect -430 7157 -396 7181
rect -430 7147 -396 7157
rect -430 7089 -396 7109
rect -430 7075 -396 7089
rect -430 7021 -396 7037
rect -430 7003 -396 7021
rect -430 6953 -396 6965
rect -430 6931 -396 6953
rect -430 6885 -396 6893
rect -430 6859 -396 6885
rect -430 6817 -396 6821
rect -430 6787 -396 6817
rect -430 6715 -396 6749
rect -430 6647 -396 6677
rect -430 6643 -396 6647
rect -430 6579 -396 6605
rect -430 6571 -396 6579
rect -430 6511 -396 6533
rect -430 6499 -396 6511
rect -430 6443 -396 6461
rect -430 6427 -396 6443
rect -430 6375 -396 6389
rect -430 6355 -396 6375
rect -430 6307 -396 6317
rect -430 6283 -396 6307
rect -430 6239 -396 6245
rect -430 6211 -396 6239
rect -430 6171 -396 6173
rect -430 6139 -396 6171
rect -430 6069 -396 6101
rect -430 6067 -396 6069
rect -430 6001 -396 6029
rect -430 5995 -396 6001
rect -430 5933 -396 5957
rect -430 5923 -396 5933
rect -430 5865 -396 5885
rect -430 5851 -396 5865
rect -430 5797 -396 5813
rect -430 5779 -396 5797
rect -430 5729 -396 5741
rect -430 5707 -396 5729
rect -430 5661 -396 5669
rect -430 5635 -396 5661
rect -430 5593 -396 5597
rect -430 5563 -396 5593
rect -430 5491 -396 5525
rect -430 5423 -396 5453
rect -430 5419 -396 5423
rect -430 5355 -396 5381
rect -430 5347 -396 5355
rect -430 5287 -396 5309
rect -430 5275 -396 5287
rect -430 5219 -396 5237
rect -430 5203 -396 5219
rect -430 5151 -396 5165
rect -430 5131 -396 5151
rect -430 5083 -396 5093
rect -430 5059 -396 5083
rect -430 5015 -396 5021
rect -430 4987 -396 5015
rect -430 4947 -396 4949
rect -430 4915 -396 4947
rect -430 4845 -396 4877
rect -430 4843 -396 4845
rect -430 4777 -396 4805
rect -430 4771 -396 4777
rect -430 4709 -396 4733
rect -430 4699 -396 4709
rect -430 4641 -396 4661
rect -430 4627 -396 4641
rect -430 4573 -396 4589
rect -430 4555 -396 4573
rect -430 4505 -396 4517
rect -430 4483 -396 4505
rect -430 4437 -396 4445
rect -430 4411 -396 4437
rect -430 4369 -396 4373
rect -430 4339 -396 4369
rect -430 4267 -396 4301
rect -430 4199 -396 4229
rect -430 4195 -396 4199
rect -430 4131 -396 4157
rect -430 4123 -396 4131
rect -430 4063 -396 4085
rect -430 4051 -396 4063
rect -430 3995 -396 4013
rect -430 3979 -396 3995
rect -430 3927 -396 3941
rect -430 3907 -396 3927
rect -430 3859 -396 3869
rect -430 3835 -396 3859
rect -430 3791 -396 3797
rect -430 3763 -396 3791
rect -430 3723 -396 3725
rect -430 3691 -396 3723
rect -430 3621 -396 3653
rect -430 3619 -396 3621
rect -430 3553 -396 3581
rect -430 3547 -396 3553
rect -430 3485 -396 3509
rect -430 3475 -396 3485
rect -430 3417 -396 3437
rect -430 3403 -396 3417
rect -430 3349 -396 3365
rect -430 3331 -396 3349
rect -430 3281 -396 3293
rect -430 3259 -396 3281
rect -430 3213 -396 3221
rect -430 3187 -396 3213
rect -430 3145 -396 3149
rect -430 3115 -396 3145
rect -430 3043 -396 3077
rect -430 2975 -396 3005
rect -430 2971 -396 2975
rect -430 2907 -396 2933
rect -430 2899 -396 2907
rect -430 2839 -396 2861
rect -430 2827 -396 2839
rect -430 2771 -396 2789
rect -430 2755 -396 2771
rect -430 2703 -396 2717
rect -430 2683 -396 2703
rect -430 2635 -396 2645
rect -430 2611 -396 2635
rect -430 2567 -396 2573
rect -430 2539 -396 2567
rect -430 2499 -396 2501
rect -430 2467 -396 2499
rect -430 2397 -396 2429
rect -430 2395 -396 2397
rect -430 2329 -396 2357
rect -430 2323 -396 2329
rect -430 2261 -396 2285
rect -430 2251 -396 2261
rect -430 2193 -396 2213
rect -430 2179 -396 2193
rect -430 2125 -396 2141
rect -430 2107 -396 2125
rect -430 2057 -396 2069
rect -430 2035 -396 2057
rect -430 1989 -396 1997
rect -430 1963 -396 1989
rect -430 1921 -396 1925
rect -430 1891 -396 1921
rect -430 1819 -396 1853
rect -430 1751 -396 1781
rect -430 1747 -396 1751
rect -430 1683 -396 1709
rect -430 1675 -396 1683
rect -430 1615 -396 1637
rect -430 1603 -396 1615
rect -430 1547 -396 1565
rect -430 1531 -396 1547
rect -430 1479 -396 1493
rect -430 1459 -396 1479
rect -430 1411 -396 1421
rect -430 1387 -396 1411
rect -430 1343 -396 1349
rect -430 1315 -396 1343
rect -430 1275 -396 1277
rect -430 1243 -396 1275
rect -430 1173 -396 1205
rect -430 1171 -396 1173
rect -430 1105 -396 1133
rect -430 1099 -396 1105
rect -430 1037 -396 1061
rect -430 1027 -396 1037
rect -430 969 -396 989
rect -430 955 -396 969
rect -430 901 -396 917
rect -430 883 -396 901
rect -430 833 -396 845
rect -430 811 -396 833
rect -430 765 -396 773
rect -430 739 -396 765
rect -430 697 -396 701
rect -430 667 -396 697
rect -430 595 -396 629
rect -430 527 -396 557
rect -430 523 -396 527
rect -430 459 -396 485
rect -430 451 -396 459
rect -430 391 -396 413
rect -430 379 -396 391
rect -430 323 -396 341
rect -430 307 -396 323
rect -430 255 -396 269
rect -430 235 -396 255
rect -430 187 -396 197
rect -430 163 -396 187
rect -430 119 -396 125
rect -430 91 -396 119
rect -430 51 -396 53
rect -430 19 -396 51
rect -430 -51 -396 -19
rect -430 -53 -396 -51
rect -430 -119 -396 -91
rect -430 -125 -396 -119
rect -430 -187 -396 -163
rect -430 -197 -396 -187
rect -430 -255 -396 -235
rect -430 -269 -396 -255
rect -430 -323 -396 -307
rect -430 -341 -396 -323
rect -430 -391 -396 -379
rect -430 -413 -396 -391
rect -430 -459 -396 -451
rect -430 -485 -396 -459
rect -430 -527 -396 -523
rect -430 -557 -396 -527
rect -430 -629 -396 -595
rect -430 -697 -396 -667
rect -430 -701 -396 -697
rect -430 -765 -396 -739
rect -430 -773 -396 -765
rect -430 -833 -396 -811
rect -430 -845 -396 -833
rect -430 -901 -396 -883
rect -430 -917 -396 -901
rect -430 -969 -396 -955
rect -430 -989 -396 -969
rect -430 -1037 -396 -1027
rect -430 -1061 -396 -1037
rect -430 -1105 -396 -1099
rect -430 -1133 -396 -1105
rect -430 -1173 -396 -1171
rect -430 -1205 -396 -1173
rect -430 -1275 -396 -1243
rect -430 -1277 -396 -1275
rect -430 -1343 -396 -1315
rect -430 -1349 -396 -1343
rect -430 -1411 -396 -1387
rect -430 -1421 -396 -1411
rect -430 -1479 -396 -1459
rect -430 -1493 -396 -1479
rect -430 -1547 -396 -1531
rect -430 -1565 -396 -1547
rect -430 -1615 -396 -1603
rect -430 -1637 -396 -1615
rect -430 -1683 -396 -1675
rect -430 -1709 -396 -1683
rect -430 -1751 -396 -1747
rect -430 -1781 -396 -1751
rect -430 -1853 -396 -1819
rect -430 -1921 -396 -1891
rect -430 -1925 -396 -1921
rect -430 -1989 -396 -1963
rect -430 -1997 -396 -1989
rect -430 -2057 -396 -2035
rect -430 -2069 -396 -2057
rect -430 -2125 -396 -2107
rect -430 -2141 -396 -2125
rect -430 -2193 -396 -2179
rect -430 -2213 -396 -2193
rect -430 -2261 -396 -2251
rect -430 -2285 -396 -2261
rect -430 -2329 -396 -2323
rect -430 -2357 -396 -2329
rect -430 -2397 -396 -2395
rect -430 -2429 -396 -2397
rect -430 -2499 -396 -2467
rect -430 -2501 -396 -2499
rect -430 -2567 -396 -2539
rect -430 -2573 -396 -2567
rect -430 -2635 -396 -2611
rect -430 -2645 -396 -2635
rect -430 -2703 -396 -2683
rect -430 -2717 -396 -2703
rect -430 -2771 -396 -2755
rect -430 -2789 -396 -2771
rect -430 -2839 -396 -2827
rect -430 -2861 -396 -2839
rect -430 -2907 -396 -2899
rect -430 -2933 -396 -2907
rect -430 -2975 -396 -2971
rect -430 -3005 -396 -2975
rect -430 -3077 -396 -3043
rect -430 -3145 -396 -3115
rect -430 -3149 -396 -3145
rect -430 -3213 -396 -3187
rect -430 -3221 -396 -3213
rect -430 -3281 -396 -3259
rect -430 -3293 -396 -3281
rect -430 -3349 -396 -3331
rect -430 -3365 -396 -3349
rect -430 -3417 -396 -3403
rect -430 -3437 -396 -3417
rect -430 -3485 -396 -3475
rect -430 -3509 -396 -3485
rect -430 -3553 -396 -3547
rect -430 -3581 -396 -3553
rect -430 -3621 -396 -3619
rect -430 -3653 -396 -3621
rect -430 -3723 -396 -3691
rect -430 -3725 -396 -3723
rect -430 -3791 -396 -3763
rect -430 -3797 -396 -3791
rect -430 -3859 -396 -3835
rect -430 -3869 -396 -3859
rect -430 -3927 -396 -3907
rect -430 -3941 -396 -3927
rect -430 -3995 -396 -3979
rect -430 -4013 -396 -3995
rect -430 -4063 -396 -4051
rect -430 -4085 -396 -4063
rect -430 -4131 -396 -4123
rect -430 -4157 -396 -4131
rect -430 -4199 -396 -4195
rect -430 -4229 -396 -4199
rect -430 -4301 -396 -4267
rect -430 -4369 -396 -4339
rect -430 -4373 -396 -4369
rect -430 -4437 -396 -4411
rect -430 -4445 -396 -4437
rect -430 -4505 -396 -4483
rect -430 -4517 -396 -4505
rect -430 -4573 -396 -4555
rect -430 -4589 -396 -4573
rect -430 -4641 -396 -4627
rect -430 -4661 -396 -4641
rect -430 -4709 -396 -4699
rect -430 -4733 -396 -4709
rect -430 -4777 -396 -4771
rect -430 -4805 -396 -4777
rect -430 -4845 -396 -4843
rect -430 -4877 -396 -4845
rect -430 -4947 -396 -4915
rect -430 -4949 -396 -4947
rect -430 -5015 -396 -4987
rect -430 -5021 -396 -5015
rect -430 -5083 -396 -5059
rect -430 -5093 -396 -5083
rect -430 -5151 -396 -5131
rect -430 -5165 -396 -5151
rect -430 -5219 -396 -5203
rect -430 -5237 -396 -5219
rect -430 -5287 -396 -5275
rect -430 -5309 -396 -5287
rect -430 -5355 -396 -5347
rect -430 -5381 -396 -5355
rect -430 -5423 -396 -5419
rect -430 -5453 -396 -5423
rect -430 -5525 -396 -5491
rect -430 -5593 -396 -5563
rect -430 -5597 -396 -5593
rect -430 -5661 -396 -5635
rect -430 -5669 -396 -5661
rect -430 -5729 -396 -5707
rect -430 -5741 -396 -5729
rect -430 -5797 -396 -5779
rect -430 -5813 -396 -5797
rect -430 -5865 -396 -5851
rect -430 -5885 -396 -5865
rect -430 -5933 -396 -5923
rect -430 -5957 -396 -5933
rect -430 -6001 -396 -5995
rect -430 -6029 -396 -6001
rect -430 -6069 -396 -6067
rect -430 -6101 -396 -6069
rect -430 -6171 -396 -6139
rect -430 -6173 -396 -6171
rect -430 -6239 -396 -6211
rect -430 -6245 -396 -6239
rect -430 -6307 -396 -6283
rect -430 -6317 -396 -6307
rect -430 -6375 -396 -6355
rect -430 -6389 -396 -6375
rect -430 -6443 -396 -6427
rect -430 -6461 -396 -6443
rect -430 -6511 -396 -6499
rect -430 -6533 -396 -6511
rect -430 -6579 -396 -6571
rect -430 -6605 -396 -6579
rect -430 -6647 -396 -6643
rect -430 -6677 -396 -6647
rect -430 -6749 -396 -6715
rect -430 -6817 -396 -6787
rect -430 -6821 -396 -6817
rect -430 -6885 -396 -6859
rect -430 -6893 -396 -6885
rect -430 -6953 -396 -6931
rect -430 -6965 -396 -6953
rect -430 -7021 -396 -7003
rect -430 -7037 -396 -7021
rect -430 -7089 -396 -7075
rect -430 -7109 -396 -7089
rect -430 -7157 -396 -7147
rect -430 -7181 -396 -7157
rect -430 -7225 -396 -7219
rect -430 -7253 -396 -7225
rect -430 -7293 -396 -7291
rect -430 -7325 -396 -7293
rect -430 -7395 -396 -7363
rect -430 -7397 -396 -7395
rect -430 -7463 -396 -7435
rect -430 -7469 -396 -7463
rect -430 -7531 -396 -7507
rect -430 -7541 -396 -7531
rect -430 -7599 -396 -7579
rect -430 -7613 -396 -7599
rect -430 -7667 -396 -7651
rect -430 -7685 -396 -7667
rect -430 -7735 -396 -7723
rect -430 -7757 -396 -7735
rect -430 -7803 -396 -7795
rect -430 -7829 -396 -7803
rect -430 -7871 -396 -7867
rect -430 -7901 -396 -7871
rect -430 -7973 -396 -7939
rect -430 -8041 -396 -8011
rect -430 -8045 -396 -8041
rect -430 -8109 -396 -8083
rect -430 -8117 -396 -8109
rect -430 -8177 -396 -8155
rect -430 -8189 -396 -8177
rect -430 -8245 -396 -8227
rect -430 -8261 -396 -8245
rect -430 -8313 -396 -8299
rect -430 -8333 -396 -8313
rect -430 -8381 -396 -8371
rect -430 -8405 -396 -8381
rect -430 -8449 -396 -8443
rect -430 -8477 -396 -8449
rect -430 -8517 -396 -8515
rect -430 -8549 -396 -8517
rect -430 -8619 -396 -8587
rect -430 -8621 -396 -8619
rect -430 -8687 -396 -8659
rect -430 -8693 -396 -8687
rect -430 -8755 -396 -8731
rect -430 -8765 -396 -8755
rect -430 -8823 -396 -8803
rect -430 -8837 -396 -8823
rect -430 -8891 -396 -8875
rect -430 -8909 -396 -8891
rect -430 -8959 -396 -8947
rect -430 -8981 -396 -8959
rect -430 -9027 -396 -9019
rect -430 -9053 -396 -9027
rect -430 -9095 -396 -9091
rect -430 -9125 -396 -9095
rect -430 -9197 -396 -9163
rect -430 -9265 -396 -9235
rect -430 -9269 -396 -9265
rect -430 -9333 -396 -9307
rect -430 -9341 -396 -9333
rect -430 -9401 -396 -9379
rect -430 -9413 -396 -9401
rect -430 -9469 -396 -9451
rect -430 -9485 -396 -9469
rect -430 -9537 -396 -9523
rect -430 -9557 -396 -9537
rect -312 9537 -278 9557
rect -312 9523 -278 9537
rect -312 9469 -278 9485
rect -312 9451 -278 9469
rect -312 9401 -278 9413
rect -312 9379 -278 9401
rect -312 9333 -278 9341
rect -312 9307 -278 9333
rect -312 9265 -278 9269
rect -312 9235 -278 9265
rect -312 9163 -278 9197
rect -312 9095 -278 9125
rect -312 9091 -278 9095
rect -312 9027 -278 9053
rect -312 9019 -278 9027
rect -312 8959 -278 8981
rect -312 8947 -278 8959
rect -312 8891 -278 8909
rect -312 8875 -278 8891
rect -312 8823 -278 8837
rect -312 8803 -278 8823
rect -312 8755 -278 8765
rect -312 8731 -278 8755
rect -312 8687 -278 8693
rect -312 8659 -278 8687
rect -312 8619 -278 8621
rect -312 8587 -278 8619
rect -312 8517 -278 8549
rect -312 8515 -278 8517
rect -312 8449 -278 8477
rect -312 8443 -278 8449
rect -312 8381 -278 8405
rect -312 8371 -278 8381
rect -312 8313 -278 8333
rect -312 8299 -278 8313
rect -312 8245 -278 8261
rect -312 8227 -278 8245
rect -312 8177 -278 8189
rect -312 8155 -278 8177
rect -312 8109 -278 8117
rect -312 8083 -278 8109
rect -312 8041 -278 8045
rect -312 8011 -278 8041
rect -312 7939 -278 7973
rect -312 7871 -278 7901
rect -312 7867 -278 7871
rect -312 7803 -278 7829
rect -312 7795 -278 7803
rect -312 7735 -278 7757
rect -312 7723 -278 7735
rect -312 7667 -278 7685
rect -312 7651 -278 7667
rect -312 7599 -278 7613
rect -312 7579 -278 7599
rect -312 7531 -278 7541
rect -312 7507 -278 7531
rect -312 7463 -278 7469
rect -312 7435 -278 7463
rect -312 7395 -278 7397
rect -312 7363 -278 7395
rect -312 7293 -278 7325
rect -312 7291 -278 7293
rect -312 7225 -278 7253
rect -312 7219 -278 7225
rect -312 7157 -278 7181
rect -312 7147 -278 7157
rect -312 7089 -278 7109
rect -312 7075 -278 7089
rect -312 7021 -278 7037
rect -312 7003 -278 7021
rect -312 6953 -278 6965
rect -312 6931 -278 6953
rect -312 6885 -278 6893
rect -312 6859 -278 6885
rect -312 6817 -278 6821
rect -312 6787 -278 6817
rect -312 6715 -278 6749
rect -312 6647 -278 6677
rect -312 6643 -278 6647
rect -312 6579 -278 6605
rect -312 6571 -278 6579
rect -312 6511 -278 6533
rect -312 6499 -278 6511
rect -312 6443 -278 6461
rect -312 6427 -278 6443
rect -312 6375 -278 6389
rect -312 6355 -278 6375
rect -312 6307 -278 6317
rect -312 6283 -278 6307
rect -312 6239 -278 6245
rect -312 6211 -278 6239
rect -312 6171 -278 6173
rect -312 6139 -278 6171
rect -312 6069 -278 6101
rect -312 6067 -278 6069
rect -312 6001 -278 6029
rect -312 5995 -278 6001
rect -312 5933 -278 5957
rect -312 5923 -278 5933
rect -312 5865 -278 5885
rect -312 5851 -278 5865
rect -312 5797 -278 5813
rect -312 5779 -278 5797
rect -312 5729 -278 5741
rect -312 5707 -278 5729
rect -312 5661 -278 5669
rect -312 5635 -278 5661
rect -312 5593 -278 5597
rect -312 5563 -278 5593
rect -312 5491 -278 5525
rect -312 5423 -278 5453
rect -312 5419 -278 5423
rect -312 5355 -278 5381
rect -312 5347 -278 5355
rect -312 5287 -278 5309
rect -312 5275 -278 5287
rect -312 5219 -278 5237
rect -312 5203 -278 5219
rect -312 5151 -278 5165
rect -312 5131 -278 5151
rect -312 5083 -278 5093
rect -312 5059 -278 5083
rect -312 5015 -278 5021
rect -312 4987 -278 5015
rect -312 4947 -278 4949
rect -312 4915 -278 4947
rect -312 4845 -278 4877
rect -312 4843 -278 4845
rect -312 4777 -278 4805
rect -312 4771 -278 4777
rect -312 4709 -278 4733
rect -312 4699 -278 4709
rect -312 4641 -278 4661
rect -312 4627 -278 4641
rect -312 4573 -278 4589
rect -312 4555 -278 4573
rect -312 4505 -278 4517
rect -312 4483 -278 4505
rect -312 4437 -278 4445
rect -312 4411 -278 4437
rect -312 4369 -278 4373
rect -312 4339 -278 4369
rect -312 4267 -278 4301
rect -312 4199 -278 4229
rect -312 4195 -278 4199
rect -312 4131 -278 4157
rect -312 4123 -278 4131
rect -312 4063 -278 4085
rect -312 4051 -278 4063
rect -312 3995 -278 4013
rect -312 3979 -278 3995
rect -312 3927 -278 3941
rect -312 3907 -278 3927
rect -312 3859 -278 3869
rect -312 3835 -278 3859
rect -312 3791 -278 3797
rect -312 3763 -278 3791
rect -312 3723 -278 3725
rect -312 3691 -278 3723
rect -312 3621 -278 3653
rect -312 3619 -278 3621
rect -312 3553 -278 3581
rect -312 3547 -278 3553
rect -312 3485 -278 3509
rect -312 3475 -278 3485
rect -312 3417 -278 3437
rect -312 3403 -278 3417
rect -312 3349 -278 3365
rect -312 3331 -278 3349
rect -312 3281 -278 3293
rect -312 3259 -278 3281
rect -312 3213 -278 3221
rect -312 3187 -278 3213
rect -312 3145 -278 3149
rect -312 3115 -278 3145
rect -312 3043 -278 3077
rect -312 2975 -278 3005
rect -312 2971 -278 2975
rect -312 2907 -278 2933
rect -312 2899 -278 2907
rect -312 2839 -278 2861
rect -312 2827 -278 2839
rect -312 2771 -278 2789
rect -312 2755 -278 2771
rect -312 2703 -278 2717
rect -312 2683 -278 2703
rect -312 2635 -278 2645
rect -312 2611 -278 2635
rect -312 2567 -278 2573
rect -312 2539 -278 2567
rect -312 2499 -278 2501
rect -312 2467 -278 2499
rect -312 2397 -278 2429
rect -312 2395 -278 2397
rect -312 2329 -278 2357
rect -312 2323 -278 2329
rect -312 2261 -278 2285
rect -312 2251 -278 2261
rect -312 2193 -278 2213
rect -312 2179 -278 2193
rect -312 2125 -278 2141
rect -312 2107 -278 2125
rect -312 2057 -278 2069
rect -312 2035 -278 2057
rect -312 1989 -278 1997
rect -312 1963 -278 1989
rect -312 1921 -278 1925
rect -312 1891 -278 1921
rect -312 1819 -278 1853
rect -312 1751 -278 1781
rect -312 1747 -278 1751
rect -312 1683 -278 1709
rect -312 1675 -278 1683
rect -312 1615 -278 1637
rect -312 1603 -278 1615
rect -312 1547 -278 1565
rect -312 1531 -278 1547
rect -312 1479 -278 1493
rect -312 1459 -278 1479
rect -312 1411 -278 1421
rect -312 1387 -278 1411
rect -312 1343 -278 1349
rect -312 1315 -278 1343
rect -312 1275 -278 1277
rect -312 1243 -278 1275
rect -312 1173 -278 1205
rect -312 1171 -278 1173
rect -312 1105 -278 1133
rect -312 1099 -278 1105
rect -312 1037 -278 1061
rect -312 1027 -278 1037
rect -312 969 -278 989
rect -312 955 -278 969
rect -312 901 -278 917
rect -312 883 -278 901
rect -312 833 -278 845
rect -312 811 -278 833
rect -312 765 -278 773
rect -312 739 -278 765
rect -312 697 -278 701
rect -312 667 -278 697
rect -312 595 -278 629
rect -312 527 -278 557
rect -312 523 -278 527
rect -312 459 -278 485
rect -312 451 -278 459
rect -312 391 -278 413
rect -312 379 -278 391
rect -312 323 -278 341
rect -312 307 -278 323
rect -312 255 -278 269
rect -312 235 -278 255
rect -312 187 -278 197
rect -312 163 -278 187
rect -312 119 -278 125
rect -312 91 -278 119
rect -312 51 -278 53
rect -312 19 -278 51
rect -312 -51 -278 -19
rect -312 -53 -278 -51
rect -312 -119 -278 -91
rect -312 -125 -278 -119
rect -312 -187 -278 -163
rect -312 -197 -278 -187
rect -312 -255 -278 -235
rect -312 -269 -278 -255
rect -312 -323 -278 -307
rect -312 -341 -278 -323
rect -312 -391 -278 -379
rect -312 -413 -278 -391
rect -312 -459 -278 -451
rect -312 -485 -278 -459
rect -312 -527 -278 -523
rect -312 -557 -278 -527
rect -312 -629 -278 -595
rect -312 -697 -278 -667
rect -312 -701 -278 -697
rect -312 -765 -278 -739
rect -312 -773 -278 -765
rect -312 -833 -278 -811
rect -312 -845 -278 -833
rect -312 -901 -278 -883
rect -312 -917 -278 -901
rect -312 -969 -278 -955
rect -312 -989 -278 -969
rect -312 -1037 -278 -1027
rect -312 -1061 -278 -1037
rect -312 -1105 -278 -1099
rect -312 -1133 -278 -1105
rect -312 -1173 -278 -1171
rect -312 -1205 -278 -1173
rect -312 -1275 -278 -1243
rect -312 -1277 -278 -1275
rect -312 -1343 -278 -1315
rect -312 -1349 -278 -1343
rect -312 -1411 -278 -1387
rect -312 -1421 -278 -1411
rect -312 -1479 -278 -1459
rect -312 -1493 -278 -1479
rect -312 -1547 -278 -1531
rect -312 -1565 -278 -1547
rect -312 -1615 -278 -1603
rect -312 -1637 -278 -1615
rect -312 -1683 -278 -1675
rect -312 -1709 -278 -1683
rect -312 -1751 -278 -1747
rect -312 -1781 -278 -1751
rect -312 -1853 -278 -1819
rect -312 -1921 -278 -1891
rect -312 -1925 -278 -1921
rect -312 -1989 -278 -1963
rect -312 -1997 -278 -1989
rect -312 -2057 -278 -2035
rect -312 -2069 -278 -2057
rect -312 -2125 -278 -2107
rect -312 -2141 -278 -2125
rect -312 -2193 -278 -2179
rect -312 -2213 -278 -2193
rect -312 -2261 -278 -2251
rect -312 -2285 -278 -2261
rect -312 -2329 -278 -2323
rect -312 -2357 -278 -2329
rect -312 -2397 -278 -2395
rect -312 -2429 -278 -2397
rect -312 -2499 -278 -2467
rect -312 -2501 -278 -2499
rect -312 -2567 -278 -2539
rect -312 -2573 -278 -2567
rect -312 -2635 -278 -2611
rect -312 -2645 -278 -2635
rect -312 -2703 -278 -2683
rect -312 -2717 -278 -2703
rect -312 -2771 -278 -2755
rect -312 -2789 -278 -2771
rect -312 -2839 -278 -2827
rect -312 -2861 -278 -2839
rect -312 -2907 -278 -2899
rect -312 -2933 -278 -2907
rect -312 -2975 -278 -2971
rect -312 -3005 -278 -2975
rect -312 -3077 -278 -3043
rect -312 -3145 -278 -3115
rect -312 -3149 -278 -3145
rect -312 -3213 -278 -3187
rect -312 -3221 -278 -3213
rect -312 -3281 -278 -3259
rect -312 -3293 -278 -3281
rect -312 -3349 -278 -3331
rect -312 -3365 -278 -3349
rect -312 -3417 -278 -3403
rect -312 -3437 -278 -3417
rect -312 -3485 -278 -3475
rect -312 -3509 -278 -3485
rect -312 -3553 -278 -3547
rect -312 -3581 -278 -3553
rect -312 -3621 -278 -3619
rect -312 -3653 -278 -3621
rect -312 -3723 -278 -3691
rect -312 -3725 -278 -3723
rect -312 -3791 -278 -3763
rect -312 -3797 -278 -3791
rect -312 -3859 -278 -3835
rect -312 -3869 -278 -3859
rect -312 -3927 -278 -3907
rect -312 -3941 -278 -3927
rect -312 -3995 -278 -3979
rect -312 -4013 -278 -3995
rect -312 -4063 -278 -4051
rect -312 -4085 -278 -4063
rect -312 -4131 -278 -4123
rect -312 -4157 -278 -4131
rect -312 -4199 -278 -4195
rect -312 -4229 -278 -4199
rect -312 -4301 -278 -4267
rect -312 -4369 -278 -4339
rect -312 -4373 -278 -4369
rect -312 -4437 -278 -4411
rect -312 -4445 -278 -4437
rect -312 -4505 -278 -4483
rect -312 -4517 -278 -4505
rect -312 -4573 -278 -4555
rect -312 -4589 -278 -4573
rect -312 -4641 -278 -4627
rect -312 -4661 -278 -4641
rect -312 -4709 -278 -4699
rect -312 -4733 -278 -4709
rect -312 -4777 -278 -4771
rect -312 -4805 -278 -4777
rect -312 -4845 -278 -4843
rect -312 -4877 -278 -4845
rect -312 -4947 -278 -4915
rect -312 -4949 -278 -4947
rect -312 -5015 -278 -4987
rect -312 -5021 -278 -5015
rect -312 -5083 -278 -5059
rect -312 -5093 -278 -5083
rect -312 -5151 -278 -5131
rect -312 -5165 -278 -5151
rect -312 -5219 -278 -5203
rect -312 -5237 -278 -5219
rect -312 -5287 -278 -5275
rect -312 -5309 -278 -5287
rect -312 -5355 -278 -5347
rect -312 -5381 -278 -5355
rect -312 -5423 -278 -5419
rect -312 -5453 -278 -5423
rect -312 -5525 -278 -5491
rect -312 -5593 -278 -5563
rect -312 -5597 -278 -5593
rect -312 -5661 -278 -5635
rect -312 -5669 -278 -5661
rect -312 -5729 -278 -5707
rect -312 -5741 -278 -5729
rect -312 -5797 -278 -5779
rect -312 -5813 -278 -5797
rect -312 -5865 -278 -5851
rect -312 -5885 -278 -5865
rect -312 -5933 -278 -5923
rect -312 -5957 -278 -5933
rect -312 -6001 -278 -5995
rect -312 -6029 -278 -6001
rect -312 -6069 -278 -6067
rect -312 -6101 -278 -6069
rect -312 -6171 -278 -6139
rect -312 -6173 -278 -6171
rect -312 -6239 -278 -6211
rect -312 -6245 -278 -6239
rect -312 -6307 -278 -6283
rect -312 -6317 -278 -6307
rect -312 -6375 -278 -6355
rect -312 -6389 -278 -6375
rect -312 -6443 -278 -6427
rect -312 -6461 -278 -6443
rect -312 -6511 -278 -6499
rect -312 -6533 -278 -6511
rect -312 -6579 -278 -6571
rect -312 -6605 -278 -6579
rect -312 -6647 -278 -6643
rect -312 -6677 -278 -6647
rect -312 -6749 -278 -6715
rect -312 -6817 -278 -6787
rect -312 -6821 -278 -6817
rect -312 -6885 -278 -6859
rect -312 -6893 -278 -6885
rect -312 -6953 -278 -6931
rect -312 -6965 -278 -6953
rect -312 -7021 -278 -7003
rect -312 -7037 -278 -7021
rect -312 -7089 -278 -7075
rect -312 -7109 -278 -7089
rect -312 -7157 -278 -7147
rect -312 -7181 -278 -7157
rect -312 -7225 -278 -7219
rect -312 -7253 -278 -7225
rect -312 -7293 -278 -7291
rect -312 -7325 -278 -7293
rect -312 -7395 -278 -7363
rect -312 -7397 -278 -7395
rect -312 -7463 -278 -7435
rect -312 -7469 -278 -7463
rect -312 -7531 -278 -7507
rect -312 -7541 -278 -7531
rect -312 -7599 -278 -7579
rect -312 -7613 -278 -7599
rect -312 -7667 -278 -7651
rect -312 -7685 -278 -7667
rect -312 -7735 -278 -7723
rect -312 -7757 -278 -7735
rect -312 -7803 -278 -7795
rect -312 -7829 -278 -7803
rect -312 -7871 -278 -7867
rect -312 -7901 -278 -7871
rect -312 -7973 -278 -7939
rect -312 -8041 -278 -8011
rect -312 -8045 -278 -8041
rect -312 -8109 -278 -8083
rect -312 -8117 -278 -8109
rect -312 -8177 -278 -8155
rect -312 -8189 -278 -8177
rect -312 -8245 -278 -8227
rect -312 -8261 -278 -8245
rect -312 -8313 -278 -8299
rect -312 -8333 -278 -8313
rect -312 -8381 -278 -8371
rect -312 -8405 -278 -8381
rect -312 -8449 -278 -8443
rect -312 -8477 -278 -8449
rect -312 -8517 -278 -8515
rect -312 -8549 -278 -8517
rect -312 -8619 -278 -8587
rect -312 -8621 -278 -8619
rect -312 -8687 -278 -8659
rect -312 -8693 -278 -8687
rect -312 -8755 -278 -8731
rect -312 -8765 -278 -8755
rect -312 -8823 -278 -8803
rect -312 -8837 -278 -8823
rect -312 -8891 -278 -8875
rect -312 -8909 -278 -8891
rect -312 -8959 -278 -8947
rect -312 -8981 -278 -8959
rect -312 -9027 -278 -9019
rect -312 -9053 -278 -9027
rect -312 -9095 -278 -9091
rect -312 -9125 -278 -9095
rect -312 -9197 -278 -9163
rect -312 -9265 -278 -9235
rect -312 -9269 -278 -9265
rect -312 -9333 -278 -9307
rect -312 -9341 -278 -9333
rect -312 -9401 -278 -9379
rect -312 -9413 -278 -9401
rect -312 -9469 -278 -9451
rect -312 -9485 -278 -9469
rect -312 -9537 -278 -9523
rect -312 -9557 -278 -9537
rect -194 9537 -160 9557
rect -194 9523 -160 9537
rect -194 9469 -160 9485
rect -194 9451 -160 9469
rect -194 9401 -160 9413
rect -194 9379 -160 9401
rect -194 9333 -160 9341
rect -194 9307 -160 9333
rect -194 9265 -160 9269
rect -194 9235 -160 9265
rect -194 9163 -160 9197
rect -194 9095 -160 9125
rect -194 9091 -160 9095
rect -194 9027 -160 9053
rect -194 9019 -160 9027
rect -194 8959 -160 8981
rect -194 8947 -160 8959
rect -194 8891 -160 8909
rect -194 8875 -160 8891
rect -194 8823 -160 8837
rect -194 8803 -160 8823
rect -194 8755 -160 8765
rect -194 8731 -160 8755
rect -194 8687 -160 8693
rect -194 8659 -160 8687
rect -194 8619 -160 8621
rect -194 8587 -160 8619
rect -194 8517 -160 8549
rect -194 8515 -160 8517
rect -194 8449 -160 8477
rect -194 8443 -160 8449
rect -194 8381 -160 8405
rect -194 8371 -160 8381
rect -194 8313 -160 8333
rect -194 8299 -160 8313
rect -194 8245 -160 8261
rect -194 8227 -160 8245
rect -194 8177 -160 8189
rect -194 8155 -160 8177
rect -194 8109 -160 8117
rect -194 8083 -160 8109
rect -194 8041 -160 8045
rect -194 8011 -160 8041
rect -194 7939 -160 7973
rect -194 7871 -160 7901
rect -194 7867 -160 7871
rect -194 7803 -160 7829
rect -194 7795 -160 7803
rect -194 7735 -160 7757
rect -194 7723 -160 7735
rect -194 7667 -160 7685
rect -194 7651 -160 7667
rect -194 7599 -160 7613
rect -194 7579 -160 7599
rect -194 7531 -160 7541
rect -194 7507 -160 7531
rect -194 7463 -160 7469
rect -194 7435 -160 7463
rect -194 7395 -160 7397
rect -194 7363 -160 7395
rect -194 7293 -160 7325
rect -194 7291 -160 7293
rect -194 7225 -160 7253
rect -194 7219 -160 7225
rect -194 7157 -160 7181
rect -194 7147 -160 7157
rect -194 7089 -160 7109
rect -194 7075 -160 7089
rect -194 7021 -160 7037
rect -194 7003 -160 7021
rect -194 6953 -160 6965
rect -194 6931 -160 6953
rect -194 6885 -160 6893
rect -194 6859 -160 6885
rect -194 6817 -160 6821
rect -194 6787 -160 6817
rect -194 6715 -160 6749
rect -194 6647 -160 6677
rect -194 6643 -160 6647
rect -194 6579 -160 6605
rect -194 6571 -160 6579
rect -194 6511 -160 6533
rect -194 6499 -160 6511
rect -194 6443 -160 6461
rect -194 6427 -160 6443
rect -194 6375 -160 6389
rect -194 6355 -160 6375
rect -194 6307 -160 6317
rect -194 6283 -160 6307
rect -194 6239 -160 6245
rect -194 6211 -160 6239
rect -194 6171 -160 6173
rect -194 6139 -160 6171
rect -194 6069 -160 6101
rect -194 6067 -160 6069
rect -194 6001 -160 6029
rect -194 5995 -160 6001
rect -194 5933 -160 5957
rect -194 5923 -160 5933
rect -194 5865 -160 5885
rect -194 5851 -160 5865
rect -194 5797 -160 5813
rect -194 5779 -160 5797
rect -194 5729 -160 5741
rect -194 5707 -160 5729
rect -194 5661 -160 5669
rect -194 5635 -160 5661
rect -194 5593 -160 5597
rect -194 5563 -160 5593
rect -194 5491 -160 5525
rect -194 5423 -160 5453
rect -194 5419 -160 5423
rect -194 5355 -160 5381
rect -194 5347 -160 5355
rect -194 5287 -160 5309
rect -194 5275 -160 5287
rect -194 5219 -160 5237
rect -194 5203 -160 5219
rect -194 5151 -160 5165
rect -194 5131 -160 5151
rect -194 5083 -160 5093
rect -194 5059 -160 5083
rect -194 5015 -160 5021
rect -194 4987 -160 5015
rect -194 4947 -160 4949
rect -194 4915 -160 4947
rect -194 4845 -160 4877
rect -194 4843 -160 4845
rect -194 4777 -160 4805
rect -194 4771 -160 4777
rect -194 4709 -160 4733
rect -194 4699 -160 4709
rect -194 4641 -160 4661
rect -194 4627 -160 4641
rect -194 4573 -160 4589
rect -194 4555 -160 4573
rect -194 4505 -160 4517
rect -194 4483 -160 4505
rect -194 4437 -160 4445
rect -194 4411 -160 4437
rect -194 4369 -160 4373
rect -194 4339 -160 4369
rect -194 4267 -160 4301
rect -194 4199 -160 4229
rect -194 4195 -160 4199
rect -194 4131 -160 4157
rect -194 4123 -160 4131
rect -194 4063 -160 4085
rect -194 4051 -160 4063
rect -194 3995 -160 4013
rect -194 3979 -160 3995
rect -194 3927 -160 3941
rect -194 3907 -160 3927
rect -194 3859 -160 3869
rect -194 3835 -160 3859
rect -194 3791 -160 3797
rect -194 3763 -160 3791
rect -194 3723 -160 3725
rect -194 3691 -160 3723
rect -194 3621 -160 3653
rect -194 3619 -160 3621
rect -194 3553 -160 3581
rect -194 3547 -160 3553
rect -194 3485 -160 3509
rect -194 3475 -160 3485
rect -194 3417 -160 3437
rect -194 3403 -160 3417
rect -194 3349 -160 3365
rect -194 3331 -160 3349
rect -194 3281 -160 3293
rect -194 3259 -160 3281
rect -194 3213 -160 3221
rect -194 3187 -160 3213
rect -194 3145 -160 3149
rect -194 3115 -160 3145
rect -194 3043 -160 3077
rect -194 2975 -160 3005
rect -194 2971 -160 2975
rect -194 2907 -160 2933
rect -194 2899 -160 2907
rect -194 2839 -160 2861
rect -194 2827 -160 2839
rect -194 2771 -160 2789
rect -194 2755 -160 2771
rect -194 2703 -160 2717
rect -194 2683 -160 2703
rect -194 2635 -160 2645
rect -194 2611 -160 2635
rect -194 2567 -160 2573
rect -194 2539 -160 2567
rect -194 2499 -160 2501
rect -194 2467 -160 2499
rect -194 2397 -160 2429
rect -194 2395 -160 2397
rect -194 2329 -160 2357
rect -194 2323 -160 2329
rect -194 2261 -160 2285
rect -194 2251 -160 2261
rect -194 2193 -160 2213
rect -194 2179 -160 2193
rect -194 2125 -160 2141
rect -194 2107 -160 2125
rect -194 2057 -160 2069
rect -194 2035 -160 2057
rect -194 1989 -160 1997
rect -194 1963 -160 1989
rect -194 1921 -160 1925
rect -194 1891 -160 1921
rect -194 1819 -160 1853
rect -194 1751 -160 1781
rect -194 1747 -160 1751
rect -194 1683 -160 1709
rect -194 1675 -160 1683
rect -194 1615 -160 1637
rect -194 1603 -160 1615
rect -194 1547 -160 1565
rect -194 1531 -160 1547
rect -194 1479 -160 1493
rect -194 1459 -160 1479
rect -194 1411 -160 1421
rect -194 1387 -160 1411
rect -194 1343 -160 1349
rect -194 1315 -160 1343
rect -194 1275 -160 1277
rect -194 1243 -160 1275
rect -194 1173 -160 1205
rect -194 1171 -160 1173
rect -194 1105 -160 1133
rect -194 1099 -160 1105
rect -194 1037 -160 1061
rect -194 1027 -160 1037
rect -194 969 -160 989
rect -194 955 -160 969
rect -194 901 -160 917
rect -194 883 -160 901
rect -194 833 -160 845
rect -194 811 -160 833
rect -194 765 -160 773
rect -194 739 -160 765
rect -194 697 -160 701
rect -194 667 -160 697
rect -194 595 -160 629
rect -194 527 -160 557
rect -194 523 -160 527
rect -194 459 -160 485
rect -194 451 -160 459
rect -194 391 -160 413
rect -194 379 -160 391
rect -194 323 -160 341
rect -194 307 -160 323
rect -194 255 -160 269
rect -194 235 -160 255
rect -194 187 -160 197
rect -194 163 -160 187
rect -194 119 -160 125
rect -194 91 -160 119
rect -194 51 -160 53
rect -194 19 -160 51
rect -194 -51 -160 -19
rect -194 -53 -160 -51
rect -194 -119 -160 -91
rect -194 -125 -160 -119
rect -194 -187 -160 -163
rect -194 -197 -160 -187
rect -194 -255 -160 -235
rect -194 -269 -160 -255
rect -194 -323 -160 -307
rect -194 -341 -160 -323
rect -194 -391 -160 -379
rect -194 -413 -160 -391
rect -194 -459 -160 -451
rect -194 -485 -160 -459
rect -194 -527 -160 -523
rect -194 -557 -160 -527
rect -194 -629 -160 -595
rect -194 -697 -160 -667
rect -194 -701 -160 -697
rect -194 -765 -160 -739
rect -194 -773 -160 -765
rect -194 -833 -160 -811
rect -194 -845 -160 -833
rect -194 -901 -160 -883
rect -194 -917 -160 -901
rect -194 -969 -160 -955
rect -194 -989 -160 -969
rect -194 -1037 -160 -1027
rect -194 -1061 -160 -1037
rect -194 -1105 -160 -1099
rect -194 -1133 -160 -1105
rect -194 -1173 -160 -1171
rect -194 -1205 -160 -1173
rect -194 -1275 -160 -1243
rect -194 -1277 -160 -1275
rect -194 -1343 -160 -1315
rect -194 -1349 -160 -1343
rect -194 -1411 -160 -1387
rect -194 -1421 -160 -1411
rect -194 -1479 -160 -1459
rect -194 -1493 -160 -1479
rect -194 -1547 -160 -1531
rect -194 -1565 -160 -1547
rect -194 -1615 -160 -1603
rect -194 -1637 -160 -1615
rect -194 -1683 -160 -1675
rect -194 -1709 -160 -1683
rect -194 -1751 -160 -1747
rect -194 -1781 -160 -1751
rect -194 -1853 -160 -1819
rect -194 -1921 -160 -1891
rect -194 -1925 -160 -1921
rect -194 -1989 -160 -1963
rect -194 -1997 -160 -1989
rect -194 -2057 -160 -2035
rect -194 -2069 -160 -2057
rect -194 -2125 -160 -2107
rect -194 -2141 -160 -2125
rect -194 -2193 -160 -2179
rect -194 -2213 -160 -2193
rect -194 -2261 -160 -2251
rect -194 -2285 -160 -2261
rect -194 -2329 -160 -2323
rect -194 -2357 -160 -2329
rect -194 -2397 -160 -2395
rect -194 -2429 -160 -2397
rect -194 -2499 -160 -2467
rect -194 -2501 -160 -2499
rect -194 -2567 -160 -2539
rect -194 -2573 -160 -2567
rect -194 -2635 -160 -2611
rect -194 -2645 -160 -2635
rect -194 -2703 -160 -2683
rect -194 -2717 -160 -2703
rect -194 -2771 -160 -2755
rect -194 -2789 -160 -2771
rect -194 -2839 -160 -2827
rect -194 -2861 -160 -2839
rect -194 -2907 -160 -2899
rect -194 -2933 -160 -2907
rect -194 -2975 -160 -2971
rect -194 -3005 -160 -2975
rect -194 -3077 -160 -3043
rect -194 -3145 -160 -3115
rect -194 -3149 -160 -3145
rect -194 -3213 -160 -3187
rect -194 -3221 -160 -3213
rect -194 -3281 -160 -3259
rect -194 -3293 -160 -3281
rect -194 -3349 -160 -3331
rect -194 -3365 -160 -3349
rect -194 -3417 -160 -3403
rect -194 -3437 -160 -3417
rect -194 -3485 -160 -3475
rect -194 -3509 -160 -3485
rect -194 -3553 -160 -3547
rect -194 -3581 -160 -3553
rect -194 -3621 -160 -3619
rect -194 -3653 -160 -3621
rect -194 -3723 -160 -3691
rect -194 -3725 -160 -3723
rect -194 -3791 -160 -3763
rect -194 -3797 -160 -3791
rect -194 -3859 -160 -3835
rect -194 -3869 -160 -3859
rect -194 -3927 -160 -3907
rect -194 -3941 -160 -3927
rect -194 -3995 -160 -3979
rect -194 -4013 -160 -3995
rect -194 -4063 -160 -4051
rect -194 -4085 -160 -4063
rect -194 -4131 -160 -4123
rect -194 -4157 -160 -4131
rect -194 -4199 -160 -4195
rect -194 -4229 -160 -4199
rect -194 -4301 -160 -4267
rect -194 -4369 -160 -4339
rect -194 -4373 -160 -4369
rect -194 -4437 -160 -4411
rect -194 -4445 -160 -4437
rect -194 -4505 -160 -4483
rect -194 -4517 -160 -4505
rect -194 -4573 -160 -4555
rect -194 -4589 -160 -4573
rect -194 -4641 -160 -4627
rect -194 -4661 -160 -4641
rect -194 -4709 -160 -4699
rect -194 -4733 -160 -4709
rect -194 -4777 -160 -4771
rect -194 -4805 -160 -4777
rect -194 -4845 -160 -4843
rect -194 -4877 -160 -4845
rect -194 -4947 -160 -4915
rect -194 -4949 -160 -4947
rect -194 -5015 -160 -4987
rect -194 -5021 -160 -5015
rect -194 -5083 -160 -5059
rect -194 -5093 -160 -5083
rect -194 -5151 -160 -5131
rect -194 -5165 -160 -5151
rect -194 -5219 -160 -5203
rect -194 -5237 -160 -5219
rect -194 -5287 -160 -5275
rect -194 -5309 -160 -5287
rect -194 -5355 -160 -5347
rect -194 -5381 -160 -5355
rect -194 -5423 -160 -5419
rect -194 -5453 -160 -5423
rect -194 -5525 -160 -5491
rect -194 -5593 -160 -5563
rect -194 -5597 -160 -5593
rect -194 -5661 -160 -5635
rect -194 -5669 -160 -5661
rect -194 -5729 -160 -5707
rect -194 -5741 -160 -5729
rect -194 -5797 -160 -5779
rect -194 -5813 -160 -5797
rect -194 -5865 -160 -5851
rect -194 -5885 -160 -5865
rect -194 -5933 -160 -5923
rect -194 -5957 -160 -5933
rect -194 -6001 -160 -5995
rect -194 -6029 -160 -6001
rect -194 -6069 -160 -6067
rect -194 -6101 -160 -6069
rect -194 -6171 -160 -6139
rect -194 -6173 -160 -6171
rect -194 -6239 -160 -6211
rect -194 -6245 -160 -6239
rect -194 -6307 -160 -6283
rect -194 -6317 -160 -6307
rect -194 -6375 -160 -6355
rect -194 -6389 -160 -6375
rect -194 -6443 -160 -6427
rect -194 -6461 -160 -6443
rect -194 -6511 -160 -6499
rect -194 -6533 -160 -6511
rect -194 -6579 -160 -6571
rect -194 -6605 -160 -6579
rect -194 -6647 -160 -6643
rect -194 -6677 -160 -6647
rect -194 -6749 -160 -6715
rect -194 -6817 -160 -6787
rect -194 -6821 -160 -6817
rect -194 -6885 -160 -6859
rect -194 -6893 -160 -6885
rect -194 -6953 -160 -6931
rect -194 -6965 -160 -6953
rect -194 -7021 -160 -7003
rect -194 -7037 -160 -7021
rect -194 -7089 -160 -7075
rect -194 -7109 -160 -7089
rect -194 -7157 -160 -7147
rect -194 -7181 -160 -7157
rect -194 -7225 -160 -7219
rect -194 -7253 -160 -7225
rect -194 -7293 -160 -7291
rect -194 -7325 -160 -7293
rect -194 -7395 -160 -7363
rect -194 -7397 -160 -7395
rect -194 -7463 -160 -7435
rect -194 -7469 -160 -7463
rect -194 -7531 -160 -7507
rect -194 -7541 -160 -7531
rect -194 -7599 -160 -7579
rect -194 -7613 -160 -7599
rect -194 -7667 -160 -7651
rect -194 -7685 -160 -7667
rect -194 -7735 -160 -7723
rect -194 -7757 -160 -7735
rect -194 -7803 -160 -7795
rect -194 -7829 -160 -7803
rect -194 -7871 -160 -7867
rect -194 -7901 -160 -7871
rect -194 -7973 -160 -7939
rect -194 -8041 -160 -8011
rect -194 -8045 -160 -8041
rect -194 -8109 -160 -8083
rect -194 -8117 -160 -8109
rect -194 -8177 -160 -8155
rect -194 -8189 -160 -8177
rect -194 -8245 -160 -8227
rect -194 -8261 -160 -8245
rect -194 -8313 -160 -8299
rect -194 -8333 -160 -8313
rect -194 -8381 -160 -8371
rect -194 -8405 -160 -8381
rect -194 -8449 -160 -8443
rect -194 -8477 -160 -8449
rect -194 -8517 -160 -8515
rect -194 -8549 -160 -8517
rect -194 -8619 -160 -8587
rect -194 -8621 -160 -8619
rect -194 -8687 -160 -8659
rect -194 -8693 -160 -8687
rect -194 -8755 -160 -8731
rect -194 -8765 -160 -8755
rect -194 -8823 -160 -8803
rect -194 -8837 -160 -8823
rect -194 -8891 -160 -8875
rect -194 -8909 -160 -8891
rect -194 -8959 -160 -8947
rect -194 -8981 -160 -8959
rect -194 -9027 -160 -9019
rect -194 -9053 -160 -9027
rect -194 -9095 -160 -9091
rect -194 -9125 -160 -9095
rect -194 -9197 -160 -9163
rect -194 -9265 -160 -9235
rect -194 -9269 -160 -9265
rect -194 -9333 -160 -9307
rect -194 -9341 -160 -9333
rect -194 -9401 -160 -9379
rect -194 -9413 -160 -9401
rect -194 -9469 -160 -9451
rect -194 -9485 -160 -9469
rect -194 -9537 -160 -9523
rect -194 -9557 -160 -9537
rect -76 9537 -42 9557
rect -76 9523 -42 9537
rect -76 9469 -42 9485
rect -76 9451 -42 9469
rect -76 9401 -42 9413
rect -76 9379 -42 9401
rect -76 9333 -42 9341
rect -76 9307 -42 9333
rect -76 9265 -42 9269
rect -76 9235 -42 9265
rect -76 9163 -42 9197
rect -76 9095 -42 9125
rect -76 9091 -42 9095
rect -76 9027 -42 9053
rect -76 9019 -42 9027
rect -76 8959 -42 8981
rect -76 8947 -42 8959
rect -76 8891 -42 8909
rect -76 8875 -42 8891
rect -76 8823 -42 8837
rect -76 8803 -42 8823
rect -76 8755 -42 8765
rect -76 8731 -42 8755
rect -76 8687 -42 8693
rect -76 8659 -42 8687
rect -76 8619 -42 8621
rect -76 8587 -42 8619
rect -76 8517 -42 8549
rect -76 8515 -42 8517
rect -76 8449 -42 8477
rect -76 8443 -42 8449
rect -76 8381 -42 8405
rect -76 8371 -42 8381
rect -76 8313 -42 8333
rect -76 8299 -42 8313
rect -76 8245 -42 8261
rect -76 8227 -42 8245
rect -76 8177 -42 8189
rect -76 8155 -42 8177
rect -76 8109 -42 8117
rect -76 8083 -42 8109
rect -76 8041 -42 8045
rect -76 8011 -42 8041
rect -76 7939 -42 7973
rect -76 7871 -42 7901
rect -76 7867 -42 7871
rect -76 7803 -42 7829
rect -76 7795 -42 7803
rect -76 7735 -42 7757
rect -76 7723 -42 7735
rect -76 7667 -42 7685
rect -76 7651 -42 7667
rect -76 7599 -42 7613
rect -76 7579 -42 7599
rect -76 7531 -42 7541
rect -76 7507 -42 7531
rect -76 7463 -42 7469
rect -76 7435 -42 7463
rect -76 7395 -42 7397
rect -76 7363 -42 7395
rect -76 7293 -42 7325
rect -76 7291 -42 7293
rect -76 7225 -42 7253
rect -76 7219 -42 7225
rect -76 7157 -42 7181
rect -76 7147 -42 7157
rect -76 7089 -42 7109
rect -76 7075 -42 7089
rect -76 7021 -42 7037
rect -76 7003 -42 7021
rect -76 6953 -42 6965
rect -76 6931 -42 6953
rect -76 6885 -42 6893
rect -76 6859 -42 6885
rect -76 6817 -42 6821
rect -76 6787 -42 6817
rect -76 6715 -42 6749
rect -76 6647 -42 6677
rect -76 6643 -42 6647
rect -76 6579 -42 6605
rect -76 6571 -42 6579
rect -76 6511 -42 6533
rect -76 6499 -42 6511
rect -76 6443 -42 6461
rect -76 6427 -42 6443
rect -76 6375 -42 6389
rect -76 6355 -42 6375
rect -76 6307 -42 6317
rect -76 6283 -42 6307
rect -76 6239 -42 6245
rect -76 6211 -42 6239
rect -76 6171 -42 6173
rect -76 6139 -42 6171
rect -76 6069 -42 6101
rect -76 6067 -42 6069
rect -76 6001 -42 6029
rect -76 5995 -42 6001
rect -76 5933 -42 5957
rect -76 5923 -42 5933
rect -76 5865 -42 5885
rect -76 5851 -42 5865
rect -76 5797 -42 5813
rect -76 5779 -42 5797
rect -76 5729 -42 5741
rect -76 5707 -42 5729
rect -76 5661 -42 5669
rect -76 5635 -42 5661
rect -76 5593 -42 5597
rect -76 5563 -42 5593
rect -76 5491 -42 5525
rect -76 5423 -42 5453
rect -76 5419 -42 5423
rect -76 5355 -42 5381
rect -76 5347 -42 5355
rect -76 5287 -42 5309
rect -76 5275 -42 5287
rect -76 5219 -42 5237
rect -76 5203 -42 5219
rect -76 5151 -42 5165
rect -76 5131 -42 5151
rect -76 5083 -42 5093
rect -76 5059 -42 5083
rect -76 5015 -42 5021
rect -76 4987 -42 5015
rect -76 4947 -42 4949
rect -76 4915 -42 4947
rect -76 4845 -42 4877
rect -76 4843 -42 4845
rect -76 4777 -42 4805
rect -76 4771 -42 4777
rect -76 4709 -42 4733
rect -76 4699 -42 4709
rect -76 4641 -42 4661
rect -76 4627 -42 4641
rect -76 4573 -42 4589
rect -76 4555 -42 4573
rect -76 4505 -42 4517
rect -76 4483 -42 4505
rect -76 4437 -42 4445
rect -76 4411 -42 4437
rect -76 4369 -42 4373
rect -76 4339 -42 4369
rect -76 4267 -42 4301
rect -76 4199 -42 4229
rect -76 4195 -42 4199
rect -76 4131 -42 4157
rect -76 4123 -42 4131
rect -76 4063 -42 4085
rect -76 4051 -42 4063
rect -76 3995 -42 4013
rect -76 3979 -42 3995
rect -76 3927 -42 3941
rect -76 3907 -42 3927
rect -76 3859 -42 3869
rect -76 3835 -42 3859
rect -76 3791 -42 3797
rect -76 3763 -42 3791
rect -76 3723 -42 3725
rect -76 3691 -42 3723
rect -76 3621 -42 3653
rect -76 3619 -42 3621
rect -76 3553 -42 3581
rect -76 3547 -42 3553
rect -76 3485 -42 3509
rect -76 3475 -42 3485
rect -76 3417 -42 3437
rect -76 3403 -42 3417
rect -76 3349 -42 3365
rect -76 3331 -42 3349
rect -76 3281 -42 3293
rect -76 3259 -42 3281
rect -76 3213 -42 3221
rect -76 3187 -42 3213
rect -76 3145 -42 3149
rect -76 3115 -42 3145
rect -76 3043 -42 3077
rect -76 2975 -42 3005
rect -76 2971 -42 2975
rect -76 2907 -42 2933
rect -76 2899 -42 2907
rect -76 2839 -42 2861
rect -76 2827 -42 2839
rect -76 2771 -42 2789
rect -76 2755 -42 2771
rect -76 2703 -42 2717
rect -76 2683 -42 2703
rect -76 2635 -42 2645
rect -76 2611 -42 2635
rect -76 2567 -42 2573
rect -76 2539 -42 2567
rect -76 2499 -42 2501
rect -76 2467 -42 2499
rect -76 2397 -42 2429
rect -76 2395 -42 2397
rect -76 2329 -42 2357
rect -76 2323 -42 2329
rect -76 2261 -42 2285
rect -76 2251 -42 2261
rect -76 2193 -42 2213
rect -76 2179 -42 2193
rect -76 2125 -42 2141
rect -76 2107 -42 2125
rect -76 2057 -42 2069
rect -76 2035 -42 2057
rect -76 1989 -42 1997
rect -76 1963 -42 1989
rect -76 1921 -42 1925
rect -76 1891 -42 1921
rect -76 1819 -42 1853
rect -76 1751 -42 1781
rect -76 1747 -42 1751
rect -76 1683 -42 1709
rect -76 1675 -42 1683
rect -76 1615 -42 1637
rect -76 1603 -42 1615
rect -76 1547 -42 1565
rect -76 1531 -42 1547
rect -76 1479 -42 1493
rect -76 1459 -42 1479
rect -76 1411 -42 1421
rect -76 1387 -42 1411
rect -76 1343 -42 1349
rect -76 1315 -42 1343
rect -76 1275 -42 1277
rect -76 1243 -42 1275
rect -76 1173 -42 1205
rect -76 1171 -42 1173
rect -76 1105 -42 1133
rect -76 1099 -42 1105
rect -76 1037 -42 1061
rect -76 1027 -42 1037
rect -76 969 -42 989
rect -76 955 -42 969
rect -76 901 -42 917
rect -76 883 -42 901
rect -76 833 -42 845
rect -76 811 -42 833
rect -76 765 -42 773
rect -76 739 -42 765
rect -76 697 -42 701
rect -76 667 -42 697
rect -76 595 -42 629
rect -76 527 -42 557
rect -76 523 -42 527
rect -76 459 -42 485
rect -76 451 -42 459
rect -76 391 -42 413
rect -76 379 -42 391
rect -76 323 -42 341
rect -76 307 -42 323
rect -76 255 -42 269
rect -76 235 -42 255
rect -76 187 -42 197
rect -76 163 -42 187
rect -76 119 -42 125
rect -76 91 -42 119
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect -76 -119 -42 -91
rect -76 -125 -42 -119
rect -76 -187 -42 -163
rect -76 -197 -42 -187
rect -76 -255 -42 -235
rect -76 -269 -42 -255
rect -76 -323 -42 -307
rect -76 -341 -42 -323
rect -76 -391 -42 -379
rect -76 -413 -42 -391
rect -76 -459 -42 -451
rect -76 -485 -42 -459
rect -76 -527 -42 -523
rect -76 -557 -42 -527
rect -76 -629 -42 -595
rect -76 -697 -42 -667
rect -76 -701 -42 -697
rect -76 -765 -42 -739
rect -76 -773 -42 -765
rect -76 -833 -42 -811
rect -76 -845 -42 -833
rect -76 -901 -42 -883
rect -76 -917 -42 -901
rect -76 -969 -42 -955
rect -76 -989 -42 -969
rect -76 -1037 -42 -1027
rect -76 -1061 -42 -1037
rect -76 -1105 -42 -1099
rect -76 -1133 -42 -1105
rect -76 -1173 -42 -1171
rect -76 -1205 -42 -1173
rect -76 -1275 -42 -1243
rect -76 -1277 -42 -1275
rect -76 -1343 -42 -1315
rect -76 -1349 -42 -1343
rect -76 -1411 -42 -1387
rect -76 -1421 -42 -1411
rect -76 -1479 -42 -1459
rect -76 -1493 -42 -1479
rect -76 -1547 -42 -1531
rect -76 -1565 -42 -1547
rect -76 -1615 -42 -1603
rect -76 -1637 -42 -1615
rect -76 -1683 -42 -1675
rect -76 -1709 -42 -1683
rect -76 -1751 -42 -1747
rect -76 -1781 -42 -1751
rect -76 -1853 -42 -1819
rect -76 -1921 -42 -1891
rect -76 -1925 -42 -1921
rect -76 -1989 -42 -1963
rect -76 -1997 -42 -1989
rect -76 -2057 -42 -2035
rect -76 -2069 -42 -2057
rect -76 -2125 -42 -2107
rect -76 -2141 -42 -2125
rect -76 -2193 -42 -2179
rect -76 -2213 -42 -2193
rect -76 -2261 -42 -2251
rect -76 -2285 -42 -2261
rect -76 -2329 -42 -2323
rect -76 -2357 -42 -2329
rect -76 -2397 -42 -2395
rect -76 -2429 -42 -2397
rect -76 -2499 -42 -2467
rect -76 -2501 -42 -2499
rect -76 -2567 -42 -2539
rect -76 -2573 -42 -2567
rect -76 -2635 -42 -2611
rect -76 -2645 -42 -2635
rect -76 -2703 -42 -2683
rect -76 -2717 -42 -2703
rect -76 -2771 -42 -2755
rect -76 -2789 -42 -2771
rect -76 -2839 -42 -2827
rect -76 -2861 -42 -2839
rect -76 -2907 -42 -2899
rect -76 -2933 -42 -2907
rect -76 -2975 -42 -2971
rect -76 -3005 -42 -2975
rect -76 -3077 -42 -3043
rect -76 -3145 -42 -3115
rect -76 -3149 -42 -3145
rect -76 -3213 -42 -3187
rect -76 -3221 -42 -3213
rect -76 -3281 -42 -3259
rect -76 -3293 -42 -3281
rect -76 -3349 -42 -3331
rect -76 -3365 -42 -3349
rect -76 -3417 -42 -3403
rect -76 -3437 -42 -3417
rect -76 -3485 -42 -3475
rect -76 -3509 -42 -3485
rect -76 -3553 -42 -3547
rect -76 -3581 -42 -3553
rect -76 -3621 -42 -3619
rect -76 -3653 -42 -3621
rect -76 -3723 -42 -3691
rect -76 -3725 -42 -3723
rect -76 -3791 -42 -3763
rect -76 -3797 -42 -3791
rect -76 -3859 -42 -3835
rect -76 -3869 -42 -3859
rect -76 -3927 -42 -3907
rect -76 -3941 -42 -3927
rect -76 -3995 -42 -3979
rect -76 -4013 -42 -3995
rect -76 -4063 -42 -4051
rect -76 -4085 -42 -4063
rect -76 -4131 -42 -4123
rect -76 -4157 -42 -4131
rect -76 -4199 -42 -4195
rect -76 -4229 -42 -4199
rect -76 -4301 -42 -4267
rect -76 -4369 -42 -4339
rect -76 -4373 -42 -4369
rect -76 -4437 -42 -4411
rect -76 -4445 -42 -4437
rect -76 -4505 -42 -4483
rect -76 -4517 -42 -4505
rect -76 -4573 -42 -4555
rect -76 -4589 -42 -4573
rect -76 -4641 -42 -4627
rect -76 -4661 -42 -4641
rect -76 -4709 -42 -4699
rect -76 -4733 -42 -4709
rect -76 -4777 -42 -4771
rect -76 -4805 -42 -4777
rect -76 -4845 -42 -4843
rect -76 -4877 -42 -4845
rect -76 -4947 -42 -4915
rect -76 -4949 -42 -4947
rect -76 -5015 -42 -4987
rect -76 -5021 -42 -5015
rect -76 -5083 -42 -5059
rect -76 -5093 -42 -5083
rect -76 -5151 -42 -5131
rect -76 -5165 -42 -5151
rect -76 -5219 -42 -5203
rect -76 -5237 -42 -5219
rect -76 -5287 -42 -5275
rect -76 -5309 -42 -5287
rect -76 -5355 -42 -5347
rect -76 -5381 -42 -5355
rect -76 -5423 -42 -5419
rect -76 -5453 -42 -5423
rect -76 -5525 -42 -5491
rect -76 -5593 -42 -5563
rect -76 -5597 -42 -5593
rect -76 -5661 -42 -5635
rect -76 -5669 -42 -5661
rect -76 -5729 -42 -5707
rect -76 -5741 -42 -5729
rect -76 -5797 -42 -5779
rect -76 -5813 -42 -5797
rect -76 -5865 -42 -5851
rect -76 -5885 -42 -5865
rect -76 -5933 -42 -5923
rect -76 -5957 -42 -5933
rect -76 -6001 -42 -5995
rect -76 -6029 -42 -6001
rect -76 -6069 -42 -6067
rect -76 -6101 -42 -6069
rect -76 -6171 -42 -6139
rect -76 -6173 -42 -6171
rect -76 -6239 -42 -6211
rect -76 -6245 -42 -6239
rect -76 -6307 -42 -6283
rect -76 -6317 -42 -6307
rect -76 -6375 -42 -6355
rect -76 -6389 -42 -6375
rect -76 -6443 -42 -6427
rect -76 -6461 -42 -6443
rect -76 -6511 -42 -6499
rect -76 -6533 -42 -6511
rect -76 -6579 -42 -6571
rect -76 -6605 -42 -6579
rect -76 -6647 -42 -6643
rect -76 -6677 -42 -6647
rect -76 -6749 -42 -6715
rect -76 -6817 -42 -6787
rect -76 -6821 -42 -6817
rect -76 -6885 -42 -6859
rect -76 -6893 -42 -6885
rect -76 -6953 -42 -6931
rect -76 -6965 -42 -6953
rect -76 -7021 -42 -7003
rect -76 -7037 -42 -7021
rect -76 -7089 -42 -7075
rect -76 -7109 -42 -7089
rect -76 -7157 -42 -7147
rect -76 -7181 -42 -7157
rect -76 -7225 -42 -7219
rect -76 -7253 -42 -7225
rect -76 -7293 -42 -7291
rect -76 -7325 -42 -7293
rect -76 -7395 -42 -7363
rect -76 -7397 -42 -7395
rect -76 -7463 -42 -7435
rect -76 -7469 -42 -7463
rect -76 -7531 -42 -7507
rect -76 -7541 -42 -7531
rect -76 -7599 -42 -7579
rect -76 -7613 -42 -7599
rect -76 -7667 -42 -7651
rect -76 -7685 -42 -7667
rect -76 -7735 -42 -7723
rect -76 -7757 -42 -7735
rect -76 -7803 -42 -7795
rect -76 -7829 -42 -7803
rect -76 -7871 -42 -7867
rect -76 -7901 -42 -7871
rect -76 -7973 -42 -7939
rect -76 -8041 -42 -8011
rect -76 -8045 -42 -8041
rect -76 -8109 -42 -8083
rect -76 -8117 -42 -8109
rect -76 -8177 -42 -8155
rect -76 -8189 -42 -8177
rect -76 -8245 -42 -8227
rect -76 -8261 -42 -8245
rect -76 -8313 -42 -8299
rect -76 -8333 -42 -8313
rect -76 -8381 -42 -8371
rect -76 -8405 -42 -8381
rect -76 -8449 -42 -8443
rect -76 -8477 -42 -8449
rect -76 -8517 -42 -8515
rect -76 -8549 -42 -8517
rect -76 -8619 -42 -8587
rect -76 -8621 -42 -8619
rect -76 -8687 -42 -8659
rect -76 -8693 -42 -8687
rect -76 -8755 -42 -8731
rect -76 -8765 -42 -8755
rect -76 -8823 -42 -8803
rect -76 -8837 -42 -8823
rect -76 -8891 -42 -8875
rect -76 -8909 -42 -8891
rect -76 -8959 -42 -8947
rect -76 -8981 -42 -8959
rect -76 -9027 -42 -9019
rect -76 -9053 -42 -9027
rect -76 -9095 -42 -9091
rect -76 -9125 -42 -9095
rect -76 -9197 -42 -9163
rect -76 -9265 -42 -9235
rect -76 -9269 -42 -9265
rect -76 -9333 -42 -9307
rect -76 -9341 -42 -9333
rect -76 -9401 -42 -9379
rect -76 -9413 -42 -9401
rect -76 -9469 -42 -9451
rect -76 -9485 -42 -9469
rect -76 -9537 -42 -9523
rect -76 -9557 -42 -9537
rect 42 9537 76 9557
rect 42 9523 76 9537
rect 42 9469 76 9485
rect 42 9451 76 9469
rect 42 9401 76 9413
rect 42 9379 76 9401
rect 42 9333 76 9341
rect 42 9307 76 9333
rect 42 9265 76 9269
rect 42 9235 76 9265
rect 42 9163 76 9197
rect 42 9095 76 9125
rect 42 9091 76 9095
rect 42 9027 76 9053
rect 42 9019 76 9027
rect 42 8959 76 8981
rect 42 8947 76 8959
rect 42 8891 76 8909
rect 42 8875 76 8891
rect 42 8823 76 8837
rect 42 8803 76 8823
rect 42 8755 76 8765
rect 42 8731 76 8755
rect 42 8687 76 8693
rect 42 8659 76 8687
rect 42 8619 76 8621
rect 42 8587 76 8619
rect 42 8517 76 8549
rect 42 8515 76 8517
rect 42 8449 76 8477
rect 42 8443 76 8449
rect 42 8381 76 8405
rect 42 8371 76 8381
rect 42 8313 76 8333
rect 42 8299 76 8313
rect 42 8245 76 8261
rect 42 8227 76 8245
rect 42 8177 76 8189
rect 42 8155 76 8177
rect 42 8109 76 8117
rect 42 8083 76 8109
rect 42 8041 76 8045
rect 42 8011 76 8041
rect 42 7939 76 7973
rect 42 7871 76 7901
rect 42 7867 76 7871
rect 42 7803 76 7829
rect 42 7795 76 7803
rect 42 7735 76 7757
rect 42 7723 76 7735
rect 42 7667 76 7685
rect 42 7651 76 7667
rect 42 7599 76 7613
rect 42 7579 76 7599
rect 42 7531 76 7541
rect 42 7507 76 7531
rect 42 7463 76 7469
rect 42 7435 76 7463
rect 42 7395 76 7397
rect 42 7363 76 7395
rect 42 7293 76 7325
rect 42 7291 76 7293
rect 42 7225 76 7253
rect 42 7219 76 7225
rect 42 7157 76 7181
rect 42 7147 76 7157
rect 42 7089 76 7109
rect 42 7075 76 7089
rect 42 7021 76 7037
rect 42 7003 76 7021
rect 42 6953 76 6965
rect 42 6931 76 6953
rect 42 6885 76 6893
rect 42 6859 76 6885
rect 42 6817 76 6821
rect 42 6787 76 6817
rect 42 6715 76 6749
rect 42 6647 76 6677
rect 42 6643 76 6647
rect 42 6579 76 6605
rect 42 6571 76 6579
rect 42 6511 76 6533
rect 42 6499 76 6511
rect 42 6443 76 6461
rect 42 6427 76 6443
rect 42 6375 76 6389
rect 42 6355 76 6375
rect 42 6307 76 6317
rect 42 6283 76 6307
rect 42 6239 76 6245
rect 42 6211 76 6239
rect 42 6171 76 6173
rect 42 6139 76 6171
rect 42 6069 76 6101
rect 42 6067 76 6069
rect 42 6001 76 6029
rect 42 5995 76 6001
rect 42 5933 76 5957
rect 42 5923 76 5933
rect 42 5865 76 5885
rect 42 5851 76 5865
rect 42 5797 76 5813
rect 42 5779 76 5797
rect 42 5729 76 5741
rect 42 5707 76 5729
rect 42 5661 76 5669
rect 42 5635 76 5661
rect 42 5593 76 5597
rect 42 5563 76 5593
rect 42 5491 76 5525
rect 42 5423 76 5453
rect 42 5419 76 5423
rect 42 5355 76 5381
rect 42 5347 76 5355
rect 42 5287 76 5309
rect 42 5275 76 5287
rect 42 5219 76 5237
rect 42 5203 76 5219
rect 42 5151 76 5165
rect 42 5131 76 5151
rect 42 5083 76 5093
rect 42 5059 76 5083
rect 42 5015 76 5021
rect 42 4987 76 5015
rect 42 4947 76 4949
rect 42 4915 76 4947
rect 42 4845 76 4877
rect 42 4843 76 4845
rect 42 4777 76 4805
rect 42 4771 76 4777
rect 42 4709 76 4733
rect 42 4699 76 4709
rect 42 4641 76 4661
rect 42 4627 76 4641
rect 42 4573 76 4589
rect 42 4555 76 4573
rect 42 4505 76 4517
rect 42 4483 76 4505
rect 42 4437 76 4445
rect 42 4411 76 4437
rect 42 4369 76 4373
rect 42 4339 76 4369
rect 42 4267 76 4301
rect 42 4199 76 4229
rect 42 4195 76 4199
rect 42 4131 76 4157
rect 42 4123 76 4131
rect 42 4063 76 4085
rect 42 4051 76 4063
rect 42 3995 76 4013
rect 42 3979 76 3995
rect 42 3927 76 3941
rect 42 3907 76 3927
rect 42 3859 76 3869
rect 42 3835 76 3859
rect 42 3791 76 3797
rect 42 3763 76 3791
rect 42 3723 76 3725
rect 42 3691 76 3723
rect 42 3621 76 3653
rect 42 3619 76 3621
rect 42 3553 76 3581
rect 42 3547 76 3553
rect 42 3485 76 3509
rect 42 3475 76 3485
rect 42 3417 76 3437
rect 42 3403 76 3417
rect 42 3349 76 3365
rect 42 3331 76 3349
rect 42 3281 76 3293
rect 42 3259 76 3281
rect 42 3213 76 3221
rect 42 3187 76 3213
rect 42 3145 76 3149
rect 42 3115 76 3145
rect 42 3043 76 3077
rect 42 2975 76 3005
rect 42 2971 76 2975
rect 42 2907 76 2933
rect 42 2899 76 2907
rect 42 2839 76 2861
rect 42 2827 76 2839
rect 42 2771 76 2789
rect 42 2755 76 2771
rect 42 2703 76 2717
rect 42 2683 76 2703
rect 42 2635 76 2645
rect 42 2611 76 2635
rect 42 2567 76 2573
rect 42 2539 76 2567
rect 42 2499 76 2501
rect 42 2467 76 2499
rect 42 2397 76 2429
rect 42 2395 76 2397
rect 42 2329 76 2357
rect 42 2323 76 2329
rect 42 2261 76 2285
rect 42 2251 76 2261
rect 42 2193 76 2213
rect 42 2179 76 2193
rect 42 2125 76 2141
rect 42 2107 76 2125
rect 42 2057 76 2069
rect 42 2035 76 2057
rect 42 1989 76 1997
rect 42 1963 76 1989
rect 42 1921 76 1925
rect 42 1891 76 1921
rect 42 1819 76 1853
rect 42 1751 76 1781
rect 42 1747 76 1751
rect 42 1683 76 1709
rect 42 1675 76 1683
rect 42 1615 76 1637
rect 42 1603 76 1615
rect 42 1547 76 1565
rect 42 1531 76 1547
rect 42 1479 76 1493
rect 42 1459 76 1479
rect 42 1411 76 1421
rect 42 1387 76 1411
rect 42 1343 76 1349
rect 42 1315 76 1343
rect 42 1275 76 1277
rect 42 1243 76 1275
rect 42 1173 76 1205
rect 42 1171 76 1173
rect 42 1105 76 1133
rect 42 1099 76 1105
rect 42 1037 76 1061
rect 42 1027 76 1037
rect 42 969 76 989
rect 42 955 76 969
rect 42 901 76 917
rect 42 883 76 901
rect 42 833 76 845
rect 42 811 76 833
rect 42 765 76 773
rect 42 739 76 765
rect 42 697 76 701
rect 42 667 76 697
rect 42 595 76 629
rect 42 527 76 557
rect 42 523 76 527
rect 42 459 76 485
rect 42 451 76 459
rect 42 391 76 413
rect 42 379 76 391
rect 42 323 76 341
rect 42 307 76 323
rect 42 255 76 269
rect 42 235 76 255
rect 42 187 76 197
rect 42 163 76 187
rect 42 119 76 125
rect 42 91 76 119
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect 42 -119 76 -91
rect 42 -125 76 -119
rect 42 -187 76 -163
rect 42 -197 76 -187
rect 42 -255 76 -235
rect 42 -269 76 -255
rect 42 -323 76 -307
rect 42 -341 76 -323
rect 42 -391 76 -379
rect 42 -413 76 -391
rect 42 -459 76 -451
rect 42 -485 76 -459
rect 42 -527 76 -523
rect 42 -557 76 -527
rect 42 -629 76 -595
rect 42 -697 76 -667
rect 42 -701 76 -697
rect 42 -765 76 -739
rect 42 -773 76 -765
rect 42 -833 76 -811
rect 42 -845 76 -833
rect 42 -901 76 -883
rect 42 -917 76 -901
rect 42 -969 76 -955
rect 42 -989 76 -969
rect 42 -1037 76 -1027
rect 42 -1061 76 -1037
rect 42 -1105 76 -1099
rect 42 -1133 76 -1105
rect 42 -1173 76 -1171
rect 42 -1205 76 -1173
rect 42 -1275 76 -1243
rect 42 -1277 76 -1275
rect 42 -1343 76 -1315
rect 42 -1349 76 -1343
rect 42 -1411 76 -1387
rect 42 -1421 76 -1411
rect 42 -1479 76 -1459
rect 42 -1493 76 -1479
rect 42 -1547 76 -1531
rect 42 -1565 76 -1547
rect 42 -1615 76 -1603
rect 42 -1637 76 -1615
rect 42 -1683 76 -1675
rect 42 -1709 76 -1683
rect 42 -1751 76 -1747
rect 42 -1781 76 -1751
rect 42 -1853 76 -1819
rect 42 -1921 76 -1891
rect 42 -1925 76 -1921
rect 42 -1989 76 -1963
rect 42 -1997 76 -1989
rect 42 -2057 76 -2035
rect 42 -2069 76 -2057
rect 42 -2125 76 -2107
rect 42 -2141 76 -2125
rect 42 -2193 76 -2179
rect 42 -2213 76 -2193
rect 42 -2261 76 -2251
rect 42 -2285 76 -2261
rect 42 -2329 76 -2323
rect 42 -2357 76 -2329
rect 42 -2397 76 -2395
rect 42 -2429 76 -2397
rect 42 -2499 76 -2467
rect 42 -2501 76 -2499
rect 42 -2567 76 -2539
rect 42 -2573 76 -2567
rect 42 -2635 76 -2611
rect 42 -2645 76 -2635
rect 42 -2703 76 -2683
rect 42 -2717 76 -2703
rect 42 -2771 76 -2755
rect 42 -2789 76 -2771
rect 42 -2839 76 -2827
rect 42 -2861 76 -2839
rect 42 -2907 76 -2899
rect 42 -2933 76 -2907
rect 42 -2975 76 -2971
rect 42 -3005 76 -2975
rect 42 -3077 76 -3043
rect 42 -3145 76 -3115
rect 42 -3149 76 -3145
rect 42 -3213 76 -3187
rect 42 -3221 76 -3213
rect 42 -3281 76 -3259
rect 42 -3293 76 -3281
rect 42 -3349 76 -3331
rect 42 -3365 76 -3349
rect 42 -3417 76 -3403
rect 42 -3437 76 -3417
rect 42 -3485 76 -3475
rect 42 -3509 76 -3485
rect 42 -3553 76 -3547
rect 42 -3581 76 -3553
rect 42 -3621 76 -3619
rect 42 -3653 76 -3621
rect 42 -3723 76 -3691
rect 42 -3725 76 -3723
rect 42 -3791 76 -3763
rect 42 -3797 76 -3791
rect 42 -3859 76 -3835
rect 42 -3869 76 -3859
rect 42 -3927 76 -3907
rect 42 -3941 76 -3927
rect 42 -3995 76 -3979
rect 42 -4013 76 -3995
rect 42 -4063 76 -4051
rect 42 -4085 76 -4063
rect 42 -4131 76 -4123
rect 42 -4157 76 -4131
rect 42 -4199 76 -4195
rect 42 -4229 76 -4199
rect 42 -4301 76 -4267
rect 42 -4369 76 -4339
rect 42 -4373 76 -4369
rect 42 -4437 76 -4411
rect 42 -4445 76 -4437
rect 42 -4505 76 -4483
rect 42 -4517 76 -4505
rect 42 -4573 76 -4555
rect 42 -4589 76 -4573
rect 42 -4641 76 -4627
rect 42 -4661 76 -4641
rect 42 -4709 76 -4699
rect 42 -4733 76 -4709
rect 42 -4777 76 -4771
rect 42 -4805 76 -4777
rect 42 -4845 76 -4843
rect 42 -4877 76 -4845
rect 42 -4947 76 -4915
rect 42 -4949 76 -4947
rect 42 -5015 76 -4987
rect 42 -5021 76 -5015
rect 42 -5083 76 -5059
rect 42 -5093 76 -5083
rect 42 -5151 76 -5131
rect 42 -5165 76 -5151
rect 42 -5219 76 -5203
rect 42 -5237 76 -5219
rect 42 -5287 76 -5275
rect 42 -5309 76 -5287
rect 42 -5355 76 -5347
rect 42 -5381 76 -5355
rect 42 -5423 76 -5419
rect 42 -5453 76 -5423
rect 42 -5525 76 -5491
rect 42 -5593 76 -5563
rect 42 -5597 76 -5593
rect 42 -5661 76 -5635
rect 42 -5669 76 -5661
rect 42 -5729 76 -5707
rect 42 -5741 76 -5729
rect 42 -5797 76 -5779
rect 42 -5813 76 -5797
rect 42 -5865 76 -5851
rect 42 -5885 76 -5865
rect 42 -5933 76 -5923
rect 42 -5957 76 -5933
rect 42 -6001 76 -5995
rect 42 -6029 76 -6001
rect 42 -6069 76 -6067
rect 42 -6101 76 -6069
rect 42 -6171 76 -6139
rect 42 -6173 76 -6171
rect 42 -6239 76 -6211
rect 42 -6245 76 -6239
rect 42 -6307 76 -6283
rect 42 -6317 76 -6307
rect 42 -6375 76 -6355
rect 42 -6389 76 -6375
rect 42 -6443 76 -6427
rect 42 -6461 76 -6443
rect 42 -6511 76 -6499
rect 42 -6533 76 -6511
rect 42 -6579 76 -6571
rect 42 -6605 76 -6579
rect 42 -6647 76 -6643
rect 42 -6677 76 -6647
rect 42 -6749 76 -6715
rect 42 -6817 76 -6787
rect 42 -6821 76 -6817
rect 42 -6885 76 -6859
rect 42 -6893 76 -6885
rect 42 -6953 76 -6931
rect 42 -6965 76 -6953
rect 42 -7021 76 -7003
rect 42 -7037 76 -7021
rect 42 -7089 76 -7075
rect 42 -7109 76 -7089
rect 42 -7157 76 -7147
rect 42 -7181 76 -7157
rect 42 -7225 76 -7219
rect 42 -7253 76 -7225
rect 42 -7293 76 -7291
rect 42 -7325 76 -7293
rect 42 -7395 76 -7363
rect 42 -7397 76 -7395
rect 42 -7463 76 -7435
rect 42 -7469 76 -7463
rect 42 -7531 76 -7507
rect 42 -7541 76 -7531
rect 42 -7599 76 -7579
rect 42 -7613 76 -7599
rect 42 -7667 76 -7651
rect 42 -7685 76 -7667
rect 42 -7735 76 -7723
rect 42 -7757 76 -7735
rect 42 -7803 76 -7795
rect 42 -7829 76 -7803
rect 42 -7871 76 -7867
rect 42 -7901 76 -7871
rect 42 -7973 76 -7939
rect 42 -8041 76 -8011
rect 42 -8045 76 -8041
rect 42 -8109 76 -8083
rect 42 -8117 76 -8109
rect 42 -8177 76 -8155
rect 42 -8189 76 -8177
rect 42 -8245 76 -8227
rect 42 -8261 76 -8245
rect 42 -8313 76 -8299
rect 42 -8333 76 -8313
rect 42 -8381 76 -8371
rect 42 -8405 76 -8381
rect 42 -8449 76 -8443
rect 42 -8477 76 -8449
rect 42 -8517 76 -8515
rect 42 -8549 76 -8517
rect 42 -8619 76 -8587
rect 42 -8621 76 -8619
rect 42 -8687 76 -8659
rect 42 -8693 76 -8687
rect 42 -8755 76 -8731
rect 42 -8765 76 -8755
rect 42 -8823 76 -8803
rect 42 -8837 76 -8823
rect 42 -8891 76 -8875
rect 42 -8909 76 -8891
rect 42 -8959 76 -8947
rect 42 -8981 76 -8959
rect 42 -9027 76 -9019
rect 42 -9053 76 -9027
rect 42 -9095 76 -9091
rect 42 -9125 76 -9095
rect 42 -9197 76 -9163
rect 42 -9265 76 -9235
rect 42 -9269 76 -9265
rect 42 -9333 76 -9307
rect 42 -9341 76 -9333
rect 42 -9401 76 -9379
rect 42 -9413 76 -9401
rect 42 -9469 76 -9451
rect 42 -9485 76 -9469
rect 42 -9537 76 -9523
rect 42 -9557 76 -9537
rect 160 9537 194 9557
rect 160 9523 194 9537
rect 160 9469 194 9485
rect 160 9451 194 9469
rect 160 9401 194 9413
rect 160 9379 194 9401
rect 160 9333 194 9341
rect 160 9307 194 9333
rect 160 9265 194 9269
rect 160 9235 194 9265
rect 160 9163 194 9197
rect 160 9095 194 9125
rect 160 9091 194 9095
rect 160 9027 194 9053
rect 160 9019 194 9027
rect 160 8959 194 8981
rect 160 8947 194 8959
rect 160 8891 194 8909
rect 160 8875 194 8891
rect 160 8823 194 8837
rect 160 8803 194 8823
rect 160 8755 194 8765
rect 160 8731 194 8755
rect 160 8687 194 8693
rect 160 8659 194 8687
rect 160 8619 194 8621
rect 160 8587 194 8619
rect 160 8517 194 8549
rect 160 8515 194 8517
rect 160 8449 194 8477
rect 160 8443 194 8449
rect 160 8381 194 8405
rect 160 8371 194 8381
rect 160 8313 194 8333
rect 160 8299 194 8313
rect 160 8245 194 8261
rect 160 8227 194 8245
rect 160 8177 194 8189
rect 160 8155 194 8177
rect 160 8109 194 8117
rect 160 8083 194 8109
rect 160 8041 194 8045
rect 160 8011 194 8041
rect 160 7939 194 7973
rect 160 7871 194 7901
rect 160 7867 194 7871
rect 160 7803 194 7829
rect 160 7795 194 7803
rect 160 7735 194 7757
rect 160 7723 194 7735
rect 160 7667 194 7685
rect 160 7651 194 7667
rect 160 7599 194 7613
rect 160 7579 194 7599
rect 160 7531 194 7541
rect 160 7507 194 7531
rect 160 7463 194 7469
rect 160 7435 194 7463
rect 160 7395 194 7397
rect 160 7363 194 7395
rect 160 7293 194 7325
rect 160 7291 194 7293
rect 160 7225 194 7253
rect 160 7219 194 7225
rect 160 7157 194 7181
rect 160 7147 194 7157
rect 160 7089 194 7109
rect 160 7075 194 7089
rect 160 7021 194 7037
rect 160 7003 194 7021
rect 160 6953 194 6965
rect 160 6931 194 6953
rect 160 6885 194 6893
rect 160 6859 194 6885
rect 160 6817 194 6821
rect 160 6787 194 6817
rect 160 6715 194 6749
rect 160 6647 194 6677
rect 160 6643 194 6647
rect 160 6579 194 6605
rect 160 6571 194 6579
rect 160 6511 194 6533
rect 160 6499 194 6511
rect 160 6443 194 6461
rect 160 6427 194 6443
rect 160 6375 194 6389
rect 160 6355 194 6375
rect 160 6307 194 6317
rect 160 6283 194 6307
rect 160 6239 194 6245
rect 160 6211 194 6239
rect 160 6171 194 6173
rect 160 6139 194 6171
rect 160 6069 194 6101
rect 160 6067 194 6069
rect 160 6001 194 6029
rect 160 5995 194 6001
rect 160 5933 194 5957
rect 160 5923 194 5933
rect 160 5865 194 5885
rect 160 5851 194 5865
rect 160 5797 194 5813
rect 160 5779 194 5797
rect 160 5729 194 5741
rect 160 5707 194 5729
rect 160 5661 194 5669
rect 160 5635 194 5661
rect 160 5593 194 5597
rect 160 5563 194 5593
rect 160 5491 194 5525
rect 160 5423 194 5453
rect 160 5419 194 5423
rect 160 5355 194 5381
rect 160 5347 194 5355
rect 160 5287 194 5309
rect 160 5275 194 5287
rect 160 5219 194 5237
rect 160 5203 194 5219
rect 160 5151 194 5165
rect 160 5131 194 5151
rect 160 5083 194 5093
rect 160 5059 194 5083
rect 160 5015 194 5021
rect 160 4987 194 5015
rect 160 4947 194 4949
rect 160 4915 194 4947
rect 160 4845 194 4877
rect 160 4843 194 4845
rect 160 4777 194 4805
rect 160 4771 194 4777
rect 160 4709 194 4733
rect 160 4699 194 4709
rect 160 4641 194 4661
rect 160 4627 194 4641
rect 160 4573 194 4589
rect 160 4555 194 4573
rect 160 4505 194 4517
rect 160 4483 194 4505
rect 160 4437 194 4445
rect 160 4411 194 4437
rect 160 4369 194 4373
rect 160 4339 194 4369
rect 160 4267 194 4301
rect 160 4199 194 4229
rect 160 4195 194 4199
rect 160 4131 194 4157
rect 160 4123 194 4131
rect 160 4063 194 4085
rect 160 4051 194 4063
rect 160 3995 194 4013
rect 160 3979 194 3995
rect 160 3927 194 3941
rect 160 3907 194 3927
rect 160 3859 194 3869
rect 160 3835 194 3859
rect 160 3791 194 3797
rect 160 3763 194 3791
rect 160 3723 194 3725
rect 160 3691 194 3723
rect 160 3621 194 3653
rect 160 3619 194 3621
rect 160 3553 194 3581
rect 160 3547 194 3553
rect 160 3485 194 3509
rect 160 3475 194 3485
rect 160 3417 194 3437
rect 160 3403 194 3417
rect 160 3349 194 3365
rect 160 3331 194 3349
rect 160 3281 194 3293
rect 160 3259 194 3281
rect 160 3213 194 3221
rect 160 3187 194 3213
rect 160 3145 194 3149
rect 160 3115 194 3145
rect 160 3043 194 3077
rect 160 2975 194 3005
rect 160 2971 194 2975
rect 160 2907 194 2933
rect 160 2899 194 2907
rect 160 2839 194 2861
rect 160 2827 194 2839
rect 160 2771 194 2789
rect 160 2755 194 2771
rect 160 2703 194 2717
rect 160 2683 194 2703
rect 160 2635 194 2645
rect 160 2611 194 2635
rect 160 2567 194 2573
rect 160 2539 194 2567
rect 160 2499 194 2501
rect 160 2467 194 2499
rect 160 2397 194 2429
rect 160 2395 194 2397
rect 160 2329 194 2357
rect 160 2323 194 2329
rect 160 2261 194 2285
rect 160 2251 194 2261
rect 160 2193 194 2213
rect 160 2179 194 2193
rect 160 2125 194 2141
rect 160 2107 194 2125
rect 160 2057 194 2069
rect 160 2035 194 2057
rect 160 1989 194 1997
rect 160 1963 194 1989
rect 160 1921 194 1925
rect 160 1891 194 1921
rect 160 1819 194 1853
rect 160 1751 194 1781
rect 160 1747 194 1751
rect 160 1683 194 1709
rect 160 1675 194 1683
rect 160 1615 194 1637
rect 160 1603 194 1615
rect 160 1547 194 1565
rect 160 1531 194 1547
rect 160 1479 194 1493
rect 160 1459 194 1479
rect 160 1411 194 1421
rect 160 1387 194 1411
rect 160 1343 194 1349
rect 160 1315 194 1343
rect 160 1275 194 1277
rect 160 1243 194 1275
rect 160 1173 194 1205
rect 160 1171 194 1173
rect 160 1105 194 1133
rect 160 1099 194 1105
rect 160 1037 194 1061
rect 160 1027 194 1037
rect 160 969 194 989
rect 160 955 194 969
rect 160 901 194 917
rect 160 883 194 901
rect 160 833 194 845
rect 160 811 194 833
rect 160 765 194 773
rect 160 739 194 765
rect 160 697 194 701
rect 160 667 194 697
rect 160 595 194 629
rect 160 527 194 557
rect 160 523 194 527
rect 160 459 194 485
rect 160 451 194 459
rect 160 391 194 413
rect 160 379 194 391
rect 160 323 194 341
rect 160 307 194 323
rect 160 255 194 269
rect 160 235 194 255
rect 160 187 194 197
rect 160 163 194 187
rect 160 119 194 125
rect 160 91 194 119
rect 160 51 194 53
rect 160 19 194 51
rect 160 -51 194 -19
rect 160 -53 194 -51
rect 160 -119 194 -91
rect 160 -125 194 -119
rect 160 -187 194 -163
rect 160 -197 194 -187
rect 160 -255 194 -235
rect 160 -269 194 -255
rect 160 -323 194 -307
rect 160 -341 194 -323
rect 160 -391 194 -379
rect 160 -413 194 -391
rect 160 -459 194 -451
rect 160 -485 194 -459
rect 160 -527 194 -523
rect 160 -557 194 -527
rect 160 -629 194 -595
rect 160 -697 194 -667
rect 160 -701 194 -697
rect 160 -765 194 -739
rect 160 -773 194 -765
rect 160 -833 194 -811
rect 160 -845 194 -833
rect 160 -901 194 -883
rect 160 -917 194 -901
rect 160 -969 194 -955
rect 160 -989 194 -969
rect 160 -1037 194 -1027
rect 160 -1061 194 -1037
rect 160 -1105 194 -1099
rect 160 -1133 194 -1105
rect 160 -1173 194 -1171
rect 160 -1205 194 -1173
rect 160 -1275 194 -1243
rect 160 -1277 194 -1275
rect 160 -1343 194 -1315
rect 160 -1349 194 -1343
rect 160 -1411 194 -1387
rect 160 -1421 194 -1411
rect 160 -1479 194 -1459
rect 160 -1493 194 -1479
rect 160 -1547 194 -1531
rect 160 -1565 194 -1547
rect 160 -1615 194 -1603
rect 160 -1637 194 -1615
rect 160 -1683 194 -1675
rect 160 -1709 194 -1683
rect 160 -1751 194 -1747
rect 160 -1781 194 -1751
rect 160 -1853 194 -1819
rect 160 -1921 194 -1891
rect 160 -1925 194 -1921
rect 160 -1989 194 -1963
rect 160 -1997 194 -1989
rect 160 -2057 194 -2035
rect 160 -2069 194 -2057
rect 160 -2125 194 -2107
rect 160 -2141 194 -2125
rect 160 -2193 194 -2179
rect 160 -2213 194 -2193
rect 160 -2261 194 -2251
rect 160 -2285 194 -2261
rect 160 -2329 194 -2323
rect 160 -2357 194 -2329
rect 160 -2397 194 -2395
rect 160 -2429 194 -2397
rect 160 -2499 194 -2467
rect 160 -2501 194 -2499
rect 160 -2567 194 -2539
rect 160 -2573 194 -2567
rect 160 -2635 194 -2611
rect 160 -2645 194 -2635
rect 160 -2703 194 -2683
rect 160 -2717 194 -2703
rect 160 -2771 194 -2755
rect 160 -2789 194 -2771
rect 160 -2839 194 -2827
rect 160 -2861 194 -2839
rect 160 -2907 194 -2899
rect 160 -2933 194 -2907
rect 160 -2975 194 -2971
rect 160 -3005 194 -2975
rect 160 -3077 194 -3043
rect 160 -3145 194 -3115
rect 160 -3149 194 -3145
rect 160 -3213 194 -3187
rect 160 -3221 194 -3213
rect 160 -3281 194 -3259
rect 160 -3293 194 -3281
rect 160 -3349 194 -3331
rect 160 -3365 194 -3349
rect 160 -3417 194 -3403
rect 160 -3437 194 -3417
rect 160 -3485 194 -3475
rect 160 -3509 194 -3485
rect 160 -3553 194 -3547
rect 160 -3581 194 -3553
rect 160 -3621 194 -3619
rect 160 -3653 194 -3621
rect 160 -3723 194 -3691
rect 160 -3725 194 -3723
rect 160 -3791 194 -3763
rect 160 -3797 194 -3791
rect 160 -3859 194 -3835
rect 160 -3869 194 -3859
rect 160 -3927 194 -3907
rect 160 -3941 194 -3927
rect 160 -3995 194 -3979
rect 160 -4013 194 -3995
rect 160 -4063 194 -4051
rect 160 -4085 194 -4063
rect 160 -4131 194 -4123
rect 160 -4157 194 -4131
rect 160 -4199 194 -4195
rect 160 -4229 194 -4199
rect 160 -4301 194 -4267
rect 160 -4369 194 -4339
rect 160 -4373 194 -4369
rect 160 -4437 194 -4411
rect 160 -4445 194 -4437
rect 160 -4505 194 -4483
rect 160 -4517 194 -4505
rect 160 -4573 194 -4555
rect 160 -4589 194 -4573
rect 160 -4641 194 -4627
rect 160 -4661 194 -4641
rect 160 -4709 194 -4699
rect 160 -4733 194 -4709
rect 160 -4777 194 -4771
rect 160 -4805 194 -4777
rect 160 -4845 194 -4843
rect 160 -4877 194 -4845
rect 160 -4947 194 -4915
rect 160 -4949 194 -4947
rect 160 -5015 194 -4987
rect 160 -5021 194 -5015
rect 160 -5083 194 -5059
rect 160 -5093 194 -5083
rect 160 -5151 194 -5131
rect 160 -5165 194 -5151
rect 160 -5219 194 -5203
rect 160 -5237 194 -5219
rect 160 -5287 194 -5275
rect 160 -5309 194 -5287
rect 160 -5355 194 -5347
rect 160 -5381 194 -5355
rect 160 -5423 194 -5419
rect 160 -5453 194 -5423
rect 160 -5525 194 -5491
rect 160 -5593 194 -5563
rect 160 -5597 194 -5593
rect 160 -5661 194 -5635
rect 160 -5669 194 -5661
rect 160 -5729 194 -5707
rect 160 -5741 194 -5729
rect 160 -5797 194 -5779
rect 160 -5813 194 -5797
rect 160 -5865 194 -5851
rect 160 -5885 194 -5865
rect 160 -5933 194 -5923
rect 160 -5957 194 -5933
rect 160 -6001 194 -5995
rect 160 -6029 194 -6001
rect 160 -6069 194 -6067
rect 160 -6101 194 -6069
rect 160 -6171 194 -6139
rect 160 -6173 194 -6171
rect 160 -6239 194 -6211
rect 160 -6245 194 -6239
rect 160 -6307 194 -6283
rect 160 -6317 194 -6307
rect 160 -6375 194 -6355
rect 160 -6389 194 -6375
rect 160 -6443 194 -6427
rect 160 -6461 194 -6443
rect 160 -6511 194 -6499
rect 160 -6533 194 -6511
rect 160 -6579 194 -6571
rect 160 -6605 194 -6579
rect 160 -6647 194 -6643
rect 160 -6677 194 -6647
rect 160 -6749 194 -6715
rect 160 -6817 194 -6787
rect 160 -6821 194 -6817
rect 160 -6885 194 -6859
rect 160 -6893 194 -6885
rect 160 -6953 194 -6931
rect 160 -6965 194 -6953
rect 160 -7021 194 -7003
rect 160 -7037 194 -7021
rect 160 -7089 194 -7075
rect 160 -7109 194 -7089
rect 160 -7157 194 -7147
rect 160 -7181 194 -7157
rect 160 -7225 194 -7219
rect 160 -7253 194 -7225
rect 160 -7293 194 -7291
rect 160 -7325 194 -7293
rect 160 -7395 194 -7363
rect 160 -7397 194 -7395
rect 160 -7463 194 -7435
rect 160 -7469 194 -7463
rect 160 -7531 194 -7507
rect 160 -7541 194 -7531
rect 160 -7599 194 -7579
rect 160 -7613 194 -7599
rect 160 -7667 194 -7651
rect 160 -7685 194 -7667
rect 160 -7735 194 -7723
rect 160 -7757 194 -7735
rect 160 -7803 194 -7795
rect 160 -7829 194 -7803
rect 160 -7871 194 -7867
rect 160 -7901 194 -7871
rect 160 -7973 194 -7939
rect 160 -8041 194 -8011
rect 160 -8045 194 -8041
rect 160 -8109 194 -8083
rect 160 -8117 194 -8109
rect 160 -8177 194 -8155
rect 160 -8189 194 -8177
rect 160 -8245 194 -8227
rect 160 -8261 194 -8245
rect 160 -8313 194 -8299
rect 160 -8333 194 -8313
rect 160 -8381 194 -8371
rect 160 -8405 194 -8381
rect 160 -8449 194 -8443
rect 160 -8477 194 -8449
rect 160 -8517 194 -8515
rect 160 -8549 194 -8517
rect 160 -8619 194 -8587
rect 160 -8621 194 -8619
rect 160 -8687 194 -8659
rect 160 -8693 194 -8687
rect 160 -8755 194 -8731
rect 160 -8765 194 -8755
rect 160 -8823 194 -8803
rect 160 -8837 194 -8823
rect 160 -8891 194 -8875
rect 160 -8909 194 -8891
rect 160 -8959 194 -8947
rect 160 -8981 194 -8959
rect 160 -9027 194 -9019
rect 160 -9053 194 -9027
rect 160 -9095 194 -9091
rect 160 -9125 194 -9095
rect 160 -9197 194 -9163
rect 160 -9265 194 -9235
rect 160 -9269 194 -9265
rect 160 -9333 194 -9307
rect 160 -9341 194 -9333
rect 160 -9401 194 -9379
rect 160 -9413 194 -9401
rect 160 -9469 194 -9451
rect 160 -9485 194 -9469
rect 160 -9537 194 -9523
rect 160 -9557 194 -9537
rect 278 9537 312 9557
rect 278 9523 312 9537
rect 278 9469 312 9485
rect 278 9451 312 9469
rect 278 9401 312 9413
rect 278 9379 312 9401
rect 278 9333 312 9341
rect 278 9307 312 9333
rect 278 9265 312 9269
rect 278 9235 312 9265
rect 278 9163 312 9197
rect 278 9095 312 9125
rect 278 9091 312 9095
rect 278 9027 312 9053
rect 278 9019 312 9027
rect 278 8959 312 8981
rect 278 8947 312 8959
rect 278 8891 312 8909
rect 278 8875 312 8891
rect 278 8823 312 8837
rect 278 8803 312 8823
rect 278 8755 312 8765
rect 278 8731 312 8755
rect 278 8687 312 8693
rect 278 8659 312 8687
rect 278 8619 312 8621
rect 278 8587 312 8619
rect 278 8517 312 8549
rect 278 8515 312 8517
rect 278 8449 312 8477
rect 278 8443 312 8449
rect 278 8381 312 8405
rect 278 8371 312 8381
rect 278 8313 312 8333
rect 278 8299 312 8313
rect 278 8245 312 8261
rect 278 8227 312 8245
rect 278 8177 312 8189
rect 278 8155 312 8177
rect 278 8109 312 8117
rect 278 8083 312 8109
rect 278 8041 312 8045
rect 278 8011 312 8041
rect 278 7939 312 7973
rect 278 7871 312 7901
rect 278 7867 312 7871
rect 278 7803 312 7829
rect 278 7795 312 7803
rect 278 7735 312 7757
rect 278 7723 312 7735
rect 278 7667 312 7685
rect 278 7651 312 7667
rect 278 7599 312 7613
rect 278 7579 312 7599
rect 278 7531 312 7541
rect 278 7507 312 7531
rect 278 7463 312 7469
rect 278 7435 312 7463
rect 278 7395 312 7397
rect 278 7363 312 7395
rect 278 7293 312 7325
rect 278 7291 312 7293
rect 278 7225 312 7253
rect 278 7219 312 7225
rect 278 7157 312 7181
rect 278 7147 312 7157
rect 278 7089 312 7109
rect 278 7075 312 7089
rect 278 7021 312 7037
rect 278 7003 312 7021
rect 278 6953 312 6965
rect 278 6931 312 6953
rect 278 6885 312 6893
rect 278 6859 312 6885
rect 278 6817 312 6821
rect 278 6787 312 6817
rect 278 6715 312 6749
rect 278 6647 312 6677
rect 278 6643 312 6647
rect 278 6579 312 6605
rect 278 6571 312 6579
rect 278 6511 312 6533
rect 278 6499 312 6511
rect 278 6443 312 6461
rect 278 6427 312 6443
rect 278 6375 312 6389
rect 278 6355 312 6375
rect 278 6307 312 6317
rect 278 6283 312 6307
rect 278 6239 312 6245
rect 278 6211 312 6239
rect 278 6171 312 6173
rect 278 6139 312 6171
rect 278 6069 312 6101
rect 278 6067 312 6069
rect 278 6001 312 6029
rect 278 5995 312 6001
rect 278 5933 312 5957
rect 278 5923 312 5933
rect 278 5865 312 5885
rect 278 5851 312 5865
rect 278 5797 312 5813
rect 278 5779 312 5797
rect 278 5729 312 5741
rect 278 5707 312 5729
rect 278 5661 312 5669
rect 278 5635 312 5661
rect 278 5593 312 5597
rect 278 5563 312 5593
rect 278 5491 312 5525
rect 278 5423 312 5453
rect 278 5419 312 5423
rect 278 5355 312 5381
rect 278 5347 312 5355
rect 278 5287 312 5309
rect 278 5275 312 5287
rect 278 5219 312 5237
rect 278 5203 312 5219
rect 278 5151 312 5165
rect 278 5131 312 5151
rect 278 5083 312 5093
rect 278 5059 312 5083
rect 278 5015 312 5021
rect 278 4987 312 5015
rect 278 4947 312 4949
rect 278 4915 312 4947
rect 278 4845 312 4877
rect 278 4843 312 4845
rect 278 4777 312 4805
rect 278 4771 312 4777
rect 278 4709 312 4733
rect 278 4699 312 4709
rect 278 4641 312 4661
rect 278 4627 312 4641
rect 278 4573 312 4589
rect 278 4555 312 4573
rect 278 4505 312 4517
rect 278 4483 312 4505
rect 278 4437 312 4445
rect 278 4411 312 4437
rect 278 4369 312 4373
rect 278 4339 312 4369
rect 278 4267 312 4301
rect 278 4199 312 4229
rect 278 4195 312 4199
rect 278 4131 312 4157
rect 278 4123 312 4131
rect 278 4063 312 4085
rect 278 4051 312 4063
rect 278 3995 312 4013
rect 278 3979 312 3995
rect 278 3927 312 3941
rect 278 3907 312 3927
rect 278 3859 312 3869
rect 278 3835 312 3859
rect 278 3791 312 3797
rect 278 3763 312 3791
rect 278 3723 312 3725
rect 278 3691 312 3723
rect 278 3621 312 3653
rect 278 3619 312 3621
rect 278 3553 312 3581
rect 278 3547 312 3553
rect 278 3485 312 3509
rect 278 3475 312 3485
rect 278 3417 312 3437
rect 278 3403 312 3417
rect 278 3349 312 3365
rect 278 3331 312 3349
rect 278 3281 312 3293
rect 278 3259 312 3281
rect 278 3213 312 3221
rect 278 3187 312 3213
rect 278 3145 312 3149
rect 278 3115 312 3145
rect 278 3043 312 3077
rect 278 2975 312 3005
rect 278 2971 312 2975
rect 278 2907 312 2933
rect 278 2899 312 2907
rect 278 2839 312 2861
rect 278 2827 312 2839
rect 278 2771 312 2789
rect 278 2755 312 2771
rect 278 2703 312 2717
rect 278 2683 312 2703
rect 278 2635 312 2645
rect 278 2611 312 2635
rect 278 2567 312 2573
rect 278 2539 312 2567
rect 278 2499 312 2501
rect 278 2467 312 2499
rect 278 2397 312 2429
rect 278 2395 312 2397
rect 278 2329 312 2357
rect 278 2323 312 2329
rect 278 2261 312 2285
rect 278 2251 312 2261
rect 278 2193 312 2213
rect 278 2179 312 2193
rect 278 2125 312 2141
rect 278 2107 312 2125
rect 278 2057 312 2069
rect 278 2035 312 2057
rect 278 1989 312 1997
rect 278 1963 312 1989
rect 278 1921 312 1925
rect 278 1891 312 1921
rect 278 1819 312 1853
rect 278 1751 312 1781
rect 278 1747 312 1751
rect 278 1683 312 1709
rect 278 1675 312 1683
rect 278 1615 312 1637
rect 278 1603 312 1615
rect 278 1547 312 1565
rect 278 1531 312 1547
rect 278 1479 312 1493
rect 278 1459 312 1479
rect 278 1411 312 1421
rect 278 1387 312 1411
rect 278 1343 312 1349
rect 278 1315 312 1343
rect 278 1275 312 1277
rect 278 1243 312 1275
rect 278 1173 312 1205
rect 278 1171 312 1173
rect 278 1105 312 1133
rect 278 1099 312 1105
rect 278 1037 312 1061
rect 278 1027 312 1037
rect 278 969 312 989
rect 278 955 312 969
rect 278 901 312 917
rect 278 883 312 901
rect 278 833 312 845
rect 278 811 312 833
rect 278 765 312 773
rect 278 739 312 765
rect 278 697 312 701
rect 278 667 312 697
rect 278 595 312 629
rect 278 527 312 557
rect 278 523 312 527
rect 278 459 312 485
rect 278 451 312 459
rect 278 391 312 413
rect 278 379 312 391
rect 278 323 312 341
rect 278 307 312 323
rect 278 255 312 269
rect 278 235 312 255
rect 278 187 312 197
rect 278 163 312 187
rect 278 119 312 125
rect 278 91 312 119
rect 278 51 312 53
rect 278 19 312 51
rect 278 -51 312 -19
rect 278 -53 312 -51
rect 278 -119 312 -91
rect 278 -125 312 -119
rect 278 -187 312 -163
rect 278 -197 312 -187
rect 278 -255 312 -235
rect 278 -269 312 -255
rect 278 -323 312 -307
rect 278 -341 312 -323
rect 278 -391 312 -379
rect 278 -413 312 -391
rect 278 -459 312 -451
rect 278 -485 312 -459
rect 278 -527 312 -523
rect 278 -557 312 -527
rect 278 -629 312 -595
rect 278 -697 312 -667
rect 278 -701 312 -697
rect 278 -765 312 -739
rect 278 -773 312 -765
rect 278 -833 312 -811
rect 278 -845 312 -833
rect 278 -901 312 -883
rect 278 -917 312 -901
rect 278 -969 312 -955
rect 278 -989 312 -969
rect 278 -1037 312 -1027
rect 278 -1061 312 -1037
rect 278 -1105 312 -1099
rect 278 -1133 312 -1105
rect 278 -1173 312 -1171
rect 278 -1205 312 -1173
rect 278 -1275 312 -1243
rect 278 -1277 312 -1275
rect 278 -1343 312 -1315
rect 278 -1349 312 -1343
rect 278 -1411 312 -1387
rect 278 -1421 312 -1411
rect 278 -1479 312 -1459
rect 278 -1493 312 -1479
rect 278 -1547 312 -1531
rect 278 -1565 312 -1547
rect 278 -1615 312 -1603
rect 278 -1637 312 -1615
rect 278 -1683 312 -1675
rect 278 -1709 312 -1683
rect 278 -1751 312 -1747
rect 278 -1781 312 -1751
rect 278 -1853 312 -1819
rect 278 -1921 312 -1891
rect 278 -1925 312 -1921
rect 278 -1989 312 -1963
rect 278 -1997 312 -1989
rect 278 -2057 312 -2035
rect 278 -2069 312 -2057
rect 278 -2125 312 -2107
rect 278 -2141 312 -2125
rect 278 -2193 312 -2179
rect 278 -2213 312 -2193
rect 278 -2261 312 -2251
rect 278 -2285 312 -2261
rect 278 -2329 312 -2323
rect 278 -2357 312 -2329
rect 278 -2397 312 -2395
rect 278 -2429 312 -2397
rect 278 -2499 312 -2467
rect 278 -2501 312 -2499
rect 278 -2567 312 -2539
rect 278 -2573 312 -2567
rect 278 -2635 312 -2611
rect 278 -2645 312 -2635
rect 278 -2703 312 -2683
rect 278 -2717 312 -2703
rect 278 -2771 312 -2755
rect 278 -2789 312 -2771
rect 278 -2839 312 -2827
rect 278 -2861 312 -2839
rect 278 -2907 312 -2899
rect 278 -2933 312 -2907
rect 278 -2975 312 -2971
rect 278 -3005 312 -2975
rect 278 -3077 312 -3043
rect 278 -3145 312 -3115
rect 278 -3149 312 -3145
rect 278 -3213 312 -3187
rect 278 -3221 312 -3213
rect 278 -3281 312 -3259
rect 278 -3293 312 -3281
rect 278 -3349 312 -3331
rect 278 -3365 312 -3349
rect 278 -3417 312 -3403
rect 278 -3437 312 -3417
rect 278 -3485 312 -3475
rect 278 -3509 312 -3485
rect 278 -3553 312 -3547
rect 278 -3581 312 -3553
rect 278 -3621 312 -3619
rect 278 -3653 312 -3621
rect 278 -3723 312 -3691
rect 278 -3725 312 -3723
rect 278 -3791 312 -3763
rect 278 -3797 312 -3791
rect 278 -3859 312 -3835
rect 278 -3869 312 -3859
rect 278 -3927 312 -3907
rect 278 -3941 312 -3927
rect 278 -3995 312 -3979
rect 278 -4013 312 -3995
rect 278 -4063 312 -4051
rect 278 -4085 312 -4063
rect 278 -4131 312 -4123
rect 278 -4157 312 -4131
rect 278 -4199 312 -4195
rect 278 -4229 312 -4199
rect 278 -4301 312 -4267
rect 278 -4369 312 -4339
rect 278 -4373 312 -4369
rect 278 -4437 312 -4411
rect 278 -4445 312 -4437
rect 278 -4505 312 -4483
rect 278 -4517 312 -4505
rect 278 -4573 312 -4555
rect 278 -4589 312 -4573
rect 278 -4641 312 -4627
rect 278 -4661 312 -4641
rect 278 -4709 312 -4699
rect 278 -4733 312 -4709
rect 278 -4777 312 -4771
rect 278 -4805 312 -4777
rect 278 -4845 312 -4843
rect 278 -4877 312 -4845
rect 278 -4947 312 -4915
rect 278 -4949 312 -4947
rect 278 -5015 312 -4987
rect 278 -5021 312 -5015
rect 278 -5083 312 -5059
rect 278 -5093 312 -5083
rect 278 -5151 312 -5131
rect 278 -5165 312 -5151
rect 278 -5219 312 -5203
rect 278 -5237 312 -5219
rect 278 -5287 312 -5275
rect 278 -5309 312 -5287
rect 278 -5355 312 -5347
rect 278 -5381 312 -5355
rect 278 -5423 312 -5419
rect 278 -5453 312 -5423
rect 278 -5525 312 -5491
rect 278 -5593 312 -5563
rect 278 -5597 312 -5593
rect 278 -5661 312 -5635
rect 278 -5669 312 -5661
rect 278 -5729 312 -5707
rect 278 -5741 312 -5729
rect 278 -5797 312 -5779
rect 278 -5813 312 -5797
rect 278 -5865 312 -5851
rect 278 -5885 312 -5865
rect 278 -5933 312 -5923
rect 278 -5957 312 -5933
rect 278 -6001 312 -5995
rect 278 -6029 312 -6001
rect 278 -6069 312 -6067
rect 278 -6101 312 -6069
rect 278 -6171 312 -6139
rect 278 -6173 312 -6171
rect 278 -6239 312 -6211
rect 278 -6245 312 -6239
rect 278 -6307 312 -6283
rect 278 -6317 312 -6307
rect 278 -6375 312 -6355
rect 278 -6389 312 -6375
rect 278 -6443 312 -6427
rect 278 -6461 312 -6443
rect 278 -6511 312 -6499
rect 278 -6533 312 -6511
rect 278 -6579 312 -6571
rect 278 -6605 312 -6579
rect 278 -6647 312 -6643
rect 278 -6677 312 -6647
rect 278 -6749 312 -6715
rect 278 -6817 312 -6787
rect 278 -6821 312 -6817
rect 278 -6885 312 -6859
rect 278 -6893 312 -6885
rect 278 -6953 312 -6931
rect 278 -6965 312 -6953
rect 278 -7021 312 -7003
rect 278 -7037 312 -7021
rect 278 -7089 312 -7075
rect 278 -7109 312 -7089
rect 278 -7157 312 -7147
rect 278 -7181 312 -7157
rect 278 -7225 312 -7219
rect 278 -7253 312 -7225
rect 278 -7293 312 -7291
rect 278 -7325 312 -7293
rect 278 -7395 312 -7363
rect 278 -7397 312 -7395
rect 278 -7463 312 -7435
rect 278 -7469 312 -7463
rect 278 -7531 312 -7507
rect 278 -7541 312 -7531
rect 278 -7599 312 -7579
rect 278 -7613 312 -7599
rect 278 -7667 312 -7651
rect 278 -7685 312 -7667
rect 278 -7735 312 -7723
rect 278 -7757 312 -7735
rect 278 -7803 312 -7795
rect 278 -7829 312 -7803
rect 278 -7871 312 -7867
rect 278 -7901 312 -7871
rect 278 -7973 312 -7939
rect 278 -8041 312 -8011
rect 278 -8045 312 -8041
rect 278 -8109 312 -8083
rect 278 -8117 312 -8109
rect 278 -8177 312 -8155
rect 278 -8189 312 -8177
rect 278 -8245 312 -8227
rect 278 -8261 312 -8245
rect 278 -8313 312 -8299
rect 278 -8333 312 -8313
rect 278 -8381 312 -8371
rect 278 -8405 312 -8381
rect 278 -8449 312 -8443
rect 278 -8477 312 -8449
rect 278 -8517 312 -8515
rect 278 -8549 312 -8517
rect 278 -8619 312 -8587
rect 278 -8621 312 -8619
rect 278 -8687 312 -8659
rect 278 -8693 312 -8687
rect 278 -8755 312 -8731
rect 278 -8765 312 -8755
rect 278 -8823 312 -8803
rect 278 -8837 312 -8823
rect 278 -8891 312 -8875
rect 278 -8909 312 -8891
rect 278 -8959 312 -8947
rect 278 -8981 312 -8959
rect 278 -9027 312 -9019
rect 278 -9053 312 -9027
rect 278 -9095 312 -9091
rect 278 -9125 312 -9095
rect 278 -9197 312 -9163
rect 278 -9265 312 -9235
rect 278 -9269 312 -9265
rect 278 -9333 312 -9307
rect 278 -9341 312 -9333
rect 278 -9401 312 -9379
rect 278 -9413 312 -9401
rect 278 -9469 312 -9451
rect 278 -9485 312 -9469
rect 278 -9537 312 -9523
rect 278 -9557 312 -9537
rect 396 9537 430 9557
rect 396 9523 430 9537
rect 396 9469 430 9485
rect 396 9451 430 9469
rect 396 9401 430 9413
rect 396 9379 430 9401
rect 396 9333 430 9341
rect 396 9307 430 9333
rect 396 9265 430 9269
rect 396 9235 430 9265
rect 396 9163 430 9197
rect 396 9095 430 9125
rect 396 9091 430 9095
rect 396 9027 430 9053
rect 396 9019 430 9027
rect 396 8959 430 8981
rect 396 8947 430 8959
rect 396 8891 430 8909
rect 396 8875 430 8891
rect 396 8823 430 8837
rect 396 8803 430 8823
rect 396 8755 430 8765
rect 396 8731 430 8755
rect 396 8687 430 8693
rect 396 8659 430 8687
rect 396 8619 430 8621
rect 396 8587 430 8619
rect 396 8517 430 8549
rect 396 8515 430 8517
rect 396 8449 430 8477
rect 396 8443 430 8449
rect 396 8381 430 8405
rect 396 8371 430 8381
rect 396 8313 430 8333
rect 396 8299 430 8313
rect 396 8245 430 8261
rect 396 8227 430 8245
rect 396 8177 430 8189
rect 396 8155 430 8177
rect 396 8109 430 8117
rect 396 8083 430 8109
rect 396 8041 430 8045
rect 396 8011 430 8041
rect 396 7939 430 7973
rect 396 7871 430 7901
rect 396 7867 430 7871
rect 396 7803 430 7829
rect 396 7795 430 7803
rect 396 7735 430 7757
rect 396 7723 430 7735
rect 396 7667 430 7685
rect 396 7651 430 7667
rect 396 7599 430 7613
rect 396 7579 430 7599
rect 396 7531 430 7541
rect 396 7507 430 7531
rect 396 7463 430 7469
rect 396 7435 430 7463
rect 396 7395 430 7397
rect 396 7363 430 7395
rect 396 7293 430 7325
rect 396 7291 430 7293
rect 396 7225 430 7253
rect 396 7219 430 7225
rect 396 7157 430 7181
rect 396 7147 430 7157
rect 396 7089 430 7109
rect 396 7075 430 7089
rect 396 7021 430 7037
rect 396 7003 430 7021
rect 396 6953 430 6965
rect 396 6931 430 6953
rect 396 6885 430 6893
rect 396 6859 430 6885
rect 396 6817 430 6821
rect 396 6787 430 6817
rect 396 6715 430 6749
rect 396 6647 430 6677
rect 396 6643 430 6647
rect 396 6579 430 6605
rect 396 6571 430 6579
rect 396 6511 430 6533
rect 396 6499 430 6511
rect 396 6443 430 6461
rect 396 6427 430 6443
rect 396 6375 430 6389
rect 396 6355 430 6375
rect 396 6307 430 6317
rect 396 6283 430 6307
rect 396 6239 430 6245
rect 396 6211 430 6239
rect 396 6171 430 6173
rect 396 6139 430 6171
rect 396 6069 430 6101
rect 396 6067 430 6069
rect 396 6001 430 6029
rect 396 5995 430 6001
rect 396 5933 430 5957
rect 396 5923 430 5933
rect 396 5865 430 5885
rect 396 5851 430 5865
rect 396 5797 430 5813
rect 396 5779 430 5797
rect 396 5729 430 5741
rect 396 5707 430 5729
rect 396 5661 430 5669
rect 396 5635 430 5661
rect 396 5593 430 5597
rect 396 5563 430 5593
rect 396 5491 430 5525
rect 396 5423 430 5453
rect 396 5419 430 5423
rect 396 5355 430 5381
rect 396 5347 430 5355
rect 396 5287 430 5309
rect 396 5275 430 5287
rect 396 5219 430 5237
rect 396 5203 430 5219
rect 396 5151 430 5165
rect 396 5131 430 5151
rect 396 5083 430 5093
rect 396 5059 430 5083
rect 396 5015 430 5021
rect 396 4987 430 5015
rect 396 4947 430 4949
rect 396 4915 430 4947
rect 396 4845 430 4877
rect 396 4843 430 4845
rect 396 4777 430 4805
rect 396 4771 430 4777
rect 396 4709 430 4733
rect 396 4699 430 4709
rect 396 4641 430 4661
rect 396 4627 430 4641
rect 396 4573 430 4589
rect 396 4555 430 4573
rect 396 4505 430 4517
rect 396 4483 430 4505
rect 396 4437 430 4445
rect 396 4411 430 4437
rect 396 4369 430 4373
rect 396 4339 430 4369
rect 396 4267 430 4301
rect 396 4199 430 4229
rect 396 4195 430 4199
rect 396 4131 430 4157
rect 396 4123 430 4131
rect 396 4063 430 4085
rect 396 4051 430 4063
rect 396 3995 430 4013
rect 396 3979 430 3995
rect 396 3927 430 3941
rect 396 3907 430 3927
rect 396 3859 430 3869
rect 396 3835 430 3859
rect 396 3791 430 3797
rect 396 3763 430 3791
rect 396 3723 430 3725
rect 396 3691 430 3723
rect 396 3621 430 3653
rect 396 3619 430 3621
rect 396 3553 430 3581
rect 396 3547 430 3553
rect 396 3485 430 3509
rect 396 3475 430 3485
rect 396 3417 430 3437
rect 396 3403 430 3417
rect 396 3349 430 3365
rect 396 3331 430 3349
rect 396 3281 430 3293
rect 396 3259 430 3281
rect 396 3213 430 3221
rect 396 3187 430 3213
rect 396 3145 430 3149
rect 396 3115 430 3145
rect 396 3043 430 3077
rect 396 2975 430 3005
rect 396 2971 430 2975
rect 396 2907 430 2933
rect 396 2899 430 2907
rect 396 2839 430 2861
rect 396 2827 430 2839
rect 396 2771 430 2789
rect 396 2755 430 2771
rect 396 2703 430 2717
rect 396 2683 430 2703
rect 396 2635 430 2645
rect 396 2611 430 2635
rect 396 2567 430 2573
rect 396 2539 430 2567
rect 396 2499 430 2501
rect 396 2467 430 2499
rect 396 2397 430 2429
rect 396 2395 430 2397
rect 396 2329 430 2357
rect 396 2323 430 2329
rect 396 2261 430 2285
rect 396 2251 430 2261
rect 396 2193 430 2213
rect 396 2179 430 2193
rect 396 2125 430 2141
rect 396 2107 430 2125
rect 396 2057 430 2069
rect 396 2035 430 2057
rect 396 1989 430 1997
rect 396 1963 430 1989
rect 396 1921 430 1925
rect 396 1891 430 1921
rect 396 1819 430 1853
rect 396 1751 430 1781
rect 396 1747 430 1751
rect 396 1683 430 1709
rect 396 1675 430 1683
rect 396 1615 430 1637
rect 396 1603 430 1615
rect 396 1547 430 1565
rect 396 1531 430 1547
rect 396 1479 430 1493
rect 396 1459 430 1479
rect 396 1411 430 1421
rect 396 1387 430 1411
rect 396 1343 430 1349
rect 396 1315 430 1343
rect 396 1275 430 1277
rect 396 1243 430 1275
rect 396 1173 430 1205
rect 396 1171 430 1173
rect 396 1105 430 1133
rect 396 1099 430 1105
rect 396 1037 430 1061
rect 396 1027 430 1037
rect 396 969 430 989
rect 396 955 430 969
rect 396 901 430 917
rect 396 883 430 901
rect 396 833 430 845
rect 396 811 430 833
rect 396 765 430 773
rect 396 739 430 765
rect 396 697 430 701
rect 396 667 430 697
rect 396 595 430 629
rect 396 527 430 557
rect 396 523 430 527
rect 396 459 430 485
rect 396 451 430 459
rect 396 391 430 413
rect 396 379 430 391
rect 396 323 430 341
rect 396 307 430 323
rect 396 255 430 269
rect 396 235 430 255
rect 396 187 430 197
rect 396 163 430 187
rect 396 119 430 125
rect 396 91 430 119
rect 396 51 430 53
rect 396 19 430 51
rect 396 -51 430 -19
rect 396 -53 430 -51
rect 396 -119 430 -91
rect 396 -125 430 -119
rect 396 -187 430 -163
rect 396 -197 430 -187
rect 396 -255 430 -235
rect 396 -269 430 -255
rect 396 -323 430 -307
rect 396 -341 430 -323
rect 396 -391 430 -379
rect 396 -413 430 -391
rect 396 -459 430 -451
rect 396 -485 430 -459
rect 396 -527 430 -523
rect 396 -557 430 -527
rect 396 -629 430 -595
rect 396 -697 430 -667
rect 396 -701 430 -697
rect 396 -765 430 -739
rect 396 -773 430 -765
rect 396 -833 430 -811
rect 396 -845 430 -833
rect 396 -901 430 -883
rect 396 -917 430 -901
rect 396 -969 430 -955
rect 396 -989 430 -969
rect 396 -1037 430 -1027
rect 396 -1061 430 -1037
rect 396 -1105 430 -1099
rect 396 -1133 430 -1105
rect 396 -1173 430 -1171
rect 396 -1205 430 -1173
rect 396 -1275 430 -1243
rect 396 -1277 430 -1275
rect 396 -1343 430 -1315
rect 396 -1349 430 -1343
rect 396 -1411 430 -1387
rect 396 -1421 430 -1411
rect 396 -1479 430 -1459
rect 396 -1493 430 -1479
rect 396 -1547 430 -1531
rect 396 -1565 430 -1547
rect 396 -1615 430 -1603
rect 396 -1637 430 -1615
rect 396 -1683 430 -1675
rect 396 -1709 430 -1683
rect 396 -1751 430 -1747
rect 396 -1781 430 -1751
rect 396 -1853 430 -1819
rect 396 -1921 430 -1891
rect 396 -1925 430 -1921
rect 396 -1989 430 -1963
rect 396 -1997 430 -1989
rect 396 -2057 430 -2035
rect 396 -2069 430 -2057
rect 396 -2125 430 -2107
rect 396 -2141 430 -2125
rect 396 -2193 430 -2179
rect 396 -2213 430 -2193
rect 396 -2261 430 -2251
rect 396 -2285 430 -2261
rect 396 -2329 430 -2323
rect 396 -2357 430 -2329
rect 396 -2397 430 -2395
rect 396 -2429 430 -2397
rect 396 -2499 430 -2467
rect 396 -2501 430 -2499
rect 396 -2567 430 -2539
rect 396 -2573 430 -2567
rect 396 -2635 430 -2611
rect 396 -2645 430 -2635
rect 396 -2703 430 -2683
rect 396 -2717 430 -2703
rect 396 -2771 430 -2755
rect 396 -2789 430 -2771
rect 396 -2839 430 -2827
rect 396 -2861 430 -2839
rect 396 -2907 430 -2899
rect 396 -2933 430 -2907
rect 396 -2975 430 -2971
rect 396 -3005 430 -2975
rect 396 -3077 430 -3043
rect 396 -3145 430 -3115
rect 396 -3149 430 -3145
rect 396 -3213 430 -3187
rect 396 -3221 430 -3213
rect 396 -3281 430 -3259
rect 396 -3293 430 -3281
rect 396 -3349 430 -3331
rect 396 -3365 430 -3349
rect 396 -3417 430 -3403
rect 396 -3437 430 -3417
rect 396 -3485 430 -3475
rect 396 -3509 430 -3485
rect 396 -3553 430 -3547
rect 396 -3581 430 -3553
rect 396 -3621 430 -3619
rect 396 -3653 430 -3621
rect 396 -3723 430 -3691
rect 396 -3725 430 -3723
rect 396 -3791 430 -3763
rect 396 -3797 430 -3791
rect 396 -3859 430 -3835
rect 396 -3869 430 -3859
rect 396 -3927 430 -3907
rect 396 -3941 430 -3927
rect 396 -3995 430 -3979
rect 396 -4013 430 -3995
rect 396 -4063 430 -4051
rect 396 -4085 430 -4063
rect 396 -4131 430 -4123
rect 396 -4157 430 -4131
rect 396 -4199 430 -4195
rect 396 -4229 430 -4199
rect 396 -4301 430 -4267
rect 396 -4369 430 -4339
rect 396 -4373 430 -4369
rect 396 -4437 430 -4411
rect 396 -4445 430 -4437
rect 396 -4505 430 -4483
rect 396 -4517 430 -4505
rect 396 -4573 430 -4555
rect 396 -4589 430 -4573
rect 396 -4641 430 -4627
rect 396 -4661 430 -4641
rect 396 -4709 430 -4699
rect 396 -4733 430 -4709
rect 396 -4777 430 -4771
rect 396 -4805 430 -4777
rect 396 -4845 430 -4843
rect 396 -4877 430 -4845
rect 396 -4947 430 -4915
rect 396 -4949 430 -4947
rect 396 -5015 430 -4987
rect 396 -5021 430 -5015
rect 396 -5083 430 -5059
rect 396 -5093 430 -5083
rect 396 -5151 430 -5131
rect 396 -5165 430 -5151
rect 396 -5219 430 -5203
rect 396 -5237 430 -5219
rect 396 -5287 430 -5275
rect 396 -5309 430 -5287
rect 396 -5355 430 -5347
rect 396 -5381 430 -5355
rect 396 -5423 430 -5419
rect 396 -5453 430 -5423
rect 396 -5525 430 -5491
rect 396 -5593 430 -5563
rect 396 -5597 430 -5593
rect 396 -5661 430 -5635
rect 396 -5669 430 -5661
rect 396 -5729 430 -5707
rect 396 -5741 430 -5729
rect 396 -5797 430 -5779
rect 396 -5813 430 -5797
rect 396 -5865 430 -5851
rect 396 -5885 430 -5865
rect 396 -5933 430 -5923
rect 396 -5957 430 -5933
rect 396 -6001 430 -5995
rect 396 -6029 430 -6001
rect 396 -6069 430 -6067
rect 396 -6101 430 -6069
rect 396 -6171 430 -6139
rect 396 -6173 430 -6171
rect 396 -6239 430 -6211
rect 396 -6245 430 -6239
rect 396 -6307 430 -6283
rect 396 -6317 430 -6307
rect 396 -6375 430 -6355
rect 396 -6389 430 -6375
rect 396 -6443 430 -6427
rect 396 -6461 430 -6443
rect 396 -6511 430 -6499
rect 396 -6533 430 -6511
rect 396 -6579 430 -6571
rect 396 -6605 430 -6579
rect 396 -6647 430 -6643
rect 396 -6677 430 -6647
rect 396 -6749 430 -6715
rect 396 -6817 430 -6787
rect 396 -6821 430 -6817
rect 396 -6885 430 -6859
rect 396 -6893 430 -6885
rect 396 -6953 430 -6931
rect 396 -6965 430 -6953
rect 396 -7021 430 -7003
rect 396 -7037 430 -7021
rect 396 -7089 430 -7075
rect 396 -7109 430 -7089
rect 396 -7157 430 -7147
rect 396 -7181 430 -7157
rect 396 -7225 430 -7219
rect 396 -7253 430 -7225
rect 396 -7293 430 -7291
rect 396 -7325 430 -7293
rect 396 -7395 430 -7363
rect 396 -7397 430 -7395
rect 396 -7463 430 -7435
rect 396 -7469 430 -7463
rect 396 -7531 430 -7507
rect 396 -7541 430 -7531
rect 396 -7599 430 -7579
rect 396 -7613 430 -7599
rect 396 -7667 430 -7651
rect 396 -7685 430 -7667
rect 396 -7735 430 -7723
rect 396 -7757 430 -7735
rect 396 -7803 430 -7795
rect 396 -7829 430 -7803
rect 396 -7871 430 -7867
rect 396 -7901 430 -7871
rect 396 -7973 430 -7939
rect 396 -8041 430 -8011
rect 396 -8045 430 -8041
rect 396 -8109 430 -8083
rect 396 -8117 430 -8109
rect 396 -8177 430 -8155
rect 396 -8189 430 -8177
rect 396 -8245 430 -8227
rect 396 -8261 430 -8245
rect 396 -8313 430 -8299
rect 396 -8333 430 -8313
rect 396 -8381 430 -8371
rect 396 -8405 430 -8381
rect 396 -8449 430 -8443
rect 396 -8477 430 -8449
rect 396 -8517 430 -8515
rect 396 -8549 430 -8517
rect 396 -8619 430 -8587
rect 396 -8621 430 -8619
rect 396 -8687 430 -8659
rect 396 -8693 430 -8687
rect 396 -8755 430 -8731
rect 396 -8765 430 -8755
rect 396 -8823 430 -8803
rect 396 -8837 430 -8823
rect 396 -8891 430 -8875
rect 396 -8909 430 -8891
rect 396 -8959 430 -8947
rect 396 -8981 430 -8959
rect 396 -9027 430 -9019
rect 396 -9053 430 -9027
rect 396 -9095 430 -9091
rect 396 -9125 430 -9095
rect 396 -9197 430 -9163
rect 396 -9265 430 -9235
rect 396 -9269 430 -9265
rect 396 -9333 430 -9307
rect 396 -9341 430 -9333
rect 396 -9401 430 -9379
rect 396 -9413 430 -9401
rect 396 -9469 430 -9451
rect 396 -9485 430 -9469
rect 396 -9537 430 -9523
rect 396 -9557 430 -9537
rect 514 9537 548 9557
rect 514 9523 548 9537
rect 514 9469 548 9485
rect 514 9451 548 9469
rect 514 9401 548 9413
rect 514 9379 548 9401
rect 514 9333 548 9341
rect 514 9307 548 9333
rect 514 9265 548 9269
rect 514 9235 548 9265
rect 514 9163 548 9197
rect 514 9095 548 9125
rect 514 9091 548 9095
rect 514 9027 548 9053
rect 514 9019 548 9027
rect 514 8959 548 8981
rect 514 8947 548 8959
rect 514 8891 548 8909
rect 514 8875 548 8891
rect 514 8823 548 8837
rect 514 8803 548 8823
rect 514 8755 548 8765
rect 514 8731 548 8755
rect 514 8687 548 8693
rect 514 8659 548 8687
rect 514 8619 548 8621
rect 514 8587 548 8619
rect 514 8517 548 8549
rect 514 8515 548 8517
rect 514 8449 548 8477
rect 514 8443 548 8449
rect 514 8381 548 8405
rect 514 8371 548 8381
rect 514 8313 548 8333
rect 514 8299 548 8313
rect 514 8245 548 8261
rect 514 8227 548 8245
rect 514 8177 548 8189
rect 514 8155 548 8177
rect 514 8109 548 8117
rect 514 8083 548 8109
rect 514 8041 548 8045
rect 514 8011 548 8041
rect 514 7939 548 7973
rect 514 7871 548 7901
rect 514 7867 548 7871
rect 514 7803 548 7829
rect 514 7795 548 7803
rect 514 7735 548 7757
rect 514 7723 548 7735
rect 514 7667 548 7685
rect 514 7651 548 7667
rect 514 7599 548 7613
rect 514 7579 548 7599
rect 514 7531 548 7541
rect 514 7507 548 7531
rect 514 7463 548 7469
rect 514 7435 548 7463
rect 514 7395 548 7397
rect 514 7363 548 7395
rect 514 7293 548 7325
rect 514 7291 548 7293
rect 514 7225 548 7253
rect 514 7219 548 7225
rect 514 7157 548 7181
rect 514 7147 548 7157
rect 514 7089 548 7109
rect 514 7075 548 7089
rect 514 7021 548 7037
rect 514 7003 548 7021
rect 514 6953 548 6965
rect 514 6931 548 6953
rect 514 6885 548 6893
rect 514 6859 548 6885
rect 514 6817 548 6821
rect 514 6787 548 6817
rect 514 6715 548 6749
rect 514 6647 548 6677
rect 514 6643 548 6647
rect 514 6579 548 6605
rect 514 6571 548 6579
rect 514 6511 548 6533
rect 514 6499 548 6511
rect 514 6443 548 6461
rect 514 6427 548 6443
rect 514 6375 548 6389
rect 514 6355 548 6375
rect 514 6307 548 6317
rect 514 6283 548 6307
rect 514 6239 548 6245
rect 514 6211 548 6239
rect 514 6171 548 6173
rect 514 6139 548 6171
rect 514 6069 548 6101
rect 514 6067 548 6069
rect 514 6001 548 6029
rect 514 5995 548 6001
rect 514 5933 548 5957
rect 514 5923 548 5933
rect 514 5865 548 5885
rect 514 5851 548 5865
rect 514 5797 548 5813
rect 514 5779 548 5797
rect 514 5729 548 5741
rect 514 5707 548 5729
rect 514 5661 548 5669
rect 514 5635 548 5661
rect 514 5593 548 5597
rect 514 5563 548 5593
rect 514 5491 548 5525
rect 514 5423 548 5453
rect 514 5419 548 5423
rect 514 5355 548 5381
rect 514 5347 548 5355
rect 514 5287 548 5309
rect 514 5275 548 5287
rect 514 5219 548 5237
rect 514 5203 548 5219
rect 514 5151 548 5165
rect 514 5131 548 5151
rect 514 5083 548 5093
rect 514 5059 548 5083
rect 514 5015 548 5021
rect 514 4987 548 5015
rect 514 4947 548 4949
rect 514 4915 548 4947
rect 514 4845 548 4877
rect 514 4843 548 4845
rect 514 4777 548 4805
rect 514 4771 548 4777
rect 514 4709 548 4733
rect 514 4699 548 4709
rect 514 4641 548 4661
rect 514 4627 548 4641
rect 514 4573 548 4589
rect 514 4555 548 4573
rect 514 4505 548 4517
rect 514 4483 548 4505
rect 514 4437 548 4445
rect 514 4411 548 4437
rect 514 4369 548 4373
rect 514 4339 548 4369
rect 514 4267 548 4301
rect 514 4199 548 4229
rect 514 4195 548 4199
rect 514 4131 548 4157
rect 514 4123 548 4131
rect 514 4063 548 4085
rect 514 4051 548 4063
rect 514 3995 548 4013
rect 514 3979 548 3995
rect 514 3927 548 3941
rect 514 3907 548 3927
rect 514 3859 548 3869
rect 514 3835 548 3859
rect 514 3791 548 3797
rect 514 3763 548 3791
rect 514 3723 548 3725
rect 514 3691 548 3723
rect 514 3621 548 3653
rect 514 3619 548 3621
rect 514 3553 548 3581
rect 514 3547 548 3553
rect 514 3485 548 3509
rect 514 3475 548 3485
rect 514 3417 548 3437
rect 514 3403 548 3417
rect 514 3349 548 3365
rect 514 3331 548 3349
rect 514 3281 548 3293
rect 514 3259 548 3281
rect 514 3213 548 3221
rect 514 3187 548 3213
rect 514 3145 548 3149
rect 514 3115 548 3145
rect 514 3043 548 3077
rect 514 2975 548 3005
rect 514 2971 548 2975
rect 514 2907 548 2933
rect 514 2899 548 2907
rect 514 2839 548 2861
rect 514 2827 548 2839
rect 514 2771 548 2789
rect 514 2755 548 2771
rect 514 2703 548 2717
rect 514 2683 548 2703
rect 514 2635 548 2645
rect 514 2611 548 2635
rect 514 2567 548 2573
rect 514 2539 548 2567
rect 514 2499 548 2501
rect 514 2467 548 2499
rect 514 2397 548 2429
rect 514 2395 548 2397
rect 514 2329 548 2357
rect 514 2323 548 2329
rect 514 2261 548 2285
rect 514 2251 548 2261
rect 514 2193 548 2213
rect 514 2179 548 2193
rect 514 2125 548 2141
rect 514 2107 548 2125
rect 514 2057 548 2069
rect 514 2035 548 2057
rect 514 1989 548 1997
rect 514 1963 548 1989
rect 514 1921 548 1925
rect 514 1891 548 1921
rect 514 1819 548 1853
rect 514 1751 548 1781
rect 514 1747 548 1751
rect 514 1683 548 1709
rect 514 1675 548 1683
rect 514 1615 548 1637
rect 514 1603 548 1615
rect 514 1547 548 1565
rect 514 1531 548 1547
rect 514 1479 548 1493
rect 514 1459 548 1479
rect 514 1411 548 1421
rect 514 1387 548 1411
rect 514 1343 548 1349
rect 514 1315 548 1343
rect 514 1275 548 1277
rect 514 1243 548 1275
rect 514 1173 548 1205
rect 514 1171 548 1173
rect 514 1105 548 1133
rect 514 1099 548 1105
rect 514 1037 548 1061
rect 514 1027 548 1037
rect 514 969 548 989
rect 514 955 548 969
rect 514 901 548 917
rect 514 883 548 901
rect 514 833 548 845
rect 514 811 548 833
rect 514 765 548 773
rect 514 739 548 765
rect 514 697 548 701
rect 514 667 548 697
rect 514 595 548 629
rect 514 527 548 557
rect 514 523 548 527
rect 514 459 548 485
rect 514 451 548 459
rect 514 391 548 413
rect 514 379 548 391
rect 514 323 548 341
rect 514 307 548 323
rect 514 255 548 269
rect 514 235 548 255
rect 514 187 548 197
rect 514 163 548 187
rect 514 119 548 125
rect 514 91 548 119
rect 514 51 548 53
rect 514 19 548 51
rect 514 -51 548 -19
rect 514 -53 548 -51
rect 514 -119 548 -91
rect 514 -125 548 -119
rect 514 -187 548 -163
rect 514 -197 548 -187
rect 514 -255 548 -235
rect 514 -269 548 -255
rect 514 -323 548 -307
rect 514 -341 548 -323
rect 514 -391 548 -379
rect 514 -413 548 -391
rect 514 -459 548 -451
rect 514 -485 548 -459
rect 514 -527 548 -523
rect 514 -557 548 -527
rect 514 -629 548 -595
rect 514 -697 548 -667
rect 514 -701 548 -697
rect 514 -765 548 -739
rect 514 -773 548 -765
rect 514 -833 548 -811
rect 514 -845 548 -833
rect 514 -901 548 -883
rect 514 -917 548 -901
rect 514 -969 548 -955
rect 514 -989 548 -969
rect 514 -1037 548 -1027
rect 514 -1061 548 -1037
rect 514 -1105 548 -1099
rect 514 -1133 548 -1105
rect 514 -1173 548 -1171
rect 514 -1205 548 -1173
rect 514 -1275 548 -1243
rect 514 -1277 548 -1275
rect 514 -1343 548 -1315
rect 514 -1349 548 -1343
rect 514 -1411 548 -1387
rect 514 -1421 548 -1411
rect 514 -1479 548 -1459
rect 514 -1493 548 -1479
rect 514 -1547 548 -1531
rect 514 -1565 548 -1547
rect 514 -1615 548 -1603
rect 514 -1637 548 -1615
rect 514 -1683 548 -1675
rect 514 -1709 548 -1683
rect 514 -1751 548 -1747
rect 514 -1781 548 -1751
rect 514 -1853 548 -1819
rect 514 -1921 548 -1891
rect 514 -1925 548 -1921
rect 514 -1989 548 -1963
rect 514 -1997 548 -1989
rect 514 -2057 548 -2035
rect 514 -2069 548 -2057
rect 514 -2125 548 -2107
rect 514 -2141 548 -2125
rect 514 -2193 548 -2179
rect 514 -2213 548 -2193
rect 514 -2261 548 -2251
rect 514 -2285 548 -2261
rect 514 -2329 548 -2323
rect 514 -2357 548 -2329
rect 514 -2397 548 -2395
rect 514 -2429 548 -2397
rect 514 -2499 548 -2467
rect 514 -2501 548 -2499
rect 514 -2567 548 -2539
rect 514 -2573 548 -2567
rect 514 -2635 548 -2611
rect 514 -2645 548 -2635
rect 514 -2703 548 -2683
rect 514 -2717 548 -2703
rect 514 -2771 548 -2755
rect 514 -2789 548 -2771
rect 514 -2839 548 -2827
rect 514 -2861 548 -2839
rect 514 -2907 548 -2899
rect 514 -2933 548 -2907
rect 514 -2975 548 -2971
rect 514 -3005 548 -2975
rect 514 -3077 548 -3043
rect 514 -3145 548 -3115
rect 514 -3149 548 -3145
rect 514 -3213 548 -3187
rect 514 -3221 548 -3213
rect 514 -3281 548 -3259
rect 514 -3293 548 -3281
rect 514 -3349 548 -3331
rect 514 -3365 548 -3349
rect 514 -3417 548 -3403
rect 514 -3437 548 -3417
rect 514 -3485 548 -3475
rect 514 -3509 548 -3485
rect 514 -3553 548 -3547
rect 514 -3581 548 -3553
rect 514 -3621 548 -3619
rect 514 -3653 548 -3621
rect 514 -3723 548 -3691
rect 514 -3725 548 -3723
rect 514 -3791 548 -3763
rect 514 -3797 548 -3791
rect 514 -3859 548 -3835
rect 514 -3869 548 -3859
rect 514 -3927 548 -3907
rect 514 -3941 548 -3927
rect 514 -3995 548 -3979
rect 514 -4013 548 -3995
rect 514 -4063 548 -4051
rect 514 -4085 548 -4063
rect 514 -4131 548 -4123
rect 514 -4157 548 -4131
rect 514 -4199 548 -4195
rect 514 -4229 548 -4199
rect 514 -4301 548 -4267
rect 514 -4369 548 -4339
rect 514 -4373 548 -4369
rect 514 -4437 548 -4411
rect 514 -4445 548 -4437
rect 514 -4505 548 -4483
rect 514 -4517 548 -4505
rect 514 -4573 548 -4555
rect 514 -4589 548 -4573
rect 514 -4641 548 -4627
rect 514 -4661 548 -4641
rect 514 -4709 548 -4699
rect 514 -4733 548 -4709
rect 514 -4777 548 -4771
rect 514 -4805 548 -4777
rect 514 -4845 548 -4843
rect 514 -4877 548 -4845
rect 514 -4947 548 -4915
rect 514 -4949 548 -4947
rect 514 -5015 548 -4987
rect 514 -5021 548 -5015
rect 514 -5083 548 -5059
rect 514 -5093 548 -5083
rect 514 -5151 548 -5131
rect 514 -5165 548 -5151
rect 514 -5219 548 -5203
rect 514 -5237 548 -5219
rect 514 -5287 548 -5275
rect 514 -5309 548 -5287
rect 514 -5355 548 -5347
rect 514 -5381 548 -5355
rect 514 -5423 548 -5419
rect 514 -5453 548 -5423
rect 514 -5525 548 -5491
rect 514 -5593 548 -5563
rect 514 -5597 548 -5593
rect 514 -5661 548 -5635
rect 514 -5669 548 -5661
rect 514 -5729 548 -5707
rect 514 -5741 548 -5729
rect 514 -5797 548 -5779
rect 514 -5813 548 -5797
rect 514 -5865 548 -5851
rect 514 -5885 548 -5865
rect 514 -5933 548 -5923
rect 514 -5957 548 -5933
rect 514 -6001 548 -5995
rect 514 -6029 548 -6001
rect 514 -6069 548 -6067
rect 514 -6101 548 -6069
rect 514 -6171 548 -6139
rect 514 -6173 548 -6171
rect 514 -6239 548 -6211
rect 514 -6245 548 -6239
rect 514 -6307 548 -6283
rect 514 -6317 548 -6307
rect 514 -6375 548 -6355
rect 514 -6389 548 -6375
rect 514 -6443 548 -6427
rect 514 -6461 548 -6443
rect 514 -6511 548 -6499
rect 514 -6533 548 -6511
rect 514 -6579 548 -6571
rect 514 -6605 548 -6579
rect 514 -6647 548 -6643
rect 514 -6677 548 -6647
rect 514 -6749 548 -6715
rect 514 -6817 548 -6787
rect 514 -6821 548 -6817
rect 514 -6885 548 -6859
rect 514 -6893 548 -6885
rect 514 -6953 548 -6931
rect 514 -6965 548 -6953
rect 514 -7021 548 -7003
rect 514 -7037 548 -7021
rect 514 -7089 548 -7075
rect 514 -7109 548 -7089
rect 514 -7157 548 -7147
rect 514 -7181 548 -7157
rect 514 -7225 548 -7219
rect 514 -7253 548 -7225
rect 514 -7293 548 -7291
rect 514 -7325 548 -7293
rect 514 -7395 548 -7363
rect 514 -7397 548 -7395
rect 514 -7463 548 -7435
rect 514 -7469 548 -7463
rect 514 -7531 548 -7507
rect 514 -7541 548 -7531
rect 514 -7599 548 -7579
rect 514 -7613 548 -7599
rect 514 -7667 548 -7651
rect 514 -7685 548 -7667
rect 514 -7735 548 -7723
rect 514 -7757 548 -7735
rect 514 -7803 548 -7795
rect 514 -7829 548 -7803
rect 514 -7871 548 -7867
rect 514 -7901 548 -7871
rect 514 -7973 548 -7939
rect 514 -8041 548 -8011
rect 514 -8045 548 -8041
rect 514 -8109 548 -8083
rect 514 -8117 548 -8109
rect 514 -8177 548 -8155
rect 514 -8189 548 -8177
rect 514 -8245 548 -8227
rect 514 -8261 548 -8245
rect 514 -8313 548 -8299
rect 514 -8333 548 -8313
rect 514 -8381 548 -8371
rect 514 -8405 548 -8381
rect 514 -8449 548 -8443
rect 514 -8477 548 -8449
rect 514 -8517 548 -8515
rect 514 -8549 548 -8517
rect 514 -8619 548 -8587
rect 514 -8621 548 -8619
rect 514 -8687 548 -8659
rect 514 -8693 548 -8687
rect 514 -8755 548 -8731
rect 514 -8765 548 -8755
rect 514 -8823 548 -8803
rect 514 -8837 548 -8823
rect 514 -8891 548 -8875
rect 514 -8909 548 -8891
rect 514 -8959 548 -8947
rect 514 -8981 548 -8959
rect 514 -9027 548 -9019
rect 514 -9053 548 -9027
rect 514 -9095 548 -9091
rect 514 -9125 548 -9095
rect 514 -9197 548 -9163
rect 514 -9265 548 -9235
rect 514 -9269 548 -9265
rect 514 -9333 548 -9307
rect 514 -9341 548 -9333
rect 514 -9401 548 -9379
rect 514 -9413 548 -9401
rect 514 -9469 548 -9451
rect 514 -9485 548 -9469
rect 514 -9537 548 -9523
rect 514 -9557 548 -9537
rect 632 9537 666 9557
rect 632 9523 666 9537
rect 632 9469 666 9485
rect 632 9451 666 9469
rect 632 9401 666 9413
rect 632 9379 666 9401
rect 632 9333 666 9341
rect 632 9307 666 9333
rect 632 9265 666 9269
rect 632 9235 666 9265
rect 632 9163 666 9197
rect 632 9095 666 9125
rect 632 9091 666 9095
rect 632 9027 666 9053
rect 632 9019 666 9027
rect 632 8959 666 8981
rect 632 8947 666 8959
rect 632 8891 666 8909
rect 632 8875 666 8891
rect 632 8823 666 8837
rect 632 8803 666 8823
rect 632 8755 666 8765
rect 632 8731 666 8755
rect 632 8687 666 8693
rect 632 8659 666 8687
rect 632 8619 666 8621
rect 632 8587 666 8619
rect 632 8517 666 8549
rect 632 8515 666 8517
rect 632 8449 666 8477
rect 632 8443 666 8449
rect 632 8381 666 8405
rect 632 8371 666 8381
rect 632 8313 666 8333
rect 632 8299 666 8313
rect 632 8245 666 8261
rect 632 8227 666 8245
rect 632 8177 666 8189
rect 632 8155 666 8177
rect 632 8109 666 8117
rect 632 8083 666 8109
rect 632 8041 666 8045
rect 632 8011 666 8041
rect 632 7939 666 7973
rect 632 7871 666 7901
rect 632 7867 666 7871
rect 632 7803 666 7829
rect 632 7795 666 7803
rect 632 7735 666 7757
rect 632 7723 666 7735
rect 632 7667 666 7685
rect 632 7651 666 7667
rect 632 7599 666 7613
rect 632 7579 666 7599
rect 632 7531 666 7541
rect 632 7507 666 7531
rect 632 7463 666 7469
rect 632 7435 666 7463
rect 632 7395 666 7397
rect 632 7363 666 7395
rect 632 7293 666 7325
rect 632 7291 666 7293
rect 632 7225 666 7253
rect 632 7219 666 7225
rect 632 7157 666 7181
rect 632 7147 666 7157
rect 632 7089 666 7109
rect 632 7075 666 7089
rect 632 7021 666 7037
rect 632 7003 666 7021
rect 632 6953 666 6965
rect 632 6931 666 6953
rect 632 6885 666 6893
rect 632 6859 666 6885
rect 632 6817 666 6821
rect 632 6787 666 6817
rect 632 6715 666 6749
rect 632 6647 666 6677
rect 632 6643 666 6647
rect 632 6579 666 6605
rect 632 6571 666 6579
rect 632 6511 666 6533
rect 632 6499 666 6511
rect 632 6443 666 6461
rect 632 6427 666 6443
rect 632 6375 666 6389
rect 632 6355 666 6375
rect 632 6307 666 6317
rect 632 6283 666 6307
rect 632 6239 666 6245
rect 632 6211 666 6239
rect 632 6171 666 6173
rect 632 6139 666 6171
rect 632 6069 666 6101
rect 632 6067 666 6069
rect 632 6001 666 6029
rect 632 5995 666 6001
rect 632 5933 666 5957
rect 632 5923 666 5933
rect 632 5865 666 5885
rect 632 5851 666 5865
rect 632 5797 666 5813
rect 632 5779 666 5797
rect 632 5729 666 5741
rect 632 5707 666 5729
rect 632 5661 666 5669
rect 632 5635 666 5661
rect 632 5593 666 5597
rect 632 5563 666 5593
rect 632 5491 666 5525
rect 632 5423 666 5453
rect 632 5419 666 5423
rect 632 5355 666 5381
rect 632 5347 666 5355
rect 632 5287 666 5309
rect 632 5275 666 5287
rect 632 5219 666 5237
rect 632 5203 666 5219
rect 632 5151 666 5165
rect 632 5131 666 5151
rect 632 5083 666 5093
rect 632 5059 666 5083
rect 632 5015 666 5021
rect 632 4987 666 5015
rect 632 4947 666 4949
rect 632 4915 666 4947
rect 632 4845 666 4877
rect 632 4843 666 4845
rect 632 4777 666 4805
rect 632 4771 666 4777
rect 632 4709 666 4733
rect 632 4699 666 4709
rect 632 4641 666 4661
rect 632 4627 666 4641
rect 632 4573 666 4589
rect 632 4555 666 4573
rect 632 4505 666 4517
rect 632 4483 666 4505
rect 632 4437 666 4445
rect 632 4411 666 4437
rect 632 4369 666 4373
rect 632 4339 666 4369
rect 632 4267 666 4301
rect 632 4199 666 4229
rect 632 4195 666 4199
rect 632 4131 666 4157
rect 632 4123 666 4131
rect 632 4063 666 4085
rect 632 4051 666 4063
rect 632 3995 666 4013
rect 632 3979 666 3995
rect 632 3927 666 3941
rect 632 3907 666 3927
rect 632 3859 666 3869
rect 632 3835 666 3859
rect 632 3791 666 3797
rect 632 3763 666 3791
rect 632 3723 666 3725
rect 632 3691 666 3723
rect 632 3621 666 3653
rect 632 3619 666 3621
rect 632 3553 666 3581
rect 632 3547 666 3553
rect 632 3485 666 3509
rect 632 3475 666 3485
rect 632 3417 666 3437
rect 632 3403 666 3417
rect 632 3349 666 3365
rect 632 3331 666 3349
rect 632 3281 666 3293
rect 632 3259 666 3281
rect 632 3213 666 3221
rect 632 3187 666 3213
rect 632 3145 666 3149
rect 632 3115 666 3145
rect 632 3043 666 3077
rect 632 2975 666 3005
rect 632 2971 666 2975
rect 632 2907 666 2933
rect 632 2899 666 2907
rect 632 2839 666 2861
rect 632 2827 666 2839
rect 632 2771 666 2789
rect 632 2755 666 2771
rect 632 2703 666 2717
rect 632 2683 666 2703
rect 632 2635 666 2645
rect 632 2611 666 2635
rect 632 2567 666 2573
rect 632 2539 666 2567
rect 632 2499 666 2501
rect 632 2467 666 2499
rect 632 2397 666 2429
rect 632 2395 666 2397
rect 632 2329 666 2357
rect 632 2323 666 2329
rect 632 2261 666 2285
rect 632 2251 666 2261
rect 632 2193 666 2213
rect 632 2179 666 2193
rect 632 2125 666 2141
rect 632 2107 666 2125
rect 632 2057 666 2069
rect 632 2035 666 2057
rect 632 1989 666 1997
rect 632 1963 666 1989
rect 632 1921 666 1925
rect 632 1891 666 1921
rect 632 1819 666 1853
rect 632 1751 666 1781
rect 632 1747 666 1751
rect 632 1683 666 1709
rect 632 1675 666 1683
rect 632 1615 666 1637
rect 632 1603 666 1615
rect 632 1547 666 1565
rect 632 1531 666 1547
rect 632 1479 666 1493
rect 632 1459 666 1479
rect 632 1411 666 1421
rect 632 1387 666 1411
rect 632 1343 666 1349
rect 632 1315 666 1343
rect 632 1275 666 1277
rect 632 1243 666 1275
rect 632 1173 666 1205
rect 632 1171 666 1173
rect 632 1105 666 1133
rect 632 1099 666 1105
rect 632 1037 666 1061
rect 632 1027 666 1037
rect 632 969 666 989
rect 632 955 666 969
rect 632 901 666 917
rect 632 883 666 901
rect 632 833 666 845
rect 632 811 666 833
rect 632 765 666 773
rect 632 739 666 765
rect 632 697 666 701
rect 632 667 666 697
rect 632 595 666 629
rect 632 527 666 557
rect 632 523 666 527
rect 632 459 666 485
rect 632 451 666 459
rect 632 391 666 413
rect 632 379 666 391
rect 632 323 666 341
rect 632 307 666 323
rect 632 255 666 269
rect 632 235 666 255
rect 632 187 666 197
rect 632 163 666 187
rect 632 119 666 125
rect 632 91 666 119
rect 632 51 666 53
rect 632 19 666 51
rect 632 -51 666 -19
rect 632 -53 666 -51
rect 632 -119 666 -91
rect 632 -125 666 -119
rect 632 -187 666 -163
rect 632 -197 666 -187
rect 632 -255 666 -235
rect 632 -269 666 -255
rect 632 -323 666 -307
rect 632 -341 666 -323
rect 632 -391 666 -379
rect 632 -413 666 -391
rect 632 -459 666 -451
rect 632 -485 666 -459
rect 632 -527 666 -523
rect 632 -557 666 -527
rect 632 -629 666 -595
rect 632 -697 666 -667
rect 632 -701 666 -697
rect 632 -765 666 -739
rect 632 -773 666 -765
rect 632 -833 666 -811
rect 632 -845 666 -833
rect 632 -901 666 -883
rect 632 -917 666 -901
rect 632 -969 666 -955
rect 632 -989 666 -969
rect 632 -1037 666 -1027
rect 632 -1061 666 -1037
rect 632 -1105 666 -1099
rect 632 -1133 666 -1105
rect 632 -1173 666 -1171
rect 632 -1205 666 -1173
rect 632 -1275 666 -1243
rect 632 -1277 666 -1275
rect 632 -1343 666 -1315
rect 632 -1349 666 -1343
rect 632 -1411 666 -1387
rect 632 -1421 666 -1411
rect 632 -1479 666 -1459
rect 632 -1493 666 -1479
rect 632 -1547 666 -1531
rect 632 -1565 666 -1547
rect 632 -1615 666 -1603
rect 632 -1637 666 -1615
rect 632 -1683 666 -1675
rect 632 -1709 666 -1683
rect 632 -1751 666 -1747
rect 632 -1781 666 -1751
rect 632 -1853 666 -1819
rect 632 -1921 666 -1891
rect 632 -1925 666 -1921
rect 632 -1989 666 -1963
rect 632 -1997 666 -1989
rect 632 -2057 666 -2035
rect 632 -2069 666 -2057
rect 632 -2125 666 -2107
rect 632 -2141 666 -2125
rect 632 -2193 666 -2179
rect 632 -2213 666 -2193
rect 632 -2261 666 -2251
rect 632 -2285 666 -2261
rect 632 -2329 666 -2323
rect 632 -2357 666 -2329
rect 632 -2397 666 -2395
rect 632 -2429 666 -2397
rect 632 -2499 666 -2467
rect 632 -2501 666 -2499
rect 632 -2567 666 -2539
rect 632 -2573 666 -2567
rect 632 -2635 666 -2611
rect 632 -2645 666 -2635
rect 632 -2703 666 -2683
rect 632 -2717 666 -2703
rect 632 -2771 666 -2755
rect 632 -2789 666 -2771
rect 632 -2839 666 -2827
rect 632 -2861 666 -2839
rect 632 -2907 666 -2899
rect 632 -2933 666 -2907
rect 632 -2975 666 -2971
rect 632 -3005 666 -2975
rect 632 -3077 666 -3043
rect 632 -3145 666 -3115
rect 632 -3149 666 -3145
rect 632 -3213 666 -3187
rect 632 -3221 666 -3213
rect 632 -3281 666 -3259
rect 632 -3293 666 -3281
rect 632 -3349 666 -3331
rect 632 -3365 666 -3349
rect 632 -3417 666 -3403
rect 632 -3437 666 -3417
rect 632 -3485 666 -3475
rect 632 -3509 666 -3485
rect 632 -3553 666 -3547
rect 632 -3581 666 -3553
rect 632 -3621 666 -3619
rect 632 -3653 666 -3621
rect 632 -3723 666 -3691
rect 632 -3725 666 -3723
rect 632 -3791 666 -3763
rect 632 -3797 666 -3791
rect 632 -3859 666 -3835
rect 632 -3869 666 -3859
rect 632 -3927 666 -3907
rect 632 -3941 666 -3927
rect 632 -3995 666 -3979
rect 632 -4013 666 -3995
rect 632 -4063 666 -4051
rect 632 -4085 666 -4063
rect 632 -4131 666 -4123
rect 632 -4157 666 -4131
rect 632 -4199 666 -4195
rect 632 -4229 666 -4199
rect 632 -4301 666 -4267
rect 632 -4369 666 -4339
rect 632 -4373 666 -4369
rect 632 -4437 666 -4411
rect 632 -4445 666 -4437
rect 632 -4505 666 -4483
rect 632 -4517 666 -4505
rect 632 -4573 666 -4555
rect 632 -4589 666 -4573
rect 632 -4641 666 -4627
rect 632 -4661 666 -4641
rect 632 -4709 666 -4699
rect 632 -4733 666 -4709
rect 632 -4777 666 -4771
rect 632 -4805 666 -4777
rect 632 -4845 666 -4843
rect 632 -4877 666 -4845
rect 632 -4947 666 -4915
rect 632 -4949 666 -4947
rect 632 -5015 666 -4987
rect 632 -5021 666 -5015
rect 632 -5083 666 -5059
rect 632 -5093 666 -5083
rect 632 -5151 666 -5131
rect 632 -5165 666 -5151
rect 632 -5219 666 -5203
rect 632 -5237 666 -5219
rect 632 -5287 666 -5275
rect 632 -5309 666 -5287
rect 632 -5355 666 -5347
rect 632 -5381 666 -5355
rect 632 -5423 666 -5419
rect 632 -5453 666 -5423
rect 632 -5525 666 -5491
rect 632 -5593 666 -5563
rect 632 -5597 666 -5593
rect 632 -5661 666 -5635
rect 632 -5669 666 -5661
rect 632 -5729 666 -5707
rect 632 -5741 666 -5729
rect 632 -5797 666 -5779
rect 632 -5813 666 -5797
rect 632 -5865 666 -5851
rect 632 -5885 666 -5865
rect 632 -5933 666 -5923
rect 632 -5957 666 -5933
rect 632 -6001 666 -5995
rect 632 -6029 666 -6001
rect 632 -6069 666 -6067
rect 632 -6101 666 -6069
rect 632 -6171 666 -6139
rect 632 -6173 666 -6171
rect 632 -6239 666 -6211
rect 632 -6245 666 -6239
rect 632 -6307 666 -6283
rect 632 -6317 666 -6307
rect 632 -6375 666 -6355
rect 632 -6389 666 -6375
rect 632 -6443 666 -6427
rect 632 -6461 666 -6443
rect 632 -6511 666 -6499
rect 632 -6533 666 -6511
rect 632 -6579 666 -6571
rect 632 -6605 666 -6579
rect 632 -6647 666 -6643
rect 632 -6677 666 -6647
rect 632 -6749 666 -6715
rect 632 -6817 666 -6787
rect 632 -6821 666 -6817
rect 632 -6885 666 -6859
rect 632 -6893 666 -6885
rect 632 -6953 666 -6931
rect 632 -6965 666 -6953
rect 632 -7021 666 -7003
rect 632 -7037 666 -7021
rect 632 -7089 666 -7075
rect 632 -7109 666 -7089
rect 632 -7157 666 -7147
rect 632 -7181 666 -7157
rect 632 -7225 666 -7219
rect 632 -7253 666 -7225
rect 632 -7293 666 -7291
rect 632 -7325 666 -7293
rect 632 -7395 666 -7363
rect 632 -7397 666 -7395
rect 632 -7463 666 -7435
rect 632 -7469 666 -7463
rect 632 -7531 666 -7507
rect 632 -7541 666 -7531
rect 632 -7599 666 -7579
rect 632 -7613 666 -7599
rect 632 -7667 666 -7651
rect 632 -7685 666 -7667
rect 632 -7735 666 -7723
rect 632 -7757 666 -7735
rect 632 -7803 666 -7795
rect 632 -7829 666 -7803
rect 632 -7871 666 -7867
rect 632 -7901 666 -7871
rect 632 -7973 666 -7939
rect 632 -8041 666 -8011
rect 632 -8045 666 -8041
rect 632 -8109 666 -8083
rect 632 -8117 666 -8109
rect 632 -8177 666 -8155
rect 632 -8189 666 -8177
rect 632 -8245 666 -8227
rect 632 -8261 666 -8245
rect 632 -8313 666 -8299
rect 632 -8333 666 -8313
rect 632 -8381 666 -8371
rect 632 -8405 666 -8381
rect 632 -8449 666 -8443
rect 632 -8477 666 -8449
rect 632 -8517 666 -8515
rect 632 -8549 666 -8517
rect 632 -8619 666 -8587
rect 632 -8621 666 -8619
rect 632 -8687 666 -8659
rect 632 -8693 666 -8687
rect 632 -8755 666 -8731
rect 632 -8765 666 -8755
rect 632 -8823 666 -8803
rect 632 -8837 666 -8823
rect 632 -8891 666 -8875
rect 632 -8909 666 -8891
rect 632 -8959 666 -8947
rect 632 -8981 666 -8959
rect 632 -9027 666 -9019
rect 632 -9053 666 -9027
rect 632 -9095 666 -9091
rect 632 -9125 666 -9095
rect 632 -9197 666 -9163
rect 632 -9265 666 -9235
rect 632 -9269 666 -9265
rect 632 -9333 666 -9307
rect 632 -9341 666 -9333
rect 632 -9401 666 -9379
rect 632 -9413 666 -9401
rect 632 -9469 666 -9451
rect 632 -9485 666 -9469
rect 632 -9537 666 -9523
rect 632 -9557 666 -9537
rect 750 9537 784 9557
rect 750 9523 784 9537
rect 750 9469 784 9485
rect 750 9451 784 9469
rect 750 9401 784 9413
rect 750 9379 784 9401
rect 750 9333 784 9341
rect 750 9307 784 9333
rect 750 9265 784 9269
rect 750 9235 784 9265
rect 750 9163 784 9197
rect 750 9095 784 9125
rect 750 9091 784 9095
rect 750 9027 784 9053
rect 750 9019 784 9027
rect 750 8959 784 8981
rect 750 8947 784 8959
rect 750 8891 784 8909
rect 750 8875 784 8891
rect 750 8823 784 8837
rect 750 8803 784 8823
rect 750 8755 784 8765
rect 750 8731 784 8755
rect 750 8687 784 8693
rect 750 8659 784 8687
rect 750 8619 784 8621
rect 750 8587 784 8619
rect 750 8517 784 8549
rect 750 8515 784 8517
rect 750 8449 784 8477
rect 750 8443 784 8449
rect 750 8381 784 8405
rect 750 8371 784 8381
rect 750 8313 784 8333
rect 750 8299 784 8313
rect 750 8245 784 8261
rect 750 8227 784 8245
rect 750 8177 784 8189
rect 750 8155 784 8177
rect 750 8109 784 8117
rect 750 8083 784 8109
rect 750 8041 784 8045
rect 750 8011 784 8041
rect 750 7939 784 7973
rect 750 7871 784 7901
rect 750 7867 784 7871
rect 750 7803 784 7829
rect 750 7795 784 7803
rect 750 7735 784 7757
rect 750 7723 784 7735
rect 750 7667 784 7685
rect 750 7651 784 7667
rect 750 7599 784 7613
rect 750 7579 784 7599
rect 750 7531 784 7541
rect 750 7507 784 7531
rect 750 7463 784 7469
rect 750 7435 784 7463
rect 750 7395 784 7397
rect 750 7363 784 7395
rect 750 7293 784 7325
rect 750 7291 784 7293
rect 750 7225 784 7253
rect 750 7219 784 7225
rect 750 7157 784 7181
rect 750 7147 784 7157
rect 750 7089 784 7109
rect 750 7075 784 7089
rect 750 7021 784 7037
rect 750 7003 784 7021
rect 750 6953 784 6965
rect 750 6931 784 6953
rect 750 6885 784 6893
rect 750 6859 784 6885
rect 750 6817 784 6821
rect 750 6787 784 6817
rect 750 6715 784 6749
rect 750 6647 784 6677
rect 750 6643 784 6647
rect 750 6579 784 6605
rect 750 6571 784 6579
rect 750 6511 784 6533
rect 750 6499 784 6511
rect 750 6443 784 6461
rect 750 6427 784 6443
rect 750 6375 784 6389
rect 750 6355 784 6375
rect 750 6307 784 6317
rect 750 6283 784 6307
rect 750 6239 784 6245
rect 750 6211 784 6239
rect 750 6171 784 6173
rect 750 6139 784 6171
rect 750 6069 784 6101
rect 750 6067 784 6069
rect 750 6001 784 6029
rect 750 5995 784 6001
rect 750 5933 784 5957
rect 750 5923 784 5933
rect 750 5865 784 5885
rect 750 5851 784 5865
rect 750 5797 784 5813
rect 750 5779 784 5797
rect 750 5729 784 5741
rect 750 5707 784 5729
rect 750 5661 784 5669
rect 750 5635 784 5661
rect 750 5593 784 5597
rect 750 5563 784 5593
rect 750 5491 784 5525
rect 750 5423 784 5453
rect 750 5419 784 5423
rect 750 5355 784 5381
rect 750 5347 784 5355
rect 750 5287 784 5309
rect 750 5275 784 5287
rect 750 5219 784 5237
rect 750 5203 784 5219
rect 750 5151 784 5165
rect 750 5131 784 5151
rect 750 5083 784 5093
rect 750 5059 784 5083
rect 750 5015 784 5021
rect 750 4987 784 5015
rect 750 4947 784 4949
rect 750 4915 784 4947
rect 750 4845 784 4877
rect 750 4843 784 4845
rect 750 4777 784 4805
rect 750 4771 784 4777
rect 750 4709 784 4733
rect 750 4699 784 4709
rect 750 4641 784 4661
rect 750 4627 784 4641
rect 750 4573 784 4589
rect 750 4555 784 4573
rect 750 4505 784 4517
rect 750 4483 784 4505
rect 750 4437 784 4445
rect 750 4411 784 4437
rect 750 4369 784 4373
rect 750 4339 784 4369
rect 750 4267 784 4301
rect 750 4199 784 4229
rect 750 4195 784 4199
rect 750 4131 784 4157
rect 750 4123 784 4131
rect 750 4063 784 4085
rect 750 4051 784 4063
rect 750 3995 784 4013
rect 750 3979 784 3995
rect 750 3927 784 3941
rect 750 3907 784 3927
rect 750 3859 784 3869
rect 750 3835 784 3859
rect 750 3791 784 3797
rect 750 3763 784 3791
rect 750 3723 784 3725
rect 750 3691 784 3723
rect 750 3621 784 3653
rect 750 3619 784 3621
rect 750 3553 784 3581
rect 750 3547 784 3553
rect 750 3485 784 3509
rect 750 3475 784 3485
rect 750 3417 784 3437
rect 750 3403 784 3417
rect 750 3349 784 3365
rect 750 3331 784 3349
rect 750 3281 784 3293
rect 750 3259 784 3281
rect 750 3213 784 3221
rect 750 3187 784 3213
rect 750 3145 784 3149
rect 750 3115 784 3145
rect 750 3043 784 3077
rect 750 2975 784 3005
rect 750 2971 784 2975
rect 750 2907 784 2933
rect 750 2899 784 2907
rect 750 2839 784 2861
rect 750 2827 784 2839
rect 750 2771 784 2789
rect 750 2755 784 2771
rect 750 2703 784 2717
rect 750 2683 784 2703
rect 750 2635 784 2645
rect 750 2611 784 2635
rect 750 2567 784 2573
rect 750 2539 784 2567
rect 750 2499 784 2501
rect 750 2467 784 2499
rect 750 2397 784 2429
rect 750 2395 784 2397
rect 750 2329 784 2357
rect 750 2323 784 2329
rect 750 2261 784 2285
rect 750 2251 784 2261
rect 750 2193 784 2213
rect 750 2179 784 2193
rect 750 2125 784 2141
rect 750 2107 784 2125
rect 750 2057 784 2069
rect 750 2035 784 2057
rect 750 1989 784 1997
rect 750 1963 784 1989
rect 750 1921 784 1925
rect 750 1891 784 1921
rect 750 1819 784 1853
rect 750 1751 784 1781
rect 750 1747 784 1751
rect 750 1683 784 1709
rect 750 1675 784 1683
rect 750 1615 784 1637
rect 750 1603 784 1615
rect 750 1547 784 1565
rect 750 1531 784 1547
rect 750 1479 784 1493
rect 750 1459 784 1479
rect 750 1411 784 1421
rect 750 1387 784 1411
rect 750 1343 784 1349
rect 750 1315 784 1343
rect 750 1275 784 1277
rect 750 1243 784 1275
rect 750 1173 784 1205
rect 750 1171 784 1173
rect 750 1105 784 1133
rect 750 1099 784 1105
rect 750 1037 784 1061
rect 750 1027 784 1037
rect 750 969 784 989
rect 750 955 784 969
rect 750 901 784 917
rect 750 883 784 901
rect 750 833 784 845
rect 750 811 784 833
rect 750 765 784 773
rect 750 739 784 765
rect 750 697 784 701
rect 750 667 784 697
rect 750 595 784 629
rect 750 527 784 557
rect 750 523 784 527
rect 750 459 784 485
rect 750 451 784 459
rect 750 391 784 413
rect 750 379 784 391
rect 750 323 784 341
rect 750 307 784 323
rect 750 255 784 269
rect 750 235 784 255
rect 750 187 784 197
rect 750 163 784 187
rect 750 119 784 125
rect 750 91 784 119
rect 750 51 784 53
rect 750 19 784 51
rect 750 -51 784 -19
rect 750 -53 784 -51
rect 750 -119 784 -91
rect 750 -125 784 -119
rect 750 -187 784 -163
rect 750 -197 784 -187
rect 750 -255 784 -235
rect 750 -269 784 -255
rect 750 -323 784 -307
rect 750 -341 784 -323
rect 750 -391 784 -379
rect 750 -413 784 -391
rect 750 -459 784 -451
rect 750 -485 784 -459
rect 750 -527 784 -523
rect 750 -557 784 -527
rect 750 -629 784 -595
rect 750 -697 784 -667
rect 750 -701 784 -697
rect 750 -765 784 -739
rect 750 -773 784 -765
rect 750 -833 784 -811
rect 750 -845 784 -833
rect 750 -901 784 -883
rect 750 -917 784 -901
rect 750 -969 784 -955
rect 750 -989 784 -969
rect 750 -1037 784 -1027
rect 750 -1061 784 -1037
rect 750 -1105 784 -1099
rect 750 -1133 784 -1105
rect 750 -1173 784 -1171
rect 750 -1205 784 -1173
rect 750 -1275 784 -1243
rect 750 -1277 784 -1275
rect 750 -1343 784 -1315
rect 750 -1349 784 -1343
rect 750 -1411 784 -1387
rect 750 -1421 784 -1411
rect 750 -1479 784 -1459
rect 750 -1493 784 -1479
rect 750 -1547 784 -1531
rect 750 -1565 784 -1547
rect 750 -1615 784 -1603
rect 750 -1637 784 -1615
rect 750 -1683 784 -1675
rect 750 -1709 784 -1683
rect 750 -1751 784 -1747
rect 750 -1781 784 -1751
rect 750 -1853 784 -1819
rect 750 -1921 784 -1891
rect 750 -1925 784 -1921
rect 750 -1989 784 -1963
rect 750 -1997 784 -1989
rect 750 -2057 784 -2035
rect 750 -2069 784 -2057
rect 750 -2125 784 -2107
rect 750 -2141 784 -2125
rect 750 -2193 784 -2179
rect 750 -2213 784 -2193
rect 750 -2261 784 -2251
rect 750 -2285 784 -2261
rect 750 -2329 784 -2323
rect 750 -2357 784 -2329
rect 750 -2397 784 -2395
rect 750 -2429 784 -2397
rect 750 -2499 784 -2467
rect 750 -2501 784 -2499
rect 750 -2567 784 -2539
rect 750 -2573 784 -2567
rect 750 -2635 784 -2611
rect 750 -2645 784 -2635
rect 750 -2703 784 -2683
rect 750 -2717 784 -2703
rect 750 -2771 784 -2755
rect 750 -2789 784 -2771
rect 750 -2839 784 -2827
rect 750 -2861 784 -2839
rect 750 -2907 784 -2899
rect 750 -2933 784 -2907
rect 750 -2975 784 -2971
rect 750 -3005 784 -2975
rect 750 -3077 784 -3043
rect 750 -3145 784 -3115
rect 750 -3149 784 -3145
rect 750 -3213 784 -3187
rect 750 -3221 784 -3213
rect 750 -3281 784 -3259
rect 750 -3293 784 -3281
rect 750 -3349 784 -3331
rect 750 -3365 784 -3349
rect 750 -3417 784 -3403
rect 750 -3437 784 -3417
rect 750 -3485 784 -3475
rect 750 -3509 784 -3485
rect 750 -3553 784 -3547
rect 750 -3581 784 -3553
rect 750 -3621 784 -3619
rect 750 -3653 784 -3621
rect 750 -3723 784 -3691
rect 750 -3725 784 -3723
rect 750 -3791 784 -3763
rect 750 -3797 784 -3791
rect 750 -3859 784 -3835
rect 750 -3869 784 -3859
rect 750 -3927 784 -3907
rect 750 -3941 784 -3927
rect 750 -3995 784 -3979
rect 750 -4013 784 -3995
rect 750 -4063 784 -4051
rect 750 -4085 784 -4063
rect 750 -4131 784 -4123
rect 750 -4157 784 -4131
rect 750 -4199 784 -4195
rect 750 -4229 784 -4199
rect 750 -4301 784 -4267
rect 750 -4369 784 -4339
rect 750 -4373 784 -4369
rect 750 -4437 784 -4411
rect 750 -4445 784 -4437
rect 750 -4505 784 -4483
rect 750 -4517 784 -4505
rect 750 -4573 784 -4555
rect 750 -4589 784 -4573
rect 750 -4641 784 -4627
rect 750 -4661 784 -4641
rect 750 -4709 784 -4699
rect 750 -4733 784 -4709
rect 750 -4777 784 -4771
rect 750 -4805 784 -4777
rect 750 -4845 784 -4843
rect 750 -4877 784 -4845
rect 750 -4947 784 -4915
rect 750 -4949 784 -4947
rect 750 -5015 784 -4987
rect 750 -5021 784 -5015
rect 750 -5083 784 -5059
rect 750 -5093 784 -5083
rect 750 -5151 784 -5131
rect 750 -5165 784 -5151
rect 750 -5219 784 -5203
rect 750 -5237 784 -5219
rect 750 -5287 784 -5275
rect 750 -5309 784 -5287
rect 750 -5355 784 -5347
rect 750 -5381 784 -5355
rect 750 -5423 784 -5419
rect 750 -5453 784 -5423
rect 750 -5525 784 -5491
rect 750 -5593 784 -5563
rect 750 -5597 784 -5593
rect 750 -5661 784 -5635
rect 750 -5669 784 -5661
rect 750 -5729 784 -5707
rect 750 -5741 784 -5729
rect 750 -5797 784 -5779
rect 750 -5813 784 -5797
rect 750 -5865 784 -5851
rect 750 -5885 784 -5865
rect 750 -5933 784 -5923
rect 750 -5957 784 -5933
rect 750 -6001 784 -5995
rect 750 -6029 784 -6001
rect 750 -6069 784 -6067
rect 750 -6101 784 -6069
rect 750 -6171 784 -6139
rect 750 -6173 784 -6171
rect 750 -6239 784 -6211
rect 750 -6245 784 -6239
rect 750 -6307 784 -6283
rect 750 -6317 784 -6307
rect 750 -6375 784 -6355
rect 750 -6389 784 -6375
rect 750 -6443 784 -6427
rect 750 -6461 784 -6443
rect 750 -6511 784 -6499
rect 750 -6533 784 -6511
rect 750 -6579 784 -6571
rect 750 -6605 784 -6579
rect 750 -6647 784 -6643
rect 750 -6677 784 -6647
rect 750 -6749 784 -6715
rect 750 -6817 784 -6787
rect 750 -6821 784 -6817
rect 750 -6885 784 -6859
rect 750 -6893 784 -6885
rect 750 -6953 784 -6931
rect 750 -6965 784 -6953
rect 750 -7021 784 -7003
rect 750 -7037 784 -7021
rect 750 -7089 784 -7075
rect 750 -7109 784 -7089
rect 750 -7157 784 -7147
rect 750 -7181 784 -7157
rect 750 -7225 784 -7219
rect 750 -7253 784 -7225
rect 750 -7293 784 -7291
rect 750 -7325 784 -7293
rect 750 -7395 784 -7363
rect 750 -7397 784 -7395
rect 750 -7463 784 -7435
rect 750 -7469 784 -7463
rect 750 -7531 784 -7507
rect 750 -7541 784 -7531
rect 750 -7599 784 -7579
rect 750 -7613 784 -7599
rect 750 -7667 784 -7651
rect 750 -7685 784 -7667
rect 750 -7735 784 -7723
rect 750 -7757 784 -7735
rect 750 -7803 784 -7795
rect 750 -7829 784 -7803
rect 750 -7871 784 -7867
rect 750 -7901 784 -7871
rect 750 -7973 784 -7939
rect 750 -8041 784 -8011
rect 750 -8045 784 -8041
rect 750 -8109 784 -8083
rect 750 -8117 784 -8109
rect 750 -8177 784 -8155
rect 750 -8189 784 -8177
rect 750 -8245 784 -8227
rect 750 -8261 784 -8245
rect 750 -8313 784 -8299
rect 750 -8333 784 -8313
rect 750 -8381 784 -8371
rect 750 -8405 784 -8381
rect 750 -8449 784 -8443
rect 750 -8477 784 -8449
rect 750 -8517 784 -8515
rect 750 -8549 784 -8517
rect 750 -8619 784 -8587
rect 750 -8621 784 -8619
rect 750 -8687 784 -8659
rect 750 -8693 784 -8687
rect 750 -8755 784 -8731
rect 750 -8765 784 -8755
rect 750 -8823 784 -8803
rect 750 -8837 784 -8823
rect 750 -8891 784 -8875
rect 750 -8909 784 -8891
rect 750 -8959 784 -8947
rect 750 -8981 784 -8959
rect 750 -9027 784 -9019
rect 750 -9053 784 -9027
rect 750 -9095 784 -9091
rect 750 -9125 784 -9095
rect 750 -9197 784 -9163
rect 750 -9265 784 -9235
rect 750 -9269 784 -9265
rect 750 -9333 784 -9307
rect 750 -9341 784 -9333
rect 750 -9401 784 -9379
rect 750 -9413 784 -9401
rect 750 -9469 784 -9451
rect 750 -9485 784 -9469
rect 750 -9537 784 -9523
rect 750 -9557 784 -9537
rect 868 9537 902 9557
rect 868 9523 902 9537
rect 868 9469 902 9485
rect 868 9451 902 9469
rect 868 9401 902 9413
rect 868 9379 902 9401
rect 868 9333 902 9341
rect 868 9307 902 9333
rect 868 9265 902 9269
rect 868 9235 902 9265
rect 868 9163 902 9197
rect 868 9095 902 9125
rect 868 9091 902 9095
rect 868 9027 902 9053
rect 868 9019 902 9027
rect 868 8959 902 8981
rect 868 8947 902 8959
rect 868 8891 902 8909
rect 868 8875 902 8891
rect 868 8823 902 8837
rect 868 8803 902 8823
rect 868 8755 902 8765
rect 868 8731 902 8755
rect 868 8687 902 8693
rect 868 8659 902 8687
rect 868 8619 902 8621
rect 868 8587 902 8619
rect 868 8517 902 8549
rect 868 8515 902 8517
rect 868 8449 902 8477
rect 868 8443 902 8449
rect 868 8381 902 8405
rect 868 8371 902 8381
rect 868 8313 902 8333
rect 868 8299 902 8313
rect 868 8245 902 8261
rect 868 8227 902 8245
rect 868 8177 902 8189
rect 868 8155 902 8177
rect 868 8109 902 8117
rect 868 8083 902 8109
rect 868 8041 902 8045
rect 868 8011 902 8041
rect 868 7939 902 7973
rect 868 7871 902 7901
rect 868 7867 902 7871
rect 868 7803 902 7829
rect 868 7795 902 7803
rect 868 7735 902 7757
rect 868 7723 902 7735
rect 868 7667 902 7685
rect 868 7651 902 7667
rect 868 7599 902 7613
rect 868 7579 902 7599
rect 868 7531 902 7541
rect 868 7507 902 7531
rect 868 7463 902 7469
rect 868 7435 902 7463
rect 868 7395 902 7397
rect 868 7363 902 7395
rect 868 7293 902 7325
rect 868 7291 902 7293
rect 868 7225 902 7253
rect 868 7219 902 7225
rect 868 7157 902 7181
rect 868 7147 902 7157
rect 868 7089 902 7109
rect 868 7075 902 7089
rect 868 7021 902 7037
rect 868 7003 902 7021
rect 868 6953 902 6965
rect 868 6931 902 6953
rect 868 6885 902 6893
rect 868 6859 902 6885
rect 868 6817 902 6821
rect 868 6787 902 6817
rect 868 6715 902 6749
rect 868 6647 902 6677
rect 868 6643 902 6647
rect 868 6579 902 6605
rect 868 6571 902 6579
rect 868 6511 902 6533
rect 868 6499 902 6511
rect 868 6443 902 6461
rect 868 6427 902 6443
rect 868 6375 902 6389
rect 868 6355 902 6375
rect 868 6307 902 6317
rect 868 6283 902 6307
rect 868 6239 902 6245
rect 868 6211 902 6239
rect 868 6171 902 6173
rect 868 6139 902 6171
rect 868 6069 902 6101
rect 868 6067 902 6069
rect 868 6001 902 6029
rect 868 5995 902 6001
rect 868 5933 902 5957
rect 868 5923 902 5933
rect 868 5865 902 5885
rect 868 5851 902 5865
rect 868 5797 902 5813
rect 868 5779 902 5797
rect 868 5729 902 5741
rect 868 5707 902 5729
rect 868 5661 902 5669
rect 868 5635 902 5661
rect 868 5593 902 5597
rect 868 5563 902 5593
rect 868 5491 902 5525
rect 868 5423 902 5453
rect 868 5419 902 5423
rect 868 5355 902 5381
rect 868 5347 902 5355
rect 868 5287 902 5309
rect 868 5275 902 5287
rect 868 5219 902 5237
rect 868 5203 902 5219
rect 868 5151 902 5165
rect 868 5131 902 5151
rect 868 5083 902 5093
rect 868 5059 902 5083
rect 868 5015 902 5021
rect 868 4987 902 5015
rect 868 4947 902 4949
rect 868 4915 902 4947
rect 868 4845 902 4877
rect 868 4843 902 4845
rect 868 4777 902 4805
rect 868 4771 902 4777
rect 868 4709 902 4733
rect 868 4699 902 4709
rect 868 4641 902 4661
rect 868 4627 902 4641
rect 868 4573 902 4589
rect 868 4555 902 4573
rect 868 4505 902 4517
rect 868 4483 902 4505
rect 868 4437 902 4445
rect 868 4411 902 4437
rect 868 4369 902 4373
rect 868 4339 902 4369
rect 868 4267 902 4301
rect 868 4199 902 4229
rect 868 4195 902 4199
rect 868 4131 902 4157
rect 868 4123 902 4131
rect 868 4063 902 4085
rect 868 4051 902 4063
rect 868 3995 902 4013
rect 868 3979 902 3995
rect 868 3927 902 3941
rect 868 3907 902 3927
rect 868 3859 902 3869
rect 868 3835 902 3859
rect 868 3791 902 3797
rect 868 3763 902 3791
rect 868 3723 902 3725
rect 868 3691 902 3723
rect 868 3621 902 3653
rect 868 3619 902 3621
rect 868 3553 902 3581
rect 868 3547 902 3553
rect 868 3485 902 3509
rect 868 3475 902 3485
rect 868 3417 902 3437
rect 868 3403 902 3417
rect 868 3349 902 3365
rect 868 3331 902 3349
rect 868 3281 902 3293
rect 868 3259 902 3281
rect 868 3213 902 3221
rect 868 3187 902 3213
rect 868 3145 902 3149
rect 868 3115 902 3145
rect 868 3043 902 3077
rect 868 2975 902 3005
rect 868 2971 902 2975
rect 868 2907 902 2933
rect 868 2899 902 2907
rect 868 2839 902 2861
rect 868 2827 902 2839
rect 868 2771 902 2789
rect 868 2755 902 2771
rect 868 2703 902 2717
rect 868 2683 902 2703
rect 868 2635 902 2645
rect 868 2611 902 2635
rect 868 2567 902 2573
rect 868 2539 902 2567
rect 868 2499 902 2501
rect 868 2467 902 2499
rect 868 2397 902 2429
rect 868 2395 902 2397
rect 868 2329 902 2357
rect 868 2323 902 2329
rect 868 2261 902 2285
rect 868 2251 902 2261
rect 868 2193 902 2213
rect 868 2179 902 2193
rect 868 2125 902 2141
rect 868 2107 902 2125
rect 868 2057 902 2069
rect 868 2035 902 2057
rect 868 1989 902 1997
rect 868 1963 902 1989
rect 868 1921 902 1925
rect 868 1891 902 1921
rect 868 1819 902 1853
rect 868 1751 902 1781
rect 868 1747 902 1751
rect 868 1683 902 1709
rect 868 1675 902 1683
rect 868 1615 902 1637
rect 868 1603 902 1615
rect 868 1547 902 1565
rect 868 1531 902 1547
rect 868 1479 902 1493
rect 868 1459 902 1479
rect 868 1411 902 1421
rect 868 1387 902 1411
rect 868 1343 902 1349
rect 868 1315 902 1343
rect 868 1275 902 1277
rect 868 1243 902 1275
rect 868 1173 902 1205
rect 868 1171 902 1173
rect 868 1105 902 1133
rect 868 1099 902 1105
rect 868 1037 902 1061
rect 868 1027 902 1037
rect 868 969 902 989
rect 868 955 902 969
rect 868 901 902 917
rect 868 883 902 901
rect 868 833 902 845
rect 868 811 902 833
rect 868 765 902 773
rect 868 739 902 765
rect 868 697 902 701
rect 868 667 902 697
rect 868 595 902 629
rect 868 527 902 557
rect 868 523 902 527
rect 868 459 902 485
rect 868 451 902 459
rect 868 391 902 413
rect 868 379 902 391
rect 868 323 902 341
rect 868 307 902 323
rect 868 255 902 269
rect 868 235 902 255
rect 868 187 902 197
rect 868 163 902 187
rect 868 119 902 125
rect 868 91 902 119
rect 868 51 902 53
rect 868 19 902 51
rect 868 -51 902 -19
rect 868 -53 902 -51
rect 868 -119 902 -91
rect 868 -125 902 -119
rect 868 -187 902 -163
rect 868 -197 902 -187
rect 868 -255 902 -235
rect 868 -269 902 -255
rect 868 -323 902 -307
rect 868 -341 902 -323
rect 868 -391 902 -379
rect 868 -413 902 -391
rect 868 -459 902 -451
rect 868 -485 902 -459
rect 868 -527 902 -523
rect 868 -557 902 -527
rect 868 -629 902 -595
rect 868 -697 902 -667
rect 868 -701 902 -697
rect 868 -765 902 -739
rect 868 -773 902 -765
rect 868 -833 902 -811
rect 868 -845 902 -833
rect 868 -901 902 -883
rect 868 -917 902 -901
rect 868 -969 902 -955
rect 868 -989 902 -969
rect 868 -1037 902 -1027
rect 868 -1061 902 -1037
rect 868 -1105 902 -1099
rect 868 -1133 902 -1105
rect 868 -1173 902 -1171
rect 868 -1205 902 -1173
rect 868 -1275 902 -1243
rect 868 -1277 902 -1275
rect 868 -1343 902 -1315
rect 868 -1349 902 -1343
rect 868 -1411 902 -1387
rect 868 -1421 902 -1411
rect 868 -1479 902 -1459
rect 868 -1493 902 -1479
rect 868 -1547 902 -1531
rect 868 -1565 902 -1547
rect 868 -1615 902 -1603
rect 868 -1637 902 -1615
rect 868 -1683 902 -1675
rect 868 -1709 902 -1683
rect 868 -1751 902 -1747
rect 868 -1781 902 -1751
rect 868 -1853 902 -1819
rect 868 -1921 902 -1891
rect 868 -1925 902 -1921
rect 868 -1989 902 -1963
rect 868 -1997 902 -1989
rect 868 -2057 902 -2035
rect 868 -2069 902 -2057
rect 868 -2125 902 -2107
rect 868 -2141 902 -2125
rect 868 -2193 902 -2179
rect 868 -2213 902 -2193
rect 868 -2261 902 -2251
rect 868 -2285 902 -2261
rect 868 -2329 902 -2323
rect 868 -2357 902 -2329
rect 868 -2397 902 -2395
rect 868 -2429 902 -2397
rect 868 -2499 902 -2467
rect 868 -2501 902 -2499
rect 868 -2567 902 -2539
rect 868 -2573 902 -2567
rect 868 -2635 902 -2611
rect 868 -2645 902 -2635
rect 868 -2703 902 -2683
rect 868 -2717 902 -2703
rect 868 -2771 902 -2755
rect 868 -2789 902 -2771
rect 868 -2839 902 -2827
rect 868 -2861 902 -2839
rect 868 -2907 902 -2899
rect 868 -2933 902 -2907
rect 868 -2975 902 -2971
rect 868 -3005 902 -2975
rect 868 -3077 902 -3043
rect 868 -3145 902 -3115
rect 868 -3149 902 -3145
rect 868 -3213 902 -3187
rect 868 -3221 902 -3213
rect 868 -3281 902 -3259
rect 868 -3293 902 -3281
rect 868 -3349 902 -3331
rect 868 -3365 902 -3349
rect 868 -3417 902 -3403
rect 868 -3437 902 -3417
rect 868 -3485 902 -3475
rect 868 -3509 902 -3485
rect 868 -3553 902 -3547
rect 868 -3581 902 -3553
rect 868 -3621 902 -3619
rect 868 -3653 902 -3621
rect 868 -3723 902 -3691
rect 868 -3725 902 -3723
rect 868 -3791 902 -3763
rect 868 -3797 902 -3791
rect 868 -3859 902 -3835
rect 868 -3869 902 -3859
rect 868 -3927 902 -3907
rect 868 -3941 902 -3927
rect 868 -3995 902 -3979
rect 868 -4013 902 -3995
rect 868 -4063 902 -4051
rect 868 -4085 902 -4063
rect 868 -4131 902 -4123
rect 868 -4157 902 -4131
rect 868 -4199 902 -4195
rect 868 -4229 902 -4199
rect 868 -4301 902 -4267
rect 868 -4369 902 -4339
rect 868 -4373 902 -4369
rect 868 -4437 902 -4411
rect 868 -4445 902 -4437
rect 868 -4505 902 -4483
rect 868 -4517 902 -4505
rect 868 -4573 902 -4555
rect 868 -4589 902 -4573
rect 868 -4641 902 -4627
rect 868 -4661 902 -4641
rect 868 -4709 902 -4699
rect 868 -4733 902 -4709
rect 868 -4777 902 -4771
rect 868 -4805 902 -4777
rect 868 -4845 902 -4843
rect 868 -4877 902 -4845
rect 868 -4947 902 -4915
rect 868 -4949 902 -4947
rect 868 -5015 902 -4987
rect 868 -5021 902 -5015
rect 868 -5083 902 -5059
rect 868 -5093 902 -5083
rect 868 -5151 902 -5131
rect 868 -5165 902 -5151
rect 868 -5219 902 -5203
rect 868 -5237 902 -5219
rect 868 -5287 902 -5275
rect 868 -5309 902 -5287
rect 868 -5355 902 -5347
rect 868 -5381 902 -5355
rect 868 -5423 902 -5419
rect 868 -5453 902 -5423
rect 868 -5525 902 -5491
rect 868 -5593 902 -5563
rect 868 -5597 902 -5593
rect 868 -5661 902 -5635
rect 868 -5669 902 -5661
rect 868 -5729 902 -5707
rect 868 -5741 902 -5729
rect 868 -5797 902 -5779
rect 868 -5813 902 -5797
rect 868 -5865 902 -5851
rect 868 -5885 902 -5865
rect 868 -5933 902 -5923
rect 868 -5957 902 -5933
rect 868 -6001 902 -5995
rect 868 -6029 902 -6001
rect 868 -6069 902 -6067
rect 868 -6101 902 -6069
rect 868 -6171 902 -6139
rect 868 -6173 902 -6171
rect 868 -6239 902 -6211
rect 868 -6245 902 -6239
rect 868 -6307 902 -6283
rect 868 -6317 902 -6307
rect 868 -6375 902 -6355
rect 868 -6389 902 -6375
rect 868 -6443 902 -6427
rect 868 -6461 902 -6443
rect 868 -6511 902 -6499
rect 868 -6533 902 -6511
rect 868 -6579 902 -6571
rect 868 -6605 902 -6579
rect 868 -6647 902 -6643
rect 868 -6677 902 -6647
rect 868 -6749 902 -6715
rect 868 -6817 902 -6787
rect 868 -6821 902 -6817
rect 868 -6885 902 -6859
rect 868 -6893 902 -6885
rect 868 -6953 902 -6931
rect 868 -6965 902 -6953
rect 868 -7021 902 -7003
rect 868 -7037 902 -7021
rect 868 -7089 902 -7075
rect 868 -7109 902 -7089
rect 868 -7157 902 -7147
rect 868 -7181 902 -7157
rect 868 -7225 902 -7219
rect 868 -7253 902 -7225
rect 868 -7293 902 -7291
rect 868 -7325 902 -7293
rect 868 -7395 902 -7363
rect 868 -7397 902 -7395
rect 868 -7463 902 -7435
rect 868 -7469 902 -7463
rect 868 -7531 902 -7507
rect 868 -7541 902 -7531
rect 868 -7599 902 -7579
rect 868 -7613 902 -7599
rect 868 -7667 902 -7651
rect 868 -7685 902 -7667
rect 868 -7735 902 -7723
rect 868 -7757 902 -7735
rect 868 -7803 902 -7795
rect 868 -7829 902 -7803
rect 868 -7871 902 -7867
rect 868 -7901 902 -7871
rect 868 -7973 902 -7939
rect 868 -8041 902 -8011
rect 868 -8045 902 -8041
rect 868 -8109 902 -8083
rect 868 -8117 902 -8109
rect 868 -8177 902 -8155
rect 868 -8189 902 -8177
rect 868 -8245 902 -8227
rect 868 -8261 902 -8245
rect 868 -8313 902 -8299
rect 868 -8333 902 -8313
rect 868 -8381 902 -8371
rect 868 -8405 902 -8381
rect 868 -8449 902 -8443
rect 868 -8477 902 -8449
rect 868 -8517 902 -8515
rect 868 -8549 902 -8517
rect 868 -8619 902 -8587
rect 868 -8621 902 -8619
rect 868 -8687 902 -8659
rect 868 -8693 902 -8687
rect 868 -8755 902 -8731
rect 868 -8765 902 -8755
rect 868 -8823 902 -8803
rect 868 -8837 902 -8823
rect 868 -8891 902 -8875
rect 868 -8909 902 -8891
rect 868 -8959 902 -8947
rect 868 -8981 902 -8959
rect 868 -9027 902 -9019
rect 868 -9053 902 -9027
rect 868 -9095 902 -9091
rect 868 -9125 902 -9095
rect 868 -9197 902 -9163
rect 868 -9265 902 -9235
rect 868 -9269 902 -9265
rect 868 -9333 902 -9307
rect 868 -9341 902 -9333
rect 868 -9401 902 -9379
rect 868 -9413 902 -9401
rect 868 -9469 902 -9451
rect 868 -9485 902 -9469
rect 868 -9537 902 -9523
rect 868 -9557 902 -9537
rect 986 9537 1020 9557
rect 986 9523 1020 9537
rect 986 9469 1020 9485
rect 986 9451 1020 9469
rect 986 9401 1020 9413
rect 986 9379 1020 9401
rect 986 9333 1020 9341
rect 986 9307 1020 9333
rect 986 9265 1020 9269
rect 986 9235 1020 9265
rect 986 9163 1020 9197
rect 986 9095 1020 9125
rect 986 9091 1020 9095
rect 986 9027 1020 9053
rect 986 9019 1020 9027
rect 986 8959 1020 8981
rect 986 8947 1020 8959
rect 986 8891 1020 8909
rect 986 8875 1020 8891
rect 986 8823 1020 8837
rect 986 8803 1020 8823
rect 986 8755 1020 8765
rect 986 8731 1020 8755
rect 986 8687 1020 8693
rect 986 8659 1020 8687
rect 986 8619 1020 8621
rect 986 8587 1020 8619
rect 986 8517 1020 8549
rect 986 8515 1020 8517
rect 986 8449 1020 8477
rect 986 8443 1020 8449
rect 986 8381 1020 8405
rect 986 8371 1020 8381
rect 986 8313 1020 8333
rect 986 8299 1020 8313
rect 986 8245 1020 8261
rect 986 8227 1020 8245
rect 986 8177 1020 8189
rect 986 8155 1020 8177
rect 986 8109 1020 8117
rect 986 8083 1020 8109
rect 986 8041 1020 8045
rect 986 8011 1020 8041
rect 986 7939 1020 7973
rect 986 7871 1020 7901
rect 986 7867 1020 7871
rect 986 7803 1020 7829
rect 986 7795 1020 7803
rect 986 7735 1020 7757
rect 986 7723 1020 7735
rect 986 7667 1020 7685
rect 986 7651 1020 7667
rect 986 7599 1020 7613
rect 986 7579 1020 7599
rect 986 7531 1020 7541
rect 986 7507 1020 7531
rect 986 7463 1020 7469
rect 986 7435 1020 7463
rect 986 7395 1020 7397
rect 986 7363 1020 7395
rect 986 7293 1020 7325
rect 986 7291 1020 7293
rect 986 7225 1020 7253
rect 986 7219 1020 7225
rect 986 7157 1020 7181
rect 986 7147 1020 7157
rect 986 7089 1020 7109
rect 986 7075 1020 7089
rect 986 7021 1020 7037
rect 986 7003 1020 7021
rect 986 6953 1020 6965
rect 986 6931 1020 6953
rect 986 6885 1020 6893
rect 986 6859 1020 6885
rect 986 6817 1020 6821
rect 986 6787 1020 6817
rect 986 6715 1020 6749
rect 986 6647 1020 6677
rect 986 6643 1020 6647
rect 986 6579 1020 6605
rect 986 6571 1020 6579
rect 986 6511 1020 6533
rect 986 6499 1020 6511
rect 986 6443 1020 6461
rect 986 6427 1020 6443
rect 986 6375 1020 6389
rect 986 6355 1020 6375
rect 986 6307 1020 6317
rect 986 6283 1020 6307
rect 986 6239 1020 6245
rect 986 6211 1020 6239
rect 986 6171 1020 6173
rect 986 6139 1020 6171
rect 986 6069 1020 6101
rect 986 6067 1020 6069
rect 986 6001 1020 6029
rect 986 5995 1020 6001
rect 986 5933 1020 5957
rect 986 5923 1020 5933
rect 986 5865 1020 5885
rect 986 5851 1020 5865
rect 986 5797 1020 5813
rect 986 5779 1020 5797
rect 986 5729 1020 5741
rect 986 5707 1020 5729
rect 986 5661 1020 5669
rect 986 5635 1020 5661
rect 986 5593 1020 5597
rect 986 5563 1020 5593
rect 986 5491 1020 5525
rect 986 5423 1020 5453
rect 986 5419 1020 5423
rect 986 5355 1020 5381
rect 986 5347 1020 5355
rect 986 5287 1020 5309
rect 986 5275 1020 5287
rect 986 5219 1020 5237
rect 986 5203 1020 5219
rect 986 5151 1020 5165
rect 986 5131 1020 5151
rect 986 5083 1020 5093
rect 986 5059 1020 5083
rect 986 5015 1020 5021
rect 986 4987 1020 5015
rect 986 4947 1020 4949
rect 986 4915 1020 4947
rect 986 4845 1020 4877
rect 986 4843 1020 4845
rect 986 4777 1020 4805
rect 986 4771 1020 4777
rect 986 4709 1020 4733
rect 986 4699 1020 4709
rect 986 4641 1020 4661
rect 986 4627 1020 4641
rect 986 4573 1020 4589
rect 986 4555 1020 4573
rect 986 4505 1020 4517
rect 986 4483 1020 4505
rect 986 4437 1020 4445
rect 986 4411 1020 4437
rect 986 4369 1020 4373
rect 986 4339 1020 4369
rect 986 4267 1020 4301
rect 986 4199 1020 4229
rect 986 4195 1020 4199
rect 986 4131 1020 4157
rect 986 4123 1020 4131
rect 986 4063 1020 4085
rect 986 4051 1020 4063
rect 986 3995 1020 4013
rect 986 3979 1020 3995
rect 986 3927 1020 3941
rect 986 3907 1020 3927
rect 986 3859 1020 3869
rect 986 3835 1020 3859
rect 986 3791 1020 3797
rect 986 3763 1020 3791
rect 986 3723 1020 3725
rect 986 3691 1020 3723
rect 986 3621 1020 3653
rect 986 3619 1020 3621
rect 986 3553 1020 3581
rect 986 3547 1020 3553
rect 986 3485 1020 3509
rect 986 3475 1020 3485
rect 986 3417 1020 3437
rect 986 3403 1020 3417
rect 986 3349 1020 3365
rect 986 3331 1020 3349
rect 986 3281 1020 3293
rect 986 3259 1020 3281
rect 986 3213 1020 3221
rect 986 3187 1020 3213
rect 986 3145 1020 3149
rect 986 3115 1020 3145
rect 986 3043 1020 3077
rect 986 2975 1020 3005
rect 986 2971 1020 2975
rect 986 2907 1020 2933
rect 986 2899 1020 2907
rect 986 2839 1020 2861
rect 986 2827 1020 2839
rect 986 2771 1020 2789
rect 986 2755 1020 2771
rect 986 2703 1020 2717
rect 986 2683 1020 2703
rect 986 2635 1020 2645
rect 986 2611 1020 2635
rect 986 2567 1020 2573
rect 986 2539 1020 2567
rect 986 2499 1020 2501
rect 986 2467 1020 2499
rect 986 2397 1020 2429
rect 986 2395 1020 2397
rect 986 2329 1020 2357
rect 986 2323 1020 2329
rect 986 2261 1020 2285
rect 986 2251 1020 2261
rect 986 2193 1020 2213
rect 986 2179 1020 2193
rect 986 2125 1020 2141
rect 986 2107 1020 2125
rect 986 2057 1020 2069
rect 986 2035 1020 2057
rect 986 1989 1020 1997
rect 986 1963 1020 1989
rect 986 1921 1020 1925
rect 986 1891 1020 1921
rect 986 1819 1020 1853
rect 986 1751 1020 1781
rect 986 1747 1020 1751
rect 986 1683 1020 1709
rect 986 1675 1020 1683
rect 986 1615 1020 1637
rect 986 1603 1020 1615
rect 986 1547 1020 1565
rect 986 1531 1020 1547
rect 986 1479 1020 1493
rect 986 1459 1020 1479
rect 986 1411 1020 1421
rect 986 1387 1020 1411
rect 986 1343 1020 1349
rect 986 1315 1020 1343
rect 986 1275 1020 1277
rect 986 1243 1020 1275
rect 986 1173 1020 1205
rect 986 1171 1020 1173
rect 986 1105 1020 1133
rect 986 1099 1020 1105
rect 986 1037 1020 1061
rect 986 1027 1020 1037
rect 986 969 1020 989
rect 986 955 1020 969
rect 986 901 1020 917
rect 986 883 1020 901
rect 986 833 1020 845
rect 986 811 1020 833
rect 986 765 1020 773
rect 986 739 1020 765
rect 986 697 1020 701
rect 986 667 1020 697
rect 986 595 1020 629
rect 986 527 1020 557
rect 986 523 1020 527
rect 986 459 1020 485
rect 986 451 1020 459
rect 986 391 1020 413
rect 986 379 1020 391
rect 986 323 1020 341
rect 986 307 1020 323
rect 986 255 1020 269
rect 986 235 1020 255
rect 986 187 1020 197
rect 986 163 1020 187
rect 986 119 1020 125
rect 986 91 1020 119
rect 986 51 1020 53
rect 986 19 1020 51
rect 986 -51 1020 -19
rect 986 -53 1020 -51
rect 986 -119 1020 -91
rect 986 -125 1020 -119
rect 986 -187 1020 -163
rect 986 -197 1020 -187
rect 986 -255 1020 -235
rect 986 -269 1020 -255
rect 986 -323 1020 -307
rect 986 -341 1020 -323
rect 986 -391 1020 -379
rect 986 -413 1020 -391
rect 986 -459 1020 -451
rect 986 -485 1020 -459
rect 986 -527 1020 -523
rect 986 -557 1020 -527
rect 986 -629 1020 -595
rect 986 -697 1020 -667
rect 986 -701 1020 -697
rect 986 -765 1020 -739
rect 986 -773 1020 -765
rect 986 -833 1020 -811
rect 986 -845 1020 -833
rect 986 -901 1020 -883
rect 986 -917 1020 -901
rect 986 -969 1020 -955
rect 986 -989 1020 -969
rect 986 -1037 1020 -1027
rect 986 -1061 1020 -1037
rect 986 -1105 1020 -1099
rect 986 -1133 1020 -1105
rect 986 -1173 1020 -1171
rect 986 -1205 1020 -1173
rect 986 -1275 1020 -1243
rect 986 -1277 1020 -1275
rect 986 -1343 1020 -1315
rect 986 -1349 1020 -1343
rect 986 -1411 1020 -1387
rect 986 -1421 1020 -1411
rect 986 -1479 1020 -1459
rect 986 -1493 1020 -1479
rect 986 -1547 1020 -1531
rect 986 -1565 1020 -1547
rect 986 -1615 1020 -1603
rect 986 -1637 1020 -1615
rect 986 -1683 1020 -1675
rect 986 -1709 1020 -1683
rect 986 -1751 1020 -1747
rect 986 -1781 1020 -1751
rect 986 -1853 1020 -1819
rect 986 -1921 1020 -1891
rect 986 -1925 1020 -1921
rect 986 -1989 1020 -1963
rect 986 -1997 1020 -1989
rect 986 -2057 1020 -2035
rect 986 -2069 1020 -2057
rect 986 -2125 1020 -2107
rect 986 -2141 1020 -2125
rect 986 -2193 1020 -2179
rect 986 -2213 1020 -2193
rect 986 -2261 1020 -2251
rect 986 -2285 1020 -2261
rect 986 -2329 1020 -2323
rect 986 -2357 1020 -2329
rect 986 -2397 1020 -2395
rect 986 -2429 1020 -2397
rect 986 -2499 1020 -2467
rect 986 -2501 1020 -2499
rect 986 -2567 1020 -2539
rect 986 -2573 1020 -2567
rect 986 -2635 1020 -2611
rect 986 -2645 1020 -2635
rect 986 -2703 1020 -2683
rect 986 -2717 1020 -2703
rect 986 -2771 1020 -2755
rect 986 -2789 1020 -2771
rect 986 -2839 1020 -2827
rect 986 -2861 1020 -2839
rect 986 -2907 1020 -2899
rect 986 -2933 1020 -2907
rect 986 -2975 1020 -2971
rect 986 -3005 1020 -2975
rect 986 -3077 1020 -3043
rect 986 -3145 1020 -3115
rect 986 -3149 1020 -3145
rect 986 -3213 1020 -3187
rect 986 -3221 1020 -3213
rect 986 -3281 1020 -3259
rect 986 -3293 1020 -3281
rect 986 -3349 1020 -3331
rect 986 -3365 1020 -3349
rect 986 -3417 1020 -3403
rect 986 -3437 1020 -3417
rect 986 -3485 1020 -3475
rect 986 -3509 1020 -3485
rect 986 -3553 1020 -3547
rect 986 -3581 1020 -3553
rect 986 -3621 1020 -3619
rect 986 -3653 1020 -3621
rect 986 -3723 1020 -3691
rect 986 -3725 1020 -3723
rect 986 -3791 1020 -3763
rect 986 -3797 1020 -3791
rect 986 -3859 1020 -3835
rect 986 -3869 1020 -3859
rect 986 -3927 1020 -3907
rect 986 -3941 1020 -3927
rect 986 -3995 1020 -3979
rect 986 -4013 1020 -3995
rect 986 -4063 1020 -4051
rect 986 -4085 1020 -4063
rect 986 -4131 1020 -4123
rect 986 -4157 1020 -4131
rect 986 -4199 1020 -4195
rect 986 -4229 1020 -4199
rect 986 -4301 1020 -4267
rect 986 -4369 1020 -4339
rect 986 -4373 1020 -4369
rect 986 -4437 1020 -4411
rect 986 -4445 1020 -4437
rect 986 -4505 1020 -4483
rect 986 -4517 1020 -4505
rect 986 -4573 1020 -4555
rect 986 -4589 1020 -4573
rect 986 -4641 1020 -4627
rect 986 -4661 1020 -4641
rect 986 -4709 1020 -4699
rect 986 -4733 1020 -4709
rect 986 -4777 1020 -4771
rect 986 -4805 1020 -4777
rect 986 -4845 1020 -4843
rect 986 -4877 1020 -4845
rect 986 -4947 1020 -4915
rect 986 -4949 1020 -4947
rect 986 -5015 1020 -4987
rect 986 -5021 1020 -5015
rect 986 -5083 1020 -5059
rect 986 -5093 1020 -5083
rect 986 -5151 1020 -5131
rect 986 -5165 1020 -5151
rect 986 -5219 1020 -5203
rect 986 -5237 1020 -5219
rect 986 -5287 1020 -5275
rect 986 -5309 1020 -5287
rect 986 -5355 1020 -5347
rect 986 -5381 1020 -5355
rect 986 -5423 1020 -5419
rect 986 -5453 1020 -5423
rect 986 -5525 1020 -5491
rect 986 -5593 1020 -5563
rect 986 -5597 1020 -5593
rect 986 -5661 1020 -5635
rect 986 -5669 1020 -5661
rect 986 -5729 1020 -5707
rect 986 -5741 1020 -5729
rect 986 -5797 1020 -5779
rect 986 -5813 1020 -5797
rect 986 -5865 1020 -5851
rect 986 -5885 1020 -5865
rect 986 -5933 1020 -5923
rect 986 -5957 1020 -5933
rect 986 -6001 1020 -5995
rect 986 -6029 1020 -6001
rect 986 -6069 1020 -6067
rect 986 -6101 1020 -6069
rect 986 -6171 1020 -6139
rect 986 -6173 1020 -6171
rect 986 -6239 1020 -6211
rect 986 -6245 1020 -6239
rect 986 -6307 1020 -6283
rect 986 -6317 1020 -6307
rect 986 -6375 1020 -6355
rect 986 -6389 1020 -6375
rect 986 -6443 1020 -6427
rect 986 -6461 1020 -6443
rect 986 -6511 1020 -6499
rect 986 -6533 1020 -6511
rect 986 -6579 1020 -6571
rect 986 -6605 1020 -6579
rect 986 -6647 1020 -6643
rect 986 -6677 1020 -6647
rect 986 -6749 1020 -6715
rect 986 -6817 1020 -6787
rect 986 -6821 1020 -6817
rect 986 -6885 1020 -6859
rect 986 -6893 1020 -6885
rect 986 -6953 1020 -6931
rect 986 -6965 1020 -6953
rect 986 -7021 1020 -7003
rect 986 -7037 1020 -7021
rect 986 -7089 1020 -7075
rect 986 -7109 1020 -7089
rect 986 -7157 1020 -7147
rect 986 -7181 1020 -7157
rect 986 -7225 1020 -7219
rect 986 -7253 1020 -7225
rect 986 -7293 1020 -7291
rect 986 -7325 1020 -7293
rect 986 -7395 1020 -7363
rect 986 -7397 1020 -7395
rect 986 -7463 1020 -7435
rect 986 -7469 1020 -7463
rect 986 -7531 1020 -7507
rect 986 -7541 1020 -7531
rect 986 -7599 1020 -7579
rect 986 -7613 1020 -7599
rect 986 -7667 1020 -7651
rect 986 -7685 1020 -7667
rect 986 -7735 1020 -7723
rect 986 -7757 1020 -7735
rect 986 -7803 1020 -7795
rect 986 -7829 1020 -7803
rect 986 -7871 1020 -7867
rect 986 -7901 1020 -7871
rect 986 -7973 1020 -7939
rect 986 -8041 1020 -8011
rect 986 -8045 1020 -8041
rect 986 -8109 1020 -8083
rect 986 -8117 1020 -8109
rect 986 -8177 1020 -8155
rect 986 -8189 1020 -8177
rect 986 -8245 1020 -8227
rect 986 -8261 1020 -8245
rect 986 -8313 1020 -8299
rect 986 -8333 1020 -8313
rect 986 -8381 1020 -8371
rect 986 -8405 1020 -8381
rect 986 -8449 1020 -8443
rect 986 -8477 1020 -8449
rect 986 -8517 1020 -8515
rect 986 -8549 1020 -8517
rect 986 -8619 1020 -8587
rect 986 -8621 1020 -8619
rect 986 -8687 1020 -8659
rect 986 -8693 1020 -8687
rect 986 -8755 1020 -8731
rect 986 -8765 1020 -8755
rect 986 -8823 1020 -8803
rect 986 -8837 1020 -8823
rect 986 -8891 1020 -8875
rect 986 -8909 1020 -8891
rect 986 -8959 1020 -8947
rect 986 -8981 1020 -8959
rect 986 -9027 1020 -9019
rect 986 -9053 1020 -9027
rect 986 -9095 1020 -9091
rect 986 -9125 1020 -9095
rect 986 -9197 1020 -9163
rect 986 -9265 1020 -9235
rect 986 -9269 1020 -9265
rect 986 -9333 1020 -9307
rect 986 -9341 1020 -9333
rect 986 -9401 1020 -9379
rect 986 -9413 1020 -9401
rect 986 -9469 1020 -9451
rect 986 -9485 1020 -9469
rect 986 -9537 1020 -9523
rect 986 -9557 1020 -9537
rect 1104 9537 1138 9557
rect 1104 9523 1138 9537
rect 1104 9469 1138 9485
rect 1104 9451 1138 9469
rect 1104 9401 1138 9413
rect 1104 9379 1138 9401
rect 1104 9333 1138 9341
rect 1104 9307 1138 9333
rect 1104 9265 1138 9269
rect 1104 9235 1138 9265
rect 1104 9163 1138 9197
rect 1104 9095 1138 9125
rect 1104 9091 1138 9095
rect 1104 9027 1138 9053
rect 1104 9019 1138 9027
rect 1104 8959 1138 8981
rect 1104 8947 1138 8959
rect 1104 8891 1138 8909
rect 1104 8875 1138 8891
rect 1104 8823 1138 8837
rect 1104 8803 1138 8823
rect 1104 8755 1138 8765
rect 1104 8731 1138 8755
rect 1104 8687 1138 8693
rect 1104 8659 1138 8687
rect 1104 8619 1138 8621
rect 1104 8587 1138 8619
rect 1104 8517 1138 8549
rect 1104 8515 1138 8517
rect 1104 8449 1138 8477
rect 1104 8443 1138 8449
rect 1104 8381 1138 8405
rect 1104 8371 1138 8381
rect 1104 8313 1138 8333
rect 1104 8299 1138 8313
rect 1104 8245 1138 8261
rect 1104 8227 1138 8245
rect 1104 8177 1138 8189
rect 1104 8155 1138 8177
rect 1104 8109 1138 8117
rect 1104 8083 1138 8109
rect 1104 8041 1138 8045
rect 1104 8011 1138 8041
rect 1104 7939 1138 7973
rect 1104 7871 1138 7901
rect 1104 7867 1138 7871
rect 1104 7803 1138 7829
rect 1104 7795 1138 7803
rect 1104 7735 1138 7757
rect 1104 7723 1138 7735
rect 1104 7667 1138 7685
rect 1104 7651 1138 7667
rect 1104 7599 1138 7613
rect 1104 7579 1138 7599
rect 1104 7531 1138 7541
rect 1104 7507 1138 7531
rect 1104 7463 1138 7469
rect 1104 7435 1138 7463
rect 1104 7395 1138 7397
rect 1104 7363 1138 7395
rect 1104 7293 1138 7325
rect 1104 7291 1138 7293
rect 1104 7225 1138 7253
rect 1104 7219 1138 7225
rect 1104 7157 1138 7181
rect 1104 7147 1138 7157
rect 1104 7089 1138 7109
rect 1104 7075 1138 7089
rect 1104 7021 1138 7037
rect 1104 7003 1138 7021
rect 1104 6953 1138 6965
rect 1104 6931 1138 6953
rect 1104 6885 1138 6893
rect 1104 6859 1138 6885
rect 1104 6817 1138 6821
rect 1104 6787 1138 6817
rect 1104 6715 1138 6749
rect 1104 6647 1138 6677
rect 1104 6643 1138 6647
rect 1104 6579 1138 6605
rect 1104 6571 1138 6579
rect 1104 6511 1138 6533
rect 1104 6499 1138 6511
rect 1104 6443 1138 6461
rect 1104 6427 1138 6443
rect 1104 6375 1138 6389
rect 1104 6355 1138 6375
rect 1104 6307 1138 6317
rect 1104 6283 1138 6307
rect 1104 6239 1138 6245
rect 1104 6211 1138 6239
rect 1104 6171 1138 6173
rect 1104 6139 1138 6171
rect 1104 6069 1138 6101
rect 1104 6067 1138 6069
rect 1104 6001 1138 6029
rect 1104 5995 1138 6001
rect 1104 5933 1138 5957
rect 1104 5923 1138 5933
rect 1104 5865 1138 5885
rect 1104 5851 1138 5865
rect 1104 5797 1138 5813
rect 1104 5779 1138 5797
rect 1104 5729 1138 5741
rect 1104 5707 1138 5729
rect 1104 5661 1138 5669
rect 1104 5635 1138 5661
rect 1104 5593 1138 5597
rect 1104 5563 1138 5593
rect 1104 5491 1138 5525
rect 1104 5423 1138 5453
rect 1104 5419 1138 5423
rect 1104 5355 1138 5381
rect 1104 5347 1138 5355
rect 1104 5287 1138 5309
rect 1104 5275 1138 5287
rect 1104 5219 1138 5237
rect 1104 5203 1138 5219
rect 1104 5151 1138 5165
rect 1104 5131 1138 5151
rect 1104 5083 1138 5093
rect 1104 5059 1138 5083
rect 1104 5015 1138 5021
rect 1104 4987 1138 5015
rect 1104 4947 1138 4949
rect 1104 4915 1138 4947
rect 1104 4845 1138 4877
rect 1104 4843 1138 4845
rect 1104 4777 1138 4805
rect 1104 4771 1138 4777
rect 1104 4709 1138 4733
rect 1104 4699 1138 4709
rect 1104 4641 1138 4661
rect 1104 4627 1138 4641
rect 1104 4573 1138 4589
rect 1104 4555 1138 4573
rect 1104 4505 1138 4517
rect 1104 4483 1138 4505
rect 1104 4437 1138 4445
rect 1104 4411 1138 4437
rect 1104 4369 1138 4373
rect 1104 4339 1138 4369
rect 1104 4267 1138 4301
rect 1104 4199 1138 4229
rect 1104 4195 1138 4199
rect 1104 4131 1138 4157
rect 1104 4123 1138 4131
rect 1104 4063 1138 4085
rect 1104 4051 1138 4063
rect 1104 3995 1138 4013
rect 1104 3979 1138 3995
rect 1104 3927 1138 3941
rect 1104 3907 1138 3927
rect 1104 3859 1138 3869
rect 1104 3835 1138 3859
rect 1104 3791 1138 3797
rect 1104 3763 1138 3791
rect 1104 3723 1138 3725
rect 1104 3691 1138 3723
rect 1104 3621 1138 3653
rect 1104 3619 1138 3621
rect 1104 3553 1138 3581
rect 1104 3547 1138 3553
rect 1104 3485 1138 3509
rect 1104 3475 1138 3485
rect 1104 3417 1138 3437
rect 1104 3403 1138 3417
rect 1104 3349 1138 3365
rect 1104 3331 1138 3349
rect 1104 3281 1138 3293
rect 1104 3259 1138 3281
rect 1104 3213 1138 3221
rect 1104 3187 1138 3213
rect 1104 3145 1138 3149
rect 1104 3115 1138 3145
rect 1104 3043 1138 3077
rect 1104 2975 1138 3005
rect 1104 2971 1138 2975
rect 1104 2907 1138 2933
rect 1104 2899 1138 2907
rect 1104 2839 1138 2861
rect 1104 2827 1138 2839
rect 1104 2771 1138 2789
rect 1104 2755 1138 2771
rect 1104 2703 1138 2717
rect 1104 2683 1138 2703
rect 1104 2635 1138 2645
rect 1104 2611 1138 2635
rect 1104 2567 1138 2573
rect 1104 2539 1138 2567
rect 1104 2499 1138 2501
rect 1104 2467 1138 2499
rect 1104 2397 1138 2429
rect 1104 2395 1138 2397
rect 1104 2329 1138 2357
rect 1104 2323 1138 2329
rect 1104 2261 1138 2285
rect 1104 2251 1138 2261
rect 1104 2193 1138 2213
rect 1104 2179 1138 2193
rect 1104 2125 1138 2141
rect 1104 2107 1138 2125
rect 1104 2057 1138 2069
rect 1104 2035 1138 2057
rect 1104 1989 1138 1997
rect 1104 1963 1138 1989
rect 1104 1921 1138 1925
rect 1104 1891 1138 1921
rect 1104 1819 1138 1853
rect 1104 1751 1138 1781
rect 1104 1747 1138 1751
rect 1104 1683 1138 1709
rect 1104 1675 1138 1683
rect 1104 1615 1138 1637
rect 1104 1603 1138 1615
rect 1104 1547 1138 1565
rect 1104 1531 1138 1547
rect 1104 1479 1138 1493
rect 1104 1459 1138 1479
rect 1104 1411 1138 1421
rect 1104 1387 1138 1411
rect 1104 1343 1138 1349
rect 1104 1315 1138 1343
rect 1104 1275 1138 1277
rect 1104 1243 1138 1275
rect 1104 1173 1138 1205
rect 1104 1171 1138 1173
rect 1104 1105 1138 1133
rect 1104 1099 1138 1105
rect 1104 1037 1138 1061
rect 1104 1027 1138 1037
rect 1104 969 1138 989
rect 1104 955 1138 969
rect 1104 901 1138 917
rect 1104 883 1138 901
rect 1104 833 1138 845
rect 1104 811 1138 833
rect 1104 765 1138 773
rect 1104 739 1138 765
rect 1104 697 1138 701
rect 1104 667 1138 697
rect 1104 595 1138 629
rect 1104 527 1138 557
rect 1104 523 1138 527
rect 1104 459 1138 485
rect 1104 451 1138 459
rect 1104 391 1138 413
rect 1104 379 1138 391
rect 1104 323 1138 341
rect 1104 307 1138 323
rect 1104 255 1138 269
rect 1104 235 1138 255
rect 1104 187 1138 197
rect 1104 163 1138 187
rect 1104 119 1138 125
rect 1104 91 1138 119
rect 1104 51 1138 53
rect 1104 19 1138 51
rect 1104 -51 1138 -19
rect 1104 -53 1138 -51
rect 1104 -119 1138 -91
rect 1104 -125 1138 -119
rect 1104 -187 1138 -163
rect 1104 -197 1138 -187
rect 1104 -255 1138 -235
rect 1104 -269 1138 -255
rect 1104 -323 1138 -307
rect 1104 -341 1138 -323
rect 1104 -391 1138 -379
rect 1104 -413 1138 -391
rect 1104 -459 1138 -451
rect 1104 -485 1138 -459
rect 1104 -527 1138 -523
rect 1104 -557 1138 -527
rect 1104 -629 1138 -595
rect 1104 -697 1138 -667
rect 1104 -701 1138 -697
rect 1104 -765 1138 -739
rect 1104 -773 1138 -765
rect 1104 -833 1138 -811
rect 1104 -845 1138 -833
rect 1104 -901 1138 -883
rect 1104 -917 1138 -901
rect 1104 -969 1138 -955
rect 1104 -989 1138 -969
rect 1104 -1037 1138 -1027
rect 1104 -1061 1138 -1037
rect 1104 -1105 1138 -1099
rect 1104 -1133 1138 -1105
rect 1104 -1173 1138 -1171
rect 1104 -1205 1138 -1173
rect 1104 -1275 1138 -1243
rect 1104 -1277 1138 -1275
rect 1104 -1343 1138 -1315
rect 1104 -1349 1138 -1343
rect 1104 -1411 1138 -1387
rect 1104 -1421 1138 -1411
rect 1104 -1479 1138 -1459
rect 1104 -1493 1138 -1479
rect 1104 -1547 1138 -1531
rect 1104 -1565 1138 -1547
rect 1104 -1615 1138 -1603
rect 1104 -1637 1138 -1615
rect 1104 -1683 1138 -1675
rect 1104 -1709 1138 -1683
rect 1104 -1751 1138 -1747
rect 1104 -1781 1138 -1751
rect 1104 -1853 1138 -1819
rect 1104 -1921 1138 -1891
rect 1104 -1925 1138 -1921
rect 1104 -1989 1138 -1963
rect 1104 -1997 1138 -1989
rect 1104 -2057 1138 -2035
rect 1104 -2069 1138 -2057
rect 1104 -2125 1138 -2107
rect 1104 -2141 1138 -2125
rect 1104 -2193 1138 -2179
rect 1104 -2213 1138 -2193
rect 1104 -2261 1138 -2251
rect 1104 -2285 1138 -2261
rect 1104 -2329 1138 -2323
rect 1104 -2357 1138 -2329
rect 1104 -2397 1138 -2395
rect 1104 -2429 1138 -2397
rect 1104 -2499 1138 -2467
rect 1104 -2501 1138 -2499
rect 1104 -2567 1138 -2539
rect 1104 -2573 1138 -2567
rect 1104 -2635 1138 -2611
rect 1104 -2645 1138 -2635
rect 1104 -2703 1138 -2683
rect 1104 -2717 1138 -2703
rect 1104 -2771 1138 -2755
rect 1104 -2789 1138 -2771
rect 1104 -2839 1138 -2827
rect 1104 -2861 1138 -2839
rect 1104 -2907 1138 -2899
rect 1104 -2933 1138 -2907
rect 1104 -2975 1138 -2971
rect 1104 -3005 1138 -2975
rect 1104 -3077 1138 -3043
rect 1104 -3145 1138 -3115
rect 1104 -3149 1138 -3145
rect 1104 -3213 1138 -3187
rect 1104 -3221 1138 -3213
rect 1104 -3281 1138 -3259
rect 1104 -3293 1138 -3281
rect 1104 -3349 1138 -3331
rect 1104 -3365 1138 -3349
rect 1104 -3417 1138 -3403
rect 1104 -3437 1138 -3417
rect 1104 -3485 1138 -3475
rect 1104 -3509 1138 -3485
rect 1104 -3553 1138 -3547
rect 1104 -3581 1138 -3553
rect 1104 -3621 1138 -3619
rect 1104 -3653 1138 -3621
rect 1104 -3723 1138 -3691
rect 1104 -3725 1138 -3723
rect 1104 -3791 1138 -3763
rect 1104 -3797 1138 -3791
rect 1104 -3859 1138 -3835
rect 1104 -3869 1138 -3859
rect 1104 -3927 1138 -3907
rect 1104 -3941 1138 -3927
rect 1104 -3995 1138 -3979
rect 1104 -4013 1138 -3995
rect 1104 -4063 1138 -4051
rect 1104 -4085 1138 -4063
rect 1104 -4131 1138 -4123
rect 1104 -4157 1138 -4131
rect 1104 -4199 1138 -4195
rect 1104 -4229 1138 -4199
rect 1104 -4301 1138 -4267
rect 1104 -4369 1138 -4339
rect 1104 -4373 1138 -4369
rect 1104 -4437 1138 -4411
rect 1104 -4445 1138 -4437
rect 1104 -4505 1138 -4483
rect 1104 -4517 1138 -4505
rect 1104 -4573 1138 -4555
rect 1104 -4589 1138 -4573
rect 1104 -4641 1138 -4627
rect 1104 -4661 1138 -4641
rect 1104 -4709 1138 -4699
rect 1104 -4733 1138 -4709
rect 1104 -4777 1138 -4771
rect 1104 -4805 1138 -4777
rect 1104 -4845 1138 -4843
rect 1104 -4877 1138 -4845
rect 1104 -4947 1138 -4915
rect 1104 -4949 1138 -4947
rect 1104 -5015 1138 -4987
rect 1104 -5021 1138 -5015
rect 1104 -5083 1138 -5059
rect 1104 -5093 1138 -5083
rect 1104 -5151 1138 -5131
rect 1104 -5165 1138 -5151
rect 1104 -5219 1138 -5203
rect 1104 -5237 1138 -5219
rect 1104 -5287 1138 -5275
rect 1104 -5309 1138 -5287
rect 1104 -5355 1138 -5347
rect 1104 -5381 1138 -5355
rect 1104 -5423 1138 -5419
rect 1104 -5453 1138 -5423
rect 1104 -5525 1138 -5491
rect 1104 -5593 1138 -5563
rect 1104 -5597 1138 -5593
rect 1104 -5661 1138 -5635
rect 1104 -5669 1138 -5661
rect 1104 -5729 1138 -5707
rect 1104 -5741 1138 -5729
rect 1104 -5797 1138 -5779
rect 1104 -5813 1138 -5797
rect 1104 -5865 1138 -5851
rect 1104 -5885 1138 -5865
rect 1104 -5933 1138 -5923
rect 1104 -5957 1138 -5933
rect 1104 -6001 1138 -5995
rect 1104 -6029 1138 -6001
rect 1104 -6069 1138 -6067
rect 1104 -6101 1138 -6069
rect 1104 -6171 1138 -6139
rect 1104 -6173 1138 -6171
rect 1104 -6239 1138 -6211
rect 1104 -6245 1138 -6239
rect 1104 -6307 1138 -6283
rect 1104 -6317 1138 -6307
rect 1104 -6375 1138 -6355
rect 1104 -6389 1138 -6375
rect 1104 -6443 1138 -6427
rect 1104 -6461 1138 -6443
rect 1104 -6511 1138 -6499
rect 1104 -6533 1138 -6511
rect 1104 -6579 1138 -6571
rect 1104 -6605 1138 -6579
rect 1104 -6647 1138 -6643
rect 1104 -6677 1138 -6647
rect 1104 -6749 1138 -6715
rect 1104 -6817 1138 -6787
rect 1104 -6821 1138 -6817
rect 1104 -6885 1138 -6859
rect 1104 -6893 1138 -6885
rect 1104 -6953 1138 -6931
rect 1104 -6965 1138 -6953
rect 1104 -7021 1138 -7003
rect 1104 -7037 1138 -7021
rect 1104 -7089 1138 -7075
rect 1104 -7109 1138 -7089
rect 1104 -7157 1138 -7147
rect 1104 -7181 1138 -7157
rect 1104 -7225 1138 -7219
rect 1104 -7253 1138 -7225
rect 1104 -7293 1138 -7291
rect 1104 -7325 1138 -7293
rect 1104 -7395 1138 -7363
rect 1104 -7397 1138 -7395
rect 1104 -7463 1138 -7435
rect 1104 -7469 1138 -7463
rect 1104 -7531 1138 -7507
rect 1104 -7541 1138 -7531
rect 1104 -7599 1138 -7579
rect 1104 -7613 1138 -7599
rect 1104 -7667 1138 -7651
rect 1104 -7685 1138 -7667
rect 1104 -7735 1138 -7723
rect 1104 -7757 1138 -7735
rect 1104 -7803 1138 -7795
rect 1104 -7829 1138 -7803
rect 1104 -7871 1138 -7867
rect 1104 -7901 1138 -7871
rect 1104 -7973 1138 -7939
rect 1104 -8041 1138 -8011
rect 1104 -8045 1138 -8041
rect 1104 -8109 1138 -8083
rect 1104 -8117 1138 -8109
rect 1104 -8177 1138 -8155
rect 1104 -8189 1138 -8177
rect 1104 -8245 1138 -8227
rect 1104 -8261 1138 -8245
rect 1104 -8313 1138 -8299
rect 1104 -8333 1138 -8313
rect 1104 -8381 1138 -8371
rect 1104 -8405 1138 -8381
rect 1104 -8449 1138 -8443
rect 1104 -8477 1138 -8449
rect 1104 -8517 1138 -8515
rect 1104 -8549 1138 -8517
rect 1104 -8619 1138 -8587
rect 1104 -8621 1138 -8619
rect 1104 -8687 1138 -8659
rect 1104 -8693 1138 -8687
rect 1104 -8755 1138 -8731
rect 1104 -8765 1138 -8755
rect 1104 -8823 1138 -8803
rect 1104 -8837 1138 -8823
rect 1104 -8891 1138 -8875
rect 1104 -8909 1138 -8891
rect 1104 -8959 1138 -8947
rect 1104 -8981 1138 -8959
rect 1104 -9027 1138 -9019
rect 1104 -9053 1138 -9027
rect 1104 -9095 1138 -9091
rect 1104 -9125 1138 -9095
rect 1104 -9197 1138 -9163
rect 1104 -9265 1138 -9235
rect 1104 -9269 1138 -9265
rect 1104 -9333 1138 -9307
rect 1104 -9341 1138 -9333
rect 1104 -9401 1138 -9379
rect 1104 -9413 1138 -9401
rect 1104 -9469 1138 -9451
rect 1104 -9485 1138 -9469
rect 1104 -9537 1138 -9523
rect 1104 -9557 1138 -9537
rect 1222 9537 1256 9557
rect 1222 9523 1256 9537
rect 1222 9469 1256 9485
rect 1222 9451 1256 9469
rect 1222 9401 1256 9413
rect 1222 9379 1256 9401
rect 1222 9333 1256 9341
rect 1222 9307 1256 9333
rect 1222 9265 1256 9269
rect 1222 9235 1256 9265
rect 1222 9163 1256 9197
rect 1222 9095 1256 9125
rect 1222 9091 1256 9095
rect 1222 9027 1256 9053
rect 1222 9019 1256 9027
rect 1222 8959 1256 8981
rect 1222 8947 1256 8959
rect 1222 8891 1256 8909
rect 1222 8875 1256 8891
rect 1222 8823 1256 8837
rect 1222 8803 1256 8823
rect 1222 8755 1256 8765
rect 1222 8731 1256 8755
rect 1222 8687 1256 8693
rect 1222 8659 1256 8687
rect 1222 8619 1256 8621
rect 1222 8587 1256 8619
rect 1222 8517 1256 8549
rect 1222 8515 1256 8517
rect 1222 8449 1256 8477
rect 1222 8443 1256 8449
rect 1222 8381 1256 8405
rect 1222 8371 1256 8381
rect 1222 8313 1256 8333
rect 1222 8299 1256 8313
rect 1222 8245 1256 8261
rect 1222 8227 1256 8245
rect 1222 8177 1256 8189
rect 1222 8155 1256 8177
rect 1222 8109 1256 8117
rect 1222 8083 1256 8109
rect 1222 8041 1256 8045
rect 1222 8011 1256 8041
rect 1222 7939 1256 7973
rect 1222 7871 1256 7901
rect 1222 7867 1256 7871
rect 1222 7803 1256 7829
rect 1222 7795 1256 7803
rect 1222 7735 1256 7757
rect 1222 7723 1256 7735
rect 1222 7667 1256 7685
rect 1222 7651 1256 7667
rect 1222 7599 1256 7613
rect 1222 7579 1256 7599
rect 1222 7531 1256 7541
rect 1222 7507 1256 7531
rect 1222 7463 1256 7469
rect 1222 7435 1256 7463
rect 1222 7395 1256 7397
rect 1222 7363 1256 7395
rect 1222 7293 1256 7325
rect 1222 7291 1256 7293
rect 1222 7225 1256 7253
rect 1222 7219 1256 7225
rect 1222 7157 1256 7181
rect 1222 7147 1256 7157
rect 1222 7089 1256 7109
rect 1222 7075 1256 7089
rect 1222 7021 1256 7037
rect 1222 7003 1256 7021
rect 1222 6953 1256 6965
rect 1222 6931 1256 6953
rect 1222 6885 1256 6893
rect 1222 6859 1256 6885
rect 1222 6817 1256 6821
rect 1222 6787 1256 6817
rect 1222 6715 1256 6749
rect 1222 6647 1256 6677
rect 1222 6643 1256 6647
rect 1222 6579 1256 6605
rect 1222 6571 1256 6579
rect 1222 6511 1256 6533
rect 1222 6499 1256 6511
rect 1222 6443 1256 6461
rect 1222 6427 1256 6443
rect 1222 6375 1256 6389
rect 1222 6355 1256 6375
rect 1222 6307 1256 6317
rect 1222 6283 1256 6307
rect 1222 6239 1256 6245
rect 1222 6211 1256 6239
rect 1222 6171 1256 6173
rect 1222 6139 1256 6171
rect 1222 6069 1256 6101
rect 1222 6067 1256 6069
rect 1222 6001 1256 6029
rect 1222 5995 1256 6001
rect 1222 5933 1256 5957
rect 1222 5923 1256 5933
rect 1222 5865 1256 5885
rect 1222 5851 1256 5865
rect 1222 5797 1256 5813
rect 1222 5779 1256 5797
rect 1222 5729 1256 5741
rect 1222 5707 1256 5729
rect 1222 5661 1256 5669
rect 1222 5635 1256 5661
rect 1222 5593 1256 5597
rect 1222 5563 1256 5593
rect 1222 5491 1256 5525
rect 1222 5423 1256 5453
rect 1222 5419 1256 5423
rect 1222 5355 1256 5381
rect 1222 5347 1256 5355
rect 1222 5287 1256 5309
rect 1222 5275 1256 5287
rect 1222 5219 1256 5237
rect 1222 5203 1256 5219
rect 1222 5151 1256 5165
rect 1222 5131 1256 5151
rect 1222 5083 1256 5093
rect 1222 5059 1256 5083
rect 1222 5015 1256 5021
rect 1222 4987 1256 5015
rect 1222 4947 1256 4949
rect 1222 4915 1256 4947
rect 1222 4845 1256 4877
rect 1222 4843 1256 4845
rect 1222 4777 1256 4805
rect 1222 4771 1256 4777
rect 1222 4709 1256 4733
rect 1222 4699 1256 4709
rect 1222 4641 1256 4661
rect 1222 4627 1256 4641
rect 1222 4573 1256 4589
rect 1222 4555 1256 4573
rect 1222 4505 1256 4517
rect 1222 4483 1256 4505
rect 1222 4437 1256 4445
rect 1222 4411 1256 4437
rect 1222 4369 1256 4373
rect 1222 4339 1256 4369
rect 1222 4267 1256 4301
rect 1222 4199 1256 4229
rect 1222 4195 1256 4199
rect 1222 4131 1256 4157
rect 1222 4123 1256 4131
rect 1222 4063 1256 4085
rect 1222 4051 1256 4063
rect 1222 3995 1256 4013
rect 1222 3979 1256 3995
rect 1222 3927 1256 3941
rect 1222 3907 1256 3927
rect 1222 3859 1256 3869
rect 1222 3835 1256 3859
rect 1222 3791 1256 3797
rect 1222 3763 1256 3791
rect 1222 3723 1256 3725
rect 1222 3691 1256 3723
rect 1222 3621 1256 3653
rect 1222 3619 1256 3621
rect 1222 3553 1256 3581
rect 1222 3547 1256 3553
rect 1222 3485 1256 3509
rect 1222 3475 1256 3485
rect 1222 3417 1256 3437
rect 1222 3403 1256 3417
rect 1222 3349 1256 3365
rect 1222 3331 1256 3349
rect 1222 3281 1256 3293
rect 1222 3259 1256 3281
rect 1222 3213 1256 3221
rect 1222 3187 1256 3213
rect 1222 3145 1256 3149
rect 1222 3115 1256 3145
rect 1222 3043 1256 3077
rect 1222 2975 1256 3005
rect 1222 2971 1256 2975
rect 1222 2907 1256 2933
rect 1222 2899 1256 2907
rect 1222 2839 1256 2861
rect 1222 2827 1256 2839
rect 1222 2771 1256 2789
rect 1222 2755 1256 2771
rect 1222 2703 1256 2717
rect 1222 2683 1256 2703
rect 1222 2635 1256 2645
rect 1222 2611 1256 2635
rect 1222 2567 1256 2573
rect 1222 2539 1256 2567
rect 1222 2499 1256 2501
rect 1222 2467 1256 2499
rect 1222 2397 1256 2429
rect 1222 2395 1256 2397
rect 1222 2329 1256 2357
rect 1222 2323 1256 2329
rect 1222 2261 1256 2285
rect 1222 2251 1256 2261
rect 1222 2193 1256 2213
rect 1222 2179 1256 2193
rect 1222 2125 1256 2141
rect 1222 2107 1256 2125
rect 1222 2057 1256 2069
rect 1222 2035 1256 2057
rect 1222 1989 1256 1997
rect 1222 1963 1256 1989
rect 1222 1921 1256 1925
rect 1222 1891 1256 1921
rect 1222 1819 1256 1853
rect 1222 1751 1256 1781
rect 1222 1747 1256 1751
rect 1222 1683 1256 1709
rect 1222 1675 1256 1683
rect 1222 1615 1256 1637
rect 1222 1603 1256 1615
rect 1222 1547 1256 1565
rect 1222 1531 1256 1547
rect 1222 1479 1256 1493
rect 1222 1459 1256 1479
rect 1222 1411 1256 1421
rect 1222 1387 1256 1411
rect 1222 1343 1256 1349
rect 1222 1315 1256 1343
rect 1222 1275 1256 1277
rect 1222 1243 1256 1275
rect 1222 1173 1256 1205
rect 1222 1171 1256 1173
rect 1222 1105 1256 1133
rect 1222 1099 1256 1105
rect 1222 1037 1256 1061
rect 1222 1027 1256 1037
rect 1222 969 1256 989
rect 1222 955 1256 969
rect 1222 901 1256 917
rect 1222 883 1256 901
rect 1222 833 1256 845
rect 1222 811 1256 833
rect 1222 765 1256 773
rect 1222 739 1256 765
rect 1222 697 1256 701
rect 1222 667 1256 697
rect 1222 595 1256 629
rect 1222 527 1256 557
rect 1222 523 1256 527
rect 1222 459 1256 485
rect 1222 451 1256 459
rect 1222 391 1256 413
rect 1222 379 1256 391
rect 1222 323 1256 341
rect 1222 307 1256 323
rect 1222 255 1256 269
rect 1222 235 1256 255
rect 1222 187 1256 197
rect 1222 163 1256 187
rect 1222 119 1256 125
rect 1222 91 1256 119
rect 1222 51 1256 53
rect 1222 19 1256 51
rect 1222 -51 1256 -19
rect 1222 -53 1256 -51
rect 1222 -119 1256 -91
rect 1222 -125 1256 -119
rect 1222 -187 1256 -163
rect 1222 -197 1256 -187
rect 1222 -255 1256 -235
rect 1222 -269 1256 -255
rect 1222 -323 1256 -307
rect 1222 -341 1256 -323
rect 1222 -391 1256 -379
rect 1222 -413 1256 -391
rect 1222 -459 1256 -451
rect 1222 -485 1256 -459
rect 1222 -527 1256 -523
rect 1222 -557 1256 -527
rect 1222 -629 1256 -595
rect 1222 -697 1256 -667
rect 1222 -701 1256 -697
rect 1222 -765 1256 -739
rect 1222 -773 1256 -765
rect 1222 -833 1256 -811
rect 1222 -845 1256 -833
rect 1222 -901 1256 -883
rect 1222 -917 1256 -901
rect 1222 -969 1256 -955
rect 1222 -989 1256 -969
rect 1222 -1037 1256 -1027
rect 1222 -1061 1256 -1037
rect 1222 -1105 1256 -1099
rect 1222 -1133 1256 -1105
rect 1222 -1173 1256 -1171
rect 1222 -1205 1256 -1173
rect 1222 -1275 1256 -1243
rect 1222 -1277 1256 -1275
rect 1222 -1343 1256 -1315
rect 1222 -1349 1256 -1343
rect 1222 -1411 1256 -1387
rect 1222 -1421 1256 -1411
rect 1222 -1479 1256 -1459
rect 1222 -1493 1256 -1479
rect 1222 -1547 1256 -1531
rect 1222 -1565 1256 -1547
rect 1222 -1615 1256 -1603
rect 1222 -1637 1256 -1615
rect 1222 -1683 1256 -1675
rect 1222 -1709 1256 -1683
rect 1222 -1751 1256 -1747
rect 1222 -1781 1256 -1751
rect 1222 -1853 1256 -1819
rect 1222 -1921 1256 -1891
rect 1222 -1925 1256 -1921
rect 1222 -1989 1256 -1963
rect 1222 -1997 1256 -1989
rect 1222 -2057 1256 -2035
rect 1222 -2069 1256 -2057
rect 1222 -2125 1256 -2107
rect 1222 -2141 1256 -2125
rect 1222 -2193 1256 -2179
rect 1222 -2213 1256 -2193
rect 1222 -2261 1256 -2251
rect 1222 -2285 1256 -2261
rect 1222 -2329 1256 -2323
rect 1222 -2357 1256 -2329
rect 1222 -2397 1256 -2395
rect 1222 -2429 1256 -2397
rect 1222 -2499 1256 -2467
rect 1222 -2501 1256 -2499
rect 1222 -2567 1256 -2539
rect 1222 -2573 1256 -2567
rect 1222 -2635 1256 -2611
rect 1222 -2645 1256 -2635
rect 1222 -2703 1256 -2683
rect 1222 -2717 1256 -2703
rect 1222 -2771 1256 -2755
rect 1222 -2789 1256 -2771
rect 1222 -2839 1256 -2827
rect 1222 -2861 1256 -2839
rect 1222 -2907 1256 -2899
rect 1222 -2933 1256 -2907
rect 1222 -2975 1256 -2971
rect 1222 -3005 1256 -2975
rect 1222 -3077 1256 -3043
rect 1222 -3145 1256 -3115
rect 1222 -3149 1256 -3145
rect 1222 -3213 1256 -3187
rect 1222 -3221 1256 -3213
rect 1222 -3281 1256 -3259
rect 1222 -3293 1256 -3281
rect 1222 -3349 1256 -3331
rect 1222 -3365 1256 -3349
rect 1222 -3417 1256 -3403
rect 1222 -3437 1256 -3417
rect 1222 -3485 1256 -3475
rect 1222 -3509 1256 -3485
rect 1222 -3553 1256 -3547
rect 1222 -3581 1256 -3553
rect 1222 -3621 1256 -3619
rect 1222 -3653 1256 -3621
rect 1222 -3723 1256 -3691
rect 1222 -3725 1256 -3723
rect 1222 -3791 1256 -3763
rect 1222 -3797 1256 -3791
rect 1222 -3859 1256 -3835
rect 1222 -3869 1256 -3859
rect 1222 -3927 1256 -3907
rect 1222 -3941 1256 -3927
rect 1222 -3995 1256 -3979
rect 1222 -4013 1256 -3995
rect 1222 -4063 1256 -4051
rect 1222 -4085 1256 -4063
rect 1222 -4131 1256 -4123
rect 1222 -4157 1256 -4131
rect 1222 -4199 1256 -4195
rect 1222 -4229 1256 -4199
rect 1222 -4301 1256 -4267
rect 1222 -4369 1256 -4339
rect 1222 -4373 1256 -4369
rect 1222 -4437 1256 -4411
rect 1222 -4445 1256 -4437
rect 1222 -4505 1256 -4483
rect 1222 -4517 1256 -4505
rect 1222 -4573 1256 -4555
rect 1222 -4589 1256 -4573
rect 1222 -4641 1256 -4627
rect 1222 -4661 1256 -4641
rect 1222 -4709 1256 -4699
rect 1222 -4733 1256 -4709
rect 1222 -4777 1256 -4771
rect 1222 -4805 1256 -4777
rect 1222 -4845 1256 -4843
rect 1222 -4877 1256 -4845
rect 1222 -4947 1256 -4915
rect 1222 -4949 1256 -4947
rect 1222 -5015 1256 -4987
rect 1222 -5021 1256 -5015
rect 1222 -5083 1256 -5059
rect 1222 -5093 1256 -5083
rect 1222 -5151 1256 -5131
rect 1222 -5165 1256 -5151
rect 1222 -5219 1256 -5203
rect 1222 -5237 1256 -5219
rect 1222 -5287 1256 -5275
rect 1222 -5309 1256 -5287
rect 1222 -5355 1256 -5347
rect 1222 -5381 1256 -5355
rect 1222 -5423 1256 -5419
rect 1222 -5453 1256 -5423
rect 1222 -5525 1256 -5491
rect 1222 -5593 1256 -5563
rect 1222 -5597 1256 -5593
rect 1222 -5661 1256 -5635
rect 1222 -5669 1256 -5661
rect 1222 -5729 1256 -5707
rect 1222 -5741 1256 -5729
rect 1222 -5797 1256 -5779
rect 1222 -5813 1256 -5797
rect 1222 -5865 1256 -5851
rect 1222 -5885 1256 -5865
rect 1222 -5933 1256 -5923
rect 1222 -5957 1256 -5933
rect 1222 -6001 1256 -5995
rect 1222 -6029 1256 -6001
rect 1222 -6069 1256 -6067
rect 1222 -6101 1256 -6069
rect 1222 -6171 1256 -6139
rect 1222 -6173 1256 -6171
rect 1222 -6239 1256 -6211
rect 1222 -6245 1256 -6239
rect 1222 -6307 1256 -6283
rect 1222 -6317 1256 -6307
rect 1222 -6375 1256 -6355
rect 1222 -6389 1256 -6375
rect 1222 -6443 1256 -6427
rect 1222 -6461 1256 -6443
rect 1222 -6511 1256 -6499
rect 1222 -6533 1256 -6511
rect 1222 -6579 1256 -6571
rect 1222 -6605 1256 -6579
rect 1222 -6647 1256 -6643
rect 1222 -6677 1256 -6647
rect 1222 -6749 1256 -6715
rect 1222 -6817 1256 -6787
rect 1222 -6821 1256 -6817
rect 1222 -6885 1256 -6859
rect 1222 -6893 1256 -6885
rect 1222 -6953 1256 -6931
rect 1222 -6965 1256 -6953
rect 1222 -7021 1256 -7003
rect 1222 -7037 1256 -7021
rect 1222 -7089 1256 -7075
rect 1222 -7109 1256 -7089
rect 1222 -7157 1256 -7147
rect 1222 -7181 1256 -7157
rect 1222 -7225 1256 -7219
rect 1222 -7253 1256 -7225
rect 1222 -7293 1256 -7291
rect 1222 -7325 1256 -7293
rect 1222 -7395 1256 -7363
rect 1222 -7397 1256 -7395
rect 1222 -7463 1256 -7435
rect 1222 -7469 1256 -7463
rect 1222 -7531 1256 -7507
rect 1222 -7541 1256 -7531
rect 1222 -7599 1256 -7579
rect 1222 -7613 1256 -7599
rect 1222 -7667 1256 -7651
rect 1222 -7685 1256 -7667
rect 1222 -7735 1256 -7723
rect 1222 -7757 1256 -7735
rect 1222 -7803 1256 -7795
rect 1222 -7829 1256 -7803
rect 1222 -7871 1256 -7867
rect 1222 -7901 1256 -7871
rect 1222 -7973 1256 -7939
rect 1222 -8041 1256 -8011
rect 1222 -8045 1256 -8041
rect 1222 -8109 1256 -8083
rect 1222 -8117 1256 -8109
rect 1222 -8177 1256 -8155
rect 1222 -8189 1256 -8177
rect 1222 -8245 1256 -8227
rect 1222 -8261 1256 -8245
rect 1222 -8313 1256 -8299
rect 1222 -8333 1256 -8313
rect 1222 -8381 1256 -8371
rect 1222 -8405 1256 -8381
rect 1222 -8449 1256 -8443
rect 1222 -8477 1256 -8449
rect 1222 -8517 1256 -8515
rect 1222 -8549 1256 -8517
rect 1222 -8619 1256 -8587
rect 1222 -8621 1256 -8619
rect 1222 -8687 1256 -8659
rect 1222 -8693 1256 -8687
rect 1222 -8755 1256 -8731
rect 1222 -8765 1256 -8755
rect 1222 -8823 1256 -8803
rect 1222 -8837 1256 -8823
rect 1222 -8891 1256 -8875
rect 1222 -8909 1256 -8891
rect 1222 -8959 1256 -8947
rect 1222 -8981 1256 -8959
rect 1222 -9027 1256 -9019
rect 1222 -9053 1256 -9027
rect 1222 -9095 1256 -9091
rect 1222 -9125 1256 -9095
rect 1222 -9197 1256 -9163
rect 1222 -9265 1256 -9235
rect 1222 -9269 1256 -9265
rect 1222 -9333 1256 -9307
rect 1222 -9341 1256 -9333
rect 1222 -9401 1256 -9379
rect 1222 -9413 1256 -9401
rect 1222 -9469 1256 -9451
rect 1222 -9485 1256 -9469
rect 1222 -9537 1256 -9523
rect 1222 -9557 1256 -9537
rect 1340 9537 1374 9557
rect 1340 9523 1374 9537
rect 1340 9469 1374 9485
rect 1340 9451 1374 9469
rect 1340 9401 1374 9413
rect 1340 9379 1374 9401
rect 1340 9333 1374 9341
rect 1340 9307 1374 9333
rect 1340 9265 1374 9269
rect 1340 9235 1374 9265
rect 1340 9163 1374 9197
rect 1340 9095 1374 9125
rect 1340 9091 1374 9095
rect 1340 9027 1374 9053
rect 1340 9019 1374 9027
rect 1340 8959 1374 8981
rect 1340 8947 1374 8959
rect 1340 8891 1374 8909
rect 1340 8875 1374 8891
rect 1340 8823 1374 8837
rect 1340 8803 1374 8823
rect 1340 8755 1374 8765
rect 1340 8731 1374 8755
rect 1340 8687 1374 8693
rect 1340 8659 1374 8687
rect 1340 8619 1374 8621
rect 1340 8587 1374 8619
rect 1340 8517 1374 8549
rect 1340 8515 1374 8517
rect 1340 8449 1374 8477
rect 1340 8443 1374 8449
rect 1340 8381 1374 8405
rect 1340 8371 1374 8381
rect 1340 8313 1374 8333
rect 1340 8299 1374 8313
rect 1340 8245 1374 8261
rect 1340 8227 1374 8245
rect 1340 8177 1374 8189
rect 1340 8155 1374 8177
rect 1340 8109 1374 8117
rect 1340 8083 1374 8109
rect 1340 8041 1374 8045
rect 1340 8011 1374 8041
rect 1340 7939 1374 7973
rect 1340 7871 1374 7901
rect 1340 7867 1374 7871
rect 1340 7803 1374 7829
rect 1340 7795 1374 7803
rect 1340 7735 1374 7757
rect 1340 7723 1374 7735
rect 1340 7667 1374 7685
rect 1340 7651 1374 7667
rect 1340 7599 1374 7613
rect 1340 7579 1374 7599
rect 1340 7531 1374 7541
rect 1340 7507 1374 7531
rect 1340 7463 1374 7469
rect 1340 7435 1374 7463
rect 1340 7395 1374 7397
rect 1340 7363 1374 7395
rect 1340 7293 1374 7325
rect 1340 7291 1374 7293
rect 1340 7225 1374 7253
rect 1340 7219 1374 7225
rect 1340 7157 1374 7181
rect 1340 7147 1374 7157
rect 1340 7089 1374 7109
rect 1340 7075 1374 7089
rect 1340 7021 1374 7037
rect 1340 7003 1374 7021
rect 1340 6953 1374 6965
rect 1340 6931 1374 6953
rect 1340 6885 1374 6893
rect 1340 6859 1374 6885
rect 1340 6817 1374 6821
rect 1340 6787 1374 6817
rect 1340 6715 1374 6749
rect 1340 6647 1374 6677
rect 1340 6643 1374 6647
rect 1340 6579 1374 6605
rect 1340 6571 1374 6579
rect 1340 6511 1374 6533
rect 1340 6499 1374 6511
rect 1340 6443 1374 6461
rect 1340 6427 1374 6443
rect 1340 6375 1374 6389
rect 1340 6355 1374 6375
rect 1340 6307 1374 6317
rect 1340 6283 1374 6307
rect 1340 6239 1374 6245
rect 1340 6211 1374 6239
rect 1340 6171 1374 6173
rect 1340 6139 1374 6171
rect 1340 6069 1374 6101
rect 1340 6067 1374 6069
rect 1340 6001 1374 6029
rect 1340 5995 1374 6001
rect 1340 5933 1374 5957
rect 1340 5923 1374 5933
rect 1340 5865 1374 5885
rect 1340 5851 1374 5865
rect 1340 5797 1374 5813
rect 1340 5779 1374 5797
rect 1340 5729 1374 5741
rect 1340 5707 1374 5729
rect 1340 5661 1374 5669
rect 1340 5635 1374 5661
rect 1340 5593 1374 5597
rect 1340 5563 1374 5593
rect 1340 5491 1374 5525
rect 1340 5423 1374 5453
rect 1340 5419 1374 5423
rect 1340 5355 1374 5381
rect 1340 5347 1374 5355
rect 1340 5287 1374 5309
rect 1340 5275 1374 5287
rect 1340 5219 1374 5237
rect 1340 5203 1374 5219
rect 1340 5151 1374 5165
rect 1340 5131 1374 5151
rect 1340 5083 1374 5093
rect 1340 5059 1374 5083
rect 1340 5015 1374 5021
rect 1340 4987 1374 5015
rect 1340 4947 1374 4949
rect 1340 4915 1374 4947
rect 1340 4845 1374 4877
rect 1340 4843 1374 4845
rect 1340 4777 1374 4805
rect 1340 4771 1374 4777
rect 1340 4709 1374 4733
rect 1340 4699 1374 4709
rect 1340 4641 1374 4661
rect 1340 4627 1374 4641
rect 1340 4573 1374 4589
rect 1340 4555 1374 4573
rect 1340 4505 1374 4517
rect 1340 4483 1374 4505
rect 1340 4437 1374 4445
rect 1340 4411 1374 4437
rect 1340 4369 1374 4373
rect 1340 4339 1374 4369
rect 1340 4267 1374 4301
rect 1340 4199 1374 4229
rect 1340 4195 1374 4199
rect 1340 4131 1374 4157
rect 1340 4123 1374 4131
rect 1340 4063 1374 4085
rect 1340 4051 1374 4063
rect 1340 3995 1374 4013
rect 1340 3979 1374 3995
rect 1340 3927 1374 3941
rect 1340 3907 1374 3927
rect 1340 3859 1374 3869
rect 1340 3835 1374 3859
rect 1340 3791 1374 3797
rect 1340 3763 1374 3791
rect 1340 3723 1374 3725
rect 1340 3691 1374 3723
rect 1340 3621 1374 3653
rect 1340 3619 1374 3621
rect 1340 3553 1374 3581
rect 1340 3547 1374 3553
rect 1340 3485 1374 3509
rect 1340 3475 1374 3485
rect 1340 3417 1374 3437
rect 1340 3403 1374 3417
rect 1340 3349 1374 3365
rect 1340 3331 1374 3349
rect 1340 3281 1374 3293
rect 1340 3259 1374 3281
rect 1340 3213 1374 3221
rect 1340 3187 1374 3213
rect 1340 3145 1374 3149
rect 1340 3115 1374 3145
rect 1340 3043 1374 3077
rect 1340 2975 1374 3005
rect 1340 2971 1374 2975
rect 1340 2907 1374 2933
rect 1340 2899 1374 2907
rect 1340 2839 1374 2861
rect 1340 2827 1374 2839
rect 1340 2771 1374 2789
rect 1340 2755 1374 2771
rect 1340 2703 1374 2717
rect 1340 2683 1374 2703
rect 1340 2635 1374 2645
rect 1340 2611 1374 2635
rect 1340 2567 1374 2573
rect 1340 2539 1374 2567
rect 1340 2499 1374 2501
rect 1340 2467 1374 2499
rect 1340 2397 1374 2429
rect 1340 2395 1374 2397
rect 1340 2329 1374 2357
rect 1340 2323 1374 2329
rect 1340 2261 1374 2285
rect 1340 2251 1374 2261
rect 1340 2193 1374 2213
rect 1340 2179 1374 2193
rect 1340 2125 1374 2141
rect 1340 2107 1374 2125
rect 1340 2057 1374 2069
rect 1340 2035 1374 2057
rect 1340 1989 1374 1997
rect 1340 1963 1374 1989
rect 1340 1921 1374 1925
rect 1340 1891 1374 1921
rect 1340 1819 1374 1853
rect 1340 1751 1374 1781
rect 1340 1747 1374 1751
rect 1340 1683 1374 1709
rect 1340 1675 1374 1683
rect 1340 1615 1374 1637
rect 1340 1603 1374 1615
rect 1340 1547 1374 1565
rect 1340 1531 1374 1547
rect 1340 1479 1374 1493
rect 1340 1459 1374 1479
rect 1340 1411 1374 1421
rect 1340 1387 1374 1411
rect 1340 1343 1374 1349
rect 1340 1315 1374 1343
rect 1340 1275 1374 1277
rect 1340 1243 1374 1275
rect 1340 1173 1374 1205
rect 1340 1171 1374 1173
rect 1340 1105 1374 1133
rect 1340 1099 1374 1105
rect 1340 1037 1374 1061
rect 1340 1027 1374 1037
rect 1340 969 1374 989
rect 1340 955 1374 969
rect 1340 901 1374 917
rect 1340 883 1374 901
rect 1340 833 1374 845
rect 1340 811 1374 833
rect 1340 765 1374 773
rect 1340 739 1374 765
rect 1340 697 1374 701
rect 1340 667 1374 697
rect 1340 595 1374 629
rect 1340 527 1374 557
rect 1340 523 1374 527
rect 1340 459 1374 485
rect 1340 451 1374 459
rect 1340 391 1374 413
rect 1340 379 1374 391
rect 1340 323 1374 341
rect 1340 307 1374 323
rect 1340 255 1374 269
rect 1340 235 1374 255
rect 1340 187 1374 197
rect 1340 163 1374 187
rect 1340 119 1374 125
rect 1340 91 1374 119
rect 1340 51 1374 53
rect 1340 19 1374 51
rect 1340 -51 1374 -19
rect 1340 -53 1374 -51
rect 1340 -119 1374 -91
rect 1340 -125 1374 -119
rect 1340 -187 1374 -163
rect 1340 -197 1374 -187
rect 1340 -255 1374 -235
rect 1340 -269 1374 -255
rect 1340 -323 1374 -307
rect 1340 -341 1374 -323
rect 1340 -391 1374 -379
rect 1340 -413 1374 -391
rect 1340 -459 1374 -451
rect 1340 -485 1374 -459
rect 1340 -527 1374 -523
rect 1340 -557 1374 -527
rect 1340 -629 1374 -595
rect 1340 -697 1374 -667
rect 1340 -701 1374 -697
rect 1340 -765 1374 -739
rect 1340 -773 1374 -765
rect 1340 -833 1374 -811
rect 1340 -845 1374 -833
rect 1340 -901 1374 -883
rect 1340 -917 1374 -901
rect 1340 -969 1374 -955
rect 1340 -989 1374 -969
rect 1340 -1037 1374 -1027
rect 1340 -1061 1374 -1037
rect 1340 -1105 1374 -1099
rect 1340 -1133 1374 -1105
rect 1340 -1173 1374 -1171
rect 1340 -1205 1374 -1173
rect 1340 -1275 1374 -1243
rect 1340 -1277 1374 -1275
rect 1340 -1343 1374 -1315
rect 1340 -1349 1374 -1343
rect 1340 -1411 1374 -1387
rect 1340 -1421 1374 -1411
rect 1340 -1479 1374 -1459
rect 1340 -1493 1374 -1479
rect 1340 -1547 1374 -1531
rect 1340 -1565 1374 -1547
rect 1340 -1615 1374 -1603
rect 1340 -1637 1374 -1615
rect 1340 -1683 1374 -1675
rect 1340 -1709 1374 -1683
rect 1340 -1751 1374 -1747
rect 1340 -1781 1374 -1751
rect 1340 -1853 1374 -1819
rect 1340 -1921 1374 -1891
rect 1340 -1925 1374 -1921
rect 1340 -1989 1374 -1963
rect 1340 -1997 1374 -1989
rect 1340 -2057 1374 -2035
rect 1340 -2069 1374 -2057
rect 1340 -2125 1374 -2107
rect 1340 -2141 1374 -2125
rect 1340 -2193 1374 -2179
rect 1340 -2213 1374 -2193
rect 1340 -2261 1374 -2251
rect 1340 -2285 1374 -2261
rect 1340 -2329 1374 -2323
rect 1340 -2357 1374 -2329
rect 1340 -2397 1374 -2395
rect 1340 -2429 1374 -2397
rect 1340 -2499 1374 -2467
rect 1340 -2501 1374 -2499
rect 1340 -2567 1374 -2539
rect 1340 -2573 1374 -2567
rect 1340 -2635 1374 -2611
rect 1340 -2645 1374 -2635
rect 1340 -2703 1374 -2683
rect 1340 -2717 1374 -2703
rect 1340 -2771 1374 -2755
rect 1340 -2789 1374 -2771
rect 1340 -2839 1374 -2827
rect 1340 -2861 1374 -2839
rect 1340 -2907 1374 -2899
rect 1340 -2933 1374 -2907
rect 1340 -2975 1374 -2971
rect 1340 -3005 1374 -2975
rect 1340 -3077 1374 -3043
rect 1340 -3145 1374 -3115
rect 1340 -3149 1374 -3145
rect 1340 -3213 1374 -3187
rect 1340 -3221 1374 -3213
rect 1340 -3281 1374 -3259
rect 1340 -3293 1374 -3281
rect 1340 -3349 1374 -3331
rect 1340 -3365 1374 -3349
rect 1340 -3417 1374 -3403
rect 1340 -3437 1374 -3417
rect 1340 -3485 1374 -3475
rect 1340 -3509 1374 -3485
rect 1340 -3553 1374 -3547
rect 1340 -3581 1374 -3553
rect 1340 -3621 1374 -3619
rect 1340 -3653 1374 -3621
rect 1340 -3723 1374 -3691
rect 1340 -3725 1374 -3723
rect 1340 -3791 1374 -3763
rect 1340 -3797 1374 -3791
rect 1340 -3859 1374 -3835
rect 1340 -3869 1374 -3859
rect 1340 -3927 1374 -3907
rect 1340 -3941 1374 -3927
rect 1340 -3995 1374 -3979
rect 1340 -4013 1374 -3995
rect 1340 -4063 1374 -4051
rect 1340 -4085 1374 -4063
rect 1340 -4131 1374 -4123
rect 1340 -4157 1374 -4131
rect 1340 -4199 1374 -4195
rect 1340 -4229 1374 -4199
rect 1340 -4301 1374 -4267
rect 1340 -4369 1374 -4339
rect 1340 -4373 1374 -4369
rect 1340 -4437 1374 -4411
rect 1340 -4445 1374 -4437
rect 1340 -4505 1374 -4483
rect 1340 -4517 1374 -4505
rect 1340 -4573 1374 -4555
rect 1340 -4589 1374 -4573
rect 1340 -4641 1374 -4627
rect 1340 -4661 1374 -4641
rect 1340 -4709 1374 -4699
rect 1340 -4733 1374 -4709
rect 1340 -4777 1374 -4771
rect 1340 -4805 1374 -4777
rect 1340 -4845 1374 -4843
rect 1340 -4877 1374 -4845
rect 1340 -4947 1374 -4915
rect 1340 -4949 1374 -4947
rect 1340 -5015 1374 -4987
rect 1340 -5021 1374 -5015
rect 1340 -5083 1374 -5059
rect 1340 -5093 1374 -5083
rect 1340 -5151 1374 -5131
rect 1340 -5165 1374 -5151
rect 1340 -5219 1374 -5203
rect 1340 -5237 1374 -5219
rect 1340 -5287 1374 -5275
rect 1340 -5309 1374 -5287
rect 1340 -5355 1374 -5347
rect 1340 -5381 1374 -5355
rect 1340 -5423 1374 -5419
rect 1340 -5453 1374 -5423
rect 1340 -5525 1374 -5491
rect 1340 -5593 1374 -5563
rect 1340 -5597 1374 -5593
rect 1340 -5661 1374 -5635
rect 1340 -5669 1374 -5661
rect 1340 -5729 1374 -5707
rect 1340 -5741 1374 -5729
rect 1340 -5797 1374 -5779
rect 1340 -5813 1374 -5797
rect 1340 -5865 1374 -5851
rect 1340 -5885 1374 -5865
rect 1340 -5933 1374 -5923
rect 1340 -5957 1374 -5933
rect 1340 -6001 1374 -5995
rect 1340 -6029 1374 -6001
rect 1340 -6069 1374 -6067
rect 1340 -6101 1374 -6069
rect 1340 -6171 1374 -6139
rect 1340 -6173 1374 -6171
rect 1340 -6239 1374 -6211
rect 1340 -6245 1374 -6239
rect 1340 -6307 1374 -6283
rect 1340 -6317 1374 -6307
rect 1340 -6375 1374 -6355
rect 1340 -6389 1374 -6375
rect 1340 -6443 1374 -6427
rect 1340 -6461 1374 -6443
rect 1340 -6511 1374 -6499
rect 1340 -6533 1374 -6511
rect 1340 -6579 1374 -6571
rect 1340 -6605 1374 -6579
rect 1340 -6647 1374 -6643
rect 1340 -6677 1374 -6647
rect 1340 -6749 1374 -6715
rect 1340 -6817 1374 -6787
rect 1340 -6821 1374 -6817
rect 1340 -6885 1374 -6859
rect 1340 -6893 1374 -6885
rect 1340 -6953 1374 -6931
rect 1340 -6965 1374 -6953
rect 1340 -7021 1374 -7003
rect 1340 -7037 1374 -7021
rect 1340 -7089 1374 -7075
rect 1340 -7109 1374 -7089
rect 1340 -7157 1374 -7147
rect 1340 -7181 1374 -7157
rect 1340 -7225 1374 -7219
rect 1340 -7253 1374 -7225
rect 1340 -7293 1374 -7291
rect 1340 -7325 1374 -7293
rect 1340 -7395 1374 -7363
rect 1340 -7397 1374 -7395
rect 1340 -7463 1374 -7435
rect 1340 -7469 1374 -7463
rect 1340 -7531 1374 -7507
rect 1340 -7541 1374 -7531
rect 1340 -7599 1374 -7579
rect 1340 -7613 1374 -7599
rect 1340 -7667 1374 -7651
rect 1340 -7685 1374 -7667
rect 1340 -7735 1374 -7723
rect 1340 -7757 1374 -7735
rect 1340 -7803 1374 -7795
rect 1340 -7829 1374 -7803
rect 1340 -7871 1374 -7867
rect 1340 -7901 1374 -7871
rect 1340 -7973 1374 -7939
rect 1340 -8041 1374 -8011
rect 1340 -8045 1374 -8041
rect 1340 -8109 1374 -8083
rect 1340 -8117 1374 -8109
rect 1340 -8177 1374 -8155
rect 1340 -8189 1374 -8177
rect 1340 -8245 1374 -8227
rect 1340 -8261 1374 -8245
rect 1340 -8313 1374 -8299
rect 1340 -8333 1374 -8313
rect 1340 -8381 1374 -8371
rect 1340 -8405 1374 -8381
rect 1340 -8449 1374 -8443
rect 1340 -8477 1374 -8449
rect 1340 -8517 1374 -8515
rect 1340 -8549 1374 -8517
rect 1340 -8619 1374 -8587
rect 1340 -8621 1374 -8619
rect 1340 -8687 1374 -8659
rect 1340 -8693 1374 -8687
rect 1340 -8755 1374 -8731
rect 1340 -8765 1374 -8755
rect 1340 -8823 1374 -8803
rect 1340 -8837 1374 -8823
rect 1340 -8891 1374 -8875
rect 1340 -8909 1374 -8891
rect 1340 -8959 1374 -8947
rect 1340 -8981 1374 -8959
rect 1340 -9027 1374 -9019
rect 1340 -9053 1374 -9027
rect 1340 -9095 1374 -9091
rect 1340 -9125 1374 -9095
rect 1340 -9197 1374 -9163
rect 1340 -9265 1374 -9235
rect 1340 -9269 1374 -9265
rect 1340 -9333 1374 -9307
rect 1340 -9341 1374 -9333
rect 1340 -9401 1374 -9379
rect 1340 -9413 1374 -9401
rect 1340 -9469 1374 -9451
rect 1340 -9485 1374 -9469
rect 1340 -9537 1374 -9523
rect 1340 -9557 1374 -9537
rect 1458 9537 1492 9557
rect 1458 9523 1492 9537
rect 1458 9469 1492 9485
rect 1458 9451 1492 9469
rect 1458 9401 1492 9413
rect 1458 9379 1492 9401
rect 1458 9333 1492 9341
rect 1458 9307 1492 9333
rect 1458 9265 1492 9269
rect 1458 9235 1492 9265
rect 1458 9163 1492 9197
rect 1458 9095 1492 9125
rect 1458 9091 1492 9095
rect 1458 9027 1492 9053
rect 1458 9019 1492 9027
rect 1458 8959 1492 8981
rect 1458 8947 1492 8959
rect 1458 8891 1492 8909
rect 1458 8875 1492 8891
rect 1458 8823 1492 8837
rect 1458 8803 1492 8823
rect 1458 8755 1492 8765
rect 1458 8731 1492 8755
rect 1458 8687 1492 8693
rect 1458 8659 1492 8687
rect 1458 8619 1492 8621
rect 1458 8587 1492 8619
rect 1458 8517 1492 8549
rect 1458 8515 1492 8517
rect 1458 8449 1492 8477
rect 1458 8443 1492 8449
rect 1458 8381 1492 8405
rect 1458 8371 1492 8381
rect 1458 8313 1492 8333
rect 1458 8299 1492 8313
rect 1458 8245 1492 8261
rect 1458 8227 1492 8245
rect 1458 8177 1492 8189
rect 1458 8155 1492 8177
rect 1458 8109 1492 8117
rect 1458 8083 1492 8109
rect 1458 8041 1492 8045
rect 1458 8011 1492 8041
rect 1458 7939 1492 7973
rect 1458 7871 1492 7901
rect 1458 7867 1492 7871
rect 1458 7803 1492 7829
rect 1458 7795 1492 7803
rect 1458 7735 1492 7757
rect 1458 7723 1492 7735
rect 1458 7667 1492 7685
rect 1458 7651 1492 7667
rect 1458 7599 1492 7613
rect 1458 7579 1492 7599
rect 1458 7531 1492 7541
rect 1458 7507 1492 7531
rect 1458 7463 1492 7469
rect 1458 7435 1492 7463
rect 1458 7395 1492 7397
rect 1458 7363 1492 7395
rect 1458 7293 1492 7325
rect 1458 7291 1492 7293
rect 1458 7225 1492 7253
rect 1458 7219 1492 7225
rect 1458 7157 1492 7181
rect 1458 7147 1492 7157
rect 1458 7089 1492 7109
rect 1458 7075 1492 7089
rect 1458 7021 1492 7037
rect 1458 7003 1492 7021
rect 1458 6953 1492 6965
rect 1458 6931 1492 6953
rect 1458 6885 1492 6893
rect 1458 6859 1492 6885
rect 1458 6817 1492 6821
rect 1458 6787 1492 6817
rect 1458 6715 1492 6749
rect 1458 6647 1492 6677
rect 1458 6643 1492 6647
rect 1458 6579 1492 6605
rect 1458 6571 1492 6579
rect 1458 6511 1492 6533
rect 1458 6499 1492 6511
rect 1458 6443 1492 6461
rect 1458 6427 1492 6443
rect 1458 6375 1492 6389
rect 1458 6355 1492 6375
rect 1458 6307 1492 6317
rect 1458 6283 1492 6307
rect 1458 6239 1492 6245
rect 1458 6211 1492 6239
rect 1458 6171 1492 6173
rect 1458 6139 1492 6171
rect 1458 6069 1492 6101
rect 1458 6067 1492 6069
rect 1458 6001 1492 6029
rect 1458 5995 1492 6001
rect 1458 5933 1492 5957
rect 1458 5923 1492 5933
rect 1458 5865 1492 5885
rect 1458 5851 1492 5865
rect 1458 5797 1492 5813
rect 1458 5779 1492 5797
rect 1458 5729 1492 5741
rect 1458 5707 1492 5729
rect 1458 5661 1492 5669
rect 1458 5635 1492 5661
rect 1458 5593 1492 5597
rect 1458 5563 1492 5593
rect 1458 5491 1492 5525
rect 1458 5423 1492 5453
rect 1458 5419 1492 5423
rect 1458 5355 1492 5381
rect 1458 5347 1492 5355
rect 1458 5287 1492 5309
rect 1458 5275 1492 5287
rect 1458 5219 1492 5237
rect 1458 5203 1492 5219
rect 1458 5151 1492 5165
rect 1458 5131 1492 5151
rect 1458 5083 1492 5093
rect 1458 5059 1492 5083
rect 1458 5015 1492 5021
rect 1458 4987 1492 5015
rect 1458 4947 1492 4949
rect 1458 4915 1492 4947
rect 1458 4845 1492 4877
rect 1458 4843 1492 4845
rect 1458 4777 1492 4805
rect 1458 4771 1492 4777
rect 1458 4709 1492 4733
rect 1458 4699 1492 4709
rect 1458 4641 1492 4661
rect 1458 4627 1492 4641
rect 1458 4573 1492 4589
rect 1458 4555 1492 4573
rect 1458 4505 1492 4517
rect 1458 4483 1492 4505
rect 1458 4437 1492 4445
rect 1458 4411 1492 4437
rect 1458 4369 1492 4373
rect 1458 4339 1492 4369
rect 1458 4267 1492 4301
rect 1458 4199 1492 4229
rect 1458 4195 1492 4199
rect 1458 4131 1492 4157
rect 1458 4123 1492 4131
rect 1458 4063 1492 4085
rect 1458 4051 1492 4063
rect 1458 3995 1492 4013
rect 1458 3979 1492 3995
rect 1458 3927 1492 3941
rect 1458 3907 1492 3927
rect 1458 3859 1492 3869
rect 1458 3835 1492 3859
rect 1458 3791 1492 3797
rect 1458 3763 1492 3791
rect 1458 3723 1492 3725
rect 1458 3691 1492 3723
rect 1458 3621 1492 3653
rect 1458 3619 1492 3621
rect 1458 3553 1492 3581
rect 1458 3547 1492 3553
rect 1458 3485 1492 3509
rect 1458 3475 1492 3485
rect 1458 3417 1492 3437
rect 1458 3403 1492 3417
rect 1458 3349 1492 3365
rect 1458 3331 1492 3349
rect 1458 3281 1492 3293
rect 1458 3259 1492 3281
rect 1458 3213 1492 3221
rect 1458 3187 1492 3213
rect 1458 3145 1492 3149
rect 1458 3115 1492 3145
rect 1458 3043 1492 3077
rect 1458 2975 1492 3005
rect 1458 2971 1492 2975
rect 1458 2907 1492 2933
rect 1458 2899 1492 2907
rect 1458 2839 1492 2861
rect 1458 2827 1492 2839
rect 1458 2771 1492 2789
rect 1458 2755 1492 2771
rect 1458 2703 1492 2717
rect 1458 2683 1492 2703
rect 1458 2635 1492 2645
rect 1458 2611 1492 2635
rect 1458 2567 1492 2573
rect 1458 2539 1492 2567
rect 1458 2499 1492 2501
rect 1458 2467 1492 2499
rect 1458 2397 1492 2429
rect 1458 2395 1492 2397
rect 1458 2329 1492 2357
rect 1458 2323 1492 2329
rect 1458 2261 1492 2285
rect 1458 2251 1492 2261
rect 1458 2193 1492 2213
rect 1458 2179 1492 2193
rect 1458 2125 1492 2141
rect 1458 2107 1492 2125
rect 1458 2057 1492 2069
rect 1458 2035 1492 2057
rect 1458 1989 1492 1997
rect 1458 1963 1492 1989
rect 1458 1921 1492 1925
rect 1458 1891 1492 1921
rect 1458 1819 1492 1853
rect 1458 1751 1492 1781
rect 1458 1747 1492 1751
rect 1458 1683 1492 1709
rect 1458 1675 1492 1683
rect 1458 1615 1492 1637
rect 1458 1603 1492 1615
rect 1458 1547 1492 1565
rect 1458 1531 1492 1547
rect 1458 1479 1492 1493
rect 1458 1459 1492 1479
rect 1458 1411 1492 1421
rect 1458 1387 1492 1411
rect 1458 1343 1492 1349
rect 1458 1315 1492 1343
rect 1458 1275 1492 1277
rect 1458 1243 1492 1275
rect 1458 1173 1492 1205
rect 1458 1171 1492 1173
rect 1458 1105 1492 1133
rect 1458 1099 1492 1105
rect 1458 1037 1492 1061
rect 1458 1027 1492 1037
rect 1458 969 1492 989
rect 1458 955 1492 969
rect 1458 901 1492 917
rect 1458 883 1492 901
rect 1458 833 1492 845
rect 1458 811 1492 833
rect 1458 765 1492 773
rect 1458 739 1492 765
rect 1458 697 1492 701
rect 1458 667 1492 697
rect 1458 595 1492 629
rect 1458 527 1492 557
rect 1458 523 1492 527
rect 1458 459 1492 485
rect 1458 451 1492 459
rect 1458 391 1492 413
rect 1458 379 1492 391
rect 1458 323 1492 341
rect 1458 307 1492 323
rect 1458 255 1492 269
rect 1458 235 1492 255
rect 1458 187 1492 197
rect 1458 163 1492 187
rect 1458 119 1492 125
rect 1458 91 1492 119
rect 1458 51 1492 53
rect 1458 19 1492 51
rect 1458 -51 1492 -19
rect 1458 -53 1492 -51
rect 1458 -119 1492 -91
rect 1458 -125 1492 -119
rect 1458 -187 1492 -163
rect 1458 -197 1492 -187
rect 1458 -255 1492 -235
rect 1458 -269 1492 -255
rect 1458 -323 1492 -307
rect 1458 -341 1492 -323
rect 1458 -391 1492 -379
rect 1458 -413 1492 -391
rect 1458 -459 1492 -451
rect 1458 -485 1492 -459
rect 1458 -527 1492 -523
rect 1458 -557 1492 -527
rect 1458 -629 1492 -595
rect 1458 -697 1492 -667
rect 1458 -701 1492 -697
rect 1458 -765 1492 -739
rect 1458 -773 1492 -765
rect 1458 -833 1492 -811
rect 1458 -845 1492 -833
rect 1458 -901 1492 -883
rect 1458 -917 1492 -901
rect 1458 -969 1492 -955
rect 1458 -989 1492 -969
rect 1458 -1037 1492 -1027
rect 1458 -1061 1492 -1037
rect 1458 -1105 1492 -1099
rect 1458 -1133 1492 -1105
rect 1458 -1173 1492 -1171
rect 1458 -1205 1492 -1173
rect 1458 -1275 1492 -1243
rect 1458 -1277 1492 -1275
rect 1458 -1343 1492 -1315
rect 1458 -1349 1492 -1343
rect 1458 -1411 1492 -1387
rect 1458 -1421 1492 -1411
rect 1458 -1479 1492 -1459
rect 1458 -1493 1492 -1479
rect 1458 -1547 1492 -1531
rect 1458 -1565 1492 -1547
rect 1458 -1615 1492 -1603
rect 1458 -1637 1492 -1615
rect 1458 -1683 1492 -1675
rect 1458 -1709 1492 -1683
rect 1458 -1751 1492 -1747
rect 1458 -1781 1492 -1751
rect 1458 -1853 1492 -1819
rect 1458 -1921 1492 -1891
rect 1458 -1925 1492 -1921
rect 1458 -1989 1492 -1963
rect 1458 -1997 1492 -1989
rect 1458 -2057 1492 -2035
rect 1458 -2069 1492 -2057
rect 1458 -2125 1492 -2107
rect 1458 -2141 1492 -2125
rect 1458 -2193 1492 -2179
rect 1458 -2213 1492 -2193
rect 1458 -2261 1492 -2251
rect 1458 -2285 1492 -2261
rect 1458 -2329 1492 -2323
rect 1458 -2357 1492 -2329
rect 1458 -2397 1492 -2395
rect 1458 -2429 1492 -2397
rect 1458 -2499 1492 -2467
rect 1458 -2501 1492 -2499
rect 1458 -2567 1492 -2539
rect 1458 -2573 1492 -2567
rect 1458 -2635 1492 -2611
rect 1458 -2645 1492 -2635
rect 1458 -2703 1492 -2683
rect 1458 -2717 1492 -2703
rect 1458 -2771 1492 -2755
rect 1458 -2789 1492 -2771
rect 1458 -2839 1492 -2827
rect 1458 -2861 1492 -2839
rect 1458 -2907 1492 -2899
rect 1458 -2933 1492 -2907
rect 1458 -2975 1492 -2971
rect 1458 -3005 1492 -2975
rect 1458 -3077 1492 -3043
rect 1458 -3145 1492 -3115
rect 1458 -3149 1492 -3145
rect 1458 -3213 1492 -3187
rect 1458 -3221 1492 -3213
rect 1458 -3281 1492 -3259
rect 1458 -3293 1492 -3281
rect 1458 -3349 1492 -3331
rect 1458 -3365 1492 -3349
rect 1458 -3417 1492 -3403
rect 1458 -3437 1492 -3417
rect 1458 -3485 1492 -3475
rect 1458 -3509 1492 -3485
rect 1458 -3553 1492 -3547
rect 1458 -3581 1492 -3553
rect 1458 -3621 1492 -3619
rect 1458 -3653 1492 -3621
rect 1458 -3723 1492 -3691
rect 1458 -3725 1492 -3723
rect 1458 -3791 1492 -3763
rect 1458 -3797 1492 -3791
rect 1458 -3859 1492 -3835
rect 1458 -3869 1492 -3859
rect 1458 -3927 1492 -3907
rect 1458 -3941 1492 -3927
rect 1458 -3995 1492 -3979
rect 1458 -4013 1492 -3995
rect 1458 -4063 1492 -4051
rect 1458 -4085 1492 -4063
rect 1458 -4131 1492 -4123
rect 1458 -4157 1492 -4131
rect 1458 -4199 1492 -4195
rect 1458 -4229 1492 -4199
rect 1458 -4301 1492 -4267
rect 1458 -4369 1492 -4339
rect 1458 -4373 1492 -4369
rect 1458 -4437 1492 -4411
rect 1458 -4445 1492 -4437
rect 1458 -4505 1492 -4483
rect 1458 -4517 1492 -4505
rect 1458 -4573 1492 -4555
rect 1458 -4589 1492 -4573
rect 1458 -4641 1492 -4627
rect 1458 -4661 1492 -4641
rect 1458 -4709 1492 -4699
rect 1458 -4733 1492 -4709
rect 1458 -4777 1492 -4771
rect 1458 -4805 1492 -4777
rect 1458 -4845 1492 -4843
rect 1458 -4877 1492 -4845
rect 1458 -4947 1492 -4915
rect 1458 -4949 1492 -4947
rect 1458 -5015 1492 -4987
rect 1458 -5021 1492 -5015
rect 1458 -5083 1492 -5059
rect 1458 -5093 1492 -5083
rect 1458 -5151 1492 -5131
rect 1458 -5165 1492 -5151
rect 1458 -5219 1492 -5203
rect 1458 -5237 1492 -5219
rect 1458 -5287 1492 -5275
rect 1458 -5309 1492 -5287
rect 1458 -5355 1492 -5347
rect 1458 -5381 1492 -5355
rect 1458 -5423 1492 -5419
rect 1458 -5453 1492 -5423
rect 1458 -5525 1492 -5491
rect 1458 -5593 1492 -5563
rect 1458 -5597 1492 -5593
rect 1458 -5661 1492 -5635
rect 1458 -5669 1492 -5661
rect 1458 -5729 1492 -5707
rect 1458 -5741 1492 -5729
rect 1458 -5797 1492 -5779
rect 1458 -5813 1492 -5797
rect 1458 -5865 1492 -5851
rect 1458 -5885 1492 -5865
rect 1458 -5933 1492 -5923
rect 1458 -5957 1492 -5933
rect 1458 -6001 1492 -5995
rect 1458 -6029 1492 -6001
rect 1458 -6069 1492 -6067
rect 1458 -6101 1492 -6069
rect 1458 -6171 1492 -6139
rect 1458 -6173 1492 -6171
rect 1458 -6239 1492 -6211
rect 1458 -6245 1492 -6239
rect 1458 -6307 1492 -6283
rect 1458 -6317 1492 -6307
rect 1458 -6375 1492 -6355
rect 1458 -6389 1492 -6375
rect 1458 -6443 1492 -6427
rect 1458 -6461 1492 -6443
rect 1458 -6511 1492 -6499
rect 1458 -6533 1492 -6511
rect 1458 -6579 1492 -6571
rect 1458 -6605 1492 -6579
rect 1458 -6647 1492 -6643
rect 1458 -6677 1492 -6647
rect 1458 -6749 1492 -6715
rect 1458 -6817 1492 -6787
rect 1458 -6821 1492 -6817
rect 1458 -6885 1492 -6859
rect 1458 -6893 1492 -6885
rect 1458 -6953 1492 -6931
rect 1458 -6965 1492 -6953
rect 1458 -7021 1492 -7003
rect 1458 -7037 1492 -7021
rect 1458 -7089 1492 -7075
rect 1458 -7109 1492 -7089
rect 1458 -7157 1492 -7147
rect 1458 -7181 1492 -7157
rect 1458 -7225 1492 -7219
rect 1458 -7253 1492 -7225
rect 1458 -7293 1492 -7291
rect 1458 -7325 1492 -7293
rect 1458 -7395 1492 -7363
rect 1458 -7397 1492 -7395
rect 1458 -7463 1492 -7435
rect 1458 -7469 1492 -7463
rect 1458 -7531 1492 -7507
rect 1458 -7541 1492 -7531
rect 1458 -7599 1492 -7579
rect 1458 -7613 1492 -7599
rect 1458 -7667 1492 -7651
rect 1458 -7685 1492 -7667
rect 1458 -7735 1492 -7723
rect 1458 -7757 1492 -7735
rect 1458 -7803 1492 -7795
rect 1458 -7829 1492 -7803
rect 1458 -7871 1492 -7867
rect 1458 -7901 1492 -7871
rect 1458 -7973 1492 -7939
rect 1458 -8041 1492 -8011
rect 1458 -8045 1492 -8041
rect 1458 -8109 1492 -8083
rect 1458 -8117 1492 -8109
rect 1458 -8177 1492 -8155
rect 1458 -8189 1492 -8177
rect 1458 -8245 1492 -8227
rect 1458 -8261 1492 -8245
rect 1458 -8313 1492 -8299
rect 1458 -8333 1492 -8313
rect 1458 -8381 1492 -8371
rect 1458 -8405 1492 -8381
rect 1458 -8449 1492 -8443
rect 1458 -8477 1492 -8449
rect 1458 -8517 1492 -8515
rect 1458 -8549 1492 -8517
rect 1458 -8619 1492 -8587
rect 1458 -8621 1492 -8619
rect 1458 -8687 1492 -8659
rect 1458 -8693 1492 -8687
rect 1458 -8755 1492 -8731
rect 1458 -8765 1492 -8755
rect 1458 -8823 1492 -8803
rect 1458 -8837 1492 -8823
rect 1458 -8891 1492 -8875
rect 1458 -8909 1492 -8891
rect 1458 -8959 1492 -8947
rect 1458 -8981 1492 -8959
rect 1458 -9027 1492 -9019
rect 1458 -9053 1492 -9027
rect 1458 -9095 1492 -9091
rect 1458 -9125 1492 -9095
rect 1458 -9197 1492 -9163
rect 1458 -9265 1492 -9235
rect 1458 -9269 1492 -9265
rect 1458 -9333 1492 -9307
rect 1458 -9341 1492 -9333
rect 1458 -9401 1492 -9379
rect 1458 -9413 1492 -9401
rect 1458 -9469 1492 -9451
rect 1458 -9485 1492 -9469
rect 1458 -9537 1492 -9523
rect 1458 -9557 1492 -9537
<< metal1 >>
rect -1498 9557 -1452 9600
rect -1498 9523 -1492 9557
rect -1458 9523 -1452 9557
rect -1498 9485 -1452 9523
rect -1498 9451 -1492 9485
rect -1458 9451 -1452 9485
rect -1498 9413 -1452 9451
rect -1498 9379 -1492 9413
rect -1458 9379 -1452 9413
rect -1498 9341 -1452 9379
rect -1498 9307 -1492 9341
rect -1458 9307 -1452 9341
rect -1498 9269 -1452 9307
rect -1498 9235 -1492 9269
rect -1458 9235 -1452 9269
rect -1498 9197 -1452 9235
rect -1498 9163 -1492 9197
rect -1458 9163 -1452 9197
rect -1498 9125 -1452 9163
rect -1498 9091 -1492 9125
rect -1458 9091 -1452 9125
rect -1498 9053 -1452 9091
rect -1498 9019 -1492 9053
rect -1458 9019 -1452 9053
rect -1498 8981 -1452 9019
rect -1498 8947 -1492 8981
rect -1458 8947 -1452 8981
rect -1498 8909 -1452 8947
rect -1498 8875 -1492 8909
rect -1458 8875 -1452 8909
rect -1498 8837 -1452 8875
rect -1498 8803 -1492 8837
rect -1458 8803 -1452 8837
rect -1498 8765 -1452 8803
rect -1498 8731 -1492 8765
rect -1458 8731 -1452 8765
rect -1498 8693 -1452 8731
rect -1498 8659 -1492 8693
rect -1458 8659 -1452 8693
rect -1498 8621 -1452 8659
rect -1498 8587 -1492 8621
rect -1458 8587 -1452 8621
rect -1498 8549 -1452 8587
rect -1498 8515 -1492 8549
rect -1458 8515 -1452 8549
rect -1498 8477 -1452 8515
rect -1498 8443 -1492 8477
rect -1458 8443 -1452 8477
rect -1498 8405 -1452 8443
rect -1498 8371 -1492 8405
rect -1458 8371 -1452 8405
rect -1498 8333 -1452 8371
rect -1498 8299 -1492 8333
rect -1458 8299 -1452 8333
rect -1498 8261 -1452 8299
rect -1498 8227 -1492 8261
rect -1458 8227 -1452 8261
rect -1498 8189 -1452 8227
rect -1498 8155 -1492 8189
rect -1458 8155 -1452 8189
rect -1498 8117 -1452 8155
rect -1498 8083 -1492 8117
rect -1458 8083 -1452 8117
rect -1498 8045 -1452 8083
rect -1498 8011 -1492 8045
rect -1458 8011 -1452 8045
rect -1498 7973 -1452 8011
rect -1498 7939 -1492 7973
rect -1458 7939 -1452 7973
rect -1498 7901 -1452 7939
rect -1498 7867 -1492 7901
rect -1458 7867 -1452 7901
rect -1498 7829 -1452 7867
rect -1498 7795 -1492 7829
rect -1458 7795 -1452 7829
rect -1498 7757 -1452 7795
rect -1498 7723 -1492 7757
rect -1458 7723 -1452 7757
rect -1498 7685 -1452 7723
rect -1498 7651 -1492 7685
rect -1458 7651 -1452 7685
rect -1498 7613 -1452 7651
rect -1498 7579 -1492 7613
rect -1458 7579 -1452 7613
rect -1498 7541 -1452 7579
rect -1498 7507 -1492 7541
rect -1458 7507 -1452 7541
rect -1498 7469 -1452 7507
rect -1498 7435 -1492 7469
rect -1458 7435 -1452 7469
rect -1498 7397 -1452 7435
rect -1498 7363 -1492 7397
rect -1458 7363 -1452 7397
rect -1498 7325 -1452 7363
rect -1498 7291 -1492 7325
rect -1458 7291 -1452 7325
rect -1498 7253 -1452 7291
rect -1498 7219 -1492 7253
rect -1458 7219 -1452 7253
rect -1498 7181 -1452 7219
rect -1498 7147 -1492 7181
rect -1458 7147 -1452 7181
rect -1498 7109 -1452 7147
rect -1498 7075 -1492 7109
rect -1458 7075 -1452 7109
rect -1498 7037 -1452 7075
rect -1498 7003 -1492 7037
rect -1458 7003 -1452 7037
rect -1498 6965 -1452 7003
rect -1498 6931 -1492 6965
rect -1458 6931 -1452 6965
rect -1498 6893 -1452 6931
rect -1498 6859 -1492 6893
rect -1458 6859 -1452 6893
rect -1498 6821 -1452 6859
rect -1498 6787 -1492 6821
rect -1458 6787 -1452 6821
rect -1498 6749 -1452 6787
rect -1498 6715 -1492 6749
rect -1458 6715 -1452 6749
rect -1498 6677 -1452 6715
rect -1498 6643 -1492 6677
rect -1458 6643 -1452 6677
rect -1498 6605 -1452 6643
rect -1498 6571 -1492 6605
rect -1458 6571 -1452 6605
rect -1498 6533 -1452 6571
rect -1498 6499 -1492 6533
rect -1458 6499 -1452 6533
rect -1498 6461 -1452 6499
rect -1498 6427 -1492 6461
rect -1458 6427 -1452 6461
rect -1498 6389 -1452 6427
rect -1498 6355 -1492 6389
rect -1458 6355 -1452 6389
rect -1498 6317 -1452 6355
rect -1498 6283 -1492 6317
rect -1458 6283 -1452 6317
rect -1498 6245 -1452 6283
rect -1498 6211 -1492 6245
rect -1458 6211 -1452 6245
rect -1498 6173 -1452 6211
rect -1498 6139 -1492 6173
rect -1458 6139 -1452 6173
rect -1498 6101 -1452 6139
rect -1498 6067 -1492 6101
rect -1458 6067 -1452 6101
rect -1498 6029 -1452 6067
rect -1498 5995 -1492 6029
rect -1458 5995 -1452 6029
rect -1498 5957 -1452 5995
rect -1498 5923 -1492 5957
rect -1458 5923 -1452 5957
rect -1498 5885 -1452 5923
rect -1498 5851 -1492 5885
rect -1458 5851 -1452 5885
rect -1498 5813 -1452 5851
rect -1498 5779 -1492 5813
rect -1458 5779 -1452 5813
rect -1498 5741 -1452 5779
rect -1498 5707 -1492 5741
rect -1458 5707 -1452 5741
rect -1498 5669 -1452 5707
rect -1498 5635 -1492 5669
rect -1458 5635 -1452 5669
rect -1498 5597 -1452 5635
rect -1498 5563 -1492 5597
rect -1458 5563 -1452 5597
rect -1498 5525 -1452 5563
rect -1498 5491 -1492 5525
rect -1458 5491 -1452 5525
rect -1498 5453 -1452 5491
rect -1498 5419 -1492 5453
rect -1458 5419 -1452 5453
rect -1498 5381 -1452 5419
rect -1498 5347 -1492 5381
rect -1458 5347 -1452 5381
rect -1498 5309 -1452 5347
rect -1498 5275 -1492 5309
rect -1458 5275 -1452 5309
rect -1498 5237 -1452 5275
rect -1498 5203 -1492 5237
rect -1458 5203 -1452 5237
rect -1498 5165 -1452 5203
rect -1498 5131 -1492 5165
rect -1458 5131 -1452 5165
rect -1498 5093 -1452 5131
rect -1498 5059 -1492 5093
rect -1458 5059 -1452 5093
rect -1498 5021 -1452 5059
rect -1498 4987 -1492 5021
rect -1458 4987 -1452 5021
rect -1498 4949 -1452 4987
rect -1498 4915 -1492 4949
rect -1458 4915 -1452 4949
rect -1498 4877 -1452 4915
rect -1498 4843 -1492 4877
rect -1458 4843 -1452 4877
rect -1498 4805 -1452 4843
rect -1498 4771 -1492 4805
rect -1458 4771 -1452 4805
rect -1498 4733 -1452 4771
rect -1498 4699 -1492 4733
rect -1458 4699 -1452 4733
rect -1498 4661 -1452 4699
rect -1498 4627 -1492 4661
rect -1458 4627 -1452 4661
rect -1498 4589 -1452 4627
rect -1498 4555 -1492 4589
rect -1458 4555 -1452 4589
rect -1498 4517 -1452 4555
rect -1498 4483 -1492 4517
rect -1458 4483 -1452 4517
rect -1498 4445 -1452 4483
rect -1498 4411 -1492 4445
rect -1458 4411 -1452 4445
rect -1498 4373 -1452 4411
rect -1498 4339 -1492 4373
rect -1458 4339 -1452 4373
rect -1498 4301 -1452 4339
rect -1498 4267 -1492 4301
rect -1458 4267 -1452 4301
rect -1498 4229 -1452 4267
rect -1498 4195 -1492 4229
rect -1458 4195 -1452 4229
rect -1498 4157 -1452 4195
rect -1498 4123 -1492 4157
rect -1458 4123 -1452 4157
rect -1498 4085 -1452 4123
rect -1498 4051 -1492 4085
rect -1458 4051 -1452 4085
rect -1498 4013 -1452 4051
rect -1498 3979 -1492 4013
rect -1458 3979 -1452 4013
rect -1498 3941 -1452 3979
rect -1498 3907 -1492 3941
rect -1458 3907 -1452 3941
rect -1498 3869 -1452 3907
rect -1498 3835 -1492 3869
rect -1458 3835 -1452 3869
rect -1498 3797 -1452 3835
rect -1498 3763 -1492 3797
rect -1458 3763 -1452 3797
rect -1498 3725 -1452 3763
rect -1498 3691 -1492 3725
rect -1458 3691 -1452 3725
rect -1498 3653 -1452 3691
rect -1498 3619 -1492 3653
rect -1458 3619 -1452 3653
rect -1498 3581 -1452 3619
rect -1498 3547 -1492 3581
rect -1458 3547 -1452 3581
rect -1498 3509 -1452 3547
rect -1498 3475 -1492 3509
rect -1458 3475 -1452 3509
rect -1498 3437 -1452 3475
rect -1498 3403 -1492 3437
rect -1458 3403 -1452 3437
rect -1498 3365 -1452 3403
rect -1498 3331 -1492 3365
rect -1458 3331 -1452 3365
rect -1498 3293 -1452 3331
rect -1498 3259 -1492 3293
rect -1458 3259 -1452 3293
rect -1498 3221 -1452 3259
rect -1498 3187 -1492 3221
rect -1458 3187 -1452 3221
rect -1498 3149 -1452 3187
rect -1498 3115 -1492 3149
rect -1458 3115 -1452 3149
rect -1498 3077 -1452 3115
rect -1498 3043 -1492 3077
rect -1458 3043 -1452 3077
rect -1498 3005 -1452 3043
rect -1498 2971 -1492 3005
rect -1458 2971 -1452 3005
rect -1498 2933 -1452 2971
rect -1498 2899 -1492 2933
rect -1458 2899 -1452 2933
rect -1498 2861 -1452 2899
rect -1498 2827 -1492 2861
rect -1458 2827 -1452 2861
rect -1498 2789 -1452 2827
rect -1498 2755 -1492 2789
rect -1458 2755 -1452 2789
rect -1498 2717 -1452 2755
rect -1498 2683 -1492 2717
rect -1458 2683 -1452 2717
rect -1498 2645 -1452 2683
rect -1498 2611 -1492 2645
rect -1458 2611 -1452 2645
rect -1498 2573 -1452 2611
rect -1498 2539 -1492 2573
rect -1458 2539 -1452 2573
rect -1498 2501 -1452 2539
rect -1498 2467 -1492 2501
rect -1458 2467 -1452 2501
rect -1498 2429 -1452 2467
rect -1498 2395 -1492 2429
rect -1458 2395 -1452 2429
rect -1498 2357 -1452 2395
rect -1498 2323 -1492 2357
rect -1458 2323 -1452 2357
rect -1498 2285 -1452 2323
rect -1498 2251 -1492 2285
rect -1458 2251 -1452 2285
rect -1498 2213 -1452 2251
rect -1498 2179 -1492 2213
rect -1458 2179 -1452 2213
rect -1498 2141 -1452 2179
rect -1498 2107 -1492 2141
rect -1458 2107 -1452 2141
rect -1498 2069 -1452 2107
rect -1498 2035 -1492 2069
rect -1458 2035 -1452 2069
rect -1498 1997 -1452 2035
rect -1498 1963 -1492 1997
rect -1458 1963 -1452 1997
rect -1498 1925 -1452 1963
rect -1498 1891 -1492 1925
rect -1458 1891 -1452 1925
rect -1498 1853 -1452 1891
rect -1498 1819 -1492 1853
rect -1458 1819 -1452 1853
rect -1498 1781 -1452 1819
rect -1498 1747 -1492 1781
rect -1458 1747 -1452 1781
rect -1498 1709 -1452 1747
rect -1498 1675 -1492 1709
rect -1458 1675 -1452 1709
rect -1498 1637 -1452 1675
rect -1498 1603 -1492 1637
rect -1458 1603 -1452 1637
rect -1498 1565 -1452 1603
rect -1498 1531 -1492 1565
rect -1458 1531 -1452 1565
rect -1498 1493 -1452 1531
rect -1498 1459 -1492 1493
rect -1458 1459 -1452 1493
rect -1498 1421 -1452 1459
rect -1498 1387 -1492 1421
rect -1458 1387 -1452 1421
rect -1498 1349 -1452 1387
rect -1498 1315 -1492 1349
rect -1458 1315 -1452 1349
rect -1498 1277 -1452 1315
rect -1498 1243 -1492 1277
rect -1458 1243 -1452 1277
rect -1498 1205 -1452 1243
rect -1498 1171 -1492 1205
rect -1458 1171 -1452 1205
rect -1498 1133 -1452 1171
rect -1498 1099 -1492 1133
rect -1458 1099 -1452 1133
rect -1498 1061 -1452 1099
rect -1498 1027 -1492 1061
rect -1458 1027 -1452 1061
rect -1498 989 -1452 1027
rect -1498 955 -1492 989
rect -1458 955 -1452 989
rect -1498 917 -1452 955
rect -1498 883 -1492 917
rect -1458 883 -1452 917
rect -1498 845 -1452 883
rect -1498 811 -1492 845
rect -1458 811 -1452 845
rect -1498 773 -1452 811
rect -1498 739 -1492 773
rect -1458 739 -1452 773
rect -1498 701 -1452 739
rect -1498 667 -1492 701
rect -1458 667 -1452 701
rect -1498 629 -1452 667
rect -1498 595 -1492 629
rect -1458 595 -1452 629
rect -1498 557 -1452 595
rect -1498 523 -1492 557
rect -1458 523 -1452 557
rect -1498 485 -1452 523
rect -1498 451 -1492 485
rect -1458 451 -1452 485
rect -1498 413 -1452 451
rect -1498 379 -1492 413
rect -1458 379 -1452 413
rect -1498 341 -1452 379
rect -1498 307 -1492 341
rect -1458 307 -1452 341
rect -1498 269 -1452 307
rect -1498 235 -1492 269
rect -1458 235 -1452 269
rect -1498 197 -1452 235
rect -1498 163 -1492 197
rect -1458 163 -1452 197
rect -1498 125 -1452 163
rect -1498 91 -1492 125
rect -1458 91 -1452 125
rect -1498 53 -1452 91
rect -1498 19 -1492 53
rect -1458 19 -1452 53
rect -1498 -19 -1452 19
rect -1498 -53 -1492 -19
rect -1458 -53 -1452 -19
rect -1498 -91 -1452 -53
rect -1498 -125 -1492 -91
rect -1458 -125 -1452 -91
rect -1498 -163 -1452 -125
rect -1498 -197 -1492 -163
rect -1458 -197 -1452 -163
rect -1498 -235 -1452 -197
rect -1498 -269 -1492 -235
rect -1458 -269 -1452 -235
rect -1498 -307 -1452 -269
rect -1498 -341 -1492 -307
rect -1458 -341 -1452 -307
rect -1498 -379 -1452 -341
rect -1498 -413 -1492 -379
rect -1458 -413 -1452 -379
rect -1498 -451 -1452 -413
rect -1498 -485 -1492 -451
rect -1458 -485 -1452 -451
rect -1498 -523 -1452 -485
rect -1498 -557 -1492 -523
rect -1458 -557 -1452 -523
rect -1498 -595 -1452 -557
rect -1498 -629 -1492 -595
rect -1458 -629 -1452 -595
rect -1498 -667 -1452 -629
rect -1498 -701 -1492 -667
rect -1458 -701 -1452 -667
rect -1498 -739 -1452 -701
rect -1498 -773 -1492 -739
rect -1458 -773 -1452 -739
rect -1498 -811 -1452 -773
rect -1498 -845 -1492 -811
rect -1458 -845 -1452 -811
rect -1498 -883 -1452 -845
rect -1498 -917 -1492 -883
rect -1458 -917 -1452 -883
rect -1498 -955 -1452 -917
rect -1498 -989 -1492 -955
rect -1458 -989 -1452 -955
rect -1498 -1027 -1452 -989
rect -1498 -1061 -1492 -1027
rect -1458 -1061 -1452 -1027
rect -1498 -1099 -1452 -1061
rect -1498 -1133 -1492 -1099
rect -1458 -1133 -1452 -1099
rect -1498 -1171 -1452 -1133
rect -1498 -1205 -1492 -1171
rect -1458 -1205 -1452 -1171
rect -1498 -1243 -1452 -1205
rect -1498 -1277 -1492 -1243
rect -1458 -1277 -1452 -1243
rect -1498 -1315 -1452 -1277
rect -1498 -1349 -1492 -1315
rect -1458 -1349 -1452 -1315
rect -1498 -1387 -1452 -1349
rect -1498 -1421 -1492 -1387
rect -1458 -1421 -1452 -1387
rect -1498 -1459 -1452 -1421
rect -1498 -1493 -1492 -1459
rect -1458 -1493 -1452 -1459
rect -1498 -1531 -1452 -1493
rect -1498 -1565 -1492 -1531
rect -1458 -1565 -1452 -1531
rect -1498 -1603 -1452 -1565
rect -1498 -1637 -1492 -1603
rect -1458 -1637 -1452 -1603
rect -1498 -1675 -1452 -1637
rect -1498 -1709 -1492 -1675
rect -1458 -1709 -1452 -1675
rect -1498 -1747 -1452 -1709
rect -1498 -1781 -1492 -1747
rect -1458 -1781 -1452 -1747
rect -1498 -1819 -1452 -1781
rect -1498 -1853 -1492 -1819
rect -1458 -1853 -1452 -1819
rect -1498 -1891 -1452 -1853
rect -1498 -1925 -1492 -1891
rect -1458 -1925 -1452 -1891
rect -1498 -1963 -1452 -1925
rect -1498 -1997 -1492 -1963
rect -1458 -1997 -1452 -1963
rect -1498 -2035 -1452 -1997
rect -1498 -2069 -1492 -2035
rect -1458 -2069 -1452 -2035
rect -1498 -2107 -1452 -2069
rect -1498 -2141 -1492 -2107
rect -1458 -2141 -1452 -2107
rect -1498 -2179 -1452 -2141
rect -1498 -2213 -1492 -2179
rect -1458 -2213 -1452 -2179
rect -1498 -2251 -1452 -2213
rect -1498 -2285 -1492 -2251
rect -1458 -2285 -1452 -2251
rect -1498 -2323 -1452 -2285
rect -1498 -2357 -1492 -2323
rect -1458 -2357 -1452 -2323
rect -1498 -2395 -1452 -2357
rect -1498 -2429 -1492 -2395
rect -1458 -2429 -1452 -2395
rect -1498 -2467 -1452 -2429
rect -1498 -2501 -1492 -2467
rect -1458 -2501 -1452 -2467
rect -1498 -2539 -1452 -2501
rect -1498 -2573 -1492 -2539
rect -1458 -2573 -1452 -2539
rect -1498 -2611 -1452 -2573
rect -1498 -2645 -1492 -2611
rect -1458 -2645 -1452 -2611
rect -1498 -2683 -1452 -2645
rect -1498 -2717 -1492 -2683
rect -1458 -2717 -1452 -2683
rect -1498 -2755 -1452 -2717
rect -1498 -2789 -1492 -2755
rect -1458 -2789 -1452 -2755
rect -1498 -2827 -1452 -2789
rect -1498 -2861 -1492 -2827
rect -1458 -2861 -1452 -2827
rect -1498 -2899 -1452 -2861
rect -1498 -2933 -1492 -2899
rect -1458 -2933 -1452 -2899
rect -1498 -2971 -1452 -2933
rect -1498 -3005 -1492 -2971
rect -1458 -3005 -1452 -2971
rect -1498 -3043 -1452 -3005
rect -1498 -3077 -1492 -3043
rect -1458 -3077 -1452 -3043
rect -1498 -3115 -1452 -3077
rect -1498 -3149 -1492 -3115
rect -1458 -3149 -1452 -3115
rect -1498 -3187 -1452 -3149
rect -1498 -3221 -1492 -3187
rect -1458 -3221 -1452 -3187
rect -1498 -3259 -1452 -3221
rect -1498 -3293 -1492 -3259
rect -1458 -3293 -1452 -3259
rect -1498 -3331 -1452 -3293
rect -1498 -3365 -1492 -3331
rect -1458 -3365 -1452 -3331
rect -1498 -3403 -1452 -3365
rect -1498 -3437 -1492 -3403
rect -1458 -3437 -1452 -3403
rect -1498 -3475 -1452 -3437
rect -1498 -3509 -1492 -3475
rect -1458 -3509 -1452 -3475
rect -1498 -3547 -1452 -3509
rect -1498 -3581 -1492 -3547
rect -1458 -3581 -1452 -3547
rect -1498 -3619 -1452 -3581
rect -1498 -3653 -1492 -3619
rect -1458 -3653 -1452 -3619
rect -1498 -3691 -1452 -3653
rect -1498 -3725 -1492 -3691
rect -1458 -3725 -1452 -3691
rect -1498 -3763 -1452 -3725
rect -1498 -3797 -1492 -3763
rect -1458 -3797 -1452 -3763
rect -1498 -3835 -1452 -3797
rect -1498 -3869 -1492 -3835
rect -1458 -3869 -1452 -3835
rect -1498 -3907 -1452 -3869
rect -1498 -3941 -1492 -3907
rect -1458 -3941 -1452 -3907
rect -1498 -3979 -1452 -3941
rect -1498 -4013 -1492 -3979
rect -1458 -4013 -1452 -3979
rect -1498 -4051 -1452 -4013
rect -1498 -4085 -1492 -4051
rect -1458 -4085 -1452 -4051
rect -1498 -4123 -1452 -4085
rect -1498 -4157 -1492 -4123
rect -1458 -4157 -1452 -4123
rect -1498 -4195 -1452 -4157
rect -1498 -4229 -1492 -4195
rect -1458 -4229 -1452 -4195
rect -1498 -4267 -1452 -4229
rect -1498 -4301 -1492 -4267
rect -1458 -4301 -1452 -4267
rect -1498 -4339 -1452 -4301
rect -1498 -4373 -1492 -4339
rect -1458 -4373 -1452 -4339
rect -1498 -4411 -1452 -4373
rect -1498 -4445 -1492 -4411
rect -1458 -4445 -1452 -4411
rect -1498 -4483 -1452 -4445
rect -1498 -4517 -1492 -4483
rect -1458 -4517 -1452 -4483
rect -1498 -4555 -1452 -4517
rect -1498 -4589 -1492 -4555
rect -1458 -4589 -1452 -4555
rect -1498 -4627 -1452 -4589
rect -1498 -4661 -1492 -4627
rect -1458 -4661 -1452 -4627
rect -1498 -4699 -1452 -4661
rect -1498 -4733 -1492 -4699
rect -1458 -4733 -1452 -4699
rect -1498 -4771 -1452 -4733
rect -1498 -4805 -1492 -4771
rect -1458 -4805 -1452 -4771
rect -1498 -4843 -1452 -4805
rect -1498 -4877 -1492 -4843
rect -1458 -4877 -1452 -4843
rect -1498 -4915 -1452 -4877
rect -1498 -4949 -1492 -4915
rect -1458 -4949 -1452 -4915
rect -1498 -4987 -1452 -4949
rect -1498 -5021 -1492 -4987
rect -1458 -5021 -1452 -4987
rect -1498 -5059 -1452 -5021
rect -1498 -5093 -1492 -5059
rect -1458 -5093 -1452 -5059
rect -1498 -5131 -1452 -5093
rect -1498 -5165 -1492 -5131
rect -1458 -5165 -1452 -5131
rect -1498 -5203 -1452 -5165
rect -1498 -5237 -1492 -5203
rect -1458 -5237 -1452 -5203
rect -1498 -5275 -1452 -5237
rect -1498 -5309 -1492 -5275
rect -1458 -5309 -1452 -5275
rect -1498 -5347 -1452 -5309
rect -1498 -5381 -1492 -5347
rect -1458 -5381 -1452 -5347
rect -1498 -5419 -1452 -5381
rect -1498 -5453 -1492 -5419
rect -1458 -5453 -1452 -5419
rect -1498 -5491 -1452 -5453
rect -1498 -5525 -1492 -5491
rect -1458 -5525 -1452 -5491
rect -1498 -5563 -1452 -5525
rect -1498 -5597 -1492 -5563
rect -1458 -5597 -1452 -5563
rect -1498 -5635 -1452 -5597
rect -1498 -5669 -1492 -5635
rect -1458 -5669 -1452 -5635
rect -1498 -5707 -1452 -5669
rect -1498 -5741 -1492 -5707
rect -1458 -5741 -1452 -5707
rect -1498 -5779 -1452 -5741
rect -1498 -5813 -1492 -5779
rect -1458 -5813 -1452 -5779
rect -1498 -5851 -1452 -5813
rect -1498 -5885 -1492 -5851
rect -1458 -5885 -1452 -5851
rect -1498 -5923 -1452 -5885
rect -1498 -5957 -1492 -5923
rect -1458 -5957 -1452 -5923
rect -1498 -5995 -1452 -5957
rect -1498 -6029 -1492 -5995
rect -1458 -6029 -1452 -5995
rect -1498 -6067 -1452 -6029
rect -1498 -6101 -1492 -6067
rect -1458 -6101 -1452 -6067
rect -1498 -6139 -1452 -6101
rect -1498 -6173 -1492 -6139
rect -1458 -6173 -1452 -6139
rect -1498 -6211 -1452 -6173
rect -1498 -6245 -1492 -6211
rect -1458 -6245 -1452 -6211
rect -1498 -6283 -1452 -6245
rect -1498 -6317 -1492 -6283
rect -1458 -6317 -1452 -6283
rect -1498 -6355 -1452 -6317
rect -1498 -6389 -1492 -6355
rect -1458 -6389 -1452 -6355
rect -1498 -6427 -1452 -6389
rect -1498 -6461 -1492 -6427
rect -1458 -6461 -1452 -6427
rect -1498 -6499 -1452 -6461
rect -1498 -6533 -1492 -6499
rect -1458 -6533 -1452 -6499
rect -1498 -6571 -1452 -6533
rect -1498 -6605 -1492 -6571
rect -1458 -6605 -1452 -6571
rect -1498 -6643 -1452 -6605
rect -1498 -6677 -1492 -6643
rect -1458 -6677 -1452 -6643
rect -1498 -6715 -1452 -6677
rect -1498 -6749 -1492 -6715
rect -1458 -6749 -1452 -6715
rect -1498 -6787 -1452 -6749
rect -1498 -6821 -1492 -6787
rect -1458 -6821 -1452 -6787
rect -1498 -6859 -1452 -6821
rect -1498 -6893 -1492 -6859
rect -1458 -6893 -1452 -6859
rect -1498 -6931 -1452 -6893
rect -1498 -6965 -1492 -6931
rect -1458 -6965 -1452 -6931
rect -1498 -7003 -1452 -6965
rect -1498 -7037 -1492 -7003
rect -1458 -7037 -1452 -7003
rect -1498 -7075 -1452 -7037
rect -1498 -7109 -1492 -7075
rect -1458 -7109 -1452 -7075
rect -1498 -7147 -1452 -7109
rect -1498 -7181 -1492 -7147
rect -1458 -7181 -1452 -7147
rect -1498 -7219 -1452 -7181
rect -1498 -7253 -1492 -7219
rect -1458 -7253 -1452 -7219
rect -1498 -7291 -1452 -7253
rect -1498 -7325 -1492 -7291
rect -1458 -7325 -1452 -7291
rect -1498 -7363 -1452 -7325
rect -1498 -7397 -1492 -7363
rect -1458 -7397 -1452 -7363
rect -1498 -7435 -1452 -7397
rect -1498 -7469 -1492 -7435
rect -1458 -7469 -1452 -7435
rect -1498 -7507 -1452 -7469
rect -1498 -7541 -1492 -7507
rect -1458 -7541 -1452 -7507
rect -1498 -7579 -1452 -7541
rect -1498 -7613 -1492 -7579
rect -1458 -7613 -1452 -7579
rect -1498 -7651 -1452 -7613
rect -1498 -7685 -1492 -7651
rect -1458 -7685 -1452 -7651
rect -1498 -7723 -1452 -7685
rect -1498 -7757 -1492 -7723
rect -1458 -7757 -1452 -7723
rect -1498 -7795 -1452 -7757
rect -1498 -7829 -1492 -7795
rect -1458 -7829 -1452 -7795
rect -1498 -7867 -1452 -7829
rect -1498 -7901 -1492 -7867
rect -1458 -7901 -1452 -7867
rect -1498 -7939 -1452 -7901
rect -1498 -7973 -1492 -7939
rect -1458 -7973 -1452 -7939
rect -1498 -8011 -1452 -7973
rect -1498 -8045 -1492 -8011
rect -1458 -8045 -1452 -8011
rect -1498 -8083 -1452 -8045
rect -1498 -8117 -1492 -8083
rect -1458 -8117 -1452 -8083
rect -1498 -8155 -1452 -8117
rect -1498 -8189 -1492 -8155
rect -1458 -8189 -1452 -8155
rect -1498 -8227 -1452 -8189
rect -1498 -8261 -1492 -8227
rect -1458 -8261 -1452 -8227
rect -1498 -8299 -1452 -8261
rect -1498 -8333 -1492 -8299
rect -1458 -8333 -1452 -8299
rect -1498 -8371 -1452 -8333
rect -1498 -8405 -1492 -8371
rect -1458 -8405 -1452 -8371
rect -1498 -8443 -1452 -8405
rect -1498 -8477 -1492 -8443
rect -1458 -8477 -1452 -8443
rect -1498 -8515 -1452 -8477
rect -1498 -8549 -1492 -8515
rect -1458 -8549 -1452 -8515
rect -1498 -8587 -1452 -8549
rect -1498 -8621 -1492 -8587
rect -1458 -8621 -1452 -8587
rect -1498 -8659 -1452 -8621
rect -1498 -8693 -1492 -8659
rect -1458 -8693 -1452 -8659
rect -1498 -8731 -1452 -8693
rect -1498 -8765 -1492 -8731
rect -1458 -8765 -1452 -8731
rect -1498 -8803 -1452 -8765
rect -1498 -8837 -1492 -8803
rect -1458 -8837 -1452 -8803
rect -1498 -8875 -1452 -8837
rect -1498 -8909 -1492 -8875
rect -1458 -8909 -1452 -8875
rect -1498 -8947 -1452 -8909
rect -1498 -8981 -1492 -8947
rect -1458 -8981 -1452 -8947
rect -1498 -9019 -1452 -8981
rect -1498 -9053 -1492 -9019
rect -1458 -9053 -1452 -9019
rect -1498 -9091 -1452 -9053
rect -1498 -9125 -1492 -9091
rect -1458 -9125 -1452 -9091
rect -1498 -9163 -1452 -9125
rect -1498 -9197 -1492 -9163
rect -1458 -9197 -1452 -9163
rect -1498 -9235 -1452 -9197
rect -1498 -9269 -1492 -9235
rect -1458 -9269 -1452 -9235
rect -1498 -9307 -1452 -9269
rect -1498 -9341 -1492 -9307
rect -1458 -9341 -1452 -9307
rect -1498 -9379 -1452 -9341
rect -1498 -9413 -1492 -9379
rect -1458 -9413 -1452 -9379
rect -1498 -9451 -1452 -9413
rect -1498 -9485 -1492 -9451
rect -1458 -9485 -1452 -9451
rect -1498 -9523 -1452 -9485
rect -1498 -9557 -1492 -9523
rect -1458 -9557 -1452 -9523
rect -1498 -9600 -1452 -9557
rect -1380 9557 -1334 9600
rect -1380 9523 -1374 9557
rect -1340 9523 -1334 9557
rect -1380 9485 -1334 9523
rect -1380 9451 -1374 9485
rect -1340 9451 -1334 9485
rect -1380 9413 -1334 9451
rect -1380 9379 -1374 9413
rect -1340 9379 -1334 9413
rect -1380 9341 -1334 9379
rect -1380 9307 -1374 9341
rect -1340 9307 -1334 9341
rect -1380 9269 -1334 9307
rect -1380 9235 -1374 9269
rect -1340 9235 -1334 9269
rect -1380 9197 -1334 9235
rect -1380 9163 -1374 9197
rect -1340 9163 -1334 9197
rect -1380 9125 -1334 9163
rect -1380 9091 -1374 9125
rect -1340 9091 -1334 9125
rect -1380 9053 -1334 9091
rect -1380 9019 -1374 9053
rect -1340 9019 -1334 9053
rect -1380 8981 -1334 9019
rect -1380 8947 -1374 8981
rect -1340 8947 -1334 8981
rect -1380 8909 -1334 8947
rect -1380 8875 -1374 8909
rect -1340 8875 -1334 8909
rect -1380 8837 -1334 8875
rect -1380 8803 -1374 8837
rect -1340 8803 -1334 8837
rect -1380 8765 -1334 8803
rect -1380 8731 -1374 8765
rect -1340 8731 -1334 8765
rect -1380 8693 -1334 8731
rect -1380 8659 -1374 8693
rect -1340 8659 -1334 8693
rect -1380 8621 -1334 8659
rect -1380 8587 -1374 8621
rect -1340 8587 -1334 8621
rect -1380 8549 -1334 8587
rect -1380 8515 -1374 8549
rect -1340 8515 -1334 8549
rect -1380 8477 -1334 8515
rect -1380 8443 -1374 8477
rect -1340 8443 -1334 8477
rect -1380 8405 -1334 8443
rect -1380 8371 -1374 8405
rect -1340 8371 -1334 8405
rect -1380 8333 -1334 8371
rect -1380 8299 -1374 8333
rect -1340 8299 -1334 8333
rect -1380 8261 -1334 8299
rect -1380 8227 -1374 8261
rect -1340 8227 -1334 8261
rect -1380 8189 -1334 8227
rect -1380 8155 -1374 8189
rect -1340 8155 -1334 8189
rect -1380 8117 -1334 8155
rect -1380 8083 -1374 8117
rect -1340 8083 -1334 8117
rect -1380 8045 -1334 8083
rect -1380 8011 -1374 8045
rect -1340 8011 -1334 8045
rect -1380 7973 -1334 8011
rect -1380 7939 -1374 7973
rect -1340 7939 -1334 7973
rect -1380 7901 -1334 7939
rect -1380 7867 -1374 7901
rect -1340 7867 -1334 7901
rect -1380 7829 -1334 7867
rect -1380 7795 -1374 7829
rect -1340 7795 -1334 7829
rect -1380 7757 -1334 7795
rect -1380 7723 -1374 7757
rect -1340 7723 -1334 7757
rect -1380 7685 -1334 7723
rect -1380 7651 -1374 7685
rect -1340 7651 -1334 7685
rect -1380 7613 -1334 7651
rect -1380 7579 -1374 7613
rect -1340 7579 -1334 7613
rect -1380 7541 -1334 7579
rect -1380 7507 -1374 7541
rect -1340 7507 -1334 7541
rect -1380 7469 -1334 7507
rect -1380 7435 -1374 7469
rect -1340 7435 -1334 7469
rect -1380 7397 -1334 7435
rect -1380 7363 -1374 7397
rect -1340 7363 -1334 7397
rect -1380 7325 -1334 7363
rect -1380 7291 -1374 7325
rect -1340 7291 -1334 7325
rect -1380 7253 -1334 7291
rect -1380 7219 -1374 7253
rect -1340 7219 -1334 7253
rect -1380 7181 -1334 7219
rect -1380 7147 -1374 7181
rect -1340 7147 -1334 7181
rect -1380 7109 -1334 7147
rect -1380 7075 -1374 7109
rect -1340 7075 -1334 7109
rect -1380 7037 -1334 7075
rect -1380 7003 -1374 7037
rect -1340 7003 -1334 7037
rect -1380 6965 -1334 7003
rect -1380 6931 -1374 6965
rect -1340 6931 -1334 6965
rect -1380 6893 -1334 6931
rect -1380 6859 -1374 6893
rect -1340 6859 -1334 6893
rect -1380 6821 -1334 6859
rect -1380 6787 -1374 6821
rect -1340 6787 -1334 6821
rect -1380 6749 -1334 6787
rect -1380 6715 -1374 6749
rect -1340 6715 -1334 6749
rect -1380 6677 -1334 6715
rect -1380 6643 -1374 6677
rect -1340 6643 -1334 6677
rect -1380 6605 -1334 6643
rect -1380 6571 -1374 6605
rect -1340 6571 -1334 6605
rect -1380 6533 -1334 6571
rect -1380 6499 -1374 6533
rect -1340 6499 -1334 6533
rect -1380 6461 -1334 6499
rect -1380 6427 -1374 6461
rect -1340 6427 -1334 6461
rect -1380 6389 -1334 6427
rect -1380 6355 -1374 6389
rect -1340 6355 -1334 6389
rect -1380 6317 -1334 6355
rect -1380 6283 -1374 6317
rect -1340 6283 -1334 6317
rect -1380 6245 -1334 6283
rect -1380 6211 -1374 6245
rect -1340 6211 -1334 6245
rect -1380 6173 -1334 6211
rect -1380 6139 -1374 6173
rect -1340 6139 -1334 6173
rect -1380 6101 -1334 6139
rect -1380 6067 -1374 6101
rect -1340 6067 -1334 6101
rect -1380 6029 -1334 6067
rect -1380 5995 -1374 6029
rect -1340 5995 -1334 6029
rect -1380 5957 -1334 5995
rect -1380 5923 -1374 5957
rect -1340 5923 -1334 5957
rect -1380 5885 -1334 5923
rect -1380 5851 -1374 5885
rect -1340 5851 -1334 5885
rect -1380 5813 -1334 5851
rect -1380 5779 -1374 5813
rect -1340 5779 -1334 5813
rect -1380 5741 -1334 5779
rect -1380 5707 -1374 5741
rect -1340 5707 -1334 5741
rect -1380 5669 -1334 5707
rect -1380 5635 -1374 5669
rect -1340 5635 -1334 5669
rect -1380 5597 -1334 5635
rect -1380 5563 -1374 5597
rect -1340 5563 -1334 5597
rect -1380 5525 -1334 5563
rect -1380 5491 -1374 5525
rect -1340 5491 -1334 5525
rect -1380 5453 -1334 5491
rect -1380 5419 -1374 5453
rect -1340 5419 -1334 5453
rect -1380 5381 -1334 5419
rect -1380 5347 -1374 5381
rect -1340 5347 -1334 5381
rect -1380 5309 -1334 5347
rect -1380 5275 -1374 5309
rect -1340 5275 -1334 5309
rect -1380 5237 -1334 5275
rect -1380 5203 -1374 5237
rect -1340 5203 -1334 5237
rect -1380 5165 -1334 5203
rect -1380 5131 -1374 5165
rect -1340 5131 -1334 5165
rect -1380 5093 -1334 5131
rect -1380 5059 -1374 5093
rect -1340 5059 -1334 5093
rect -1380 5021 -1334 5059
rect -1380 4987 -1374 5021
rect -1340 4987 -1334 5021
rect -1380 4949 -1334 4987
rect -1380 4915 -1374 4949
rect -1340 4915 -1334 4949
rect -1380 4877 -1334 4915
rect -1380 4843 -1374 4877
rect -1340 4843 -1334 4877
rect -1380 4805 -1334 4843
rect -1380 4771 -1374 4805
rect -1340 4771 -1334 4805
rect -1380 4733 -1334 4771
rect -1380 4699 -1374 4733
rect -1340 4699 -1334 4733
rect -1380 4661 -1334 4699
rect -1380 4627 -1374 4661
rect -1340 4627 -1334 4661
rect -1380 4589 -1334 4627
rect -1380 4555 -1374 4589
rect -1340 4555 -1334 4589
rect -1380 4517 -1334 4555
rect -1380 4483 -1374 4517
rect -1340 4483 -1334 4517
rect -1380 4445 -1334 4483
rect -1380 4411 -1374 4445
rect -1340 4411 -1334 4445
rect -1380 4373 -1334 4411
rect -1380 4339 -1374 4373
rect -1340 4339 -1334 4373
rect -1380 4301 -1334 4339
rect -1380 4267 -1374 4301
rect -1340 4267 -1334 4301
rect -1380 4229 -1334 4267
rect -1380 4195 -1374 4229
rect -1340 4195 -1334 4229
rect -1380 4157 -1334 4195
rect -1380 4123 -1374 4157
rect -1340 4123 -1334 4157
rect -1380 4085 -1334 4123
rect -1380 4051 -1374 4085
rect -1340 4051 -1334 4085
rect -1380 4013 -1334 4051
rect -1380 3979 -1374 4013
rect -1340 3979 -1334 4013
rect -1380 3941 -1334 3979
rect -1380 3907 -1374 3941
rect -1340 3907 -1334 3941
rect -1380 3869 -1334 3907
rect -1380 3835 -1374 3869
rect -1340 3835 -1334 3869
rect -1380 3797 -1334 3835
rect -1380 3763 -1374 3797
rect -1340 3763 -1334 3797
rect -1380 3725 -1334 3763
rect -1380 3691 -1374 3725
rect -1340 3691 -1334 3725
rect -1380 3653 -1334 3691
rect -1380 3619 -1374 3653
rect -1340 3619 -1334 3653
rect -1380 3581 -1334 3619
rect -1380 3547 -1374 3581
rect -1340 3547 -1334 3581
rect -1380 3509 -1334 3547
rect -1380 3475 -1374 3509
rect -1340 3475 -1334 3509
rect -1380 3437 -1334 3475
rect -1380 3403 -1374 3437
rect -1340 3403 -1334 3437
rect -1380 3365 -1334 3403
rect -1380 3331 -1374 3365
rect -1340 3331 -1334 3365
rect -1380 3293 -1334 3331
rect -1380 3259 -1374 3293
rect -1340 3259 -1334 3293
rect -1380 3221 -1334 3259
rect -1380 3187 -1374 3221
rect -1340 3187 -1334 3221
rect -1380 3149 -1334 3187
rect -1380 3115 -1374 3149
rect -1340 3115 -1334 3149
rect -1380 3077 -1334 3115
rect -1380 3043 -1374 3077
rect -1340 3043 -1334 3077
rect -1380 3005 -1334 3043
rect -1380 2971 -1374 3005
rect -1340 2971 -1334 3005
rect -1380 2933 -1334 2971
rect -1380 2899 -1374 2933
rect -1340 2899 -1334 2933
rect -1380 2861 -1334 2899
rect -1380 2827 -1374 2861
rect -1340 2827 -1334 2861
rect -1380 2789 -1334 2827
rect -1380 2755 -1374 2789
rect -1340 2755 -1334 2789
rect -1380 2717 -1334 2755
rect -1380 2683 -1374 2717
rect -1340 2683 -1334 2717
rect -1380 2645 -1334 2683
rect -1380 2611 -1374 2645
rect -1340 2611 -1334 2645
rect -1380 2573 -1334 2611
rect -1380 2539 -1374 2573
rect -1340 2539 -1334 2573
rect -1380 2501 -1334 2539
rect -1380 2467 -1374 2501
rect -1340 2467 -1334 2501
rect -1380 2429 -1334 2467
rect -1380 2395 -1374 2429
rect -1340 2395 -1334 2429
rect -1380 2357 -1334 2395
rect -1380 2323 -1374 2357
rect -1340 2323 -1334 2357
rect -1380 2285 -1334 2323
rect -1380 2251 -1374 2285
rect -1340 2251 -1334 2285
rect -1380 2213 -1334 2251
rect -1380 2179 -1374 2213
rect -1340 2179 -1334 2213
rect -1380 2141 -1334 2179
rect -1380 2107 -1374 2141
rect -1340 2107 -1334 2141
rect -1380 2069 -1334 2107
rect -1380 2035 -1374 2069
rect -1340 2035 -1334 2069
rect -1380 1997 -1334 2035
rect -1380 1963 -1374 1997
rect -1340 1963 -1334 1997
rect -1380 1925 -1334 1963
rect -1380 1891 -1374 1925
rect -1340 1891 -1334 1925
rect -1380 1853 -1334 1891
rect -1380 1819 -1374 1853
rect -1340 1819 -1334 1853
rect -1380 1781 -1334 1819
rect -1380 1747 -1374 1781
rect -1340 1747 -1334 1781
rect -1380 1709 -1334 1747
rect -1380 1675 -1374 1709
rect -1340 1675 -1334 1709
rect -1380 1637 -1334 1675
rect -1380 1603 -1374 1637
rect -1340 1603 -1334 1637
rect -1380 1565 -1334 1603
rect -1380 1531 -1374 1565
rect -1340 1531 -1334 1565
rect -1380 1493 -1334 1531
rect -1380 1459 -1374 1493
rect -1340 1459 -1334 1493
rect -1380 1421 -1334 1459
rect -1380 1387 -1374 1421
rect -1340 1387 -1334 1421
rect -1380 1349 -1334 1387
rect -1380 1315 -1374 1349
rect -1340 1315 -1334 1349
rect -1380 1277 -1334 1315
rect -1380 1243 -1374 1277
rect -1340 1243 -1334 1277
rect -1380 1205 -1334 1243
rect -1380 1171 -1374 1205
rect -1340 1171 -1334 1205
rect -1380 1133 -1334 1171
rect -1380 1099 -1374 1133
rect -1340 1099 -1334 1133
rect -1380 1061 -1334 1099
rect -1380 1027 -1374 1061
rect -1340 1027 -1334 1061
rect -1380 989 -1334 1027
rect -1380 955 -1374 989
rect -1340 955 -1334 989
rect -1380 917 -1334 955
rect -1380 883 -1374 917
rect -1340 883 -1334 917
rect -1380 845 -1334 883
rect -1380 811 -1374 845
rect -1340 811 -1334 845
rect -1380 773 -1334 811
rect -1380 739 -1374 773
rect -1340 739 -1334 773
rect -1380 701 -1334 739
rect -1380 667 -1374 701
rect -1340 667 -1334 701
rect -1380 629 -1334 667
rect -1380 595 -1374 629
rect -1340 595 -1334 629
rect -1380 557 -1334 595
rect -1380 523 -1374 557
rect -1340 523 -1334 557
rect -1380 485 -1334 523
rect -1380 451 -1374 485
rect -1340 451 -1334 485
rect -1380 413 -1334 451
rect -1380 379 -1374 413
rect -1340 379 -1334 413
rect -1380 341 -1334 379
rect -1380 307 -1374 341
rect -1340 307 -1334 341
rect -1380 269 -1334 307
rect -1380 235 -1374 269
rect -1340 235 -1334 269
rect -1380 197 -1334 235
rect -1380 163 -1374 197
rect -1340 163 -1334 197
rect -1380 125 -1334 163
rect -1380 91 -1374 125
rect -1340 91 -1334 125
rect -1380 53 -1334 91
rect -1380 19 -1374 53
rect -1340 19 -1334 53
rect -1380 -19 -1334 19
rect -1380 -53 -1374 -19
rect -1340 -53 -1334 -19
rect -1380 -91 -1334 -53
rect -1380 -125 -1374 -91
rect -1340 -125 -1334 -91
rect -1380 -163 -1334 -125
rect -1380 -197 -1374 -163
rect -1340 -197 -1334 -163
rect -1380 -235 -1334 -197
rect -1380 -269 -1374 -235
rect -1340 -269 -1334 -235
rect -1380 -307 -1334 -269
rect -1380 -341 -1374 -307
rect -1340 -341 -1334 -307
rect -1380 -379 -1334 -341
rect -1380 -413 -1374 -379
rect -1340 -413 -1334 -379
rect -1380 -451 -1334 -413
rect -1380 -485 -1374 -451
rect -1340 -485 -1334 -451
rect -1380 -523 -1334 -485
rect -1380 -557 -1374 -523
rect -1340 -557 -1334 -523
rect -1380 -595 -1334 -557
rect -1380 -629 -1374 -595
rect -1340 -629 -1334 -595
rect -1380 -667 -1334 -629
rect -1380 -701 -1374 -667
rect -1340 -701 -1334 -667
rect -1380 -739 -1334 -701
rect -1380 -773 -1374 -739
rect -1340 -773 -1334 -739
rect -1380 -811 -1334 -773
rect -1380 -845 -1374 -811
rect -1340 -845 -1334 -811
rect -1380 -883 -1334 -845
rect -1380 -917 -1374 -883
rect -1340 -917 -1334 -883
rect -1380 -955 -1334 -917
rect -1380 -989 -1374 -955
rect -1340 -989 -1334 -955
rect -1380 -1027 -1334 -989
rect -1380 -1061 -1374 -1027
rect -1340 -1061 -1334 -1027
rect -1380 -1099 -1334 -1061
rect -1380 -1133 -1374 -1099
rect -1340 -1133 -1334 -1099
rect -1380 -1171 -1334 -1133
rect -1380 -1205 -1374 -1171
rect -1340 -1205 -1334 -1171
rect -1380 -1243 -1334 -1205
rect -1380 -1277 -1374 -1243
rect -1340 -1277 -1334 -1243
rect -1380 -1315 -1334 -1277
rect -1380 -1349 -1374 -1315
rect -1340 -1349 -1334 -1315
rect -1380 -1387 -1334 -1349
rect -1380 -1421 -1374 -1387
rect -1340 -1421 -1334 -1387
rect -1380 -1459 -1334 -1421
rect -1380 -1493 -1374 -1459
rect -1340 -1493 -1334 -1459
rect -1380 -1531 -1334 -1493
rect -1380 -1565 -1374 -1531
rect -1340 -1565 -1334 -1531
rect -1380 -1603 -1334 -1565
rect -1380 -1637 -1374 -1603
rect -1340 -1637 -1334 -1603
rect -1380 -1675 -1334 -1637
rect -1380 -1709 -1374 -1675
rect -1340 -1709 -1334 -1675
rect -1380 -1747 -1334 -1709
rect -1380 -1781 -1374 -1747
rect -1340 -1781 -1334 -1747
rect -1380 -1819 -1334 -1781
rect -1380 -1853 -1374 -1819
rect -1340 -1853 -1334 -1819
rect -1380 -1891 -1334 -1853
rect -1380 -1925 -1374 -1891
rect -1340 -1925 -1334 -1891
rect -1380 -1963 -1334 -1925
rect -1380 -1997 -1374 -1963
rect -1340 -1997 -1334 -1963
rect -1380 -2035 -1334 -1997
rect -1380 -2069 -1374 -2035
rect -1340 -2069 -1334 -2035
rect -1380 -2107 -1334 -2069
rect -1380 -2141 -1374 -2107
rect -1340 -2141 -1334 -2107
rect -1380 -2179 -1334 -2141
rect -1380 -2213 -1374 -2179
rect -1340 -2213 -1334 -2179
rect -1380 -2251 -1334 -2213
rect -1380 -2285 -1374 -2251
rect -1340 -2285 -1334 -2251
rect -1380 -2323 -1334 -2285
rect -1380 -2357 -1374 -2323
rect -1340 -2357 -1334 -2323
rect -1380 -2395 -1334 -2357
rect -1380 -2429 -1374 -2395
rect -1340 -2429 -1334 -2395
rect -1380 -2467 -1334 -2429
rect -1380 -2501 -1374 -2467
rect -1340 -2501 -1334 -2467
rect -1380 -2539 -1334 -2501
rect -1380 -2573 -1374 -2539
rect -1340 -2573 -1334 -2539
rect -1380 -2611 -1334 -2573
rect -1380 -2645 -1374 -2611
rect -1340 -2645 -1334 -2611
rect -1380 -2683 -1334 -2645
rect -1380 -2717 -1374 -2683
rect -1340 -2717 -1334 -2683
rect -1380 -2755 -1334 -2717
rect -1380 -2789 -1374 -2755
rect -1340 -2789 -1334 -2755
rect -1380 -2827 -1334 -2789
rect -1380 -2861 -1374 -2827
rect -1340 -2861 -1334 -2827
rect -1380 -2899 -1334 -2861
rect -1380 -2933 -1374 -2899
rect -1340 -2933 -1334 -2899
rect -1380 -2971 -1334 -2933
rect -1380 -3005 -1374 -2971
rect -1340 -3005 -1334 -2971
rect -1380 -3043 -1334 -3005
rect -1380 -3077 -1374 -3043
rect -1340 -3077 -1334 -3043
rect -1380 -3115 -1334 -3077
rect -1380 -3149 -1374 -3115
rect -1340 -3149 -1334 -3115
rect -1380 -3187 -1334 -3149
rect -1380 -3221 -1374 -3187
rect -1340 -3221 -1334 -3187
rect -1380 -3259 -1334 -3221
rect -1380 -3293 -1374 -3259
rect -1340 -3293 -1334 -3259
rect -1380 -3331 -1334 -3293
rect -1380 -3365 -1374 -3331
rect -1340 -3365 -1334 -3331
rect -1380 -3403 -1334 -3365
rect -1380 -3437 -1374 -3403
rect -1340 -3437 -1334 -3403
rect -1380 -3475 -1334 -3437
rect -1380 -3509 -1374 -3475
rect -1340 -3509 -1334 -3475
rect -1380 -3547 -1334 -3509
rect -1380 -3581 -1374 -3547
rect -1340 -3581 -1334 -3547
rect -1380 -3619 -1334 -3581
rect -1380 -3653 -1374 -3619
rect -1340 -3653 -1334 -3619
rect -1380 -3691 -1334 -3653
rect -1380 -3725 -1374 -3691
rect -1340 -3725 -1334 -3691
rect -1380 -3763 -1334 -3725
rect -1380 -3797 -1374 -3763
rect -1340 -3797 -1334 -3763
rect -1380 -3835 -1334 -3797
rect -1380 -3869 -1374 -3835
rect -1340 -3869 -1334 -3835
rect -1380 -3907 -1334 -3869
rect -1380 -3941 -1374 -3907
rect -1340 -3941 -1334 -3907
rect -1380 -3979 -1334 -3941
rect -1380 -4013 -1374 -3979
rect -1340 -4013 -1334 -3979
rect -1380 -4051 -1334 -4013
rect -1380 -4085 -1374 -4051
rect -1340 -4085 -1334 -4051
rect -1380 -4123 -1334 -4085
rect -1380 -4157 -1374 -4123
rect -1340 -4157 -1334 -4123
rect -1380 -4195 -1334 -4157
rect -1380 -4229 -1374 -4195
rect -1340 -4229 -1334 -4195
rect -1380 -4267 -1334 -4229
rect -1380 -4301 -1374 -4267
rect -1340 -4301 -1334 -4267
rect -1380 -4339 -1334 -4301
rect -1380 -4373 -1374 -4339
rect -1340 -4373 -1334 -4339
rect -1380 -4411 -1334 -4373
rect -1380 -4445 -1374 -4411
rect -1340 -4445 -1334 -4411
rect -1380 -4483 -1334 -4445
rect -1380 -4517 -1374 -4483
rect -1340 -4517 -1334 -4483
rect -1380 -4555 -1334 -4517
rect -1380 -4589 -1374 -4555
rect -1340 -4589 -1334 -4555
rect -1380 -4627 -1334 -4589
rect -1380 -4661 -1374 -4627
rect -1340 -4661 -1334 -4627
rect -1380 -4699 -1334 -4661
rect -1380 -4733 -1374 -4699
rect -1340 -4733 -1334 -4699
rect -1380 -4771 -1334 -4733
rect -1380 -4805 -1374 -4771
rect -1340 -4805 -1334 -4771
rect -1380 -4843 -1334 -4805
rect -1380 -4877 -1374 -4843
rect -1340 -4877 -1334 -4843
rect -1380 -4915 -1334 -4877
rect -1380 -4949 -1374 -4915
rect -1340 -4949 -1334 -4915
rect -1380 -4987 -1334 -4949
rect -1380 -5021 -1374 -4987
rect -1340 -5021 -1334 -4987
rect -1380 -5059 -1334 -5021
rect -1380 -5093 -1374 -5059
rect -1340 -5093 -1334 -5059
rect -1380 -5131 -1334 -5093
rect -1380 -5165 -1374 -5131
rect -1340 -5165 -1334 -5131
rect -1380 -5203 -1334 -5165
rect -1380 -5237 -1374 -5203
rect -1340 -5237 -1334 -5203
rect -1380 -5275 -1334 -5237
rect -1380 -5309 -1374 -5275
rect -1340 -5309 -1334 -5275
rect -1380 -5347 -1334 -5309
rect -1380 -5381 -1374 -5347
rect -1340 -5381 -1334 -5347
rect -1380 -5419 -1334 -5381
rect -1380 -5453 -1374 -5419
rect -1340 -5453 -1334 -5419
rect -1380 -5491 -1334 -5453
rect -1380 -5525 -1374 -5491
rect -1340 -5525 -1334 -5491
rect -1380 -5563 -1334 -5525
rect -1380 -5597 -1374 -5563
rect -1340 -5597 -1334 -5563
rect -1380 -5635 -1334 -5597
rect -1380 -5669 -1374 -5635
rect -1340 -5669 -1334 -5635
rect -1380 -5707 -1334 -5669
rect -1380 -5741 -1374 -5707
rect -1340 -5741 -1334 -5707
rect -1380 -5779 -1334 -5741
rect -1380 -5813 -1374 -5779
rect -1340 -5813 -1334 -5779
rect -1380 -5851 -1334 -5813
rect -1380 -5885 -1374 -5851
rect -1340 -5885 -1334 -5851
rect -1380 -5923 -1334 -5885
rect -1380 -5957 -1374 -5923
rect -1340 -5957 -1334 -5923
rect -1380 -5995 -1334 -5957
rect -1380 -6029 -1374 -5995
rect -1340 -6029 -1334 -5995
rect -1380 -6067 -1334 -6029
rect -1380 -6101 -1374 -6067
rect -1340 -6101 -1334 -6067
rect -1380 -6139 -1334 -6101
rect -1380 -6173 -1374 -6139
rect -1340 -6173 -1334 -6139
rect -1380 -6211 -1334 -6173
rect -1380 -6245 -1374 -6211
rect -1340 -6245 -1334 -6211
rect -1380 -6283 -1334 -6245
rect -1380 -6317 -1374 -6283
rect -1340 -6317 -1334 -6283
rect -1380 -6355 -1334 -6317
rect -1380 -6389 -1374 -6355
rect -1340 -6389 -1334 -6355
rect -1380 -6427 -1334 -6389
rect -1380 -6461 -1374 -6427
rect -1340 -6461 -1334 -6427
rect -1380 -6499 -1334 -6461
rect -1380 -6533 -1374 -6499
rect -1340 -6533 -1334 -6499
rect -1380 -6571 -1334 -6533
rect -1380 -6605 -1374 -6571
rect -1340 -6605 -1334 -6571
rect -1380 -6643 -1334 -6605
rect -1380 -6677 -1374 -6643
rect -1340 -6677 -1334 -6643
rect -1380 -6715 -1334 -6677
rect -1380 -6749 -1374 -6715
rect -1340 -6749 -1334 -6715
rect -1380 -6787 -1334 -6749
rect -1380 -6821 -1374 -6787
rect -1340 -6821 -1334 -6787
rect -1380 -6859 -1334 -6821
rect -1380 -6893 -1374 -6859
rect -1340 -6893 -1334 -6859
rect -1380 -6931 -1334 -6893
rect -1380 -6965 -1374 -6931
rect -1340 -6965 -1334 -6931
rect -1380 -7003 -1334 -6965
rect -1380 -7037 -1374 -7003
rect -1340 -7037 -1334 -7003
rect -1380 -7075 -1334 -7037
rect -1380 -7109 -1374 -7075
rect -1340 -7109 -1334 -7075
rect -1380 -7147 -1334 -7109
rect -1380 -7181 -1374 -7147
rect -1340 -7181 -1334 -7147
rect -1380 -7219 -1334 -7181
rect -1380 -7253 -1374 -7219
rect -1340 -7253 -1334 -7219
rect -1380 -7291 -1334 -7253
rect -1380 -7325 -1374 -7291
rect -1340 -7325 -1334 -7291
rect -1380 -7363 -1334 -7325
rect -1380 -7397 -1374 -7363
rect -1340 -7397 -1334 -7363
rect -1380 -7435 -1334 -7397
rect -1380 -7469 -1374 -7435
rect -1340 -7469 -1334 -7435
rect -1380 -7507 -1334 -7469
rect -1380 -7541 -1374 -7507
rect -1340 -7541 -1334 -7507
rect -1380 -7579 -1334 -7541
rect -1380 -7613 -1374 -7579
rect -1340 -7613 -1334 -7579
rect -1380 -7651 -1334 -7613
rect -1380 -7685 -1374 -7651
rect -1340 -7685 -1334 -7651
rect -1380 -7723 -1334 -7685
rect -1380 -7757 -1374 -7723
rect -1340 -7757 -1334 -7723
rect -1380 -7795 -1334 -7757
rect -1380 -7829 -1374 -7795
rect -1340 -7829 -1334 -7795
rect -1380 -7867 -1334 -7829
rect -1380 -7901 -1374 -7867
rect -1340 -7901 -1334 -7867
rect -1380 -7939 -1334 -7901
rect -1380 -7973 -1374 -7939
rect -1340 -7973 -1334 -7939
rect -1380 -8011 -1334 -7973
rect -1380 -8045 -1374 -8011
rect -1340 -8045 -1334 -8011
rect -1380 -8083 -1334 -8045
rect -1380 -8117 -1374 -8083
rect -1340 -8117 -1334 -8083
rect -1380 -8155 -1334 -8117
rect -1380 -8189 -1374 -8155
rect -1340 -8189 -1334 -8155
rect -1380 -8227 -1334 -8189
rect -1380 -8261 -1374 -8227
rect -1340 -8261 -1334 -8227
rect -1380 -8299 -1334 -8261
rect -1380 -8333 -1374 -8299
rect -1340 -8333 -1334 -8299
rect -1380 -8371 -1334 -8333
rect -1380 -8405 -1374 -8371
rect -1340 -8405 -1334 -8371
rect -1380 -8443 -1334 -8405
rect -1380 -8477 -1374 -8443
rect -1340 -8477 -1334 -8443
rect -1380 -8515 -1334 -8477
rect -1380 -8549 -1374 -8515
rect -1340 -8549 -1334 -8515
rect -1380 -8587 -1334 -8549
rect -1380 -8621 -1374 -8587
rect -1340 -8621 -1334 -8587
rect -1380 -8659 -1334 -8621
rect -1380 -8693 -1374 -8659
rect -1340 -8693 -1334 -8659
rect -1380 -8731 -1334 -8693
rect -1380 -8765 -1374 -8731
rect -1340 -8765 -1334 -8731
rect -1380 -8803 -1334 -8765
rect -1380 -8837 -1374 -8803
rect -1340 -8837 -1334 -8803
rect -1380 -8875 -1334 -8837
rect -1380 -8909 -1374 -8875
rect -1340 -8909 -1334 -8875
rect -1380 -8947 -1334 -8909
rect -1380 -8981 -1374 -8947
rect -1340 -8981 -1334 -8947
rect -1380 -9019 -1334 -8981
rect -1380 -9053 -1374 -9019
rect -1340 -9053 -1334 -9019
rect -1380 -9091 -1334 -9053
rect -1380 -9125 -1374 -9091
rect -1340 -9125 -1334 -9091
rect -1380 -9163 -1334 -9125
rect -1380 -9197 -1374 -9163
rect -1340 -9197 -1334 -9163
rect -1380 -9235 -1334 -9197
rect -1380 -9269 -1374 -9235
rect -1340 -9269 -1334 -9235
rect -1380 -9307 -1334 -9269
rect -1380 -9341 -1374 -9307
rect -1340 -9341 -1334 -9307
rect -1380 -9379 -1334 -9341
rect -1380 -9413 -1374 -9379
rect -1340 -9413 -1334 -9379
rect -1380 -9451 -1334 -9413
rect -1380 -9485 -1374 -9451
rect -1340 -9485 -1334 -9451
rect -1380 -9523 -1334 -9485
rect -1380 -9557 -1374 -9523
rect -1340 -9557 -1334 -9523
rect -1380 -9600 -1334 -9557
rect -1262 9557 -1216 9600
rect -1262 9523 -1256 9557
rect -1222 9523 -1216 9557
rect -1262 9485 -1216 9523
rect -1262 9451 -1256 9485
rect -1222 9451 -1216 9485
rect -1262 9413 -1216 9451
rect -1262 9379 -1256 9413
rect -1222 9379 -1216 9413
rect -1262 9341 -1216 9379
rect -1262 9307 -1256 9341
rect -1222 9307 -1216 9341
rect -1262 9269 -1216 9307
rect -1262 9235 -1256 9269
rect -1222 9235 -1216 9269
rect -1262 9197 -1216 9235
rect -1262 9163 -1256 9197
rect -1222 9163 -1216 9197
rect -1262 9125 -1216 9163
rect -1262 9091 -1256 9125
rect -1222 9091 -1216 9125
rect -1262 9053 -1216 9091
rect -1262 9019 -1256 9053
rect -1222 9019 -1216 9053
rect -1262 8981 -1216 9019
rect -1262 8947 -1256 8981
rect -1222 8947 -1216 8981
rect -1262 8909 -1216 8947
rect -1262 8875 -1256 8909
rect -1222 8875 -1216 8909
rect -1262 8837 -1216 8875
rect -1262 8803 -1256 8837
rect -1222 8803 -1216 8837
rect -1262 8765 -1216 8803
rect -1262 8731 -1256 8765
rect -1222 8731 -1216 8765
rect -1262 8693 -1216 8731
rect -1262 8659 -1256 8693
rect -1222 8659 -1216 8693
rect -1262 8621 -1216 8659
rect -1262 8587 -1256 8621
rect -1222 8587 -1216 8621
rect -1262 8549 -1216 8587
rect -1262 8515 -1256 8549
rect -1222 8515 -1216 8549
rect -1262 8477 -1216 8515
rect -1262 8443 -1256 8477
rect -1222 8443 -1216 8477
rect -1262 8405 -1216 8443
rect -1262 8371 -1256 8405
rect -1222 8371 -1216 8405
rect -1262 8333 -1216 8371
rect -1262 8299 -1256 8333
rect -1222 8299 -1216 8333
rect -1262 8261 -1216 8299
rect -1262 8227 -1256 8261
rect -1222 8227 -1216 8261
rect -1262 8189 -1216 8227
rect -1262 8155 -1256 8189
rect -1222 8155 -1216 8189
rect -1262 8117 -1216 8155
rect -1262 8083 -1256 8117
rect -1222 8083 -1216 8117
rect -1262 8045 -1216 8083
rect -1262 8011 -1256 8045
rect -1222 8011 -1216 8045
rect -1262 7973 -1216 8011
rect -1262 7939 -1256 7973
rect -1222 7939 -1216 7973
rect -1262 7901 -1216 7939
rect -1262 7867 -1256 7901
rect -1222 7867 -1216 7901
rect -1262 7829 -1216 7867
rect -1262 7795 -1256 7829
rect -1222 7795 -1216 7829
rect -1262 7757 -1216 7795
rect -1262 7723 -1256 7757
rect -1222 7723 -1216 7757
rect -1262 7685 -1216 7723
rect -1262 7651 -1256 7685
rect -1222 7651 -1216 7685
rect -1262 7613 -1216 7651
rect -1262 7579 -1256 7613
rect -1222 7579 -1216 7613
rect -1262 7541 -1216 7579
rect -1262 7507 -1256 7541
rect -1222 7507 -1216 7541
rect -1262 7469 -1216 7507
rect -1262 7435 -1256 7469
rect -1222 7435 -1216 7469
rect -1262 7397 -1216 7435
rect -1262 7363 -1256 7397
rect -1222 7363 -1216 7397
rect -1262 7325 -1216 7363
rect -1262 7291 -1256 7325
rect -1222 7291 -1216 7325
rect -1262 7253 -1216 7291
rect -1262 7219 -1256 7253
rect -1222 7219 -1216 7253
rect -1262 7181 -1216 7219
rect -1262 7147 -1256 7181
rect -1222 7147 -1216 7181
rect -1262 7109 -1216 7147
rect -1262 7075 -1256 7109
rect -1222 7075 -1216 7109
rect -1262 7037 -1216 7075
rect -1262 7003 -1256 7037
rect -1222 7003 -1216 7037
rect -1262 6965 -1216 7003
rect -1262 6931 -1256 6965
rect -1222 6931 -1216 6965
rect -1262 6893 -1216 6931
rect -1262 6859 -1256 6893
rect -1222 6859 -1216 6893
rect -1262 6821 -1216 6859
rect -1262 6787 -1256 6821
rect -1222 6787 -1216 6821
rect -1262 6749 -1216 6787
rect -1262 6715 -1256 6749
rect -1222 6715 -1216 6749
rect -1262 6677 -1216 6715
rect -1262 6643 -1256 6677
rect -1222 6643 -1216 6677
rect -1262 6605 -1216 6643
rect -1262 6571 -1256 6605
rect -1222 6571 -1216 6605
rect -1262 6533 -1216 6571
rect -1262 6499 -1256 6533
rect -1222 6499 -1216 6533
rect -1262 6461 -1216 6499
rect -1262 6427 -1256 6461
rect -1222 6427 -1216 6461
rect -1262 6389 -1216 6427
rect -1262 6355 -1256 6389
rect -1222 6355 -1216 6389
rect -1262 6317 -1216 6355
rect -1262 6283 -1256 6317
rect -1222 6283 -1216 6317
rect -1262 6245 -1216 6283
rect -1262 6211 -1256 6245
rect -1222 6211 -1216 6245
rect -1262 6173 -1216 6211
rect -1262 6139 -1256 6173
rect -1222 6139 -1216 6173
rect -1262 6101 -1216 6139
rect -1262 6067 -1256 6101
rect -1222 6067 -1216 6101
rect -1262 6029 -1216 6067
rect -1262 5995 -1256 6029
rect -1222 5995 -1216 6029
rect -1262 5957 -1216 5995
rect -1262 5923 -1256 5957
rect -1222 5923 -1216 5957
rect -1262 5885 -1216 5923
rect -1262 5851 -1256 5885
rect -1222 5851 -1216 5885
rect -1262 5813 -1216 5851
rect -1262 5779 -1256 5813
rect -1222 5779 -1216 5813
rect -1262 5741 -1216 5779
rect -1262 5707 -1256 5741
rect -1222 5707 -1216 5741
rect -1262 5669 -1216 5707
rect -1262 5635 -1256 5669
rect -1222 5635 -1216 5669
rect -1262 5597 -1216 5635
rect -1262 5563 -1256 5597
rect -1222 5563 -1216 5597
rect -1262 5525 -1216 5563
rect -1262 5491 -1256 5525
rect -1222 5491 -1216 5525
rect -1262 5453 -1216 5491
rect -1262 5419 -1256 5453
rect -1222 5419 -1216 5453
rect -1262 5381 -1216 5419
rect -1262 5347 -1256 5381
rect -1222 5347 -1216 5381
rect -1262 5309 -1216 5347
rect -1262 5275 -1256 5309
rect -1222 5275 -1216 5309
rect -1262 5237 -1216 5275
rect -1262 5203 -1256 5237
rect -1222 5203 -1216 5237
rect -1262 5165 -1216 5203
rect -1262 5131 -1256 5165
rect -1222 5131 -1216 5165
rect -1262 5093 -1216 5131
rect -1262 5059 -1256 5093
rect -1222 5059 -1216 5093
rect -1262 5021 -1216 5059
rect -1262 4987 -1256 5021
rect -1222 4987 -1216 5021
rect -1262 4949 -1216 4987
rect -1262 4915 -1256 4949
rect -1222 4915 -1216 4949
rect -1262 4877 -1216 4915
rect -1262 4843 -1256 4877
rect -1222 4843 -1216 4877
rect -1262 4805 -1216 4843
rect -1262 4771 -1256 4805
rect -1222 4771 -1216 4805
rect -1262 4733 -1216 4771
rect -1262 4699 -1256 4733
rect -1222 4699 -1216 4733
rect -1262 4661 -1216 4699
rect -1262 4627 -1256 4661
rect -1222 4627 -1216 4661
rect -1262 4589 -1216 4627
rect -1262 4555 -1256 4589
rect -1222 4555 -1216 4589
rect -1262 4517 -1216 4555
rect -1262 4483 -1256 4517
rect -1222 4483 -1216 4517
rect -1262 4445 -1216 4483
rect -1262 4411 -1256 4445
rect -1222 4411 -1216 4445
rect -1262 4373 -1216 4411
rect -1262 4339 -1256 4373
rect -1222 4339 -1216 4373
rect -1262 4301 -1216 4339
rect -1262 4267 -1256 4301
rect -1222 4267 -1216 4301
rect -1262 4229 -1216 4267
rect -1262 4195 -1256 4229
rect -1222 4195 -1216 4229
rect -1262 4157 -1216 4195
rect -1262 4123 -1256 4157
rect -1222 4123 -1216 4157
rect -1262 4085 -1216 4123
rect -1262 4051 -1256 4085
rect -1222 4051 -1216 4085
rect -1262 4013 -1216 4051
rect -1262 3979 -1256 4013
rect -1222 3979 -1216 4013
rect -1262 3941 -1216 3979
rect -1262 3907 -1256 3941
rect -1222 3907 -1216 3941
rect -1262 3869 -1216 3907
rect -1262 3835 -1256 3869
rect -1222 3835 -1216 3869
rect -1262 3797 -1216 3835
rect -1262 3763 -1256 3797
rect -1222 3763 -1216 3797
rect -1262 3725 -1216 3763
rect -1262 3691 -1256 3725
rect -1222 3691 -1216 3725
rect -1262 3653 -1216 3691
rect -1262 3619 -1256 3653
rect -1222 3619 -1216 3653
rect -1262 3581 -1216 3619
rect -1262 3547 -1256 3581
rect -1222 3547 -1216 3581
rect -1262 3509 -1216 3547
rect -1262 3475 -1256 3509
rect -1222 3475 -1216 3509
rect -1262 3437 -1216 3475
rect -1262 3403 -1256 3437
rect -1222 3403 -1216 3437
rect -1262 3365 -1216 3403
rect -1262 3331 -1256 3365
rect -1222 3331 -1216 3365
rect -1262 3293 -1216 3331
rect -1262 3259 -1256 3293
rect -1222 3259 -1216 3293
rect -1262 3221 -1216 3259
rect -1262 3187 -1256 3221
rect -1222 3187 -1216 3221
rect -1262 3149 -1216 3187
rect -1262 3115 -1256 3149
rect -1222 3115 -1216 3149
rect -1262 3077 -1216 3115
rect -1262 3043 -1256 3077
rect -1222 3043 -1216 3077
rect -1262 3005 -1216 3043
rect -1262 2971 -1256 3005
rect -1222 2971 -1216 3005
rect -1262 2933 -1216 2971
rect -1262 2899 -1256 2933
rect -1222 2899 -1216 2933
rect -1262 2861 -1216 2899
rect -1262 2827 -1256 2861
rect -1222 2827 -1216 2861
rect -1262 2789 -1216 2827
rect -1262 2755 -1256 2789
rect -1222 2755 -1216 2789
rect -1262 2717 -1216 2755
rect -1262 2683 -1256 2717
rect -1222 2683 -1216 2717
rect -1262 2645 -1216 2683
rect -1262 2611 -1256 2645
rect -1222 2611 -1216 2645
rect -1262 2573 -1216 2611
rect -1262 2539 -1256 2573
rect -1222 2539 -1216 2573
rect -1262 2501 -1216 2539
rect -1262 2467 -1256 2501
rect -1222 2467 -1216 2501
rect -1262 2429 -1216 2467
rect -1262 2395 -1256 2429
rect -1222 2395 -1216 2429
rect -1262 2357 -1216 2395
rect -1262 2323 -1256 2357
rect -1222 2323 -1216 2357
rect -1262 2285 -1216 2323
rect -1262 2251 -1256 2285
rect -1222 2251 -1216 2285
rect -1262 2213 -1216 2251
rect -1262 2179 -1256 2213
rect -1222 2179 -1216 2213
rect -1262 2141 -1216 2179
rect -1262 2107 -1256 2141
rect -1222 2107 -1216 2141
rect -1262 2069 -1216 2107
rect -1262 2035 -1256 2069
rect -1222 2035 -1216 2069
rect -1262 1997 -1216 2035
rect -1262 1963 -1256 1997
rect -1222 1963 -1216 1997
rect -1262 1925 -1216 1963
rect -1262 1891 -1256 1925
rect -1222 1891 -1216 1925
rect -1262 1853 -1216 1891
rect -1262 1819 -1256 1853
rect -1222 1819 -1216 1853
rect -1262 1781 -1216 1819
rect -1262 1747 -1256 1781
rect -1222 1747 -1216 1781
rect -1262 1709 -1216 1747
rect -1262 1675 -1256 1709
rect -1222 1675 -1216 1709
rect -1262 1637 -1216 1675
rect -1262 1603 -1256 1637
rect -1222 1603 -1216 1637
rect -1262 1565 -1216 1603
rect -1262 1531 -1256 1565
rect -1222 1531 -1216 1565
rect -1262 1493 -1216 1531
rect -1262 1459 -1256 1493
rect -1222 1459 -1216 1493
rect -1262 1421 -1216 1459
rect -1262 1387 -1256 1421
rect -1222 1387 -1216 1421
rect -1262 1349 -1216 1387
rect -1262 1315 -1256 1349
rect -1222 1315 -1216 1349
rect -1262 1277 -1216 1315
rect -1262 1243 -1256 1277
rect -1222 1243 -1216 1277
rect -1262 1205 -1216 1243
rect -1262 1171 -1256 1205
rect -1222 1171 -1216 1205
rect -1262 1133 -1216 1171
rect -1262 1099 -1256 1133
rect -1222 1099 -1216 1133
rect -1262 1061 -1216 1099
rect -1262 1027 -1256 1061
rect -1222 1027 -1216 1061
rect -1262 989 -1216 1027
rect -1262 955 -1256 989
rect -1222 955 -1216 989
rect -1262 917 -1216 955
rect -1262 883 -1256 917
rect -1222 883 -1216 917
rect -1262 845 -1216 883
rect -1262 811 -1256 845
rect -1222 811 -1216 845
rect -1262 773 -1216 811
rect -1262 739 -1256 773
rect -1222 739 -1216 773
rect -1262 701 -1216 739
rect -1262 667 -1256 701
rect -1222 667 -1216 701
rect -1262 629 -1216 667
rect -1262 595 -1256 629
rect -1222 595 -1216 629
rect -1262 557 -1216 595
rect -1262 523 -1256 557
rect -1222 523 -1216 557
rect -1262 485 -1216 523
rect -1262 451 -1256 485
rect -1222 451 -1216 485
rect -1262 413 -1216 451
rect -1262 379 -1256 413
rect -1222 379 -1216 413
rect -1262 341 -1216 379
rect -1262 307 -1256 341
rect -1222 307 -1216 341
rect -1262 269 -1216 307
rect -1262 235 -1256 269
rect -1222 235 -1216 269
rect -1262 197 -1216 235
rect -1262 163 -1256 197
rect -1222 163 -1216 197
rect -1262 125 -1216 163
rect -1262 91 -1256 125
rect -1222 91 -1216 125
rect -1262 53 -1216 91
rect -1262 19 -1256 53
rect -1222 19 -1216 53
rect -1262 -19 -1216 19
rect -1262 -53 -1256 -19
rect -1222 -53 -1216 -19
rect -1262 -91 -1216 -53
rect -1262 -125 -1256 -91
rect -1222 -125 -1216 -91
rect -1262 -163 -1216 -125
rect -1262 -197 -1256 -163
rect -1222 -197 -1216 -163
rect -1262 -235 -1216 -197
rect -1262 -269 -1256 -235
rect -1222 -269 -1216 -235
rect -1262 -307 -1216 -269
rect -1262 -341 -1256 -307
rect -1222 -341 -1216 -307
rect -1262 -379 -1216 -341
rect -1262 -413 -1256 -379
rect -1222 -413 -1216 -379
rect -1262 -451 -1216 -413
rect -1262 -485 -1256 -451
rect -1222 -485 -1216 -451
rect -1262 -523 -1216 -485
rect -1262 -557 -1256 -523
rect -1222 -557 -1216 -523
rect -1262 -595 -1216 -557
rect -1262 -629 -1256 -595
rect -1222 -629 -1216 -595
rect -1262 -667 -1216 -629
rect -1262 -701 -1256 -667
rect -1222 -701 -1216 -667
rect -1262 -739 -1216 -701
rect -1262 -773 -1256 -739
rect -1222 -773 -1216 -739
rect -1262 -811 -1216 -773
rect -1262 -845 -1256 -811
rect -1222 -845 -1216 -811
rect -1262 -883 -1216 -845
rect -1262 -917 -1256 -883
rect -1222 -917 -1216 -883
rect -1262 -955 -1216 -917
rect -1262 -989 -1256 -955
rect -1222 -989 -1216 -955
rect -1262 -1027 -1216 -989
rect -1262 -1061 -1256 -1027
rect -1222 -1061 -1216 -1027
rect -1262 -1099 -1216 -1061
rect -1262 -1133 -1256 -1099
rect -1222 -1133 -1216 -1099
rect -1262 -1171 -1216 -1133
rect -1262 -1205 -1256 -1171
rect -1222 -1205 -1216 -1171
rect -1262 -1243 -1216 -1205
rect -1262 -1277 -1256 -1243
rect -1222 -1277 -1216 -1243
rect -1262 -1315 -1216 -1277
rect -1262 -1349 -1256 -1315
rect -1222 -1349 -1216 -1315
rect -1262 -1387 -1216 -1349
rect -1262 -1421 -1256 -1387
rect -1222 -1421 -1216 -1387
rect -1262 -1459 -1216 -1421
rect -1262 -1493 -1256 -1459
rect -1222 -1493 -1216 -1459
rect -1262 -1531 -1216 -1493
rect -1262 -1565 -1256 -1531
rect -1222 -1565 -1216 -1531
rect -1262 -1603 -1216 -1565
rect -1262 -1637 -1256 -1603
rect -1222 -1637 -1216 -1603
rect -1262 -1675 -1216 -1637
rect -1262 -1709 -1256 -1675
rect -1222 -1709 -1216 -1675
rect -1262 -1747 -1216 -1709
rect -1262 -1781 -1256 -1747
rect -1222 -1781 -1216 -1747
rect -1262 -1819 -1216 -1781
rect -1262 -1853 -1256 -1819
rect -1222 -1853 -1216 -1819
rect -1262 -1891 -1216 -1853
rect -1262 -1925 -1256 -1891
rect -1222 -1925 -1216 -1891
rect -1262 -1963 -1216 -1925
rect -1262 -1997 -1256 -1963
rect -1222 -1997 -1216 -1963
rect -1262 -2035 -1216 -1997
rect -1262 -2069 -1256 -2035
rect -1222 -2069 -1216 -2035
rect -1262 -2107 -1216 -2069
rect -1262 -2141 -1256 -2107
rect -1222 -2141 -1216 -2107
rect -1262 -2179 -1216 -2141
rect -1262 -2213 -1256 -2179
rect -1222 -2213 -1216 -2179
rect -1262 -2251 -1216 -2213
rect -1262 -2285 -1256 -2251
rect -1222 -2285 -1216 -2251
rect -1262 -2323 -1216 -2285
rect -1262 -2357 -1256 -2323
rect -1222 -2357 -1216 -2323
rect -1262 -2395 -1216 -2357
rect -1262 -2429 -1256 -2395
rect -1222 -2429 -1216 -2395
rect -1262 -2467 -1216 -2429
rect -1262 -2501 -1256 -2467
rect -1222 -2501 -1216 -2467
rect -1262 -2539 -1216 -2501
rect -1262 -2573 -1256 -2539
rect -1222 -2573 -1216 -2539
rect -1262 -2611 -1216 -2573
rect -1262 -2645 -1256 -2611
rect -1222 -2645 -1216 -2611
rect -1262 -2683 -1216 -2645
rect -1262 -2717 -1256 -2683
rect -1222 -2717 -1216 -2683
rect -1262 -2755 -1216 -2717
rect -1262 -2789 -1256 -2755
rect -1222 -2789 -1216 -2755
rect -1262 -2827 -1216 -2789
rect -1262 -2861 -1256 -2827
rect -1222 -2861 -1216 -2827
rect -1262 -2899 -1216 -2861
rect -1262 -2933 -1256 -2899
rect -1222 -2933 -1216 -2899
rect -1262 -2971 -1216 -2933
rect -1262 -3005 -1256 -2971
rect -1222 -3005 -1216 -2971
rect -1262 -3043 -1216 -3005
rect -1262 -3077 -1256 -3043
rect -1222 -3077 -1216 -3043
rect -1262 -3115 -1216 -3077
rect -1262 -3149 -1256 -3115
rect -1222 -3149 -1216 -3115
rect -1262 -3187 -1216 -3149
rect -1262 -3221 -1256 -3187
rect -1222 -3221 -1216 -3187
rect -1262 -3259 -1216 -3221
rect -1262 -3293 -1256 -3259
rect -1222 -3293 -1216 -3259
rect -1262 -3331 -1216 -3293
rect -1262 -3365 -1256 -3331
rect -1222 -3365 -1216 -3331
rect -1262 -3403 -1216 -3365
rect -1262 -3437 -1256 -3403
rect -1222 -3437 -1216 -3403
rect -1262 -3475 -1216 -3437
rect -1262 -3509 -1256 -3475
rect -1222 -3509 -1216 -3475
rect -1262 -3547 -1216 -3509
rect -1262 -3581 -1256 -3547
rect -1222 -3581 -1216 -3547
rect -1262 -3619 -1216 -3581
rect -1262 -3653 -1256 -3619
rect -1222 -3653 -1216 -3619
rect -1262 -3691 -1216 -3653
rect -1262 -3725 -1256 -3691
rect -1222 -3725 -1216 -3691
rect -1262 -3763 -1216 -3725
rect -1262 -3797 -1256 -3763
rect -1222 -3797 -1216 -3763
rect -1262 -3835 -1216 -3797
rect -1262 -3869 -1256 -3835
rect -1222 -3869 -1216 -3835
rect -1262 -3907 -1216 -3869
rect -1262 -3941 -1256 -3907
rect -1222 -3941 -1216 -3907
rect -1262 -3979 -1216 -3941
rect -1262 -4013 -1256 -3979
rect -1222 -4013 -1216 -3979
rect -1262 -4051 -1216 -4013
rect -1262 -4085 -1256 -4051
rect -1222 -4085 -1216 -4051
rect -1262 -4123 -1216 -4085
rect -1262 -4157 -1256 -4123
rect -1222 -4157 -1216 -4123
rect -1262 -4195 -1216 -4157
rect -1262 -4229 -1256 -4195
rect -1222 -4229 -1216 -4195
rect -1262 -4267 -1216 -4229
rect -1262 -4301 -1256 -4267
rect -1222 -4301 -1216 -4267
rect -1262 -4339 -1216 -4301
rect -1262 -4373 -1256 -4339
rect -1222 -4373 -1216 -4339
rect -1262 -4411 -1216 -4373
rect -1262 -4445 -1256 -4411
rect -1222 -4445 -1216 -4411
rect -1262 -4483 -1216 -4445
rect -1262 -4517 -1256 -4483
rect -1222 -4517 -1216 -4483
rect -1262 -4555 -1216 -4517
rect -1262 -4589 -1256 -4555
rect -1222 -4589 -1216 -4555
rect -1262 -4627 -1216 -4589
rect -1262 -4661 -1256 -4627
rect -1222 -4661 -1216 -4627
rect -1262 -4699 -1216 -4661
rect -1262 -4733 -1256 -4699
rect -1222 -4733 -1216 -4699
rect -1262 -4771 -1216 -4733
rect -1262 -4805 -1256 -4771
rect -1222 -4805 -1216 -4771
rect -1262 -4843 -1216 -4805
rect -1262 -4877 -1256 -4843
rect -1222 -4877 -1216 -4843
rect -1262 -4915 -1216 -4877
rect -1262 -4949 -1256 -4915
rect -1222 -4949 -1216 -4915
rect -1262 -4987 -1216 -4949
rect -1262 -5021 -1256 -4987
rect -1222 -5021 -1216 -4987
rect -1262 -5059 -1216 -5021
rect -1262 -5093 -1256 -5059
rect -1222 -5093 -1216 -5059
rect -1262 -5131 -1216 -5093
rect -1262 -5165 -1256 -5131
rect -1222 -5165 -1216 -5131
rect -1262 -5203 -1216 -5165
rect -1262 -5237 -1256 -5203
rect -1222 -5237 -1216 -5203
rect -1262 -5275 -1216 -5237
rect -1262 -5309 -1256 -5275
rect -1222 -5309 -1216 -5275
rect -1262 -5347 -1216 -5309
rect -1262 -5381 -1256 -5347
rect -1222 -5381 -1216 -5347
rect -1262 -5419 -1216 -5381
rect -1262 -5453 -1256 -5419
rect -1222 -5453 -1216 -5419
rect -1262 -5491 -1216 -5453
rect -1262 -5525 -1256 -5491
rect -1222 -5525 -1216 -5491
rect -1262 -5563 -1216 -5525
rect -1262 -5597 -1256 -5563
rect -1222 -5597 -1216 -5563
rect -1262 -5635 -1216 -5597
rect -1262 -5669 -1256 -5635
rect -1222 -5669 -1216 -5635
rect -1262 -5707 -1216 -5669
rect -1262 -5741 -1256 -5707
rect -1222 -5741 -1216 -5707
rect -1262 -5779 -1216 -5741
rect -1262 -5813 -1256 -5779
rect -1222 -5813 -1216 -5779
rect -1262 -5851 -1216 -5813
rect -1262 -5885 -1256 -5851
rect -1222 -5885 -1216 -5851
rect -1262 -5923 -1216 -5885
rect -1262 -5957 -1256 -5923
rect -1222 -5957 -1216 -5923
rect -1262 -5995 -1216 -5957
rect -1262 -6029 -1256 -5995
rect -1222 -6029 -1216 -5995
rect -1262 -6067 -1216 -6029
rect -1262 -6101 -1256 -6067
rect -1222 -6101 -1216 -6067
rect -1262 -6139 -1216 -6101
rect -1262 -6173 -1256 -6139
rect -1222 -6173 -1216 -6139
rect -1262 -6211 -1216 -6173
rect -1262 -6245 -1256 -6211
rect -1222 -6245 -1216 -6211
rect -1262 -6283 -1216 -6245
rect -1262 -6317 -1256 -6283
rect -1222 -6317 -1216 -6283
rect -1262 -6355 -1216 -6317
rect -1262 -6389 -1256 -6355
rect -1222 -6389 -1216 -6355
rect -1262 -6427 -1216 -6389
rect -1262 -6461 -1256 -6427
rect -1222 -6461 -1216 -6427
rect -1262 -6499 -1216 -6461
rect -1262 -6533 -1256 -6499
rect -1222 -6533 -1216 -6499
rect -1262 -6571 -1216 -6533
rect -1262 -6605 -1256 -6571
rect -1222 -6605 -1216 -6571
rect -1262 -6643 -1216 -6605
rect -1262 -6677 -1256 -6643
rect -1222 -6677 -1216 -6643
rect -1262 -6715 -1216 -6677
rect -1262 -6749 -1256 -6715
rect -1222 -6749 -1216 -6715
rect -1262 -6787 -1216 -6749
rect -1262 -6821 -1256 -6787
rect -1222 -6821 -1216 -6787
rect -1262 -6859 -1216 -6821
rect -1262 -6893 -1256 -6859
rect -1222 -6893 -1216 -6859
rect -1262 -6931 -1216 -6893
rect -1262 -6965 -1256 -6931
rect -1222 -6965 -1216 -6931
rect -1262 -7003 -1216 -6965
rect -1262 -7037 -1256 -7003
rect -1222 -7037 -1216 -7003
rect -1262 -7075 -1216 -7037
rect -1262 -7109 -1256 -7075
rect -1222 -7109 -1216 -7075
rect -1262 -7147 -1216 -7109
rect -1262 -7181 -1256 -7147
rect -1222 -7181 -1216 -7147
rect -1262 -7219 -1216 -7181
rect -1262 -7253 -1256 -7219
rect -1222 -7253 -1216 -7219
rect -1262 -7291 -1216 -7253
rect -1262 -7325 -1256 -7291
rect -1222 -7325 -1216 -7291
rect -1262 -7363 -1216 -7325
rect -1262 -7397 -1256 -7363
rect -1222 -7397 -1216 -7363
rect -1262 -7435 -1216 -7397
rect -1262 -7469 -1256 -7435
rect -1222 -7469 -1216 -7435
rect -1262 -7507 -1216 -7469
rect -1262 -7541 -1256 -7507
rect -1222 -7541 -1216 -7507
rect -1262 -7579 -1216 -7541
rect -1262 -7613 -1256 -7579
rect -1222 -7613 -1216 -7579
rect -1262 -7651 -1216 -7613
rect -1262 -7685 -1256 -7651
rect -1222 -7685 -1216 -7651
rect -1262 -7723 -1216 -7685
rect -1262 -7757 -1256 -7723
rect -1222 -7757 -1216 -7723
rect -1262 -7795 -1216 -7757
rect -1262 -7829 -1256 -7795
rect -1222 -7829 -1216 -7795
rect -1262 -7867 -1216 -7829
rect -1262 -7901 -1256 -7867
rect -1222 -7901 -1216 -7867
rect -1262 -7939 -1216 -7901
rect -1262 -7973 -1256 -7939
rect -1222 -7973 -1216 -7939
rect -1262 -8011 -1216 -7973
rect -1262 -8045 -1256 -8011
rect -1222 -8045 -1216 -8011
rect -1262 -8083 -1216 -8045
rect -1262 -8117 -1256 -8083
rect -1222 -8117 -1216 -8083
rect -1262 -8155 -1216 -8117
rect -1262 -8189 -1256 -8155
rect -1222 -8189 -1216 -8155
rect -1262 -8227 -1216 -8189
rect -1262 -8261 -1256 -8227
rect -1222 -8261 -1216 -8227
rect -1262 -8299 -1216 -8261
rect -1262 -8333 -1256 -8299
rect -1222 -8333 -1216 -8299
rect -1262 -8371 -1216 -8333
rect -1262 -8405 -1256 -8371
rect -1222 -8405 -1216 -8371
rect -1262 -8443 -1216 -8405
rect -1262 -8477 -1256 -8443
rect -1222 -8477 -1216 -8443
rect -1262 -8515 -1216 -8477
rect -1262 -8549 -1256 -8515
rect -1222 -8549 -1216 -8515
rect -1262 -8587 -1216 -8549
rect -1262 -8621 -1256 -8587
rect -1222 -8621 -1216 -8587
rect -1262 -8659 -1216 -8621
rect -1262 -8693 -1256 -8659
rect -1222 -8693 -1216 -8659
rect -1262 -8731 -1216 -8693
rect -1262 -8765 -1256 -8731
rect -1222 -8765 -1216 -8731
rect -1262 -8803 -1216 -8765
rect -1262 -8837 -1256 -8803
rect -1222 -8837 -1216 -8803
rect -1262 -8875 -1216 -8837
rect -1262 -8909 -1256 -8875
rect -1222 -8909 -1216 -8875
rect -1262 -8947 -1216 -8909
rect -1262 -8981 -1256 -8947
rect -1222 -8981 -1216 -8947
rect -1262 -9019 -1216 -8981
rect -1262 -9053 -1256 -9019
rect -1222 -9053 -1216 -9019
rect -1262 -9091 -1216 -9053
rect -1262 -9125 -1256 -9091
rect -1222 -9125 -1216 -9091
rect -1262 -9163 -1216 -9125
rect -1262 -9197 -1256 -9163
rect -1222 -9197 -1216 -9163
rect -1262 -9235 -1216 -9197
rect -1262 -9269 -1256 -9235
rect -1222 -9269 -1216 -9235
rect -1262 -9307 -1216 -9269
rect -1262 -9341 -1256 -9307
rect -1222 -9341 -1216 -9307
rect -1262 -9379 -1216 -9341
rect -1262 -9413 -1256 -9379
rect -1222 -9413 -1216 -9379
rect -1262 -9451 -1216 -9413
rect -1262 -9485 -1256 -9451
rect -1222 -9485 -1216 -9451
rect -1262 -9523 -1216 -9485
rect -1262 -9557 -1256 -9523
rect -1222 -9557 -1216 -9523
rect -1262 -9600 -1216 -9557
rect -1144 9557 -1098 9600
rect -1144 9523 -1138 9557
rect -1104 9523 -1098 9557
rect -1144 9485 -1098 9523
rect -1144 9451 -1138 9485
rect -1104 9451 -1098 9485
rect -1144 9413 -1098 9451
rect -1144 9379 -1138 9413
rect -1104 9379 -1098 9413
rect -1144 9341 -1098 9379
rect -1144 9307 -1138 9341
rect -1104 9307 -1098 9341
rect -1144 9269 -1098 9307
rect -1144 9235 -1138 9269
rect -1104 9235 -1098 9269
rect -1144 9197 -1098 9235
rect -1144 9163 -1138 9197
rect -1104 9163 -1098 9197
rect -1144 9125 -1098 9163
rect -1144 9091 -1138 9125
rect -1104 9091 -1098 9125
rect -1144 9053 -1098 9091
rect -1144 9019 -1138 9053
rect -1104 9019 -1098 9053
rect -1144 8981 -1098 9019
rect -1144 8947 -1138 8981
rect -1104 8947 -1098 8981
rect -1144 8909 -1098 8947
rect -1144 8875 -1138 8909
rect -1104 8875 -1098 8909
rect -1144 8837 -1098 8875
rect -1144 8803 -1138 8837
rect -1104 8803 -1098 8837
rect -1144 8765 -1098 8803
rect -1144 8731 -1138 8765
rect -1104 8731 -1098 8765
rect -1144 8693 -1098 8731
rect -1144 8659 -1138 8693
rect -1104 8659 -1098 8693
rect -1144 8621 -1098 8659
rect -1144 8587 -1138 8621
rect -1104 8587 -1098 8621
rect -1144 8549 -1098 8587
rect -1144 8515 -1138 8549
rect -1104 8515 -1098 8549
rect -1144 8477 -1098 8515
rect -1144 8443 -1138 8477
rect -1104 8443 -1098 8477
rect -1144 8405 -1098 8443
rect -1144 8371 -1138 8405
rect -1104 8371 -1098 8405
rect -1144 8333 -1098 8371
rect -1144 8299 -1138 8333
rect -1104 8299 -1098 8333
rect -1144 8261 -1098 8299
rect -1144 8227 -1138 8261
rect -1104 8227 -1098 8261
rect -1144 8189 -1098 8227
rect -1144 8155 -1138 8189
rect -1104 8155 -1098 8189
rect -1144 8117 -1098 8155
rect -1144 8083 -1138 8117
rect -1104 8083 -1098 8117
rect -1144 8045 -1098 8083
rect -1144 8011 -1138 8045
rect -1104 8011 -1098 8045
rect -1144 7973 -1098 8011
rect -1144 7939 -1138 7973
rect -1104 7939 -1098 7973
rect -1144 7901 -1098 7939
rect -1144 7867 -1138 7901
rect -1104 7867 -1098 7901
rect -1144 7829 -1098 7867
rect -1144 7795 -1138 7829
rect -1104 7795 -1098 7829
rect -1144 7757 -1098 7795
rect -1144 7723 -1138 7757
rect -1104 7723 -1098 7757
rect -1144 7685 -1098 7723
rect -1144 7651 -1138 7685
rect -1104 7651 -1098 7685
rect -1144 7613 -1098 7651
rect -1144 7579 -1138 7613
rect -1104 7579 -1098 7613
rect -1144 7541 -1098 7579
rect -1144 7507 -1138 7541
rect -1104 7507 -1098 7541
rect -1144 7469 -1098 7507
rect -1144 7435 -1138 7469
rect -1104 7435 -1098 7469
rect -1144 7397 -1098 7435
rect -1144 7363 -1138 7397
rect -1104 7363 -1098 7397
rect -1144 7325 -1098 7363
rect -1144 7291 -1138 7325
rect -1104 7291 -1098 7325
rect -1144 7253 -1098 7291
rect -1144 7219 -1138 7253
rect -1104 7219 -1098 7253
rect -1144 7181 -1098 7219
rect -1144 7147 -1138 7181
rect -1104 7147 -1098 7181
rect -1144 7109 -1098 7147
rect -1144 7075 -1138 7109
rect -1104 7075 -1098 7109
rect -1144 7037 -1098 7075
rect -1144 7003 -1138 7037
rect -1104 7003 -1098 7037
rect -1144 6965 -1098 7003
rect -1144 6931 -1138 6965
rect -1104 6931 -1098 6965
rect -1144 6893 -1098 6931
rect -1144 6859 -1138 6893
rect -1104 6859 -1098 6893
rect -1144 6821 -1098 6859
rect -1144 6787 -1138 6821
rect -1104 6787 -1098 6821
rect -1144 6749 -1098 6787
rect -1144 6715 -1138 6749
rect -1104 6715 -1098 6749
rect -1144 6677 -1098 6715
rect -1144 6643 -1138 6677
rect -1104 6643 -1098 6677
rect -1144 6605 -1098 6643
rect -1144 6571 -1138 6605
rect -1104 6571 -1098 6605
rect -1144 6533 -1098 6571
rect -1144 6499 -1138 6533
rect -1104 6499 -1098 6533
rect -1144 6461 -1098 6499
rect -1144 6427 -1138 6461
rect -1104 6427 -1098 6461
rect -1144 6389 -1098 6427
rect -1144 6355 -1138 6389
rect -1104 6355 -1098 6389
rect -1144 6317 -1098 6355
rect -1144 6283 -1138 6317
rect -1104 6283 -1098 6317
rect -1144 6245 -1098 6283
rect -1144 6211 -1138 6245
rect -1104 6211 -1098 6245
rect -1144 6173 -1098 6211
rect -1144 6139 -1138 6173
rect -1104 6139 -1098 6173
rect -1144 6101 -1098 6139
rect -1144 6067 -1138 6101
rect -1104 6067 -1098 6101
rect -1144 6029 -1098 6067
rect -1144 5995 -1138 6029
rect -1104 5995 -1098 6029
rect -1144 5957 -1098 5995
rect -1144 5923 -1138 5957
rect -1104 5923 -1098 5957
rect -1144 5885 -1098 5923
rect -1144 5851 -1138 5885
rect -1104 5851 -1098 5885
rect -1144 5813 -1098 5851
rect -1144 5779 -1138 5813
rect -1104 5779 -1098 5813
rect -1144 5741 -1098 5779
rect -1144 5707 -1138 5741
rect -1104 5707 -1098 5741
rect -1144 5669 -1098 5707
rect -1144 5635 -1138 5669
rect -1104 5635 -1098 5669
rect -1144 5597 -1098 5635
rect -1144 5563 -1138 5597
rect -1104 5563 -1098 5597
rect -1144 5525 -1098 5563
rect -1144 5491 -1138 5525
rect -1104 5491 -1098 5525
rect -1144 5453 -1098 5491
rect -1144 5419 -1138 5453
rect -1104 5419 -1098 5453
rect -1144 5381 -1098 5419
rect -1144 5347 -1138 5381
rect -1104 5347 -1098 5381
rect -1144 5309 -1098 5347
rect -1144 5275 -1138 5309
rect -1104 5275 -1098 5309
rect -1144 5237 -1098 5275
rect -1144 5203 -1138 5237
rect -1104 5203 -1098 5237
rect -1144 5165 -1098 5203
rect -1144 5131 -1138 5165
rect -1104 5131 -1098 5165
rect -1144 5093 -1098 5131
rect -1144 5059 -1138 5093
rect -1104 5059 -1098 5093
rect -1144 5021 -1098 5059
rect -1144 4987 -1138 5021
rect -1104 4987 -1098 5021
rect -1144 4949 -1098 4987
rect -1144 4915 -1138 4949
rect -1104 4915 -1098 4949
rect -1144 4877 -1098 4915
rect -1144 4843 -1138 4877
rect -1104 4843 -1098 4877
rect -1144 4805 -1098 4843
rect -1144 4771 -1138 4805
rect -1104 4771 -1098 4805
rect -1144 4733 -1098 4771
rect -1144 4699 -1138 4733
rect -1104 4699 -1098 4733
rect -1144 4661 -1098 4699
rect -1144 4627 -1138 4661
rect -1104 4627 -1098 4661
rect -1144 4589 -1098 4627
rect -1144 4555 -1138 4589
rect -1104 4555 -1098 4589
rect -1144 4517 -1098 4555
rect -1144 4483 -1138 4517
rect -1104 4483 -1098 4517
rect -1144 4445 -1098 4483
rect -1144 4411 -1138 4445
rect -1104 4411 -1098 4445
rect -1144 4373 -1098 4411
rect -1144 4339 -1138 4373
rect -1104 4339 -1098 4373
rect -1144 4301 -1098 4339
rect -1144 4267 -1138 4301
rect -1104 4267 -1098 4301
rect -1144 4229 -1098 4267
rect -1144 4195 -1138 4229
rect -1104 4195 -1098 4229
rect -1144 4157 -1098 4195
rect -1144 4123 -1138 4157
rect -1104 4123 -1098 4157
rect -1144 4085 -1098 4123
rect -1144 4051 -1138 4085
rect -1104 4051 -1098 4085
rect -1144 4013 -1098 4051
rect -1144 3979 -1138 4013
rect -1104 3979 -1098 4013
rect -1144 3941 -1098 3979
rect -1144 3907 -1138 3941
rect -1104 3907 -1098 3941
rect -1144 3869 -1098 3907
rect -1144 3835 -1138 3869
rect -1104 3835 -1098 3869
rect -1144 3797 -1098 3835
rect -1144 3763 -1138 3797
rect -1104 3763 -1098 3797
rect -1144 3725 -1098 3763
rect -1144 3691 -1138 3725
rect -1104 3691 -1098 3725
rect -1144 3653 -1098 3691
rect -1144 3619 -1138 3653
rect -1104 3619 -1098 3653
rect -1144 3581 -1098 3619
rect -1144 3547 -1138 3581
rect -1104 3547 -1098 3581
rect -1144 3509 -1098 3547
rect -1144 3475 -1138 3509
rect -1104 3475 -1098 3509
rect -1144 3437 -1098 3475
rect -1144 3403 -1138 3437
rect -1104 3403 -1098 3437
rect -1144 3365 -1098 3403
rect -1144 3331 -1138 3365
rect -1104 3331 -1098 3365
rect -1144 3293 -1098 3331
rect -1144 3259 -1138 3293
rect -1104 3259 -1098 3293
rect -1144 3221 -1098 3259
rect -1144 3187 -1138 3221
rect -1104 3187 -1098 3221
rect -1144 3149 -1098 3187
rect -1144 3115 -1138 3149
rect -1104 3115 -1098 3149
rect -1144 3077 -1098 3115
rect -1144 3043 -1138 3077
rect -1104 3043 -1098 3077
rect -1144 3005 -1098 3043
rect -1144 2971 -1138 3005
rect -1104 2971 -1098 3005
rect -1144 2933 -1098 2971
rect -1144 2899 -1138 2933
rect -1104 2899 -1098 2933
rect -1144 2861 -1098 2899
rect -1144 2827 -1138 2861
rect -1104 2827 -1098 2861
rect -1144 2789 -1098 2827
rect -1144 2755 -1138 2789
rect -1104 2755 -1098 2789
rect -1144 2717 -1098 2755
rect -1144 2683 -1138 2717
rect -1104 2683 -1098 2717
rect -1144 2645 -1098 2683
rect -1144 2611 -1138 2645
rect -1104 2611 -1098 2645
rect -1144 2573 -1098 2611
rect -1144 2539 -1138 2573
rect -1104 2539 -1098 2573
rect -1144 2501 -1098 2539
rect -1144 2467 -1138 2501
rect -1104 2467 -1098 2501
rect -1144 2429 -1098 2467
rect -1144 2395 -1138 2429
rect -1104 2395 -1098 2429
rect -1144 2357 -1098 2395
rect -1144 2323 -1138 2357
rect -1104 2323 -1098 2357
rect -1144 2285 -1098 2323
rect -1144 2251 -1138 2285
rect -1104 2251 -1098 2285
rect -1144 2213 -1098 2251
rect -1144 2179 -1138 2213
rect -1104 2179 -1098 2213
rect -1144 2141 -1098 2179
rect -1144 2107 -1138 2141
rect -1104 2107 -1098 2141
rect -1144 2069 -1098 2107
rect -1144 2035 -1138 2069
rect -1104 2035 -1098 2069
rect -1144 1997 -1098 2035
rect -1144 1963 -1138 1997
rect -1104 1963 -1098 1997
rect -1144 1925 -1098 1963
rect -1144 1891 -1138 1925
rect -1104 1891 -1098 1925
rect -1144 1853 -1098 1891
rect -1144 1819 -1138 1853
rect -1104 1819 -1098 1853
rect -1144 1781 -1098 1819
rect -1144 1747 -1138 1781
rect -1104 1747 -1098 1781
rect -1144 1709 -1098 1747
rect -1144 1675 -1138 1709
rect -1104 1675 -1098 1709
rect -1144 1637 -1098 1675
rect -1144 1603 -1138 1637
rect -1104 1603 -1098 1637
rect -1144 1565 -1098 1603
rect -1144 1531 -1138 1565
rect -1104 1531 -1098 1565
rect -1144 1493 -1098 1531
rect -1144 1459 -1138 1493
rect -1104 1459 -1098 1493
rect -1144 1421 -1098 1459
rect -1144 1387 -1138 1421
rect -1104 1387 -1098 1421
rect -1144 1349 -1098 1387
rect -1144 1315 -1138 1349
rect -1104 1315 -1098 1349
rect -1144 1277 -1098 1315
rect -1144 1243 -1138 1277
rect -1104 1243 -1098 1277
rect -1144 1205 -1098 1243
rect -1144 1171 -1138 1205
rect -1104 1171 -1098 1205
rect -1144 1133 -1098 1171
rect -1144 1099 -1138 1133
rect -1104 1099 -1098 1133
rect -1144 1061 -1098 1099
rect -1144 1027 -1138 1061
rect -1104 1027 -1098 1061
rect -1144 989 -1098 1027
rect -1144 955 -1138 989
rect -1104 955 -1098 989
rect -1144 917 -1098 955
rect -1144 883 -1138 917
rect -1104 883 -1098 917
rect -1144 845 -1098 883
rect -1144 811 -1138 845
rect -1104 811 -1098 845
rect -1144 773 -1098 811
rect -1144 739 -1138 773
rect -1104 739 -1098 773
rect -1144 701 -1098 739
rect -1144 667 -1138 701
rect -1104 667 -1098 701
rect -1144 629 -1098 667
rect -1144 595 -1138 629
rect -1104 595 -1098 629
rect -1144 557 -1098 595
rect -1144 523 -1138 557
rect -1104 523 -1098 557
rect -1144 485 -1098 523
rect -1144 451 -1138 485
rect -1104 451 -1098 485
rect -1144 413 -1098 451
rect -1144 379 -1138 413
rect -1104 379 -1098 413
rect -1144 341 -1098 379
rect -1144 307 -1138 341
rect -1104 307 -1098 341
rect -1144 269 -1098 307
rect -1144 235 -1138 269
rect -1104 235 -1098 269
rect -1144 197 -1098 235
rect -1144 163 -1138 197
rect -1104 163 -1098 197
rect -1144 125 -1098 163
rect -1144 91 -1138 125
rect -1104 91 -1098 125
rect -1144 53 -1098 91
rect -1144 19 -1138 53
rect -1104 19 -1098 53
rect -1144 -19 -1098 19
rect -1144 -53 -1138 -19
rect -1104 -53 -1098 -19
rect -1144 -91 -1098 -53
rect -1144 -125 -1138 -91
rect -1104 -125 -1098 -91
rect -1144 -163 -1098 -125
rect -1144 -197 -1138 -163
rect -1104 -197 -1098 -163
rect -1144 -235 -1098 -197
rect -1144 -269 -1138 -235
rect -1104 -269 -1098 -235
rect -1144 -307 -1098 -269
rect -1144 -341 -1138 -307
rect -1104 -341 -1098 -307
rect -1144 -379 -1098 -341
rect -1144 -413 -1138 -379
rect -1104 -413 -1098 -379
rect -1144 -451 -1098 -413
rect -1144 -485 -1138 -451
rect -1104 -485 -1098 -451
rect -1144 -523 -1098 -485
rect -1144 -557 -1138 -523
rect -1104 -557 -1098 -523
rect -1144 -595 -1098 -557
rect -1144 -629 -1138 -595
rect -1104 -629 -1098 -595
rect -1144 -667 -1098 -629
rect -1144 -701 -1138 -667
rect -1104 -701 -1098 -667
rect -1144 -739 -1098 -701
rect -1144 -773 -1138 -739
rect -1104 -773 -1098 -739
rect -1144 -811 -1098 -773
rect -1144 -845 -1138 -811
rect -1104 -845 -1098 -811
rect -1144 -883 -1098 -845
rect -1144 -917 -1138 -883
rect -1104 -917 -1098 -883
rect -1144 -955 -1098 -917
rect -1144 -989 -1138 -955
rect -1104 -989 -1098 -955
rect -1144 -1027 -1098 -989
rect -1144 -1061 -1138 -1027
rect -1104 -1061 -1098 -1027
rect -1144 -1099 -1098 -1061
rect -1144 -1133 -1138 -1099
rect -1104 -1133 -1098 -1099
rect -1144 -1171 -1098 -1133
rect -1144 -1205 -1138 -1171
rect -1104 -1205 -1098 -1171
rect -1144 -1243 -1098 -1205
rect -1144 -1277 -1138 -1243
rect -1104 -1277 -1098 -1243
rect -1144 -1315 -1098 -1277
rect -1144 -1349 -1138 -1315
rect -1104 -1349 -1098 -1315
rect -1144 -1387 -1098 -1349
rect -1144 -1421 -1138 -1387
rect -1104 -1421 -1098 -1387
rect -1144 -1459 -1098 -1421
rect -1144 -1493 -1138 -1459
rect -1104 -1493 -1098 -1459
rect -1144 -1531 -1098 -1493
rect -1144 -1565 -1138 -1531
rect -1104 -1565 -1098 -1531
rect -1144 -1603 -1098 -1565
rect -1144 -1637 -1138 -1603
rect -1104 -1637 -1098 -1603
rect -1144 -1675 -1098 -1637
rect -1144 -1709 -1138 -1675
rect -1104 -1709 -1098 -1675
rect -1144 -1747 -1098 -1709
rect -1144 -1781 -1138 -1747
rect -1104 -1781 -1098 -1747
rect -1144 -1819 -1098 -1781
rect -1144 -1853 -1138 -1819
rect -1104 -1853 -1098 -1819
rect -1144 -1891 -1098 -1853
rect -1144 -1925 -1138 -1891
rect -1104 -1925 -1098 -1891
rect -1144 -1963 -1098 -1925
rect -1144 -1997 -1138 -1963
rect -1104 -1997 -1098 -1963
rect -1144 -2035 -1098 -1997
rect -1144 -2069 -1138 -2035
rect -1104 -2069 -1098 -2035
rect -1144 -2107 -1098 -2069
rect -1144 -2141 -1138 -2107
rect -1104 -2141 -1098 -2107
rect -1144 -2179 -1098 -2141
rect -1144 -2213 -1138 -2179
rect -1104 -2213 -1098 -2179
rect -1144 -2251 -1098 -2213
rect -1144 -2285 -1138 -2251
rect -1104 -2285 -1098 -2251
rect -1144 -2323 -1098 -2285
rect -1144 -2357 -1138 -2323
rect -1104 -2357 -1098 -2323
rect -1144 -2395 -1098 -2357
rect -1144 -2429 -1138 -2395
rect -1104 -2429 -1098 -2395
rect -1144 -2467 -1098 -2429
rect -1144 -2501 -1138 -2467
rect -1104 -2501 -1098 -2467
rect -1144 -2539 -1098 -2501
rect -1144 -2573 -1138 -2539
rect -1104 -2573 -1098 -2539
rect -1144 -2611 -1098 -2573
rect -1144 -2645 -1138 -2611
rect -1104 -2645 -1098 -2611
rect -1144 -2683 -1098 -2645
rect -1144 -2717 -1138 -2683
rect -1104 -2717 -1098 -2683
rect -1144 -2755 -1098 -2717
rect -1144 -2789 -1138 -2755
rect -1104 -2789 -1098 -2755
rect -1144 -2827 -1098 -2789
rect -1144 -2861 -1138 -2827
rect -1104 -2861 -1098 -2827
rect -1144 -2899 -1098 -2861
rect -1144 -2933 -1138 -2899
rect -1104 -2933 -1098 -2899
rect -1144 -2971 -1098 -2933
rect -1144 -3005 -1138 -2971
rect -1104 -3005 -1098 -2971
rect -1144 -3043 -1098 -3005
rect -1144 -3077 -1138 -3043
rect -1104 -3077 -1098 -3043
rect -1144 -3115 -1098 -3077
rect -1144 -3149 -1138 -3115
rect -1104 -3149 -1098 -3115
rect -1144 -3187 -1098 -3149
rect -1144 -3221 -1138 -3187
rect -1104 -3221 -1098 -3187
rect -1144 -3259 -1098 -3221
rect -1144 -3293 -1138 -3259
rect -1104 -3293 -1098 -3259
rect -1144 -3331 -1098 -3293
rect -1144 -3365 -1138 -3331
rect -1104 -3365 -1098 -3331
rect -1144 -3403 -1098 -3365
rect -1144 -3437 -1138 -3403
rect -1104 -3437 -1098 -3403
rect -1144 -3475 -1098 -3437
rect -1144 -3509 -1138 -3475
rect -1104 -3509 -1098 -3475
rect -1144 -3547 -1098 -3509
rect -1144 -3581 -1138 -3547
rect -1104 -3581 -1098 -3547
rect -1144 -3619 -1098 -3581
rect -1144 -3653 -1138 -3619
rect -1104 -3653 -1098 -3619
rect -1144 -3691 -1098 -3653
rect -1144 -3725 -1138 -3691
rect -1104 -3725 -1098 -3691
rect -1144 -3763 -1098 -3725
rect -1144 -3797 -1138 -3763
rect -1104 -3797 -1098 -3763
rect -1144 -3835 -1098 -3797
rect -1144 -3869 -1138 -3835
rect -1104 -3869 -1098 -3835
rect -1144 -3907 -1098 -3869
rect -1144 -3941 -1138 -3907
rect -1104 -3941 -1098 -3907
rect -1144 -3979 -1098 -3941
rect -1144 -4013 -1138 -3979
rect -1104 -4013 -1098 -3979
rect -1144 -4051 -1098 -4013
rect -1144 -4085 -1138 -4051
rect -1104 -4085 -1098 -4051
rect -1144 -4123 -1098 -4085
rect -1144 -4157 -1138 -4123
rect -1104 -4157 -1098 -4123
rect -1144 -4195 -1098 -4157
rect -1144 -4229 -1138 -4195
rect -1104 -4229 -1098 -4195
rect -1144 -4267 -1098 -4229
rect -1144 -4301 -1138 -4267
rect -1104 -4301 -1098 -4267
rect -1144 -4339 -1098 -4301
rect -1144 -4373 -1138 -4339
rect -1104 -4373 -1098 -4339
rect -1144 -4411 -1098 -4373
rect -1144 -4445 -1138 -4411
rect -1104 -4445 -1098 -4411
rect -1144 -4483 -1098 -4445
rect -1144 -4517 -1138 -4483
rect -1104 -4517 -1098 -4483
rect -1144 -4555 -1098 -4517
rect -1144 -4589 -1138 -4555
rect -1104 -4589 -1098 -4555
rect -1144 -4627 -1098 -4589
rect -1144 -4661 -1138 -4627
rect -1104 -4661 -1098 -4627
rect -1144 -4699 -1098 -4661
rect -1144 -4733 -1138 -4699
rect -1104 -4733 -1098 -4699
rect -1144 -4771 -1098 -4733
rect -1144 -4805 -1138 -4771
rect -1104 -4805 -1098 -4771
rect -1144 -4843 -1098 -4805
rect -1144 -4877 -1138 -4843
rect -1104 -4877 -1098 -4843
rect -1144 -4915 -1098 -4877
rect -1144 -4949 -1138 -4915
rect -1104 -4949 -1098 -4915
rect -1144 -4987 -1098 -4949
rect -1144 -5021 -1138 -4987
rect -1104 -5021 -1098 -4987
rect -1144 -5059 -1098 -5021
rect -1144 -5093 -1138 -5059
rect -1104 -5093 -1098 -5059
rect -1144 -5131 -1098 -5093
rect -1144 -5165 -1138 -5131
rect -1104 -5165 -1098 -5131
rect -1144 -5203 -1098 -5165
rect -1144 -5237 -1138 -5203
rect -1104 -5237 -1098 -5203
rect -1144 -5275 -1098 -5237
rect -1144 -5309 -1138 -5275
rect -1104 -5309 -1098 -5275
rect -1144 -5347 -1098 -5309
rect -1144 -5381 -1138 -5347
rect -1104 -5381 -1098 -5347
rect -1144 -5419 -1098 -5381
rect -1144 -5453 -1138 -5419
rect -1104 -5453 -1098 -5419
rect -1144 -5491 -1098 -5453
rect -1144 -5525 -1138 -5491
rect -1104 -5525 -1098 -5491
rect -1144 -5563 -1098 -5525
rect -1144 -5597 -1138 -5563
rect -1104 -5597 -1098 -5563
rect -1144 -5635 -1098 -5597
rect -1144 -5669 -1138 -5635
rect -1104 -5669 -1098 -5635
rect -1144 -5707 -1098 -5669
rect -1144 -5741 -1138 -5707
rect -1104 -5741 -1098 -5707
rect -1144 -5779 -1098 -5741
rect -1144 -5813 -1138 -5779
rect -1104 -5813 -1098 -5779
rect -1144 -5851 -1098 -5813
rect -1144 -5885 -1138 -5851
rect -1104 -5885 -1098 -5851
rect -1144 -5923 -1098 -5885
rect -1144 -5957 -1138 -5923
rect -1104 -5957 -1098 -5923
rect -1144 -5995 -1098 -5957
rect -1144 -6029 -1138 -5995
rect -1104 -6029 -1098 -5995
rect -1144 -6067 -1098 -6029
rect -1144 -6101 -1138 -6067
rect -1104 -6101 -1098 -6067
rect -1144 -6139 -1098 -6101
rect -1144 -6173 -1138 -6139
rect -1104 -6173 -1098 -6139
rect -1144 -6211 -1098 -6173
rect -1144 -6245 -1138 -6211
rect -1104 -6245 -1098 -6211
rect -1144 -6283 -1098 -6245
rect -1144 -6317 -1138 -6283
rect -1104 -6317 -1098 -6283
rect -1144 -6355 -1098 -6317
rect -1144 -6389 -1138 -6355
rect -1104 -6389 -1098 -6355
rect -1144 -6427 -1098 -6389
rect -1144 -6461 -1138 -6427
rect -1104 -6461 -1098 -6427
rect -1144 -6499 -1098 -6461
rect -1144 -6533 -1138 -6499
rect -1104 -6533 -1098 -6499
rect -1144 -6571 -1098 -6533
rect -1144 -6605 -1138 -6571
rect -1104 -6605 -1098 -6571
rect -1144 -6643 -1098 -6605
rect -1144 -6677 -1138 -6643
rect -1104 -6677 -1098 -6643
rect -1144 -6715 -1098 -6677
rect -1144 -6749 -1138 -6715
rect -1104 -6749 -1098 -6715
rect -1144 -6787 -1098 -6749
rect -1144 -6821 -1138 -6787
rect -1104 -6821 -1098 -6787
rect -1144 -6859 -1098 -6821
rect -1144 -6893 -1138 -6859
rect -1104 -6893 -1098 -6859
rect -1144 -6931 -1098 -6893
rect -1144 -6965 -1138 -6931
rect -1104 -6965 -1098 -6931
rect -1144 -7003 -1098 -6965
rect -1144 -7037 -1138 -7003
rect -1104 -7037 -1098 -7003
rect -1144 -7075 -1098 -7037
rect -1144 -7109 -1138 -7075
rect -1104 -7109 -1098 -7075
rect -1144 -7147 -1098 -7109
rect -1144 -7181 -1138 -7147
rect -1104 -7181 -1098 -7147
rect -1144 -7219 -1098 -7181
rect -1144 -7253 -1138 -7219
rect -1104 -7253 -1098 -7219
rect -1144 -7291 -1098 -7253
rect -1144 -7325 -1138 -7291
rect -1104 -7325 -1098 -7291
rect -1144 -7363 -1098 -7325
rect -1144 -7397 -1138 -7363
rect -1104 -7397 -1098 -7363
rect -1144 -7435 -1098 -7397
rect -1144 -7469 -1138 -7435
rect -1104 -7469 -1098 -7435
rect -1144 -7507 -1098 -7469
rect -1144 -7541 -1138 -7507
rect -1104 -7541 -1098 -7507
rect -1144 -7579 -1098 -7541
rect -1144 -7613 -1138 -7579
rect -1104 -7613 -1098 -7579
rect -1144 -7651 -1098 -7613
rect -1144 -7685 -1138 -7651
rect -1104 -7685 -1098 -7651
rect -1144 -7723 -1098 -7685
rect -1144 -7757 -1138 -7723
rect -1104 -7757 -1098 -7723
rect -1144 -7795 -1098 -7757
rect -1144 -7829 -1138 -7795
rect -1104 -7829 -1098 -7795
rect -1144 -7867 -1098 -7829
rect -1144 -7901 -1138 -7867
rect -1104 -7901 -1098 -7867
rect -1144 -7939 -1098 -7901
rect -1144 -7973 -1138 -7939
rect -1104 -7973 -1098 -7939
rect -1144 -8011 -1098 -7973
rect -1144 -8045 -1138 -8011
rect -1104 -8045 -1098 -8011
rect -1144 -8083 -1098 -8045
rect -1144 -8117 -1138 -8083
rect -1104 -8117 -1098 -8083
rect -1144 -8155 -1098 -8117
rect -1144 -8189 -1138 -8155
rect -1104 -8189 -1098 -8155
rect -1144 -8227 -1098 -8189
rect -1144 -8261 -1138 -8227
rect -1104 -8261 -1098 -8227
rect -1144 -8299 -1098 -8261
rect -1144 -8333 -1138 -8299
rect -1104 -8333 -1098 -8299
rect -1144 -8371 -1098 -8333
rect -1144 -8405 -1138 -8371
rect -1104 -8405 -1098 -8371
rect -1144 -8443 -1098 -8405
rect -1144 -8477 -1138 -8443
rect -1104 -8477 -1098 -8443
rect -1144 -8515 -1098 -8477
rect -1144 -8549 -1138 -8515
rect -1104 -8549 -1098 -8515
rect -1144 -8587 -1098 -8549
rect -1144 -8621 -1138 -8587
rect -1104 -8621 -1098 -8587
rect -1144 -8659 -1098 -8621
rect -1144 -8693 -1138 -8659
rect -1104 -8693 -1098 -8659
rect -1144 -8731 -1098 -8693
rect -1144 -8765 -1138 -8731
rect -1104 -8765 -1098 -8731
rect -1144 -8803 -1098 -8765
rect -1144 -8837 -1138 -8803
rect -1104 -8837 -1098 -8803
rect -1144 -8875 -1098 -8837
rect -1144 -8909 -1138 -8875
rect -1104 -8909 -1098 -8875
rect -1144 -8947 -1098 -8909
rect -1144 -8981 -1138 -8947
rect -1104 -8981 -1098 -8947
rect -1144 -9019 -1098 -8981
rect -1144 -9053 -1138 -9019
rect -1104 -9053 -1098 -9019
rect -1144 -9091 -1098 -9053
rect -1144 -9125 -1138 -9091
rect -1104 -9125 -1098 -9091
rect -1144 -9163 -1098 -9125
rect -1144 -9197 -1138 -9163
rect -1104 -9197 -1098 -9163
rect -1144 -9235 -1098 -9197
rect -1144 -9269 -1138 -9235
rect -1104 -9269 -1098 -9235
rect -1144 -9307 -1098 -9269
rect -1144 -9341 -1138 -9307
rect -1104 -9341 -1098 -9307
rect -1144 -9379 -1098 -9341
rect -1144 -9413 -1138 -9379
rect -1104 -9413 -1098 -9379
rect -1144 -9451 -1098 -9413
rect -1144 -9485 -1138 -9451
rect -1104 -9485 -1098 -9451
rect -1144 -9523 -1098 -9485
rect -1144 -9557 -1138 -9523
rect -1104 -9557 -1098 -9523
rect -1144 -9600 -1098 -9557
rect -1026 9557 -980 9600
rect -1026 9523 -1020 9557
rect -986 9523 -980 9557
rect -1026 9485 -980 9523
rect -1026 9451 -1020 9485
rect -986 9451 -980 9485
rect -1026 9413 -980 9451
rect -1026 9379 -1020 9413
rect -986 9379 -980 9413
rect -1026 9341 -980 9379
rect -1026 9307 -1020 9341
rect -986 9307 -980 9341
rect -1026 9269 -980 9307
rect -1026 9235 -1020 9269
rect -986 9235 -980 9269
rect -1026 9197 -980 9235
rect -1026 9163 -1020 9197
rect -986 9163 -980 9197
rect -1026 9125 -980 9163
rect -1026 9091 -1020 9125
rect -986 9091 -980 9125
rect -1026 9053 -980 9091
rect -1026 9019 -1020 9053
rect -986 9019 -980 9053
rect -1026 8981 -980 9019
rect -1026 8947 -1020 8981
rect -986 8947 -980 8981
rect -1026 8909 -980 8947
rect -1026 8875 -1020 8909
rect -986 8875 -980 8909
rect -1026 8837 -980 8875
rect -1026 8803 -1020 8837
rect -986 8803 -980 8837
rect -1026 8765 -980 8803
rect -1026 8731 -1020 8765
rect -986 8731 -980 8765
rect -1026 8693 -980 8731
rect -1026 8659 -1020 8693
rect -986 8659 -980 8693
rect -1026 8621 -980 8659
rect -1026 8587 -1020 8621
rect -986 8587 -980 8621
rect -1026 8549 -980 8587
rect -1026 8515 -1020 8549
rect -986 8515 -980 8549
rect -1026 8477 -980 8515
rect -1026 8443 -1020 8477
rect -986 8443 -980 8477
rect -1026 8405 -980 8443
rect -1026 8371 -1020 8405
rect -986 8371 -980 8405
rect -1026 8333 -980 8371
rect -1026 8299 -1020 8333
rect -986 8299 -980 8333
rect -1026 8261 -980 8299
rect -1026 8227 -1020 8261
rect -986 8227 -980 8261
rect -1026 8189 -980 8227
rect -1026 8155 -1020 8189
rect -986 8155 -980 8189
rect -1026 8117 -980 8155
rect -1026 8083 -1020 8117
rect -986 8083 -980 8117
rect -1026 8045 -980 8083
rect -1026 8011 -1020 8045
rect -986 8011 -980 8045
rect -1026 7973 -980 8011
rect -1026 7939 -1020 7973
rect -986 7939 -980 7973
rect -1026 7901 -980 7939
rect -1026 7867 -1020 7901
rect -986 7867 -980 7901
rect -1026 7829 -980 7867
rect -1026 7795 -1020 7829
rect -986 7795 -980 7829
rect -1026 7757 -980 7795
rect -1026 7723 -1020 7757
rect -986 7723 -980 7757
rect -1026 7685 -980 7723
rect -1026 7651 -1020 7685
rect -986 7651 -980 7685
rect -1026 7613 -980 7651
rect -1026 7579 -1020 7613
rect -986 7579 -980 7613
rect -1026 7541 -980 7579
rect -1026 7507 -1020 7541
rect -986 7507 -980 7541
rect -1026 7469 -980 7507
rect -1026 7435 -1020 7469
rect -986 7435 -980 7469
rect -1026 7397 -980 7435
rect -1026 7363 -1020 7397
rect -986 7363 -980 7397
rect -1026 7325 -980 7363
rect -1026 7291 -1020 7325
rect -986 7291 -980 7325
rect -1026 7253 -980 7291
rect -1026 7219 -1020 7253
rect -986 7219 -980 7253
rect -1026 7181 -980 7219
rect -1026 7147 -1020 7181
rect -986 7147 -980 7181
rect -1026 7109 -980 7147
rect -1026 7075 -1020 7109
rect -986 7075 -980 7109
rect -1026 7037 -980 7075
rect -1026 7003 -1020 7037
rect -986 7003 -980 7037
rect -1026 6965 -980 7003
rect -1026 6931 -1020 6965
rect -986 6931 -980 6965
rect -1026 6893 -980 6931
rect -1026 6859 -1020 6893
rect -986 6859 -980 6893
rect -1026 6821 -980 6859
rect -1026 6787 -1020 6821
rect -986 6787 -980 6821
rect -1026 6749 -980 6787
rect -1026 6715 -1020 6749
rect -986 6715 -980 6749
rect -1026 6677 -980 6715
rect -1026 6643 -1020 6677
rect -986 6643 -980 6677
rect -1026 6605 -980 6643
rect -1026 6571 -1020 6605
rect -986 6571 -980 6605
rect -1026 6533 -980 6571
rect -1026 6499 -1020 6533
rect -986 6499 -980 6533
rect -1026 6461 -980 6499
rect -1026 6427 -1020 6461
rect -986 6427 -980 6461
rect -1026 6389 -980 6427
rect -1026 6355 -1020 6389
rect -986 6355 -980 6389
rect -1026 6317 -980 6355
rect -1026 6283 -1020 6317
rect -986 6283 -980 6317
rect -1026 6245 -980 6283
rect -1026 6211 -1020 6245
rect -986 6211 -980 6245
rect -1026 6173 -980 6211
rect -1026 6139 -1020 6173
rect -986 6139 -980 6173
rect -1026 6101 -980 6139
rect -1026 6067 -1020 6101
rect -986 6067 -980 6101
rect -1026 6029 -980 6067
rect -1026 5995 -1020 6029
rect -986 5995 -980 6029
rect -1026 5957 -980 5995
rect -1026 5923 -1020 5957
rect -986 5923 -980 5957
rect -1026 5885 -980 5923
rect -1026 5851 -1020 5885
rect -986 5851 -980 5885
rect -1026 5813 -980 5851
rect -1026 5779 -1020 5813
rect -986 5779 -980 5813
rect -1026 5741 -980 5779
rect -1026 5707 -1020 5741
rect -986 5707 -980 5741
rect -1026 5669 -980 5707
rect -1026 5635 -1020 5669
rect -986 5635 -980 5669
rect -1026 5597 -980 5635
rect -1026 5563 -1020 5597
rect -986 5563 -980 5597
rect -1026 5525 -980 5563
rect -1026 5491 -1020 5525
rect -986 5491 -980 5525
rect -1026 5453 -980 5491
rect -1026 5419 -1020 5453
rect -986 5419 -980 5453
rect -1026 5381 -980 5419
rect -1026 5347 -1020 5381
rect -986 5347 -980 5381
rect -1026 5309 -980 5347
rect -1026 5275 -1020 5309
rect -986 5275 -980 5309
rect -1026 5237 -980 5275
rect -1026 5203 -1020 5237
rect -986 5203 -980 5237
rect -1026 5165 -980 5203
rect -1026 5131 -1020 5165
rect -986 5131 -980 5165
rect -1026 5093 -980 5131
rect -1026 5059 -1020 5093
rect -986 5059 -980 5093
rect -1026 5021 -980 5059
rect -1026 4987 -1020 5021
rect -986 4987 -980 5021
rect -1026 4949 -980 4987
rect -1026 4915 -1020 4949
rect -986 4915 -980 4949
rect -1026 4877 -980 4915
rect -1026 4843 -1020 4877
rect -986 4843 -980 4877
rect -1026 4805 -980 4843
rect -1026 4771 -1020 4805
rect -986 4771 -980 4805
rect -1026 4733 -980 4771
rect -1026 4699 -1020 4733
rect -986 4699 -980 4733
rect -1026 4661 -980 4699
rect -1026 4627 -1020 4661
rect -986 4627 -980 4661
rect -1026 4589 -980 4627
rect -1026 4555 -1020 4589
rect -986 4555 -980 4589
rect -1026 4517 -980 4555
rect -1026 4483 -1020 4517
rect -986 4483 -980 4517
rect -1026 4445 -980 4483
rect -1026 4411 -1020 4445
rect -986 4411 -980 4445
rect -1026 4373 -980 4411
rect -1026 4339 -1020 4373
rect -986 4339 -980 4373
rect -1026 4301 -980 4339
rect -1026 4267 -1020 4301
rect -986 4267 -980 4301
rect -1026 4229 -980 4267
rect -1026 4195 -1020 4229
rect -986 4195 -980 4229
rect -1026 4157 -980 4195
rect -1026 4123 -1020 4157
rect -986 4123 -980 4157
rect -1026 4085 -980 4123
rect -1026 4051 -1020 4085
rect -986 4051 -980 4085
rect -1026 4013 -980 4051
rect -1026 3979 -1020 4013
rect -986 3979 -980 4013
rect -1026 3941 -980 3979
rect -1026 3907 -1020 3941
rect -986 3907 -980 3941
rect -1026 3869 -980 3907
rect -1026 3835 -1020 3869
rect -986 3835 -980 3869
rect -1026 3797 -980 3835
rect -1026 3763 -1020 3797
rect -986 3763 -980 3797
rect -1026 3725 -980 3763
rect -1026 3691 -1020 3725
rect -986 3691 -980 3725
rect -1026 3653 -980 3691
rect -1026 3619 -1020 3653
rect -986 3619 -980 3653
rect -1026 3581 -980 3619
rect -1026 3547 -1020 3581
rect -986 3547 -980 3581
rect -1026 3509 -980 3547
rect -1026 3475 -1020 3509
rect -986 3475 -980 3509
rect -1026 3437 -980 3475
rect -1026 3403 -1020 3437
rect -986 3403 -980 3437
rect -1026 3365 -980 3403
rect -1026 3331 -1020 3365
rect -986 3331 -980 3365
rect -1026 3293 -980 3331
rect -1026 3259 -1020 3293
rect -986 3259 -980 3293
rect -1026 3221 -980 3259
rect -1026 3187 -1020 3221
rect -986 3187 -980 3221
rect -1026 3149 -980 3187
rect -1026 3115 -1020 3149
rect -986 3115 -980 3149
rect -1026 3077 -980 3115
rect -1026 3043 -1020 3077
rect -986 3043 -980 3077
rect -1026 3005 -980 3043
rect -1026 2971 -1020 3005
rect -986 2971 -980 3005
rect -1026 2933 -980 2971
rect -1026 2899 -1020 2933
rect -986 2899 -980 2933
rect -1026 2861 -980 2899
rect -1026 2827 -1020 2861
rect -986 2827 -980 2861
rect -1026 2789 -980 2827
rect -1026 2755 -1020 2789
rect -986 2755 -980 2789
rect -1026 2717 -980 2755
rect -1026 2683 -1020 2717
rect -986 2683 -980 2717
rect -1026 2645 -980 2683
rect -1026 2611 -1020 2645
rect -986 2611 -980 2645
rect -1026 2573 -980 2611
rect -1026 2539 -1020 2573
rect -986 2539 -980 2573
rect -1026 2501 -980 2539
rect -1026 2467 -1020 2501
rect -986 2467 -980 2501
rect -1026 2429 -980 2467
rect -1026 2395 -1020 2429
rect -986 2395 -980 2429
rect -1026 2357 -980 2395
rect -1026 2323 -1020 2357
rect -986 2323 -980 2357
rect -1026 2285 -980 2323
rect -1026 2251 -1020 2285
rect -986 2251 -980 2285
rect -1026 2213 -980 2251
rect -1026 2179 -1020 2213
rect -986 2179 -980 2213
rect -1026 2141 -980 2179
rect -1026 2107 -1020 2141
rect -986 2107 -980 2141
rect -1026 2069 -980 2107
rect -1026 2035 -1020 2069
rect -986 2035 -980 2069
rect -1026 1997 -980 2035
rect -1026 1963 -1020 1997
rect -986 1963 -980 1997
rect -1026 1925 -980 1963
rect -1026 1891 -1020 1925
rect -986 1891 -980 1925
rect -1026 1853 -980 1891
rect -1026 1819 -1020 1853
rect -986 1819 -980 1853
rect -1026 1781 -980 1819
rect -1026 1747 -1020 1781
rect -986 1747 -980 1781
rect -1026 1709 -980 1747
rect -1026 1675 -1020 1709
rect -986 1675 -980 1709
rect -1026 1637 -980 1675
rect -1026 1603 -1020 1637
rect -986 1603 -980 1637
rect -1026 1565 -980 1603
rect -1026 1531 -1020 1565
rect -986 1531 -980 1565
rect -1026 1493 -980 1531
rect -1026 1459 -1020 1493
rect -986 1459 -980 1493
rect -1026 1421 -980 1459
rect -1026 1387 -1020 1421
rect -986 1387 -980 1421
rect -1026 1349 -980 1387
rect -1026 1315 -1020 1349
rect -986 1315 -980 1349
rect -1026 1277 -980 1315
rect -1026 1243 -1020 1277
rect -986 1243 -980 1277
rect -1026 1205 -980 1243
rect -1026 1171 -1020 1205
rect -986 1171 -980 1205
rect -1026 1133 -980 1171
rect -1026 1099 -1020 1133
rect -986 1099 -980 1133
rect -1026 1061 -980 1099
rect -1026 1027 -1020 1061
rect -986 1027 -980 1061
rect -1026 989 -980 1027
rect -1026 955 -1020 989
rect -986 955 -980 989
rect -1026 917 -980 955
rect -1026 883 -1020 917
rect -986 883 -980 917
rect -1026 845 -980 883
rect -1026 811 -1020 845
rect -986 811 -980 845
rect -1026 773 -980 811
rect -1026 739 -1020 773
rect -986 739 -980 773
rect -1026 701 -980 739
rect -1026 667 -1020 701
rect -986 667 -980 701
rect -1026 629 -980 667
rect -1026 595 -1020 629
rect -986 595 -980 629
rect -1026 557 -980 595
rect -1026 523 -1020 557
rect -986 523 -980 557
rect -1026 485 -980 523
rect -1026 451 -1020 485
rect -986 451 -980 485
rect -1026 413 -980 451
rect -1026 379 -1020 413
rect -986 379 -980 413
rect -1026 341 -980 379
rect -1026 307 -1020 341
rect -986 307 -980 341
rect -1026 269 -980 307
rect -1026 235 -1020 269
rect -986 235 -980 269
rect -1026 197 -980 235
rect -1026 163 -1020 197
rect -986 163 -980 197
rect -1026 125 -980 163
rect -1026 91 -1020 125
rect -986 91 -980 125
rect -1026 53 -980 91
rect -1026 19 -1020 53
rect -986 19 -980 53
rect -1026 -19 -980 19
rect -1026 -53 -1020 -19
rect -986 -53 -980 -19
rect -1026 -91 -980 -53
rect -1026 -125 -1020 -91
rect -986 -125 -980 -91
rect -1026 -163 -980 -125
rect -1026 -197 -1020 -163
rect -986 -197 -980 -163
rect -1026 -235 -980 -197
rect -1026 -269 -1020 -235
rect -986 -269 -980 -235
rect -1026 -307 -980 -269
rect -1026 -341 -1020 -307
rect -986 -341 -980 -307
rect -1026 -379 -980 -341
rect -1026 -413 -1020 -379
rect -986 -413 -980 -379
rect -1026 -451 -980 -413
rect -1026 -485 -1020 -451
rect -986 -485 -980 -451
rect -1026 -523 -980 -485
rect -1026 -557 -1020 -523
rect -986 -557 -980 -523
rect -1026 -595 -980 -557
rect -1026 -629 -1020 -595
rect -986 -629 -980 -595
rect -1026 -667 -980 -629
rect -1026 -701 -1020 -667
rect -986 -701 -980 -667
rect -1026 -739 -980 -701
rect -1026 -773 -1020 -739
rect -986 -773 -980 -739
rect -1026 -811 -980 -773
rect -1026 -845 -1020 -811
rect -986 -845 -980 -811
rect -1026 -883 -980 -845
rect -1026 -917 -1020 -883
rect -986 -917 -980 -883
rect -1026 -955 -980 -917
rect -1026 -989 -1020 -955
rect -986 -989 -980 -955
rect -1026 -1027 -980 -989
rect -1026 -1061 -1020 -1027
rect -986 -1061 -980 -1027
rect -1026 -1099 -980 -1061
rect -1026 -1133 -1020 -1099
rect -986 -1133 -980 -1099
rect -1026 -1171 -980 -1133
rect -1026 -1205 -1020 -1171
rect -986 -1205 -980 -1171
rect -1026 -1243 -980 -1205
rect -1026 -1277 -1020 -1243
rect -986 -1277 -980 -1243
rect -1026 -1315 -980 -1277
rect -1026 -1349 -1020 -1315
rect -986 -1349 -980 -1315
rect -1026 -1387 -980 -1349
rect -1026 -1421 -1020 -1387
rect -986 -1421 -980 -1387
rect -1026 -1459 -980 -1421
rect -1026 -1493 -1020 -1459
rect -986 -1493 -980 -1459
rect -1026 -1531 -980 -1493
rect -1026 -1565 -1020 -1531
rect -986 -1565 -980 -1531
rect -1026 -1603 -980 -1565
rect -1026 -1637 -1020 -1603
rect -986 -1637 -980 -1603
rect -1026 -1675 -980 -1637
rect -1026 -1709 -1020 -1675
rect -986 -1709 -980 -1675
rect -1026 -1747 -980 -1709
rect -1026 -1781 -1020 -1747
rect -986 -1781 -980 -1747
rect -1026 -1819 -980 -1781
rect -1026 -1853 -1020 -1819
rect -986 -1853 -980 -1819
rect -1026 -1891 -980 -1853
rect -1026 -1925 -1020 -1891
rect -986 -1925 -980 -1891
rect -1026 -1963 -980 -1925
rect -1026 -1997 -1020 -1963
rect -986 -1997 -980 -1963
rect -1026 -2035 -980 -1997
rect -1026 -2069 -1020 -2035
rect -986 -2069 -980 -2035
rect -1026 -2107 -980 -2069
rect -1026 -2141 -1020 -2107
rect -986 -2141 -980 -2107
rect -1026 -2179 -980 -2141
rect -1026 -2213 -1020 -2179
rect -986 -2213 -980 -2179
rect -1026 -2251 -980 -2213
rect -1026 -2285 -1020 -2251
rect -986 -2285 -980 -2251
rect -1026 -2323 -980 -2285
rect -1026 -2357 -1020 -2323
rect -986 -2357 -980 -2323
rect -1026 -2395 -980 -2357
rect -1026 -2429 -1020 -2395
rect -986 -2429 -980 -2395
rect -1026 -2467 -980 -2429
rect -1026 -2501 -1020 -2467
rect -986 -2501 -980 -2467
rect -1026 -2539 -980 -2501
rect -1026 -2573 -1020 -2539
rect -986 -2573 -980 -2539
rect -1026 -2611 -980 -2573
rect -1026 -2645 -1020 -2611
rect -986 -2645 -980 -2611
rect -1026 -2683 -980 -2645
rect -1026 -2717 -1020 -2683
rect -986 -2717 -980 -2683
rect -1026 -2755 -980 -2717
rect -1026 -2789 -1020 -2755
rect -986 -2789 -980 -2755
rect -1026 -2827 -980 -2789
rect -1026 -2861 -1020 -2827
rect -986 -2861 -980 -2827
rect -1026 -2899 -980 -2861
rect -1026 -2933 -1020 -2899
rect -986 -2933 -980 -2899
rect -1026 -2971 -980 -2933
rect -1026 -3005 -1020 -2971
rect -986 -3005 -980 -2971
rect -1026 -3043 -980 -3005
rect -1026 -3077 -1020 -3043
rect -986 -3077 -980 -3043
rect -1026 -3115 -980 -3077
rect -1026 -3149 -1020 -3115
rect -986 -3149 -980 -3115
rect -1026 -3187 -980 -3149
rect -1026 -3221 -1020 -3187
rect -986 -3221 -980 -3187
rect -1026 -3259 -980 -3221
rect -1026 -3293 -1020 -3259
rect -986 -3293 -980 -3259
rect -1026 -3331 -980 -3293
rect -1026 -3365 -1020 -3331
rect -986 -3365 -980 -3331
rect -1026 -3403 -980 -3365
rect -1026 -3437 -1020 -3403
rect -986 -3437 -980 -3403
rect -1026 -3475 -980 -3437
rect -1026 -3509 -1020 -3475
rect -986 -3509 -980 -3475
rect -1026 -3547 -980 -3509
rect -1026 -3581 -1020 -3547
rect -986 -3581 -980 -3547
rect -1026 -3619 -980 -3581
rect -1026 -3653 -1020 -3619
rect -986 -3653 -980 -3619
rect -1026 -3691 -980 -3653
rect -1026 -3725 -1020 -3691
rect -986 -3725 -980 -3691
rect -1026 -3763 -980 -3725
rect -1026 -3797 -1020 -3763
rect -986 -3797 -980 -3763
rect -1026 -3835 -980 -3797
rect -1026 -3869 -1020 -3835
rect -986 -3869 -980 -3835
rect -1026 -3907 -980 -3869
rect -1026 -3941 -1020 -3907
rect -986 -3941 -980 -3907
rect -1026 -3979 -980 -3941
rect -1026 -4013 -1020 -3979
rect -986 -4013 -980 -3979
rect -1026 -4051 -980 -4013
rect -1026 -4085 -1020 -4051
rect -986 -4085 -980 -4051
rect -1026 -4123 -980 -4085
rect -1026 -4157 -1020 -4123
rect -986 -4157 -980 -4123
rect -1026 -4195 -980 -4157
rect -1026 -4229 -1020 -4195
rect -986 -4229 -980 -4195
rect -1026 -4267 -980 -4229
rect -1026 -4301 -1020 -4267
rect -986 -4301 -980 -4267
rect -1026 -4339 -980 -4301
rect -1026 -4373 -1020 -4339
rect -986 -4373 -980 -4339
rect -1026 -4411 -980 -4373
rect -1026 -4445 -1020 -4411
rect -986 -4445 -980 -4411
rect -1026 -4483 -980 -4445
rect -1026 -4517 -1020 -4483
rect -986 -4517 -980 -4483
rect -1026 -4555 -980 -4517
rect -1026 -4589 -1020 -4555
rect -986 -4589 -980 -4555
rect -1026 -4627 -980 -4589
rect -1026 -4661 -1020 -4627
rect -986 -4661 -980 -4627
rect -1026 -4699 -980 -4661
rect -1026 -4733 -1020 -4699
rect -986 -4733 -980 -4699
rect -1026 -4771 -980 -4733
rect -1026 -4805 -1020 -4771
rect -986 -4805 -980 -4771
rect -1026 -4843 -980 -4805
rect -1026 -4877 -1020 -4843
rect -986 -4877 -980 -4843
rect -1026 -4915 -980 -4877
rect -1026 -4949 -1020 -4915
rect -986 -4949 -980 -4915
rect -1026 -4987 -980 -4949
rect -1026 -5021 -1020 -4987
rect -986 -5021 -980 -4987
rect -1026 -5059 -980 -5021
rect -1026 -5093 -1020 -5059
rect -986 -5093 -980 -5059
rect -1026 -5131 -980 -5093
rect -1026 -5165 -1020 -5131
rect -986 -5165 -980 -5131
rect -1026 -5203 -980 -5165
rect -1026 -5237 -1020 -5203
rect -986 -5237 -980 -5203
rect -1026 -5275 -980 -5237
rect -1026 -5309 -1020 -5275
rect -986 -5309 -980 -5275
rect -1026 -5347 -980 -5309
rect -1026 -5381 -1020 -5347
rect -986 -5381 -980 -5347
rect -1026 -5419 -980 -5381
rect -1026 -5453 -1020 -5419
rect -986 -5453 -980 -5419
rect -1026 -5491 -980 -5453
rect -1026 -5525 -1020 -5491
rect -986 -5525 -980 -5491
rect -1026 -5563 -980 -5525
rect -1026 -5597 -1020 -5563
rect -986 -5597 -980 -5563
rect -1026 -5635 -980 -5597
rect -1026 -5669 -1020 -5635
rect -986 -5669 -980 -5635
rect -1026 -5707 -980 -5669
rect -1026 -5741 -1020 -5707
rect -986 -5741 -980 -5707
rect -1026 -5779 -980 -5741
rect -1026 -5813 -1020 -5779
rect -986 -5813 -980 -5779
rect -1026 -5851 -980 -5813
rect -1026 -5885 -1020 -5851
rect -986 -5885 -980 -5851
rect -1026 -5923 -980 -5885
rect -1026 -5957 -1020 -5923
rect -986 -5957 -980 -5923
rect -1026 -5995 -980 -5957
rect -1026 -6029 -1020 -5995
rect -986 -6029 -980 -5995
rect -1026 -6067 -980 -6029
rect -1026 -6101 -1020 -6067
rect -986 -6101 -980 -6067
rect -1026 -6139 -980 -6101
rect -1026 -6173 -1020 -6139
rect -986 -6173 -980 -6139
rect -1026 -6211 -980 -6173
rect -1026 -6245 -1020 -6211
rect -986 -6245 -980 -6211
rect -1026 -6283 -980 -6245
rect -1026 -6317 -1020 -6283
rect -986 -6317 -980 -6283
rect -1026 -6355 -980 -6317
rect -1026 -6389 -1020 -6355
rect -986 -6389 -980 -6355
rect -1026 -6427 -980 -6389
rect -1026 -6461 -1020 -6427
rect -986 -6461 -980 -6427
rect -1026 -6499 -980 -6461
rect -1026 -6533 -1020 -6499
rect -986 -6533 -980 -6499
rect -1026 -6571 -980 -6533
rect -1026 -6605 -1020 -6571
rect -986 -6605 -980 -6571
rect -1026 -6643 -980 -6605
rect -1026 -6677 -1020 -6643
rect -986 -6677 -980 -6643
rect -1026 -6715 -980 -6677
rect -1026 -6749 -1020 -6715
rect -986 -6749 -980 -6715
rect -1026 -6787 -980 -6749
rect -1026 -6821 -1020 -6787
rect -986 -6821 -980 -6787
rect -1026 -6859 -980 -6821
rect -1026 -6893 -1020 -6859
rect -986 -6893 -980 -6859
rect -1026 -6931 -980 -6893
rect -1026 -6965 -1020 -6931
rect -986 -6965 -980 -6931
rect -1026 -7003 -980 -6965
rect -1026 -7037 -1020 -7003
rect -986 -7037 -980 -7003
rect -1026 -7075 -980 -7037
rect -1026 -7109 -1020 -7075
rect -986 -7109 -980 -7075
rect -1026 -7147 -980 -7109
rect -1026 -7181 -1020 -7147
rect -986 -7181 -980 -7147
rect -1026 -7219 -980 -7181
rect -1026 -7253 -1020 -7219
rect -986 -7253 -980 -7219
rect -1026 -7291 -980 -7253
rect -1026 -7325 -1020 -7291
rect -986 -7325 -980 -7291
rect -1026 -7363 -980 -7325
rect -1026 -7397 -1020 -7363
rect -986 -7397 -980 -7363
rect -1026 -7435 -980 -7397
rect -1026 -7469 -1020 -7435
rect -986 -7469 -980 -7435
rect -1026 -7507 -980 -7469
rect -1026 -7541 -1020 -7507
rect -986 -7541 -980 -7507
rect -1026 -7579 -980 -7541
rect -1026 -7613 -1020 -7579
rect -986 -7613 -980 -7579
rect -1026 -7651 -980 -7613
rect -1026 -7685 -1020 -7651
rect -986 -7685 -980 -7651
rect -1026 -7723 -980 -7685
rect -1026 -7757 -1020 -7723
rect -986 -7757 -980 -7723
rect -1026 -7795 -980 -7757
rect -1026 -7829 -1020 -7795
rect -986 -7829 -980 -7795
rect -1026 -7867 -980 -7829
rect -1026 -7901 -1020 -7867
rect -986 -7901 -980 -7867
rect -1026 -7939 -980 -7901
rect -1026 -7973 -1020 -7939
rect -986 -7973 -980 -7939
rect -1026 -8011 -980 -7973
rect -1026 -8045 -1020 -8011
rect -986 -8045 -980 -8011
rect -1026 -8083 -980 -8045
rect -1026 -8117 -1020 -8083
rect -986 -8117 -980 -8083
rect -1026 -8155 -980 -8117
rect -1026 -8189 -1020 -8155
rect -986 -8189 -980 -8155
rect -1026 -8227 -980 -8189
rect -1026 -8261 -1020 -8227
rect -986 -8261 -980 -8227
rect -1026 -8299 -980 -8261
rect -1026 -8333 -1020 -8299
rect -986 -8333 -980 -8299
rect -1026 -8371 -980 -8333
rect -1026 -8405 -1020 -8371
rect -986 -8405 -980 -8371
rect -1026 -8443 -980 -8405
rect -1026 -8477 -1020 -8443
rect -986 -8477 -980 -8443
rect -1026 -8515 -980 -8477
rect -1026 -8549 -1020 -8515
rect -986 -8549 -980 -8515
rect -1026 -8587 -980 -8549
rect -1026 -8621 -1020 -8587
rect -986 -8621 -980 -8587
rect -1026 -8659 -980 -8621
rect -1026 -8693 -1020 -8659
rect -986 -8693 -980 -8659
rect -1026 -8731 -980 -8693
rect -1026 -8765 -1020 -8731
rect -986 -8765 -980 -8731
rect -1026 -8803 -980 -8765
rect -1026 -8837 -1020 -8803
rect -986 -8837 -980 -8803
rect -1026 -8875 -980 -8837
rect -1026 -8909 -1020 -8875
rect -986 -8909 -980 -8875
rect -1026 -8947 -980 -8909
rect -1026 -8981 -1020 -8947
rect -986 -8981 -980 -8947
rect -1026 -9019 -980 -8981
rect -1026 -9053 -1020 -9019
rect -986 -9053 -980 -9019
rect -1026 -9091 -980 -9053
rect -1026 -9125 -1020 -9091
rect -986 -9125 -980 -9091
rect -1026 -9163 -980 -9125
rect -1026 -9197 -1020 -9163
rect -986 -9197 -980 -9163
rect -1026 -9235 -980 -9197
rect -1026 -9269 -1020 -9235
rect -986 -9269 -980 -9235
rect -1026 -9307 -980 -9269
rect -1026 -9341 -1020 -9307
rect -986 -9341 -980 -9307
rect -1026 -9379 -980 -9341
rect -1026 -9413 -1020 -9379
rect -986 -9413 -980 -9379
rect -1026 -9451 -980 -9413
rect -1026 -9485 -1020 -9451
rect -986 -9485 -980 -9451
rect -1026 -9523 -980 -9485
rect -1026 -9557 -1020 -9523
rect -986 -9557 -980 -9523
rect -1026 -9600 -980 -9557
rect -908 9557 -862 9600
rect -908 9523 -902 9557
rect -868 9523 -862 9557
rect -908 9485 -862 9523
rect -908 9451 -902 9485
rect -868 9451 -862 9485
rect -908 9413 -862 9451
rect -908 9379 -902 9413
rect -868 9379 -862 9413
rect -908 9341 -862 9379
rect -908 9307 -902 9341
rect -868 9307 -862 9341
rect -908 9269 -862 9307
rect -908 9235 -902 9269
rect -868 9235 -862 9269
rect -908 9197 -862 9235
rect -908 9163 -902 9197
rect -868 9163 -862 9197
rect -908 9125 -862 9163
rect -908 9091 -902 9125
rect -868 9091 -862 9125
rect -908 9053 -862 9091
rect -908 9019 -902 9053
rect -868 9019 -862 9053
rect -908 8981 -862 9019
rect -908 8947 -902 8981
rect -868 8947 -862 8981
rect -908 8909 -862 8947
rect -908 8875 -902 8909
rect -868 8875 -862 8909
rect -908 8837 -862 8875
rect -908 8803 -902 8837
rect -868 8803 -862 8837
rect -908 8765 -862 8803
rect -908 8731 -902 8765
rect -868 8731 -862 8765
rect -908 8693 -862 8731
rect -908 8659 -902 8693
rect -868 8659 -862 8693
rect -908 8621 -862 8659
rect -908 8587 -902 8621
rect -868 8587 -862 8621
rect -908 8549 -862 8587
rect -908 8515 -902 8549
rect -868 8515 -862 8549
rect -908 8477 -862 8515
rect -908 8443 -902 8477
rect -868 8443 -862 8477
rect -908 8405 -862 8443
rect -908 8371 -902 8405
rect -868 8371 -862 8405
rect -908 8333 -862 8371
rect -908 8299 -902 8333
rect -868 8299 -862 8333
rect -908 8261 -862 8299
rect -908 8227 -902 8261
rect -868 8227 -862 8261
rect -908 8189 -862 8227
rect -908 8155 -902 8189
rect -868 8155 -862 8189
rect -908 8117 -862 8155
rect -908 8083 -902 8117
rect -868 8083 -862 8117
rect -908 8045 -862 8083
rect -908 8011 -902 8045
rect -868 8011 -862 8045
rect -908 7973 -862 8011
rect -908 7939 -902 7973
rect -868 7939 -862 7973
rect -908 7901 -862 7939
rect -908 7867 -902 7901
rect -868 7867 -862 7901
rect -908 7829 -862 7867
rect -908 7795 -902 7829
rect -868 7795 -862 7829
rect -908 7757 -862 7795
rect -908 7723 -902 7757
rect -868 7723 -862 7757
rect -908 7685 -862 7723
rect -908 7651 -902 7685
rect -868 7651 -862 7685
rect -908 7613 -862 7651
rect -908 7579 -902 7613
rect -868 7579 -862 7613
rect -908 7541 -862 7579
rect -908 7507 -902 7541
rect -868 7507 -862 7541
rect -908 7469 -862 7507
rect -908 7435 -902 7469
rect -868 7435 -862 7469
rect -908 7397 -862 7435
rect -908 7363 -902 7397
rect -868 7363 -862 7397
rect -908 7325 -862 7363
rect -908 7291 -902 7325
rect -868 7291 -862 7325
rect -908 7253 -862 7291
rect -908 7219 -902 7253
rect -868 7219 -862 7253
rect -908 7181 -862 7219
rect -908 7147 -902 7181
rect -868 7147 -862 7181
rect -908 7109 -862 7147
rect -908 7075 -902 7109
rect -868 7075 -862 7109
rect -908 7037 -862 7075
rect -908 7003 -902 7037
rect -868 7003 -862 7037
rect -908 6965 -862 7003
rect -908 6931 -902 6965
rect -868 6931 -862 6965
rect -908 6893 -862 6931
rect -908 6859 -902 6893
rect -868 6859 -862 6893
rect -908 6821 -862 6859
rect -908 6787 -902 6821
rect -868 6787 -862 6821
rect -908 6749 -862 6787
rect -908 6715 -902 6749
rect -868 6715 -862 6749
rect -908 6677 -862 6715
rect -908 6643 -902 6677
rect -868 6643 -862 6677
rect -908 6605 -862 6643
rect -908 6571 -902 6605
rect -868 6571 -862 6605
rect -908 6533 -862 6571
rect -908 6499 -902 6533
rect -868 6499 -862 6533
rect -908 6461 -862 6499
rect -908 6427 -902 6461
rect -868 6427 -862 6461
rect -908 6389 -862 6427
rect -908 6355 -902 6389
rect -868 6355 -862 6389
rect -908 6317 -862 6355
rect -908 6283 -902 6317
rect -868 6283 -862 6317
rect -908 6245 -862 6283
rect -908 6211 -902 6245
rect -868 6211 -862 6245
rect -908 6173 -862 6211
rect -908 6139 -902 6173
rect -868 6139 -862 6173
rect -908 6101 -862 6139
rect -908 6067 -902 6101
rect -868 6067 -862 6101
rect -908 6029 -862 6067
rect -908 5995 -902 6029
rect -868 5995 -862 6029
rect -908 5957 -862 5995
rect -908 5923 -902 5957
rect -868 5923 -862 5957
rect -908 5885 -862 5923
rect -908 5851 -902 5885
rect -868 5851 -862 5885
rect -908 5813 -862 5851
rect -908 5779 -902 5813
rect -868 5779 -862 5813
rect -908 5741 -862 5779
rect -908 5707 -902 5741
rect -868 5707 -862 5741
rect -908 5669 -862 5707
rect -908 5635 -902 5669
rect -868 5635 -862 5669
rect -908 5597 -862 5635
rect -908 5563 -902 5597
rect -868 5563 -862 5597
rect -908 5525 -862 5563
rect -908 5491 -902 5525
rect -868 5491 -862 5525
rect -908 5453 -862 5491
rect -908 5419 -902 5453
rect -868 5419 -862 5453
rect -908 5381 -862 5419
rect -908 5347 -902 5381
rect -868 5347 -862 5381
rect -908 5309 -862 5347
rect -908 5275 -902 5309
rect -868 5275 -862 5309
rect -908 5237 -862 5275
rect -908 5203 -902 5237
rect -868 5203 -862 5237
rect -908 5165 -862 5203
rect -908 5131 -902 5165
rect -868 5131 -862 5165
rect -908 5093 -862 5131
rect -908 5059 -902 5093
rect -868 5059 -862 5093
rect -908 5021 -862 5059
rect -908 4987 -902 5021
rect -868 4987 -862 5021
rect -908 4949 -862 4987
rect -908 4915 -902 4949
rect -868 4915 -862 4949
rect -908 4877 -862 4915
rect -908 4843 -902 4877
rect -868 4843 -862 4877
rect -908 4805 -862 4843
rect -908 4771 -902 4805
rect -868 4771 -862 4805
rect -908 4733 -862 4771
rect -908 4699 -902 4733
rect -868 4699 -862 4733
rect -908 4661 -862 4699
rect -908 4627 -902 4661
rect -868 4627 -862 4661
rect -908 4589 -862 4627
rect -908 4555 -902 4589
rect -868 4555 -862 4589
rect -908 4517 -862 4555
rect -908 4483 -902 4517
rect -868 4483 -862 4517
rect -908 4445 -862 4483
rect -908 4411 -902 4445
rect -868 4411 -862 4445
rect -908 4373 -862 4411
rect -908 4339 -902 4373
rect -868 4339 -862 4373
rect -908 4301 -862 4339
rect -908 4267 -902 4301
rect -868 4267 -862 4301
rect -908 4229 -862 4267
rect -908 4195 -902 4229
rect -868 4195 -862 4229
rect -908 4157 -862 4195
rect -908 4123 -902 4157
rect -868 4123 -862 4157
rect -908 4085 -862 4123
rect -908 4051 -902 4085
rect -868 4051 -862 4085
rect -908 4013 -862 4051
rect -908 3979 -902 4013
rect -868 3979 -862 4013
rect -908 3941 -862 3979
rect -908 3907 -902 3941
rect -868 3907 -862 3941
rect -908 3869 -862 3907
rect -908 3835 -902 3869
rect -868 3835 -862 3869
rect -908 3797 -862 3835
rect -908 3763 -902 3797
rect -868 3763 -862 3797
rect -908 3725 -862 3763
rect -908 3691 -902 3725
rect -868 3691 -862 3725
rect -908 3653 -862 3691
rect -908 3619 -902 3653
rect -868 3619 -862 3653
rect -908 3581 -862 3619
rect -908 3547 -902 3581
rect -868 3547 -862 3581
rect -908 3509 -862 3547
rect -908 3475 -902 3509
rect -868 3475 -862 3509
rect -908 3437 -862 3475
rect -908 3403 -902 3437
rect -868 3403 -862 3437
rect -908 3365 -862 3403
rect -908 3331 -902 3365
rect -868 3331 -862 3365
rect -908 3293 -862 3331
rect -908 3259 -902 3293
rect -868 3259 -862 3293
rect -908 3221 -862 3259
rect -908 3187 -902 3221
rect -868 3187 -862 3221
rect -908 3149 -862 3187
rect -908 3115 -902 3149
rect -868 3115 -862 3149
rect -908 3077 -862 3115
rect -908 3043 -902 3077
rect -868 3043 -862 3077
rect -908 3005 -862 3043
rect -908 2971 -902 3005
rect -868 2971 -862 3005
rect -908 2933 -862 2971
rect -908 2899 -902 2933
rect -868 2899 -862 2933
rect -908 2861 -862 2899
rect -908 2827 -902 2861
rect -868 2827 -862 2861
rect -908 2789 -862 2827
rect -908 2755 -902 2789
rect -868 2755 -862 2789
rect -908 2717 -862 2755
rect -908 2683 -902 2717
rect -868 2683 -862 2717
rect -908 2645 -862 2683
rect -908 2611 -902 2645
rect -868 2611 -862 2645
rect -908 2573 -862 2611
rect -908 2539 -902 2573
rect -868 2539 -862 2573
rect -908 2501 -862 2539
rect -908 2467 -902 2501
rect -868 2467 -862 2501
rect -908 2429 -862 2467
rect -908 2395 -902 2429
rect -868 2395 -862 2429
rect -908 2357 -862 2395
rect -908 2323 -902 2357
rect -868 2323 -862 2357
rect -908 2285 -862 2323
rect -908 2251 -902 2285
rect -868 2251 -862 2285
rect -908 2213 -862 2251
rect -908 2179 -902 2213
rect -868 2179 -862 2213
rect -908 2141 -862 2179
rect -908 2107 -902 2141
rect -868 2107 -862 2141
rect -908 2069 -862 2107
rect -908 2035 -902 2069
rect -868 2035 -862 2069
rect -908 1997 -862 2035
rect -908 1963 -902 1997
rect -868 1963 -862 1997
rect -908 1925 -862 1963
rect -908 1891 -902 1925
rect -868 1891 -862 1925
rect -908 1853 -862 1891
rect -908 1819 -902 1853
rect -868 1819 -862 1853
rect -908 1781 -862 1819
rect -908 1747 -902 1781
rect -868 1747 -862 1781
rect -908 1709 -862 1747
rect -908 1675 -902 1709
rect -868 1675 -862 1709
rect -908 1637 -862 1675
rect -908 1603 -902 1637
rect -868 1603 -862 1637
rect -908 1565 -862 1603
rect -908 1531 -902 1565
rect -868 1531 -862 1565
rect -908 1493 -862 1531
rect -908 1459 -902 1493
rect -868 1459 -862 1493
rect -908 1421 -862 1459
rect -908 1387 -902 1421
rect -868 1387 -862 1421
rect -908 1349 -862 1387
rect -908 1315 -902 1349
rect -868 1315 -862 1349
rect -908 1277 -862 1315
rect -908 1243 -902 1277
rect -868 1243 -862 1277
rect -908 1205 -862 1243
rect -908 1171 -902 1205
rect -868 1171 -862 1205
rect -908 1133 -862 1171
rect -908 1099 -902 1133
rect -868 1099 -862 1133
rect -908 1061 -862 1099
rect -908 1027 -902 1061
rect -868 1027 -862 1061
rect -908 989 -862 1027
rect -908 955 -902 989
rect -868 955 -862 989
rect -908 917 -862 955
rect -908 883 -902 917
rect -868 883 -862 917
rect -908 845 -862 883
rect -908 811 -902 845
rect -868 811 -862 845
rect -908 773 -862 811
rect -908 739 -902 773
rect -868 739 -862 773
rect -908 701 -862 739
rect -908 667 -902 701
rect -868 667 -862 701
rect -908 629 -862 667
rect -908 595 -902 629
rect -868 595 -862 629
rect -908 557 -862 595
rect -908 523 -902 557
rect -868 523 -862 557
rect -908 485 -862 523
rect -908 451 -902 485
rect -868 451 -862 485
rect -908 413 -862 451
rect -908 379 -902 413
rect -868 379 -862 413
rect -908 341 -862 379
rect -908 307 -902 341
rect -868 307 -862 341
rect -908 269 -862 307
rect -908 235 -902 269
rect -868 235 -862 269
rect -908 197 -862 235
rect -908 163 -902 197
rect -868 163 -862 197
rect -908 125 -862 163
rect -908 91 -902 125
rect -868 91 -862 125
rect -908 53 -862 91
rect -908 19 -902 53
rect -868 19 -862 53
rect -908 -19 -862 19
rect -908 -53 -902 -19
rect -868 -53 -862 -19
rect -908 -91 -862 -53
rect -908 -125 -902 -91
rect -868 -125 -862 -91
rect -908 -163 -862 -125
rect -908 -197 -902 -163
rect -868 -197 -862 -163
rect -908 -235 -862 -197
rect -908 -269 -902 -235
rect -868 -269 -862 -235
rect -908 -307 -862 -269
rect -908 -341 -902 -307
rect -868 -341 -862 -307
rect -908 -379 -862 -341
rect -908 -413 -902 -379
rect -868 -413 -862 -379
rect -908 -451 -862 -413
rect -908 -485 -902 -451
rect -868 -485 -862 -451
rect -908 -523 -862 -485
rect -908 -557 -902 -523
rect -868 -557 -862 -523
rect -908 -595 -862 -557
rect -908 -629 -902 -595
rect -868 -629 -862 -595
rect -908 -667 -862 -629
rect -908 -701 -902 -667
rect -868 -701 -862 -667
rect -908 -739 -862 -701
rect -908 -773 -902 -739
rect -868 -773 -862 -739
rect -908 -811 -862 -773
rect -908 -845 -902 -811
rect -868 -845 -862 -811
rect -908 -883 -862 -845
rect -908 -917 -902 -883
rect -868 -917 -862 -883
rect -908 -955 -862 -917
rect -908 -989 -902 -955
rect -868 -989 -862 -955
rect -908 -1027 -862 -989
rect -908 -1061 -902 -1027
rect -868 -1061 -862 -1027
rect -908 -1099 -862 -1061
rect -908 -1133 -902 -1099
rect -868 -1133 -862 -1099
rect -908 -1171 -862 -1133
rect -908 -1205 -902 -1171
rect -868 -1205 -862 -1171
rect -908 -1243 -862 -1205
rect -908 -1277 -902 -1243
rect -868 -1277 -862 -1243
rect -908 -1315 -862 -1277
rect -908 -1349 -902 -1315
rect -868 -1349 -862 -1315
rect -908 -1387 -862 -1349
rect -908 -1421 -902 -1387
rect -868 -1421 -862 -1387
rect -908 -1459 -862 -1421
rect -908 -1493 -902 -1459
rect -868 -1493 -862 -1459
rect -908 -1531 -862 -1493
rect -908 -1565 -902 -1531
rect -868 -1565 -862 -1531
rect -908 -1603 -862 -1565
rect -908 -1637 -902 -1603
rect -868 -1637 -862 -1603
rect -908 -1675 -862 -1637
rect -908 -1709 -902 -1675
rect -868 -1709 -862 -1675
rect -908 -1747 -862 -1709
rect -908 -1781 -902 -1747
rect -868 -1781 -862 -1747
rect -908 -1819 -862 -1781
rect -908 -1853 -902 -1819
rect -868 -1853 -862 -1819
rect -908 -1891 -862 -1853
rect -908 -1925 -902 -1891
rect -868 -1925 -862 -1891
rect -908 -1963 -862 -1925
rect -908 -1997 -902 -1963
rect -868 -1997 -862 -1963
rect -908 -2035 -862 -1997
rect -908 -2069 -902 -2035
rect -868 -2069 -862 -2035
rect -908 -2107 -862 -2069
rect -908 -2141 -902 -2107
rect -868 -2141 -862 -2107
rect -908 -2179 -862 -2141
rect -908 -2213 -902 -2179
rect -868 -2213 -862 -2179
rect -908 -2251 -862 -2213
rect -908 -2285 -902 -2251
rect -868 -2285 -862 -2251
rect -908 -2323 -862 -2285
rect -908 -2357 -902 -2323
rect -868 -2357 -862 -2323
rect -908 -2395 -862 -2357
rect -908 -2429 -902 -2395
rect -868 -2429 -862 -2395
rect -908 -2467 -862 -2429
rect -908 -2501 -902 -2467
rect -868 -2501 -862 -2467
rect -908 -2539 -862 -2501
rect -908 -2573 -902 -2539
rect -868 -2573 -862 -2539
rect -908 -2611 -862 -2573
rect -908 -2645 -902 -2611
rect -868 -2645 -862 -2611
rect -908 -2683 -862 -2645
rect -908 -2717 -902 -2683
rect -868 -2717 -862 -2683
rect -908 -2755 -862 -2717
rect -908 -2789 -902 -2755
rect -868 -2789 -862 -2755
rect -908 -2827 -862 -2789
rect -908 -2861 -902 -2827
rect -868 -2861 -862 -2827
rect -908 -2899 -862 -2861
rect -908 -2933 -902 -2899
rect -868 -2933 -862 -2899
rect -908 -2971 -862 -2933
rect -908 -3005 -902 -2971
rect -868 -3005 -862 -2971
rect -908 -3043 -862 -3005
rect -908 -3077 -902 -3043
rect -868 -3077 -862 -3043
rect -908 -3115 -862 -3077
rect -908 -3149 -902 -3115
rect -868 -3149 -862 -3115
rect -908 -3187 -862 -3149
rect -908 -3221 -902 -3187
rect -868 -3221 -862 -3187
rect -908 -3259 -862 -3221
rect -908 -3293 -902 -3259
rect -868 -3293 -862 -3259
rect -908 -3331 -862 -3293
rect -908 -3365 -902 -3331
rect -868 -3365 -862 -3331
rect -908 -3403 -862 -3365
rect -908 -3437 -902 -3403
rect -868 -3437 -862 -3403
rect -908 -3475 -862 -3437
rect -908 -3509 -902 -3475
rect -868 -3509 -862 -3475
rect -908 -3547 -862 -3509
rect -908 -3581 -902 -3547
rect -868 -3581 -862 -3547
rect -908 -3619 -862 -3581
rect -908 -3653 -902 -3619
rect -868 -3653 -862 -3619
rect -908 -3691 -862 -3653
rect -908 -3725 -902 -3691
rect -868 -3725 -862 -3691
rect -908 -3763 -862 -3725
rect -908 -3797 -902 -3763
rect -868 -3797 -862 -3763
rect -908 -3835 -862 -3797
rect -908 -3869 -902 -3835
rect -868 -3869 -862 -3835
rect -908 -3907 -862 -3869
rect -908 -3941 -902 -3907
rect -868 -3941 -862 -3907
rect -908 -3979 -862 -3941
rect -908 -4013 -902 -3979
rect -868 -4013 -862 -3979
rect -908 -4051 -862 -4013
rect -908 -4085 -902 -4051
rect -868 -4085 -862 -4051
rect -908 -4123 -862 -4085
rect -908 -4157 -902 -4123
rect -868 -4157 -862 -4123
rect -908 -4195 -862 -4157
rect -908 -4229 -902 -4195
rect -868 -4229 -862 -4195
rect -908 -4267 -862 -4229
rect -908 -4301 -902 -4267
rect -868 -4301 -862 -4267
rect -908 -4339 -862 -4301
rect -908 -4373 -902 -4339
rect -868 -4373 -862 -4339
rect -908 -4411 -862 -4373
rect -908 -4445 -902 -4411
rect -868 -4445 -862 -4411
rect -908 -4483 -862 -4445
rect -908 -4517 -902 -4483
rect -868 -4517 -862 -4483
rect -908 -4555 -862 -4517
rect -908 -4589 -902 -4555
rect -868 -4589 -862 -4555
rect -908 -4627 -862 -4589
rect -908 -4661 -902 -4627
rect -868 -4661 -862 -4627
rect -908 -4699 -862 -4661
rect -908 -4733 -902 -4699
rect -868 -4733 -862 -4699
rect -908 -4771 -862 -4733
rect -908 -4805 -902 -4771
rect -868 -4805 -862 -4771
rect -908 -4843 -862 -4805
rect -908 -4877 -902 -4843
rect -868 -4877 -862 -4843
rect -908 -4915 -862 -4877
rect -908 -4949 -902 -4915
rect -868 -4949 -862 -4915
rect -908 -4987 -862 -4949
rect -908 -5021 -902 -4987
rect -868 -5021 -862 -4987
rect -908 -5059 -862 -5021
rect -908 -5093 -902 -5059
rect -868 -5093 -862 -5059
rect -908 -5131 -862 -5093
rect -908 -5165 -902 -5131
rect -868 -5165 -862 -5131
rect -908 -5203 -862 -5165
rect -908 -5237 -902 -5203
rect -868 -5237 -862 -5203
rect -908 -5275 -862 -5237
rect -908 -5309 -902 -5275
rect -868 -5309 -862 -5275
rect -908 -5347 -862 -5309
rect -908 -5381 -902 -5347
rect -868 -5381 -862 -5347
rect -908 -5419 -862 -5381
rect -908 -5453 -902 -5419
rect -868 -5453 -862 -5419
rect -908 -5491 -862 -5453
rect -908 -5525 -902 -5491
rect -868 -5525 -862 -5491
rect -908 -5563 -862 -5525
rect -908 -5597 -902 -5563
rect -868 -5597 -862 -5563
rect -908 -5635 -862 -5597
rect -908 -5669 -902 -5635
rect -868 -5669 -862 -5635
rect -908 -5707 -862 -5669
rect -908 -5741 -902 -5707
rect -868 -5741 -862 -5707
rect -908 -5779 -862 -5741
rect -908 -5813 -902 -5779
rect -868 -5813 -862 -5779
rect -908 -5851 -862 -5813
rect -908 -5885 -902 -5851
rect -868 -5885 -862 -5851
rect -908 -5923 -862 -5885
rect -908 -5957 -902 -5923
rect -868 -5957 -862 -5923
rect -908 -5995 -862 -5957
rect -908 -6029 -902 -5995
rect -868 -6029 -862 -5995
rect -908 -6067 -862 -6029
rect -908 -6101 -902 -6067
rect -868 -6101 -862 -6067
rect -908 -6139 -862 -6101
rect -908 -6173 -902 -6139
rect -868 -6173 -862 -6139
rect -908 -6211 -862 -6173
rect -908 -6245 -902 -6211
rect -868 -6245 -862 -6211
rect -908 -6283 -862 -6245
rect -908 -6317 -902 -6283
rect -868 -6317 -862 -6283
rect -908 -6355 -862 -6317
rect -908 -6389 -902 -6355
rect -868 -6389 -862 -6355
rect -908 -6427 -862 -6389
rect -908 -6461 -902 -6427
rect -868 -6461 -862 -6427
rect -908 -6499 -862 -6461
rect -908 -6533 -902 -6499
rect -868 -6533 -862 -6499
rect -908 -6571 -862 -6533
rect -908 -6605 -902 -6571
rect -868 -6605 -862 -6571
rect -908 -6643 -862 -6605
rect -908 -6677 -902 -6643
rect -868 -6677 -862 -6643
rect -908 -6715 -862 -6677
rect -908 -6749 -902 -6715
rect -868 -6749 -862 -6715
rect -908 -6787 -862 -6749
rect -908 -6821 -902 -6787
rect -868 -6821 -862 -6787
rect -908 -6859 -862 -6821
rect -908 -6893 -902 -6859
rect -868 -6893 -862 -6859
rect -908 -6931 -862 -6893
rect -908 -6965 -902 -6931
rect -868 -6965 -862 -6931
rect -908 -7003 -862 -6965
rect -908 -7037 -902 -7003
rect -868 -7037 -862 -7003
rect -908 -7075 -862 -7037
rect -908 -7109 -902 -7075
rect -868 -7109 -862 -7075
rect -908 -7147 -862 -7109
rect -908 -7181 -902 -7147
rect -868 -7181 -862 -7147
rect -908 -7219 -862 -7181
rect -908 -7253 -902 -7219
rect -868 -7253 -862 -7219
rect -908 -7291 -862 -7253
rect -908 -7325 -902 -7291
rect -868 -7325 -862 -7291
rect -908 -7363 -862 -7325
rect -908 -7397 -902 -7363
rect -868 -7397 -862 -7363
rect -908 -7435 -862 -7397
rect -908 -7469 -902 -7435
rect -868 -7469 -862 -7435
rect -908 -7507 -862 -7469
rect -908 -7541 -902 -7507
rect -868 -7541 -862 -7507
rect -908 -7579 -862 -7541
rect -908 -7613 -902 -7579
rect -868 -7613 -862 -7579
rect -908 -7651 -862 -7613
rect -908 -7685 -902 -7651
rect -868 -7685 -862 -7651
rect -908 -7723 -862 -7685
rect -908 -7757 -902 -7723
rect -868 -7757 -862 -7723
rect -908 -7795 -862 -7757
rect -908 -7829 -902 -7795
rect -868 -7829 -862 -7795
rect -908 -7867 -862 -7829
rect -908 -7901 -902 -7867
rect -868 -7901 -862 -7867
rect -908 -7939 -862 -7901
rect -908 -7973 -902 -7939
rect -868 -7973 -862 -7939
rect -908 -8011 -862 -7973
rect -908 -8045 -902 -8011
rect -868 -8045 -862 -8011
rect -908 -8083 -862 -8045
rect -908 -8117 -902 -8083
rect -868 -8117 -862 -8083
rect -908 -8155 -862 -8117
rect -908 -8189 -902 -8155
rect -868 -8189 -862 -8155
rect -908 -8227 -862 -8189
rect -908 -8261 -902 -8227
rect -868 -8261 -862 -8227
rect -908 -8299 -862 -8261
rect -908 -8333 -902 -8299
rect -868 -8333 -862 -8299
rect -908 -8371 -862 -8333
rect -908 -8405 -902 -8371
rect -868 -8405 -862 -8371
rect -908 -8443 -862 -8405
rect -908 -8477 -902 -8443
rect -868 -8477 -862 -8443
rect -908 -8515 -862 -8477
rect -908 -8549 -902 -8515
rect -868 -8549 -862 -8515
rect -908 -8587 -862 -8549
rect -908 -8621 -902 -8587
rect -868 -8621 -862 -8587
rect -908 -8659 -862 -8621
rect -908 -8693 -902 -8659
rect -868 -8693 -862 -8659
rect -908 -8731 -862 -8693
rect -908 -8765 -902 -8731
rect -868 -8765 -862 -8731
rect -908 -8803 -862 -8765
rect -908 -8837 -902 -8803
rect -868 -8837 -862 -8803
rect -908 -8875 -862 -8837
rect -908 -8909 -902 -8875
rect -868 -8909 -862 -8875
rect -908 -8947 -862 -8909
rect -908 -8981 -902 -8947
rect -868 -8981 -862 -8947
rect -908 -9019 -862 -8981
rect -908 -9053 -902 -9019
rect -868 -9053 -862 -9019
rect -908 -9091 -862 -9053
rect -908 -9125 -902 -9091
rect -868 -9125 -862 -9091
rect -908 -9163 -862 -9125
rect -908 -9197 -902 -9163
rect -868 -9197 -862 -9163
rect -908 -9235 -862 -9197
rect -908 -9269 -902 -9235
rect -868 -9269 -862 -9235
rect -908 -9307 -862 -9269
rect -908 -9341 -902 -9307
rect -868 -9341 -862 -9307
rect -908 -9379 -862 -9341
rect -908 -9413 -902 -9379
rect -868 -9413 -862 -9379
rect -908 -9451 -862 -9413
rect -908 -9485 -902 -9451
rect -868 -9485 -862 -9451
rect -908 -9523 -862 -9485
rect -908 -9557 -902 -9523
rect -868 -9557 -862 -9523
rect -908 -9600 -862 -9557
rect -790 9557 -744 9600
rect -790 9523 -784 9557
rect -750 9523 -744 9557
rect -790 9485 -744 9523
rect -790 9451 -784 9485
rect -750 9451 -744 9485
rect -790 9413 -744 9451
rect -790 9379 -784 9413
rect -750 9379 -744 9413
rect -790 9341 -744 9379
rect -790 9307 -784 9341
rect -750 9307 -744 9341
rect -790 9269 -744 9307
rect -790 9235 -784 9269
rect -750 9235 -744 9269
rect -790 9197 -744 9235
rect -790 9163 -784 9197
rect -750 9163 -744 9197
rect -790 9125 -744 9163
rect -790 9091 -784 9125
rect -750 9091 -744 9125
rect -790 9053 -744 9091
rect -790 9019 -784 9053
rect -750 9019 -744 9053
rect -790 8981 -744 9019
rect -790 8947 -784 8981
rect -750 8947 -744 8981
rect -790 8909 -744 8947
rect -790 8875 -784 8909
rect -750 8875 -744 8909
rect -790 8837 -744 8875
rect -790 8803 -784 8837
rect -750 8803 -744 8837
rect -790 8765 -744 8803
rect -790 8731 -784 8765
rect -750 8731 -744 8765
rect -790 8693 -744 8731
rect -790 8659 -784 8693
rect -750 8659 -744 8693
rect -790 8621 -744 8659
rect -790 8587 -784 8621
rect -750 8587 -744 8621
rect -790 8549 -744 8587
rect -790 8515 -784 8549
rect -750 8515 -744 8549
rect -790 8477 -744 8515
rect -790 8443 -784 8477
rect -750 8443 -744 8477
rect -790 8405 -744 8443
rect -790 8371 -784 8405
rect -750 8371 -744 8405
rect -790 8333 -744 8371
rect -790 8299 -784 8333
rect -750 8299 -744 8333
rect -790 8261 -744 8299
rect -790 8227 -784 8261
rect -750 8227 -744 8261
rect -790 8189 -744 8227
rect -790 8155 -784 8189
rect -750 8155 -744 8189
rect -790 8117 -744 8155
rect -790 8083 -784 8117
rect -750 8083 -744 8117
rect -790 8045 -744 8083
rect -790 8011 -784 8045
rect -750 8011 -744 8045
rect -790 7973 -744 8011
rect -790 7939 -784 7973
rect -750 7939 -744 7973
rect -790 7901 -744 7939
rect -790 7867 -784 7901
rect -750 7867 -744 7901
rect -790 7829 -744 7867
rect -790 7795 -784 7829
rect -750 7795 -744 7829
rect -790 7757 -744 7795
rect -790 7723 -784 7757
rect -750 7723 -744 7757
rect -790 7685 -744 7723
rect -790 7651 -784 7685
rect -750 7651 -744 7685
rect -790 7613 -744 7651
rect -790 7579 -784 7613
rect -750 7579 -744 7613
rect -790 7541 -744 7579
rect -790 7507 -784 7541
rect -750 7507 -744 7541
rect -790 7469 -744 7507
rect -790 7435 -784 7469
rect -750 7435 -744 7469
rect -790 7397 -744 7435
rect -790 7363 -784 7397
rect -750 7363 -744 7397
rect -790 7325 -744 7363
rect -790 7291 -784 7325
rect -750 7291 -744 7325
rect -790 7253 -744 7291
rect -790 7219 -784 7253
rect -750 7219 -744 7253
rect -790 7181 -744 7219
rect -790 7147 -784 7181
rect -750 7147 -744 7181
rect -790 7109 -744 7147
rect -790 7075 -784 7109
rect -750 7075 -744 7109
rect -790 7037 -744 7075
rect -790 7003 -784 7037
rect -750 7003 -744 7037
rect -790 6965 -744 7003
rect -790 6931 -784 6965
rect -750 6931 -744 6965
rect -790 6893 -744 6931
rect -790 6859 -784 6893
rect -750 6859 -744 6893
rect -790 6821 -744 6859
rect -790 6787 -784 6821
rect -750 6787 -744 6821
rect -790 6749 -744 6787
rect -790 6715 -784 6749
rect -750 6715 -744 6749
rect -790 6677 -744 6715
rect -790 6643 -784 6677
rect -750 6643 -744 6677
rect -790 6605 -744 6643
rect -790 6571 -784 6605
rect -750 6571 -744 6605
rect -790 6533 -744 6571
rect -790 6499 -784 6533
rect -750 6499 -744 6533
rect -790 6461 -744 6499
rect -790 6427 -784 6461
rect -750 6427 -744 6461
rect -790 6389 -744 6427
rect -790 6355 -784 6389
rect -750 6355 -744 6389
rect -790 6317 -744 6355
rect -790 6283 -784 6317
rect -750 6283 -744 6317
rect -790 6245 -744 6283
rect -790 6211 -784 6245
rect -750 6211 -744 6245
rect -790 6173 -744 6211
rect -790 6139 -784 6173
rect -750 6139 -744 6173
rect -790 6101 -744 6139
rect -790 6067 -784 6101
rect -750 6067 -744 6101
rect -790 6029 -744 6067
rect -790 5995 -784 6029
rect -750 5995 -744 6029
rect -790 5957 -744 5995
rect -790 5923 -784 5957
rect -750 5923 -744 5957
rect -790 5885 -744 5923
rect -790 5851 -784 5885
rect -750 5851 -744 5885
rect -790 5813 -744 5851
rect -790 5779 -784 5813
rect -750 5779 -744 5813
rect -790 5741 -744 5779
rect -790 5707 -784 5741
rect -750 5707 -744 5741
rect -790 5669 -744 5707
rect -790 5635 -784 5669
rect -750 5635 -744 5669
rect -790 5597 -744 5635
rect -790 5563 -784 5597
rect -750 5563 -744 5597
rect -790 5525 -744 5563
rect -790 5491 -784 5525
rect -750 5491 -744 5525
rect -790 5453 -744 5491
rect -790 5419 -784 5453
rect -750 5419 -744 5453
rect -790 5381 -744 5419
rect -790 5347 -784 5381
rect -750 5347 -744 5381
rect -790 5309 -744 5347
rect -790 5275 -784 5309
rect -750 5275 -744 5309
rect -790 5237 -744 5275
rect -790 5203 -784 5237
rect -750 5203 -744 5237
rect -790 5165 -744 5203
rect -790 5131 -784 5165
rect -750 5131 -744 5165
rect -790 5093 -744 5131
rect -790 5059 -784 5093
rect -750 5059 -744 5093
rect -790 5021 -744 5059
rect -790 4987 -784 5021
rect -750 4987 -744 5021
rect -790 4949 -744 4987
rect -790 4915 -784 4949
rect -750 4915 -744 4949
rect -790 4877 -744 4915
rect -790 4843 -784 4877
rect -750 4843 -744 4877
rect -790 4805 -744 4843
rect -790 4771 -784 4805
rect -750 4771 -744 4805
rect -790 4733 -744 4771
rect -790 4699 -784 4733
rect -750 4699 -744 4733
rect -790 4661 -744 4699
rect -790 4627 -784 4661
rect -750 4627 -744 4661
rect -790 4589 -744 4627
rect -790 4555 -784 4589
rect -750 4555 -744 4589
rect -790 4517 -744 4555
rect -790 4483 -784 4517
rect -750 4483 -744 4517
rect -790 4445 -744 4483
rect -790 4411 -784 4445
rect -750 4411 -744 4445
rect -790 4373 -744 4411
rect -790 4339 -784 4373
rect -750 4339 -744 4373
rect -790 4301 -744 4339
rect -790 4267 -784 4301
rect -750 4267 -744 4301
rect -790 4229 -744 4267
rect -790 4195 -784 4229
rect -750 4195 -744 4229
rect -790 4157 -744 4195
rect -790 4123 -784 4157
rect -750 4123 -744 4157
rect -790 4085 -744 4123
rect -790 4051 -784 4085
rect -750 4051 -744 4085
rect -790 4013 -744 4051
rect -790 3979 -784 4013
rect -750 3979 -744 4013
rect -790 3941 -744 3979
rect -790 3907 -784 3941
rect -750 3907 -744 3941
rect -790 3869 -744 3907
rect -790 3835 -784 3869
rect -750 3835 -744 3869
rect -790 3797 -744 3835
rect -790 3763 -784 3797
rect -750 3763 -744 3797
rect -790 3725 -744 3763
rect -790 3691 -784 3725
rect -750 3691 -744 3725
rect -790 3653 -744 3691
rect -790 3619 -784 3653
rect -750 3619 -744 3653
rect -790 3581 -744 3619
rect -790 3547 -784 3581
rect -750 3547 -744 3581
rect -790 3509 -744 3547
rect -790 3475 -784 3509
rect -750 3475 -744 3509
rect -790 3437 -744 3475
rect -790 3403 -784 3437
rect -750 3403 -744 3437
rect -790 3365 -744 3403
rect -790 3331 -784 3365
rect -750 3331 -744 3365
rect -790 3293 -744 3331
rect -790 3259 -784 3293
rect -750 3259 -744 3293
rect -790 3221 -744 3259
rect -790 3187 -784 3221
rect -750 3187 -744 3221
rect -790 3149 -744 3187
rect -790 3115 -784 3149
rect -750 3115 -744 3149
rect -790 3077 -744 3115
rect -790 3043 -784 3077
rect -750 3043 -744 3077
rect -790 3005 -744 3043
rect -790 2971 -784 3005
rect -750 2971 -744 3005
rect -790 2933 -744 2971
rect -790 2899 -784 2933
rect -750 2899 -744 2933
rect -790 2861 -744 2899
rect -790 2827 -784 2861
rect -750 2827 -744 2861
rect -790 2789 -744 2827
rect -790 2755 -784 2789
rect -750 2755 -744 2789
rect -790 2717 -744 2755
rect -790 2683 -784 2717
rect -750 2683 -744 2717
rect -790 2645 -744 2683
rect -790 2611 -784 2645
rect -750 2611 -744 2645
rect -790 2573 -744 2611
rect -790 2539 -784 2573
rect -750 2539 -744 2573
rect -790 2501 -744 2539
rect -790 2467 -784 2501
rect -750 2467 -744 2501
rect -790 2429 -744 2467
rect -790 2395 -784 2429
rect -750 2395 -744 2429
rect -790 2357 -744 2395
rect -790 2323 -784 2357
rect -750 2323 -744 2357
rect -790 2285 -744 2323
rect -790 2251 -784 2285
rect -750 2251 -744 2285
rect -790 2213 -744 2251
rect -790 2179 -784 2213
rect -750 2179 -744 2213
rect -790 2141 -744 2179
rect -790 2107 -784 2141
rect -750 2107 -744 2141
rect -790 2069 -744 2107
rect -790 2035 -784 2069
rect -750 2035 -744 2069
rect -790 1997 -744 2035
rect -790 1963 -784 1997
rect -750 1963 -744 1997
rect -790 1925 -744 1963
rect -790 1891 -784 1925
rect -750 1891 -744 1925
rect -790 1853 -744 1891
rect -790 1819 -784 1853
rect -750 1819 -744 1853
rect -790 1781 -744 1819
rect -790 1747 -784 1781
rect -750 1747 -744 1781
rect -790 1709 -744 1747
rect -790 1675 -784 1709
rect -750 1675 -744 1709
rect -790 1637 -744 1675
rect -790 1603 -784 1637
rect -750 1603 -744 1637
rect -790 1565 -744 1603
rect -790 1531 -784 1565
rect -750 1531 -744 1565
rect -790 1493 -744 1531
rect -790 1459 -784 1493
rect -750 1459 -744 1493
rect -790 1421 -744 1459
rect -790 1387 -784 1421
rect -750 1387 -744 1421
rect -790 1349 -744 1387
rect -790 1315 -784 1349
rect -750 1315 -744 1349
rect -790 1277 -744 1315
rect -790 1243 -784 1277
rect -750 1243 -744 1277
rect -790 1205 -744 1243
rect -790 1171 -784 1205
rect -750 1171 -744 1205
rect -790 1133 -744 1171
rect -790 1099 -784 1133
rect -750 1099 -744 1133
rect -790 1061 -744 1099
rect -790 1027 -784 1061
rect -750 1027 -744 1061
rect -790 989 -744 1027
rect -790 955 -784 989
rect -750 955 -744 989
rect -790 917 -744 955
rect -790 883 -784 917
rect -750 883 -744 917
rect -790 845 -744 883
rect -790 811 -784 845
rect -750 811 -744 845
rect -790 773 -744 811
rect -790 739 -784 773
rect -750 739 -744 773
rect -790 701 -744 739
rect -790 667 -784 701
rect -750 667 -744 701
rect -790 629 -744 667
rect -790 595 -784 629
rect -750 595 -744 629
rect -790 557 -744 595
rect -790 523 -784 557
rect -750 523 -744 557
rect -790 485 -744 523
rect -790 451 -784 485
rect -750 451 -744 485
rect -790 413 -744 451
rect -790 379 -784 413
rect -750 379 -744 413
rect -790 341 -744 379
rect -790 307 -784 341
rect -750 307 -744 341
rect -790 269 -744 307
rect -790 235 -784 269
rect -750 235 -744 269
rect -790 197 -744 235
rect -790 163 -784 197
rect -750 163 -744 197
rect -790 125 -744 163
rect -790 91 -784 125
rect -750 91 -744 125
rect -790 53 -744 91
rect -790 19 -784 53
rect -750 19 -744 53
rect -790 -19 -744 19
rect -790 -53 -784 -19
rect -750 -53 -744 -19
rect -790 -91 -744 -53
rect -790 -125 -784 -91
rect -750 -125 -744 -91
rect -790 -163 -744 -125
rect -790 -197 -784 -163
rect -750 -197 -744 -163
rect -790 -235 -744 -197
rect -790 -269 -784 -235
rect -750 -269 -744 -235
rect -790 -307 -744 -269
rect -790 -341 -784 -307
rect -750 -341 -744 -307
rect -790 -379 -744 -341
rect -790 -413 -784 -379
rect -750 -413 -744 -379
rect -790 -451 -744 -413
rect -790 -485 -784 -451
rect -750 -485 -744 -451
rect -790 -523 -744 -485
rect -790 -557 -784 -523
rect -750 -557 -744 -523
rect -790 -595 -744 -557
rect -790 -629 -784 -595
rect -750 -629 -744 -595
rect -790 -667 -744 -629
rect -790 -701 -784 -667
rect -750 -701 -744 -667
rect -790 -739 -744 -701
rect -790 -773 -784 -739
rect -750 -773 -744 -739
rect -790 -811 -744 -773
rect -790 -845 -784 -811
rect -750 -845 -744 -811
rect -790 -883 -744 -845
rect -790 -917 -784 -883
rect -750 -917 -744 -883
rect -790 -955 -744 -917
rect -790 -989 -784 -955
rect -750 -989 -744 -955
rect -790 -1027 -744 -989
rect -790 -1061 -784 -1027
rect -750 -1061 -744 -1027
rect -790 -1099 -744 -1061
rect -790 -1133 -784 -1099
rect -750 -1133 -744 -1099
rect -790 -1171 -744 -1133
rect -790 -1205 -784 -1171
rect -750 -1205 -744 -1171
rect -790 -1243 -744 -1205
rect -790 -1277 -784 -1243
rect -750 -1277 -744 -1243
rect -790 -1315 -744 -1277
rect -790 -1349 -784 -1315
rect -750 -1349 -744 -1315
rect -790 -1387 -744 -1349
rect -790 -1421 -784 -1387
rect -750 -1421 -744 -1387
rect -790 -1459 -744 -1421
rect -790 -1493 -784 -1459
rect -750 -1493 -744 -1459
rect -790 -1531 -744 -1493
rect -790 -1565 -784 -1531
rect -750 -1565 -744 -1531
rect -790 -1603 -744 -1565
rect -790 -1637 -784 -1603
rect -750 -1637 -744 -1603
rect -790 -1675 -744 -1637
rect -790 -1709 -784 -1675
rect -750 -1709 -744 -1675
rect -790 -1747 -744 -1709
rect -790 -1781 -784 -1747
rect -750 -1781 -744 -1747
rect -790 -1819 -744 -1781
rect -790 -1853 -784 -1819
rect -750 -1853 -744 -1819
rect -790 -1891 -744 -1853
rect -790 -1925 -784 -1891
rect -750 -1925 -744 -1891
rect -790 -1963 -744 -1925
rect -790 -1997 -784 -1963
rect -750 -1997 -744 -1963
rect -790 -2035 -744 -1997
rect -790 -2069 -784 -2035
rect -750 -2069 -744 -2035
rect -790 -2107 -744 -2069
rect -790 -2141 -784 -2107
rect -750 -2141 -744 -2107
rect -790 -2179 -744 -2141
rect -790 -2213 -784 -2179
rect -750 -2213 -744 -2179
rect -790 -2251 -744 -2213
rect -790 -2285 -784 -2251
rect -750 -2285 -744 -2251
rect -790 -2323 -744 -2285
rect -790 -2357 -784 -2323
rect -750 -2357 -744 -2323
rect -790 -2395 -744 -2357
rect -790 -2429 -784 -2395
rect -750 -2429 -744 -2395
rect -790 -2467 -744 -2429
rect -790 -2501 -784 -2467
rect -750 -2501 -744 -2467
rect -790 -2539 -744 -2501
rect -790 -2573 -784 -2539
rect -750 -2573 -744 -2539
rect -790 -2611 -744 -2573
rect -790 -2645 -784 -2611
rect -750 -2645 -744 -2611
rect -790 -2683 -744 -2645
rect -790 -2717 -784 -2683
rect -750 -2717 -744 -2683
rect -790 -2755 -744 -2717
rect -790 -2789 -784 -2755
rect -750 -2789 -744 -2755
rect -790 -2827 -744 -2789
rect -790 -2861 -784 -2827
rect -750 -2861 -744 -2827
rect -790 -2899 -744 -2861
rect -790 -2933 -784 -2899
rect -750 -2933 -744 -2899
rect -790 -2971 -744 -2933
rect -790 -3005 -784 -2971
rect -750 -3005 -744 -2971
rect -790 -3043 -744 -3005
rect -790 -3077 -784 -3043
rect -750 -3077 -744 -3043
rect -790 -3115 -744 -3077
rect -790 -3149 -784 -3115
rect -750 -3149 -744 -3115
rect -790 -3187 -744 -3149
rect -790 -3221 -784 -3187
rect -750 -3221 -744 -3187
rect -790 -3259 -744 -3221
rect -790 -3293 -784 -3259
rect -750 -3293 -744 -3259
rect -790 -3331 -744 -3293
rect -790 -3365 -784 -3331
rect -750 -3365 -744 -3331
rect -790 -3403 -744 -3365
rect -790 -3437 -784 -3403
rect -750 -3437 -744 -3403
rect -790 -3475 -744 -3437
rect -790 -3509 -784 -3475
rect -750 -3509 -744 -3475
rect -790 -3547 -744 -3509
rect -790 -3581 -784 -3547
rect -750 -3581 -744 -3547
rect -790 -3619 -744 -3581
rect -790 -3653 -784 -3619
rect -750 -3653 -744 -3619
rect -790 -3691 -744 -3653
rect -790 -3725 -784 -3691
rect -750 -3725 -744 -3691
rect -790 -3763 -744 -3725
rect -790 -3797 -784 -3763
rect -750 -3797 -744 -3763
rect -790 -3835 -744 -3797
rect -790 -3869 -784 -3835
rect -750 -3869 -744 -3835
rect -790 -3907 -744 -3869
rect -790 -3941 -784 -3907
rect -750 -3941 -744 -3907
rect -790 -3979 -744 -3941
rect -790 -4013 -784 -3979
rect -750 -4013 -744 -3979
rect -790 -4051 -744 -4013
rect -790 -4085 -784 -4051
rect -750 -4085 -744 -4051
rect -790 -4123 -744 -4085
rect -790 -4157 -784 -4123
rect -750 -4157 -744 -4123
rect -790 -4195 -744 -4157
rect -790 -4229 -784 -4195
rect -750 -4229 -744 -4195
rect -790 -4267 -744 -4229
rect -790 -4301 -784 -4267
rect -750 -4301 -744 -4267
rect -790 -4339 -744 -4301
rect -790 -4373 -784 -4339
rect -750 -4373 -744 -4339
rect -790 -4411 -744 -4373
rect -790 -4445 -784 -4411
rect -750 -4445 -744 -4411
rect -790 -4483 -744 -4445
rect -790 -4517 -784 -4483
rect -750 -4517 -744 -4483
rect -790 -4555 -744 -4517
rect -790 -4589 -784 -4555
rect -750 -4589 -744 -4555
rect -790 -4627 -744 -4589
rect -790 -4661 -784 -4627
rect -750 -4661 -744 -4627
rect -790 -4699 -744 -4661
rect -790 -4733 -784 -4699
rect -750 -4733 -744 -4699
rect -790 -4771 -744 -4733
rect -790 -4805 -784 -4771
rect -750 -4805 -744 -4771
rect -790 -4843 -744 -4805
rect -790 -4877 -784 -4843
rect -750 -4877 -744 -4843
rect -790 -4915 -744 -4877
rect -790 -4949 -784 -4915
rect -750 -4949 -744 -4915
rect -790 -4987 -744 -4949
rect -790 -5021 -784 -4987
rect -750 -5021 -744 -4987
rect -790 -5059 -744 -5021
rect -790 -5093 -784 -5059
rect -750 -5093 -744 -5059
rect -790 -5131 -744 -5093
rect -790 -5165 -784 -5131
rect -750 -5165 -744 -5131
rect -790 -5203 -744 -5165
rect -790 -5237 -784 -5203
rect -750 -5237 -744 -5203
rect -790 -5275 -744 -5237
rect -790 -5309 -784 -5275
rect -750 -5309 -744 -5275
rect -790 -5347 -744 -5309
rect -790 -5381 -784 -5347
rect -750 -5381 -744 -5347
rect -790 -5419 -744 -5381
rect -790 -5453 -784 -5419
rect -750 -5453 -744 -5419
rect -790 -5491 -744 -5453
rect -790 -5525 -784 -5491
rect -750 -5525 -744 -5491
rect -790 -5563 -744 -5525
rect -790 -5597 -784 -5563
rect -750 -5597 -744 -5563
rect -790 -5635 -744 -5597
rect -790 -5669 -784 -5635
rect -750 -5669 -744 -5635
rect -790 -5707 -744 -5669
rect -790 -5741 -784 -5707
rect -750 -5741 -744 -5707
rect -790 -5779 -744 -5741
rect -790 -5813 -784 -5779
rect -750 -5813 -744 -5779
rect -790 -5851 -744 -5813
rect -790 -5885 -784 -5851
rect -750 -5885 -744 -5851
rect -790 -5923 -744 -5885
rect -790 -5957 -784 -5923
rect -750 -5957 -744 -5923
rect -790 -5995 -744 -5957
rect -790 -6029 -784 -5995
rect -750 -6029 -744 -5995
rect -790 -6067 -744 -6029
rect -790 -6101 -784 -6067
rect -750 -6101 -744 -6067
rect -790 -6139 -744 -6101
rect -790 -6173 -784 -6139
rect -750 -6173 -744 -6139
rect -790 -6211 -744 -6173
rect -790 -6245 -784 -6211
rect -750 -6245 -744 -6211
rect -790 -6283 -744 -6245
rect -790 -6317 -784 -6283
rect -750 -6317 -744 -6283
rect -790 -6355 -744 -6317
rect -790 -6389 -784 -6355
rect -750 -6389 -744 -6355
rect -790 -6427 -744 -6389
rect -790 -6461 -784 -6427
rect -750 -6461 -744 -6427
rect -790 -6499 -744 -6461
rect -790 -6533 -784 -6499
rect -750 -6533 -744 -6499
rect -790 -6571 -744 -6533
rect -790 -6605 -784 -6571
rect -750 -6605 -744 -6571
rect -790 -6643 -744 -6605
rect -790 -6677 -784 -6643
rect -750 -6677 -744 -6643
rect -790 -6715 -744 -6677
rect -790 -6749 -784 -6715
rect -750 -6749 -744 -6715
rect -790 -6787 -744 -6749
rect -790 -6821 -784 -6787
rect -750 -6821 -744 -6787
rect -790 -6859 -744 -6821
rect -790 -6893 -784 -6859
rect -750 -6893 -744 -6859
rect -790 -6931 -744 -6893
rect -790 -6965 -784 -6931
rect -750 -6965 -744 -6931
rect -790 -7003 -744 -6965
rect -790 -7037 -784 -7003
rect -750 -7037 -744 -7003
rect -790 -7075 -744 -7037
rect -790 -7109 -784 -7075
rect -750 -7109 -744 -7075
rect -790 -7147 -744 -7109
rect -790 -7181 -784 -7147
rect -750 -7181 -744 -7147
rect -790 -7219 -744 -7181
rect -790 -7253 -784 -7219
rect -750 -7253 -744 -7219
rect -790 -7291 -744 -7253
rect -790 -7325 -784 -7291
rect -750 -7325 -744 -7291
rect -790 -7363 -744 -7325
rect -790 -7397 -784 -7363
rect -750 -7397 -744 -7363
rect -790 -7435 -744 -7397
rect -790 -7469 -784 -7435
rect -750 -7469 -744 -7435
rect -790 -7507 -744 -7469
rect -790 -7541 -784 -7507
rect -750 -7541 -744 -7507
rect -790 -7579 -744 -7541
rect -790 -7613 -784 -7579
rect -750 -7613 -744 -7579
rect -790 -7651 -744 -7613
rect -790 -7685 -784 -7651
rect -750 -7685 -744 -7651
rect -790 -7723 -744 -7685
rect -790 -7757 -784 -7723
rect -750 -7757 -744 -7723
rect -790 -7795 -744 -7757
rect -790 -7829 -784 -7795
rect -750 -7829 -744 -7795
rect -790 -7867 -744 -7829
rect -790 -7901 -784 -7867
rect -750 -7901 -744 -7867
rect -790 -7939 -744 -7901
rect -790 -7973 -784 -7939
rect -750 -7973 -744 -7939
rect -790 -8011 -744 -7973
rect -790 -8045 -784 -8011
rect -750 -8045 -744 -8011
rect -790 -8083 -744 -8045
rect -790 -8117 -784 -8083
rect -750 -8117 -744 -8083
rect -790 -8155 -744 -8117
rect -790 -8189 -784 -8155
rect -750 -8189 -744 -8155
rect -790 -8227 -744 -8189
rect -790 -8261 -784 -8227
rect -750 -8261 -744 -8227
rect -790 -8299 -744 -8261
rect -790 -8333 -784 -8299
rect -750 -8333 -744 -8299
rect -790 -8371 -744 -8333
rect -790 -8405 -784 -8371
rect -750 -8405 -744 -8371
rect -790 -8443 -744 -8405
rect -790 -8477 -784 -8443
rect -750 -8477 -744 -8443
rect -790 -8515 -744 -8477
rect -790 -8549 -784 -8515
rect -750 -8549 -744 -8515
rect -790 -8587 -744 -8549
rect -790 -8621 -784 -8587
rect -750 -8621 -744 -8587
rect -790 -8659 -744 -8621
rect -790 -8693 -784 -8659
rect -750 -8693 -744 -8659
rect -790 -8731 -744 -8693
rect -790 -8765 -784 -8731
rect -750 -8765 -744 -8731
rect -790 -8803 -744 -8765
rect -790 -8837 -784 -8803
rect -750 -8837 -744 -8803
rect -790 -8875 -744 -8837
rect -790 -8909 -784 -8875
rect -750 -8909 -744 -8875
rect -790 -8947 -744 -8909
rect -790 -8981 -784 -8947
rect -750 -8981 -744 -8947
rect -790 -9019 -744 -8981
rect -790 -9053 -784 -9019
rect -750 -9053 -744 -9019
rect -790 -9091 -744 -9053
rect -790 -9125 -784 -9091
rect -750 -9125 -744 -9091
rect -790 -9163 -744 -9125
rect -790 -9197 -784 -9163
rect -750 -9197 -744 -9163
rect -790 -9235 -744 -9197
rect -790 -9269 -784 -9235
rect -750 -9269 -744 -9235
rect -790 -9307 -744 -9269
rect -790 -9341 -784 -9307
rect -750 -9341 -744 -9307
rect -790 -9379 -744 -9341
rect -790 -9413 -784 -9379
rect -750 -9413 -744 -9379
rect -790 -9451 -744 -9413
rect -790 -9485 -784 -9451
rect -750 -9485 -744 -9451
rect -790 -9523 -744 -9485
rect -790 -9557 -784 -9523
rect -750 -9557 -744 -9523
rect -790 -9600 -744 -9557
rect -672 9557 -626 9600
rect -672 9523 -666 9557
rect -632 9523 -626 9557
rect -672 9485 -626 9523
rect -672 9451 -666 9485
rect -632 9451 -626 9485
rect -672 9413 -626 9451
rect -672 9379 -666 9413
rect -632 9379 -626 9413
rect -672 9341 -626 9379
rect -672 9307 -666 9341
rect -632 9307 -626 9341
rect -672 9269 -626 9307
rect -672 9235 -666 9269
rect -632 9235 -626 9269
rect -672 9197 -626 9235
rect -672 9163 -666 9197
rect -632 9163 -626 9197
rect -672 9125 -626 9163
rect -672 9091 -666 9125
rect -632 9091 -626 9125
rect -672 9053 -626 9091
rect -672 9019 -666 9053
rect -632 9019 -626 9053
rect -672 8981 -626 9019
rect -672 8947 -666 8981
rect -632 8947 -626 8981
rect -672 8909 -626 8947
rect -672 8875 -666 8909
rect -632 8875 -626 8909
rect -672 8837 -626 8875
rect -672 8803 -666 8837
rect -632 8803 -626 8837
rect -672 8765 -626 8803
rect -672 8731 -666 8765
rect -632 8731 -626 8765
rect -672 8693 -626 8731
rect -672 8659 -666 8693
rect -632 8659 -626 8693
rect -672 8621 -626 8659
rect -672 8587 -666 8621
rect -632 8587 -626 8621
rect -672 8549 -626 8587
rect -672 8515 -666 8549
rect -632 8515 -626 8549
rect -672 8477 -626 8515
rect -672 8443 -666 8477
rect -632 8443 -626 8477
rect -672 8405 -626 8443
rect -672 8371 -666 8405
rect -632 8371 -626 8405
rect -672 8333 -626 8371
rect -672 8299 -666 8333
rect -632 8299 -626 8333
rect -672 8261 -626 8299
rect -672 8227 -666 8261
rect -632 8227 -626 8261
rect -672 8189 -626 8227
rect -672 8155 -666 8189
rect -632 8155 -626 8189
rect -672 8117 -626 8155
rect -672 8083 -666 8117
rect -632 8083 -626 8117
rect -672 8045 -626 8083
rect -672 8011 -666 8045
rect -632 8011 -626 8045
rect -672 7973 -626 8011
rect -672 7939 -666 7973
rect -632 7939 -626 7973
rect -672 7901 -626 7939
rect -672 7867 -666 7901
rect -632 7867 -626 7901
rect -672 7829 -626 7867
rect -672 7795 -666 7829
rect -632 7795 -626 7829
rect -672 7757 -626 7795
rect -672 7723 -666 7757
rect -632 7723 -626 7757
rect -672 7685 -626 7723
rect -672 7651 -666 7685
rect -632 7651 -626 7685
rect -672 7613 -626 7651
rect -672 7579 -666 7613
rect -632 7579 -626 7613
rect -672 7541 -626 7579
rect -672 7507 -666 7541
rect -632 7507 -626 7541
rect -672 7469 -626 7507
rect -672 7435 -666 7469
rect -632 7435 -626 7469
rect -672 7397 -626 7435
rect -672 7363 -666 7397
rect -632 7363 -626 7397
rect -672 7325 -626 7363
rect -672 7291 -666 7325
rect -632 7291 -626 7325
rect -672 7253 -626 7291
rect -672 7219 -666 7253
rect -632 7219 -626 7253
rect -672 7181 -626 7219
rect -672 7147 -666 7181
rect -632 7147 -626 7181
rect -672 7109 -626 7147
rect -672 7075 -666 7109
rect -632 7075 -626 7109
rect -672 7037 -626 7075
rect -672 7003 -666 7037
rect -632 7003 -626 7037
rect -672 6965 -626 7003
rect -672 6931 -666 6965
rect -632 6931 -626 6965
rect -672 6893 -626 6931
rect -672 6859 -666 6893
rect -632 6859 -626 6893
rect -672 6821 -626 6859
rect -672 6787 -666 6821
rect -632 6787 -626 6821
rect -672 6749 -626 6787
rect -672 6715 -666 6749
rect -632 6715 -626 6749
rect -672 6677 -626 6715
rect -672 6643 -666 6677
rect -632 6643 -626 6677
rect -672 6605 -626 6643
rect -672 6571 -666 6605
rect -632 6571 -626 6605
rect -672 6533 -626 6571
rect -672 6499 -666 6533
rect -632 6499 -626 6533
rect -672 6461 -626 6499
rect -672 6427 -666 6461
rect -632 6427 -626 6461
rect -672 6389 -626 6427
rect -672 6355 -666 6389
rect -632 6355 -626 6389
rect -672 6317 -626 6355
rect -672 6283 -666 6317
rect -632 6283 -626 6317
rect -672 6245 -626 6283
rect -672 6211 -666 6245
rect -632 6211 -626 6245
rect -672 6173 -626 6211
rect -672 6139 -666 6173
rect -632 6139 -626 6173
rect -672 6101 -626 6139
rect -672 6067 -666 6101
rect -632 6067 -626 6101
rect -672 6029 -626 6067
rect -672 5995 -666 6029
rect -632 5995 -626 6029
rect -672 5957 -626 5995
rect -672 5923 -666 5957
rect -632 5923 -626 5957
rect -672 5885 -626 5923
rect -672 5851 -666 5885
rect -632 5851 -626 5885
rect -672 5813 -626 5851
rect -672 5779 -666 5813
rect -632 5779 -626 5813
rect -672 5741 -626 5779
rect -672 5707 -666 5741
rect -632 5707 -626 5741
rect -672 5669 -626 5707
rect -672 5635 -666 5669
rect -632 5635 -626 5669
rect -672 5597 -626 5635
rect -672 5563 -666 5597
rect -632 5563 -626 5597
rect -672 5525 -626 5563
rect -672 5491 -666 5525
rect -632 5491 -626 5525
rect -672 5453 -626 5491
rect -672 5419 -666 5453
rect -632 5419 -626 5453
rect -672 5381 -626 5419
rect -672 5347 -666 5381
rect -632 5347 -626 5381
rect -672 5309 -626 5347
rect -672 5275 -666 5309
rect -632 5275 -626 5309
rect -672 5237 -626 5275
rect -672 5203 -666 5237
rect -632 5203 -626 5237
rect -672 5165 -626 5203
rect -672 5131 -666 5165
rect -632 5131 -626 5165
rect -672 5093 -626 5131
rect -672 5059 -666 5093
rect -632 5059 -626 5093
rect -672 5021 -626 5059
rect -672 4987 -666 5021
rect -632 4987 -626 5021
rect -672 4949 -626 4987
rect -672 4915 -666 4949
rect -632 4915 -626 4949
rect -672 4877 -626 4915
rect -672 4843 -666 4877
rect -632 4843 -626 4877
rect -672 4805 -626 4843
rect -672 4771 -666 4805
rect -632 4771 -626 4805
rect -672 4733 -626 4771
rect -672 4699 -666 4733
rect -632 4699 -626 4733
rect -672 4661 -626 4699
rect -672 4627 -666 4661
rect -632 4627 -626 4661
rect -672 4589 -626 4627
rect -672 4555 -666 4589
rect -632 4555 -626 4589
rect -672 4517 -626 4555
rect -672 4483 -666 4517
rect -632 4483 -626 4517
rect -672 4445 -626 4483
rect -672 4411 -666 4445
rect -632 4411 -626 4445
rect -672 4373 -626 4411
rect -672 4339 -666 4373
rect -632 4339 -626 4373
rect -672 4301 -626 4339
rect -672 4267 -666 4301
rect -632 4267 -626 4301
rect -672 4229 -626 4267
rect -672 4195 -666 4229
rect -632 4195 -626 4229
rect -672 4157 -626 4195
rect -672 4123 -666 4157
rect -632 4123 -626 4157
rect -672 4085 -626 4123
rect -672 4051 -666 4085
rect -632 4051 -626 4085
rect -672 4013 -626 4051
rect -672 3979 -666 4013
rect -632 3979 -626 4013
rect -672 3941 -626 3979
rect -672 3907 -666 3941
rect -632 3907 -626 3941
rect -672 3869 -626 3907
rect -672 3835 -666 3869
rect -632 3835 -626 3869
rect -672 3797 -626 3835
rect -672 3763 -666 3797
rect -632 3763 -626 3797
rect -672 3725 -626 3763
rect -672 3691 -666 3725
rect -632 3691 -626 3725
rect -672 3653 -626 3691
rect -672 3619 -666 3653
rect -632 3619 -626 3653
rect -672 3581 -626 3619
rect -672 3547 -666 3581
rect -632 3547 -626 3581
rect -672 3509 -626 3547
rect -672 3475 -666 3509
rect -632 3475 -626 3509
rect -672 3437 -626 3475
rect -672 3403 -666 3437
rect -632 3403 -626 3437
rect -672 3365 -626 3403
rect -672 3331 -666 3365
rect -632 3331 -626 3365
rect -672 3293 -626 3331
rect -672 3259 -666 3293
rect -632 3259 -626 3293
rect -672 3221 -626 3259
rect -672 3187 -666 3221
rect -632 3187 -626 3221
rect -672 3149 -626 3187
rect -672 3115 -666 3149
rect -632 3115 -626 3149
rect -672 3077 -626 3115
rect -672 3043 -666 3077
rect -632 3043 -626 3077
rect -672 3005 -626 3043
rect -672 2971 -666 3005
rect -632 2971 -626 3005
rect -672 2933 -626 2971
rect -672 2899 -666 2933
rect -632 2899 -626 2933
rect -672 2861 -626 2899
rect -672 2827 -666 2861
rect -632 2827 -626 2861
rect -672 2789 -626 2827
rect -672 2755 -666 2789
rect -632 2755 -626 2789
rect -672 2717 -626 2755
rect -672 2683 -666 2717
rect -632 2683 -626 2717
rect -672 2645 -626 2683
rect -672 2611 -666 2645
rect -632 2611 -626 2645
rect -672 2573 -626 2611
rect -672 2539 -666 2573
rect -632 2539 -626 2573
rect -672 2501 -626 2539
rect -672 2467 -666 2501
rect -632 2467 -626 2501
rect -672 2429 -626 2467
rect -672 2395 -666 2429
rect -632 2395 -626 2429
rect -672 2357 -626 2395
rect -672 2323 -666 2357
rect -632 2323 -626 2357
rect -672 2285 -626 2323
rect -672 2251 -666 2285
rect -632 2251 -626 2285
rect -672 2213 -626 2251
rect -672 2179 -666 2213
rect -632 2179 -626 2213
rect -672 2141 -626 2179
rect -672 2107 -666 2141
rect -632 2107 -626 2141
rect -672 2069 -626 2107
rect -672 2035 -666 2069
rect -632 2035 -626 2069
rect -672 1997 -626 2035
rect -672 1963 -666 1997
rect -632 1963 -626 1997
rect -672 1925 -626 1963
rect -672 1891 -666 1925
rect -632 1891 -626 1925
rect -672 1853 -626 1891
rect -672 1819 -666 1853
rect -632 1819 -626 1853
rect -672 1781 -626 1819
rect -672 1747 -666 1781
rect -632 1747 -626 1781
rect -672 1709 -626 1747
rect -672 1675 -666 1709
rect -632 1675 -626 1709
rect -672 1637 -626 1675
rect -672 1603 -666 1637
rect -632 1603 -626 1637
rect -672 1565 -626 1603
rect -672 1531 -666 1565
rect -632 1531 -626 1565
rect -672 1493 -626 1531
rect -672 1459 -666 1493
rect -632 1459 -626 1493
rect -672 1421 -626 1459
rect -672 1387 -666 1421
rect -632 1387 -626 1421
rect -672 1349 -626 1387
rect -672 1315 -666 1349
rect -632 1315 -626 1349
rect -672 1277 -626 1315
rect -672 1243 -666 1277
rect -632 1243 -626 1277
rect -672 1205 -626 1243
rect -672 1171 -666 1205
rect -632 1171 -626 1205
rect -672 1133 -626 1171
rect -672 1099 -666 1133
rect -632 1099 -626 1133
rect -672 1061 -626 1099
rect -672 1027 -666 1061
rect -632 1027 -626 1061
rect -672 989 -626 1027
rect -672 955 -666 989
rect -632 955 -626 989
rect -672 917 -626 955
rect -672 883 -666 917
rect -632 883 -626 917
rect -672 845 -626 883
rect -672 811 -666 845
rect -632 811 -626 845
rect -672 773 -626 811
rect -672 739 -666 773
rect -632 739 -626 773
rect -672 701 -626 739
rect -672 667 -666 701
rect -632 667 -626 701
rect -672 629 -626 667
rect -672 595 -666 629
rect -632 595 -626 629
rect -672 557 -626 595
rect -672 523 -666 557
rect -632 523 -626 557
rect -672 485 -626 523
rect -672 451 -666 485
rect -632 451 -626 485
rect -672 413 -626 451
rect -672 379 -666 413
rect -632 379 -626 413
rect -672 341 -626 379
rect -672 307 -666 341
rect -632 307 -626 341
rect -672 269 -626 307
rect -672 235 -666 269
rect -632 235 -626 269
rect -672 197 -626 235
rect -672 163 -666 197
rect -632 163 -626 197
rect -672 125 -626 163
rect -672 91 -666 125
rect -632 91 -626 125
rect -672 53 -626 91
rect -672 19 -666 53
rect -632 19 -626 53
rect -672 -19 -626 19
rect -672 -53 -666 -19
rect -632 -53 -626 -19
rect -672 -91 -626 -53
rect -672 -125 -666 -91
rect -632 -125 -626 -91
rect -672 -163 -626 -125
rect -672 -197 -666 -163
rect -632 -197 -626 -163
rect -672 -235 -626 -197
rect -672 -269 -666 -235
rect -632 -269 -626 -235
rect -672 -307 -626 -269
rect -672 -341 -666 -307
rect -632 -341 -626 -307
rect -672 -379 -626 -341
rect -672 -413 -666 -379
rect -632 -413 -626 -379
rect -672 -451 -626 -413
rect -672 -485 -666 -451
rect -632 -485 -626 -451
rect -672 -523 -626 -485
rect -672 -557 -666 -523
rect -632 -557 -626 -523
rect -672 -595 -626 -557
rect -672 -629 -666 -595
rect -632 -629 -626 -595
rect -672 -667 -626 -629
rect -672 -701 -666 -667
rect -632 -701 -626 -667
rect -672 -739 -626 -701
rect -672 -773 -666 -739
rect -632 -773 -626 -739
rect -672 -811 -626 -773
rect -672 -845 -666 -811
rect -632 -845 -626 -811
rect -672 -883 -626 -845
rect -672 -917 -666 -883
rect -632 -917 -626 -883
rect -672 -955 -626 -917
rect -672 -989 -666 -955
rect -632 -989 -626 -955
rect -672 -1027 -626 -989
rect -672 -1061 -666 -1027
rect -632 -1061 -626 -1027
rect -672 -1099 -626 -1061
rect -672 -1133 -666 -1099
rect -632 -1133 -626 -1099
rect -672 -1171 -626 -1133
rect -672 -1205 -666 -1171
rect -632 -1205 -626 -1171
rect -672 -1243 -626 -1205
rect -672 -1277 -666 -1243
rect -632 -1277 -626 -1243
rect -672 -1315 -626 -1277
rect -672 -1349 -666 -1315
rect -632 -1349 -626 -1315
rect -672 -1387 -626 -1349
rect -672 -1421 -666 -1387
rect -632 -1421 -626 -1387
rect -672 -1459 -626 -1421
rect -672 -1493 -666 -1459
rect -632 -1493 -626 -1459
rect -672 -1531 -626 -1493
rect -672 -1565 -666 -1531
rect -632 -1565 -626 -1531
rect -672 -1603 -626 -1565
rect -672 -1637 -666 -1603
rect -632 -1637 -626 -1603
rect -672 -1675 -626 -1637
rect -672 -1709 -666 -1675
rect -632 -1709 -626 -1675
rect -672 -1747 -626 -1709
rect -672 -1781 -666 -1747
rect -632 -1781 -626 -1747
rect -672 -1819 -626 -1781
rect -672 -1853 -666 -1819
rect -632 -1853 -626 -1819
rect -672 -1891 -626 -1853
rect -672 -1925 -666 -1891
rect -632 -1925 -626 -1891
rect -672 -1963 -626 -1925
rect -672 -1997 -666 -1963
rect -632 -1997 -626 -1963
rect -672 -2035 -626 -1997
rect -672 -2069 -666 -2035
rect -632 -2069 -626 -2035
rect -672 -2107 -626 -2069
rect -672 -2141 -666 -2107
rect -632 -2141 -626 -2107
rect -672 -2179 -626 -2141
rect -672 -2213 -666 -2179
rect -632 -2213 -626 -2179
rect -672 -2251 -626 -2213
rect -672 -2285 -666 -2251
rect -632 -2285 -626 -2251
rect -672 -2323 -626 -2285
rect -672 -2357 -666 -2323
rect -632 -2357 -626 -2323
rect -672 -2395 -626 -2357
rect -672 -2429 -666 -2395
rect -632 -2429 -626 -2395
rect -672 -2467 -626 -2429
rect -672 -2501 -666 -2467
rect -632 -2501 -626 -2467
rect -672 -2539 -626 -2501
rect -672 -2573 -666 -2539
rect -632 -2573 -626 -2539
rect -672 -2611 -626 -2573
rect -672 -2645 -666 -2611
rect -632 -2645 -626 -2611
rect -672 -2683 -626 -2645
rect -672 -2717 -666 -2683
rect -632 -2717 -626 -2683
rect -672 -2755 -626 -2717
rect -672 -2789 -666 -2755
rect -632 -2789 -626 -2755
rect -672 -2827 -626 -2789
rect -672 -2861 -666 -2827
rect -632 -2861 -626 -2827
rect -672 -2899 -626 -2861
rect -672 -2933 -666 -2899
rect -632 -2933 -626 -2899
rect -672 -2971 -626 -2933
rect -672 -3005 -666 -2971
rect -632 -3005 -626 -2971
rect -672 -3043 -626 -3005
rect -672 -3077 -666 -3043
rect -632 -3077 -626 -3043
rect -672 -3115 -626 -3077
rect -672 -3149 -666 -3115
rect -632 -3149 -626 -3115
rect -672 -3187 -626 -3149
rect -672 -3221 -666 -3187
rect -632 -3221 -626 -3187
rect -672 -3259 -626 -3221
rect -672 -3293 -666 -3259
rect -632 -3293 -626 -3259
rect -672 -3331 -626 -3293
rect -672 -3365 -666 -3331
rect -632 -3365 -626 -3331
rect -672 -3403 -626 -3365
rect -672 -3437 -666 -3403
rect -632 -3437 -626 -3403
rect -672 -3475 -626 -3437
rect -672 -3509 -666 -3475
rect -632 -3509 -626 -3475
rect -672 -3547 -626 -3509
rect -672 -3581 -666 -3547
rect -632 -3581 -626 -3547
rect -672 -3619 -626 -3581
rect -672 -3653 -666 -3619
rect -632 -3653 -626 -3619
rect -672 -3691 -626 -3653
rect -672 -3725 -666 -3691
rect -632 -3725 -626 -3691
rect -672 -3763 -626 -3725
rect -672 -3797 -666 -3763
rect -632 -3797 -626 -3763
rect -672 -3835 -626 -3797
rect -672 -3869 -666 -3835
rect -632 -3869 -626 -3835
rect -672 -3907 -626 -3869
rect -672 -3941 -666 -3907
rect -632 -3941 -626 -3907
rect -672 -3979 -626 -3941
rect -672 -4013 -666 -3979
rect -632 -4013 -626 -3979
rect -672 -4051 -626 -4013
rect -672 -4085 -666 -4051
rect -632 -4085 -626 -4051
rect -672 -4123 -626 -4085
rect -672 -4157 -666 -4123
rect -632 -4157 -626 -4123
rect -672 -4195 -626 -4157
rect -672 -4229 -666 -4195
rect -632 -4229 -626 -4195
rect -672 -4267 -626 -4229
rect -672 -4301 -666 -4267
rect -632 -4301 -626 -4267
rect -672 -4339 -626 -4301
rect -672 -4373 -666 -4339
rect -632 -4373 -626 -4339
rect -672 -4411 -626 -4373
rect -672 -4445 -666 -4411
rect -632 -4445 -626 -4411
rect -672 -4483 -626 -4445
rect -672 -4517 -666 -4483
rect -632 -4517 -626 -4483
rect -672 -4555 -626 -4517
rect -672 -4589 -666 -4555
rect -632 -4589 -626 -4555
rect -672 -4627 -626 -4589
rect -672 -4661 -666 -4627
rect -632 -4661 -626 -4627
rect -672 -4699 -626 -4661
rect -672 -4733 -666 -4699
rect -632 -4733 -626 -4699
rect -672 -4771 -626 -4733
rect -672 -4805 -666 -4771
rect -632 -4805 -626 -4771
rect -672 -4843 -626 -4805
rect -672 -4877 -666 -4843
rect -632 -4877 -626 -4843
rect -672 -4915 -626 -4877
rect -672 -4949 -666 -4915
rect -632 -4949 -626 -4915
rect -672 -4987 -626 -4949
rect -672 -5021 -666 -4987
rect -632 -5021 -626 -4987
rect -672 -5059 -626 -5021
rect -672 -5093 -666 -5059
rect -632 -5093 -626 -5059
rect -672 -5131 -626 -5093
rect -672 -5165 -666 -5131
rect -632 -5165 -626 -5131
rect -672 -5203 -626 -5165
rect -672 -5237 -666 -5203
rect -632 -5237 -626 -5203
rect -672 -5275 -626 -5237
rect -672 -5309 -666 -5275
rect -632 -5309 -626 -5275
rect -672 -5347 -626 -5309
rect -672 -5381 -666 -5347
rect -632 -5381 -626 -5347
rect -672 -5419 -626 -5381
rect -672 -5453 -666 -5419
rect -632 -5453 -626 -5419
rect -672 -5491 -626 -5453
rect -672 -5525 -666 -5491
rect -632 -5525 -626 -5491
rect -672 -5563 -626 -5525
rect -672 -5597 -666 -5563
rect -632 -5597 -626 -5563
rect -672 -5635 -626 -5597
rect -672 -5669 -666 -5635
rect -632 -5669 -626 -5635
rect -672 -5707 -626 -5669
rect -672 -5741 -666 -5707
rect -632 -5741 -626 -5707
rect -672 -5779 -626 -5741
rect -672 -5813 -666 -5779
rect -632 -5813 -626 -5779
rect -672 -5851 -626 -5813
rect -672 -5885 -666 -5851
rect -632 -5885 -626 -5851
rect -672 -5923 -626 -5885
rect -672 -5957 -666 -5923
rect -632 -5957 -626 -5923
rect -672 -5995 -626 -5957
rect -672 -6029 -666 -5995
rect -632 -6029 -626 -5995
rect -672 -6067 -626 -6029
rect -672 -6101 -666 -6067
rect -632 -6101 -626 -6067
rect -672 -6139 -626 -6101
rect -672 -6173 -666 -6139
rect -632 -6173 -626 -6139
rect -672 -6211 -626 -6173
rect -672 -6245 -666 -6211
rect -632 -6245 -626 -6211
rect -672 -6283 -626 -6245
rect -672 -6317 -666 -6283
rect -632 -6317 -626 -6283
rect -672 -6355 -626 -6317
rect -672 -6389 -666 -6355
rect -632 -6389 -626 -6355
rect -672 -6427 -626 -6389
rect -672 -6461 -666 -6427
rect -632 -6461 -626 -6427
rect -672 -6499 -626 -6461
rect -672 -6533 -666 -6499
rect -632 -6533 -626 -6499
rect -672 -6571 -626 -6533
rect -672 -6605 -666 -6571
rect -632 -6605 -626 -6571
rect -672 -6643 -626 -6605
rect -672 -6677 -666 -6643
rect -632 -6677 -626 -6643
rect -672 -6715 -626 -6677
rect -672 -6749 -666 -6715
rect -632 -6749 -626 -6715
rect -672 -6787 -626 -6749
rect -672 -6821 -666 -6787
rect -632 -6821 -626 -6787
rect -672 -6859 -626 -6821
rect -672 -6893 -666 -6859
rect -632 -6893 -626 -6859
rect -672 -6931 -626 -6893
rect -672 -6965 -666 -6931
rect -632 -6965 -626 -6931
rect -672 -7003 -626 -6965
rect -672 -7037 -666 -7003
rect -632 -7037 -626 -7003
rect -672 -7075 -626 -7037
rect -672 -7109 -666 -7075
rect -632 -7109 -626 -7075
rect -672 -7147 -626 -7109
rect -672 -7181 -666 -7147
rect -632 -7181 -626 -7147
rect -672 -7219 -626 -7181
rect -672 -7253 -666 -7219
rect -632 -7253 -626 -7219
rect -672 -7291 -626 -7253
rect -672 -7325 -666 -7291
rect -632 -7325 -626 -7291
rect -672 -7363 -626 -7325
rect -672 -7397 -666 -7363
rect -632 -7397 -626 -7363
rect -672 -7435 -626 -7397
rect -672 -7469 -666 -7435
rect -632 -7469 -626 -7435
rect -672 -7507 -626 -7469
rect -672 -7541 -666 -7507
rect -632 -7541 -626 -7507
rect -672 -7579 -626 -7541
rect -672 -7613 -666 -7579
rect -632 -7613 -626 -7579
rect -672 -7651 -626 -7613
rect -672 -7685 -666 -7651
rect -632 -7685 -626 -7651
rect -672 -7723 -626 -7685
rect -672 -7757 -666 -7723
rect -632 -7757 -626 -7723
rect -672 -7795 -626 -7757
rect -672 -7829 -666 -7795
rect -632 -7829 -626 -7795
rect -672 -7867 -626 -7829
rect -672 -7901 -666 -7867
rect -632 -7901 -626 -7867
rect -672 -7939 -626 -7901
rect -672 -7973 -666 -7939
rect -632 -7973 -626 -7939
rect -672 -8011 -626 -7973
rect -672 -8045 -666 -8011
rect -632 -8045 -626 -8011
rect -672 -8083 -626 -8045
rect -672 -8117 -666 -8083
rect -632 -8117 -626 -8083
rect -672 -8155 -626 -8117
rect -672 -8189 -666 -8155
rect -632 -8189 -626 -8155
rect -672 -8227 -626 -8189
rect -672 -8261 -666 -8227
rect -632 -8261 -626 -8227
rect -672 -8299 -626 -8261
rect -672 -8333 -666 -8299
rect -632 -8333 -626 -8299
rect -672 -8371 -626 -8333
rect -672 -8405 -666 -8371
rect -632 -8405 -626 -8371
rect -672 -8443 -626 -8405
rect -672 -8477 -666 -8443
rect -632 -8477 -626 -8443
rect -672 -8515 -626 -8477
rect -672 -8549 -666 -8515
rect -632 -8549 -626 -8515
rect -672 -8587 -626 -8549
rect -672 -8621 -666 -8587
rect -632 -8621 -626 -8587
rect -672 -8659 -626 -8621
rect -672 -8693 -666 -8659
rect -632 -8693 -626 -8659
rect -672 -8731 -626 -8693
rect -672 -8765 -666 -8731
rect -632 -8765 -626 -8731
rect -672 -8803 -626 -8765
rect -672 -8837 -666 -8803
rect -632 -8837 -626 -8803
rect -672 -8875 -626 -8837
rect -672 -8909 -666 -8875
rect -632 -8909 -626 -8875
rect -672 -8947 -626 -8909
rect -672 -8981 -666 -8947
rect -632 -8981 -626 -8947
rect -672 -9019 -626 -8981
rect -672 -9053 -666 -9019
rect -632 -9053 -626 -9019
rect -672 -9091 -626 -9053
rect -672 -9125 -666 -9091
rect -632 -9125 -626 -9091
rect -672 -9163 -626 -9125
rect -672 -9197 -666 -9163
rect -632 -9197 -626 -9163
rect -672 -9235 -626 -9197
rect -672 -9269 -666 -9235
rect -632 -9269 -626 -9235
rect -672 -9307 -626 -9269
rect -672 -9341 -666 -9307
rect -632 -9341 -626 -9307
rect -672 -9379 -626 -9341
rect -672 -9413 -666 -9379
rect -632 -9413 -626 -9379
rect -672 -9451 -626 -9413
rect -672 -9485 -666 -9451
rect -632 -9485 -626 -9451
rect -672 -9523 -626 -9485
rect -672 -9557 -666 -9523
rect -632 -9557 -626 -9523
rect -672 -9600 -626 -9557
rect -554 9557 -508 9600
rect -554 9523 -548 9557
rect -514 9523 -508 9557
rect -554 9485 -508 9523
rect -554 9451 -548 9485
rect -514 9451 -508 9485
rect -554 9413 -508 9451
rect -554 9379 -548 9413
rect -514 9379 -508 9413
rect -554 9341 -508 9379
rect -554 9307 -548 9341
rect -514 9307 -508 9341
rect -554 9269 -508 9307
rect -554 9235 -548 9269
rect -514 9235 -508 9269
rect -554 9197 -508 9235
rect -554 9163 -548 9197
rect -514 9163 -508 9197
rect -554 9125 -508 9163
rect -554 9091 -548 9125
rect -514 9091 -508 9125
rect -554 9053 -508 9091
rect -554 9019 -548 9053
rect -514 9019 -508 9053
rect -554 8981 -508 9019
rect -554 8947 -548 8981
rect -514 8947 -508 8981
rect -554 8909 -508 8947
rect -554 8875 -548 8909
rect -514 8875 -508 8909
rect -554 8837 -508 8875
rect -554 8803 -548 8837
rect -514 8803 -508 8837
rect -554 8765 -508 8803
rect -554 8731 -548 8765
rect -514 8731 -508 8765
rect -554 8693 -508 8731
rect -554 8659 -548 8693
rect -514 8659 -508 8693
rect -554 8621 -508 8659
rect -554 8587 -548 8621
rect -514 8587 -508 8621
rect -554 8549 -508 8587
rect -554 8515 -548 8549
rect -514 8515 -508 8549
rect -554 8477 -508 8515
rect -554 8443 -548 8477
rect -514 8443 -508 8477
rect -554 8405 -508 8443
rect -554 8371 -548 8405
rect -514 8371 -508 8405
rect -554 8333 -508 8371
rect -554 8299 -548 8333
rect -514 8299 -508 8333
rect -554 8261 -508 8299
rect -554 8227 -548 8261
rect -514 8227 -508 8261
rect -554 8189 -508 8227
rect -554 8155 -548 8189
rect -514 8155 -508 8189
rect -554 8117 -508 8155
rect -554 8083 -548 8117
rect -514 8083 -508 8117
rect -554 8045 -508 8083
rect -554 8011 -548 8045
rect -514 8011 -508 8045
rect -554 7973 -508 8011
rect -554 7939 -548 7973
rect -514 7939 -508 7973
rect -554 7901 -508 7939
rect -554 7867 -548 7901
rect -514 7867 -508 7901
rect -554 7829 -508 7867
rect -554 7795 -548 7829
rect -514 7795 -508 7829
rect -554 7757 -508 7795
rect -554 7723 -548 7757
rect -514 7723 -508 7757
rect -554 7685 -508 7723
rect -554 7651 -548 7685
rect -514 7651 -508 7685
rect -554 7613 -508 7651
rect -554 7579 -548 7613
rect -514 7579 -508 7613
rect -554 7541 -508 7579
rect -554 7507 -548 7541
rect -514 7507 -508 7541
rect -554 7469 -508 7507
rect -554 7435 -548 7469
rect -514 7435 -508 7469
rect -554 7397 -508 7435
rect -554 7363 -548 7397
rect -514 7363 -508 7397
rect -554 7325 -508 7363
rect -554 7291 -548 7325
rect -514 7291 -508 7325
rect -554 7253 -508 7291
rect -554 7219 -548 7253
rect -514 7219 -508 7253
rect -554 7181 -508 7219
rect -554 7147 -548 7181
rect -514 7147 -508 7181
rect -554 7109 -508 7147
rect -554 7075 -548 7109
rect -514 7075 -508 7109
rect -554 7037 -508 7075
rect -554 7003 -548 7037
rect -514 7003 -508 7037
rect -554 6965 -508 7003
rect -554 6931 -548 6965
rect -514 6931 -508 6965
rect -554 6893 -508 6931
rect -554 6859 -548 6893
rect -514 6859 -508 6893
rect -554 6821 -508 6859
rect -554 6787 -548 6821
rect -514 6787 -508 6821
rect -554 6749 -508 6787
rect -554 6715 -548 6749
rect -514 6715 -508 6749
rect -554 6677 -508 6715
rect -554 6643 -548 6677
rect -514 6643 -508 6677
rect -554 6605 -508 6643
rect -554 6571 -548 6605
rect -514 6571 -508 6605
rect -554 6533 -508 6571
rect -554 6499 -548 6533
rect -514 6499 -508 6533
rect -554 6461 -508 6499
rect -554 6427 -548 6461
rect -514 6427 -508 6461
rect -554 6389 -508 6427
rect -554 6355 -548 6389
rect -514 6355 -508 6389
rect -554 6317 -508 6355
rect -554 6283 -548 6317
rect -514 6283 -508 6317
rect -554 6245 -508 6283
rect -554 6211 -548 6245
rect -514 6211 -508 6245
rect -554 6173 -508 6211
rect -554 6139 -548 6173
rect -514 6139 -508 6173
rect -554 6101 -508 6139
rect -554 6067 -548 6101
rect -514 6067 -508 6101
rect -554 6029 -508 6067
rect -554 5995 -548 6029
rect -514 5995 -508 6029
rect -554 5957 -508 5995
rect -554 5923 -548 5957
rect -514 5923 -508 5957
rect -554 5885 -508 5923
rect -554 5851 -548 5885
rect -514 5851 -508 5885
rect -554 5813 -508 5851
rect -554 5779 -548 5813
rect -514 5779 -508 5813
rect -554 5741 -508 5779
rect -554 5707 -548 5741
rect -514 5707 -508 5741
rect -554 5669 -508 5707
rect -554 5635 -548 5669
rect -514 5635 -508 5669
rect -554 5597 -508 5635
rect -554 5563 -548 5597
rect -514 5563 -508 5597
rect -554 5525 -508 5563
rect -554 5491 -548 5525
rect -514 5491 -508 5525
rect -554 5453 -508 5491
rect -554 5419 -548 5453
rect -514 5419 -508 5453
rect -554 5381 -508 5419
rect -554 5347 -548 5381
rect -514 5347 -508 5381
rect -554 5309 -508 5347
rect -554 5275 -548 5309
rect -514 5275 -508 5309
rect -554 5237 -508 5275
rect -554 5203 -548 5237
rect -514 5203 -508 5237
rect -554 5165 -508 5203
rect -554 5131 -548 5165
rect -514 5131 -508 5165
rect -554 5093 -508 5131
rect -554 5059 -548 5093
rect -514 5059 -508 5093
rect -554 5021 -508 5059
rect -554 4987 -548 5021
rect -514 4987 -508 5021
rect -554 4949 -508 4987
rect -554 4915 -548 4949
rect -514 4915 -508 4949
rect -554 4877 -508 4915
rect -554 4843 -548 4877
rect -514 4843 -508 4877
rect -554 4805 -508 4843
rect -554 4771 -548 4805
rect -514 4771 -508 4805
rect -554 4733 -508 4771
rect -554 4699 -548 4733
rect -514 4699 -508 4733
rect -554 4661 -508 4699
rect -554 4627 -548 4661
rect -514 4627 -508 4661
rect -554 4589 -508 4627
rect -554 4555 -548 4589
rect -514 4555 -508 4589
rect -554 4517 -508 4555
rect -554 4483 -548 4517
rect -514 4483 -508 4517
rect -554 4445 -508 4483
rect -554 4411 -548 4445
rect -514 4411 -508 4445
rect -554 4373 -508 4411
rect -554 4339 -548 4373
rect -514 4339 -508 4373
rect -554 4301 -508 4339
rect -554 4267 -548 4301
rect -514 4267 -508 4301
rect -554 4229 -508 4267
rect -554 4195 -548 4229
rect -514 4195 -508 4229
rect -554 4157 -508 4195
rect -554 4123 -548 4157
rect -514 4123 -508 4157
rect -554 4085 -508 4123
rect -554 4051 -548 4085
rect -514 4051 -508 4085
rect -554 4013 -508 4051
rect -554 3979 -548 4013
rect -514 3979 -508 4013
rect -554 3941 -508 3979
rect -554 3907 -548 3941
rect -514 3907 -508 3941
rect -554 3869 -508 3907
rect -554 3835 -548 3869
rect -514 3835 -508 3869
rect -554 3797 -508 3835
rect -554 3763 -548 3797
rect -514 3763 -508 3797
rect -554 3725 -508 3763
rect -554 3691 -548 3725
rect -514 3691 -508 3725
rect -554 3653 -508 3691
rect -554 3619 -548 3653
rect -514 3619 -508 3653
rect -554 3581 -508 3619
rect -554 3547 -548 3581
rect -514 3547 -508 3581
rect -554 3509 -508 3547
rect -554 3475 -548 3509
rect -514 3475 -508 3509
rect -554 3437 -508 3475
rect -554 3403 -548 3437
rect -514 3403 -508 3437
rect -554 3365 -508 3403
rect -554 3331 -548 3365
rect -514 3331 -508 3365
rect -554 3293 -508 3331
rect -554 3259 -548 3293
rect -514 3259 -508 3293
rect -554 3221 -508 3259
rect -554 3187 -548 3221
rect -514 3187 -508 3221
rect -554 3149 -508 3187
rect -554 3115 -548 3149
rect -514 3115 -508 3149
rect -554 3077 -508 3115
rect -554 3043 -548 3077
rect -514 3043 -508 3077
rect -554 3005 -508 3043
rect -554 2971 -548 3005
rect -514 2971 -508 3005
rect -554 2933 -508 2971
rect -554 2899 -548 2933
rect -514 2899 -508 2933
rect -554 2861 -508 2899
rect -554 2827 -548 2861
rect -514 2827 -508 2861
rect -554 2789 -508 2827
rect -554 2755 -548 2789
rect -514 2755 -508 2789
rect -554 2717 -508 2755
rect -554 2683 -548 2717
rect -514 2683 -508 2717
rect -554 2645 -508 2683
rect -554 2611 -548 2645
rect -514 2611 -508 2645
rect -554 2573 -508 2611
rect -554 2539 -548 2573
rect -514 2539 -508 2573
rect -554 2501 -508 2539
rect -554 2467 -548 2501
rect -514 2467 -508 2501
rect -554 2429 -508 2467
rect -554 2395 -548 2429
rect -514 2395 -508 2429
rect -554 2357 -508 2395
rect -554 2323 -548 2357
rect -514 2323 -508 2357
rect -554 2285 -508 2323
rect -554 2251 -548 2285
rect -514 2251 -508 2285
rect -554 2213 -508 2251
rect -554 2179 -548 2213
rect -514 2179 -508 2213
rect -554 2141 -508 2179
rect -554 2107 -548 2141
rect -514 2107 -508 2141
rect -554 2069 -508 2107
rect -554 2035 -548 2069
rect -514 2035 -508 2069
rect -554 1997 -508 2035
rect -554 1963 -548 1997
rect -514 1963 -508 1997
rect -554 1925 -508 1963
rect -554 1891 -548 1925
rect -514 1891 -508 1925
rect -554 1853 -508 1891
rect -554 1819 -548 1853
rect -514 1819 -508 1853
rect -554 1781 -508 1819
rect -554 1747 -548 1781
rect -514 1747 -508 1781
rect -554 1709 -508 1747
rect -554 1675 -548 1709
rect -514 1675 -508 1709
rect -554 1637 -508 1675
rect -554 1603 -548 1637
rect -514 1603 -508 1637
rect -554 1565 -508 1603
rect -554 1531 -548 1565
rect -514 1531 -508 1565
rect -554 1493 -508 1531
rect -554 1459 -548 1493
rect -514 1459 -508 1493
rect -554 1421 -508 1459
rect -554 1387 -548 1421
rect -514 1387 -508 1421
rect -554 1349 -508 1387
rect -554 1315 -548 1349
rect -514 1315 -508 1349
rect -554 1277 -508 1315
rect -554 1243 -548 1277
rect -514 1243 -508 1277
rect -554 1205 -508 1243
rect -554 1171 -548 1205
rect -514 1171 -508 1205
rect -554 1133 -508 1171
rect -554 1099 -548 1133
rect -514 1099 -508 1133
rect -554 1061 -508 1099
rect -554 1027 -548 1061
rect -514 1027 -508 1061
rect -554 989 -508 1027
rect -554 955 -548 989
rect -514 955 -508 989
rect -554 917 -508 955
rect -554 883 -548 917
rect -514 883 -508 917
rect -554 845 -508 883
rect -554 811 -548 845
rect -514 811 -508 845
rect -554 773 -508 811
rect -554 739 -548 773
rect -514 739 -508 773
rect -554 701 -508 739
rect -554 667 -548 701
rect -514 667 -508 701
rect -554 629 -508 667
rect -554 595 -548 629
rect -514 595 -508 629
rect -554 557 -508 595
rect -554 523 -548 557
rect -514 523 -508 557
rect -554 485 -508 523
rect -554 451 -548 485
rect -514 451 -508 485
rect -554 413 -508 451
rect -554 379 -548 413
rect -514 379 -508 413
rect -554 341 -508 379
rect -554 307 -548 341
rect -514 307 -508 341
rect -554 269 -508 307
rect -554 235 -548 269
rect -514 235 -508 269
rect -554 197 -508 235
rect -554 163 -548 197
rect -514 163 -508 197
rect -554 125 -508 163
rect -554 91 -548 125
rect -514 91 -508 125
rect -554 53 -508 91
rect -554 19 -548 53
rect -514 19 -508 53
rect -554 -19 -508 19
rect -554 -53 -548 -19
rect -514 -53 -508 -19
rect -554 -91 -508 -53
rect -554 -125 -548 -91
rect -514 -125 -508 -91
rect -554 -163 -508 -125
rect -554 -197 -548 -163
rect -514 -197 -508 -163
rect -554 -235 -508 -197
rect -554 -269 -548 -235
rect -514 -269 -508 -235
rect -554 -307 -508 -269
rect -554 -341 -548 -307
rect -514 -341 -508 -307
rect -554 -379 -508 -341
rect -554 -413 -548 -379
rect -514 -413 -508 -379
rect -554 -451 -508 -413
rect -554 -485 -548 -451
rect -514 -485 -508 -451
rect -554 -523 -508 -485
rect -554 -557 -548 -523
rect -514 -557 -508 -523
rect -554 -595 -508 -557
rect -554 -629 -548 -595
rect -514 -629 -508 -595
rect -554 -667 -508 -629
rect -554 -701 -548 -667
rect -514 -701 -508 -667
rect -554 -739 -508 -701
rect -554 -773 -548 -739
rect -514 -773 -508 -739
rect -554 -811 -508 -773
rect -554 -845 -548 -811
rect -514 -845 -508 -811
rect -554 -883 -508 -845
rect -554 -917 -548 -883
rect -514 -917 -508 -883
rect -554 -955 -508 -917
rect -554 -989 -548 -955
rect -514 -989 -508 -955
rect -554 -1027 -508 -989
rect -554 -1061 -548 -1027
rect -514 -1061 -508 -1027
rect -554 -1099 -508 -1061
rect -554 -1133 -548 -1099
rect -514 -1133 -508 -1099
rect -554 -1171 -508 -1133
rect -554 -1205 -548 -1171
rect -514 -1205 -508 -1171
rect -554 -1243 -508 -1205
rect -554 -1277 -548 -1243
rect -514 -1277 -508 -1243
rect -554 -1315 -508 -1277
rect -554 -1349 -548 -1315
rect -514 -1349 -508 -1315
rect -554 -1387 -508 -1349
rect -554 -1421 -548 -1387
rect -514 -1421 -508 -1387
rect -554 -1459 -508 -1421
rect -554 -1493 -548 -1459
rect -514 -1493 -508 -1459
rect -554 -1531 -508 -1493
rect -554 -1565 -548 -1531
rect -514 -1565 -508 -1531
rect -554 -1603 -508 -1565
rect -554 -1637 -548 -1603
rect -514 -1637 -508 -1603
rect -554 -1675 -508 -1637
rect -554 -1709 -548 -1675
rect -514 -1709 -508 -1675
rect -554 -1747 -508 -1709
rect -554 -1781 -548 -1747
rect -514 -1781 -508 -1747
rect -554 -1819 -508 -1781
rect -554 -1853 -548 -1819
rect -514 -1853 -508 -1819
rect -554 -1891 -508 -1853
rect -554 -1925 -548 -1891
rect -514 -1925 -508 -1891
rect -554 -1963 -508 -1925
rect -554 -1997 -548 -1963
rect -514 -1997 -508 -1963
rect -554 -2035 -508 -1997
rect -554 -2069 -548 -2035
rect -514 -2069 -508 -2035
rect -554 -2107 -508 -2069
rect -554 -2141 -548 -2107
rect -514 -2141 -508 -2107
rect -554 -2179 -508 -2141
rect -554 -2213 -548 -2179
rect -514 -2213 -508 -2179
rect -554 -2251 -508 -2213
rect -554 -2285 -548 -2251
rect -514 -2285 -508 -2251
rect -554 -2323 -508 -2285
rect -554 -2357 -548 -2323
rect -514 -2357 -508 -2323
rect -554 -2395 -508 -2357
rect -554 -2429 -548 -2395
rect -514 -2429 -508 -2395
rect -554 -2467 -508 -2429
rect -554 -2501 -548 -2467
rect -514 -2501 -508 -2467
rect -554 -2539 -508 -2501
rect -554 -2573 -548 -2539
rect -514 -2573 -508 -2539
rect -554 -2611 -508 -2573
rect -554 -2645 -548 -2611
rect -514 -2645 -508 -2611
rect -554 -2683 -508 -2645
rect -554 -2717 -548 -2683
rect -514 -2717 -508 -2683
rect -554 -2755 -508 -2717
rect -554 -2789 -548 -2755
rect -514 -2789 -508 -2755
rect -554 -2827 -508 -2789
rect -554 -2861 -548 -2827
rect -514 -2861 -508 -2827
rect -554 -2899 -508 -2861
rect -554 -2933 -548 -2899
rect -514 -2933 -508 -2899
rect -554 -2971 -508 -2933
rect -554 -3005 -548 -2971
rect -514 -3005 -508 -2971
rect -554 -3043 -508 -3005
rect -554 -3077 -548 -3043
rect -514 -3077 -508 -3043
rect -554 -3115 -508 -3077
rect -554 -3149 -548 -3115
rect -514 -3149 -508 -3115
rect -554 -3187 -508 -3149
rect -554 -3221 -548 -3187
rect -514 -3221 -508 -3187
rect -554 -3259 -508 -3221
rect -554 -3293 -548 -3259
rect -514 -3293 -508 -3259
rect -554 -3331 -508 -3293
rect -554 -3365 -548 -3331
rect -514 -3365 -508 -3331
rect -554 -3403 -508 -3365
rect -554 -3437 -548 -3403
rect -514 -3437 -508 -3403
rect -554 -3475 -508 -3437
rect -554 -3509 -548 -3475
rect -514 -3509 -508 -3475
rect -554 -3547 -508 -3509
rect -554 -3581 -548 -3547
rect -514 -3581 -508 -3547
rect -554 -3619 -508 -3581
rect -554 -3653 -548 -3619
rect -514 -3653 -508 -3619
rect -554 -3691 -508 -3653
rect -554 -3725 -548 -3691
rect -514 -3725 -508 -3691
rect -554 -3763 -508 -3725
rect -554 -3797 -548 -3763
rect -514 -3797 -508 -3763
rect -554 -3835 -508 -3797
rect -554 -3869 -548 -3835
rect -514 -3869 -508 -3835
rect -554 -3907 -508 -3869
rect -554 -3941 -548 -3907
rect -514 -3941 -508 -3907
rect -554 -3979 -508 -3941
rect -554 -4013 -548 -3979
rect -514 -4013 -508 -3979
rect -554 -4051 -508 -4013
rect -554 -4085 -548 -4051
rect -514 -4085 -508 -4051
rect -554 -4123 -508 -4085
rect -554 -4157 -548 -4123
rect -514 -4157 -508 -4123
rect -554 -4195 -508 -4157
rect -554 -4229 -548 -4195
rect -514 -4229 -508 -4195
rect -554 -4267 -508 -4229
rect -554 -4301 -548 -4267
rect -514 -4301 -508 -4267
rect -554 -4339 -508 -4301
rect -554 -4373 -548 -4339
rect -514 -4373 -508 -4339
rect -554 -4411 -508 -4373
rect -554 -4445 -548 -4411
rect -514 -4445 -508 -4411
rect -554 -4483 -508 -4445
rect -554 -4517 -548 -4483
rect -514 -4517 -508 -4483
rect -554 -4555 -508 -4517
rect -554 -4589 -548 -4555
rect -514 -4589 -508 -4555
rect -554 -4627 -508 -4589
rect -554 -4661 -548 -4627
rect -514 -4661 -508 -4627
rect -554 -4699 -508 -4661
rect -554 -4733 -548 -4699
rect -514 -4733 -508 -4699
rect -554 -4771 -508 -4733
rect -554 -4805 -548 -4771
rect -514 -4805 -508 -4771
rect -554 -4843 -508 -4805
rect -554 -4877 -548 -4843
rect -514 -4877 -508 -4843
rect -554 -4915 -508 -4877
rect -554 -4949 -548 -4915
rect -514 -4949 -508 -4915
rect -554 -4987 -508 -4949
rect -554 -5021 -548 -4987
rect -514 -5021 -508 -4987
rect -554 -5059 -508 -5021
rect -554 -5093 -548 -5059
rect -514 -5093 -508 -5059
rect -554 -5131 -508 -5093
rect -554 -5165 -548 -5131
rect -514 -5165 -508 -5131
rect -554 -5203 -508 -5165
rect -554 -5237 -548 -5203
rect -514 -5237 -508 -5203
rect -554 -5275 -508 -5237
rect -554 -5309 -548 -5275
rect -514 -5309 -508 -5275
rect -554 -5347 -508 -5309
rect -554 -5381 -548 -5347
rect -514 -5381 -508 -5347
rect -554 -5419 -508 -5381
rect -554 -5453 -548 -5419
rect -514 -5453 -508 -5419
rect -554 -5491 -508 -5453
rect -554 -5525 -548 -5491
rect -514 -5525 -508 -5491
rect -554 -5563 -508 -5525
rect -554 -5597 -548 -5563
rect -514 -5597 -508 -5563
rect -554 -5635 -508 -5597
rect -554 -5669 -548 -5635
rect -514 -5669 -508 -5635
rect -554 -5707 -508 -5669
rect -554 -5741 -548 -5707
rect -514 -5741 -508 -5707
rect -554 -5779 -508 -5741
rect -554 -5813 -548 -5779
rect -514 -5813 -508 -5779
rect -554 -5851 -508 -5813
rect -554 -5885 -548 -5851
rect -514 -5885 -508 -5851
rect -554 -5923 -508 -5885
rect -554 -5957 -548 -5923
rect -514 -5957 -508 -5923
rect -554 -5995 -508 -5957
rect -554 -6029 -548 -5995
rect -514 -6029 -508 -5995
rect -554 -6067 -508 -6029
rect -554 -6101 -548 -6067
rect -514 -6101 -508 -6067
rect -554 -6139 -508 -6101
rect -554 -6173 -548 -6139
rect -514 -6173 -508 -6139
rect -554 -6211 -508 -6173
rect -554 -6245 -548 -6211
rect -514 -6245 -508 -6211
rect -554 -6283 -508 -6245
rect -554 -6317 -548 -6283
rect -514 -6317 -508 -6283
rect -554 -6355 -508 -6317
rect -554 -6389 -548 -6355
rect -514 -6389 -508 -6355
rect -554 -6427 -508 -6389
rect -554 -6461 -548 -6427
rect -514 -6461 -508 -6427
rect -554 -6499 -508 -6461
rect -554 -6533 -548 -6499
rect -514 -6533 -508 -6499
rect -554 -6571 -508 -6533
rect -554 -6605 -548 -6571
rect -514 -6605 -508 -6571
rect -554 -6643 -508 -6605
rect -554 -6677 -548 -6643
rect -514 -6677 -508 -6643
rect -554 -6715 -508 -6677
rect -554 -6749 -548 -6715
rect -514 -6749 -508 -6715
rect -554 -6787 -508 -6749
rect -554 -6821 -548 -6787
rect -514 -6821 -508 -6787
rect -554 -6859 -508 -6821
rect -554 -6893 -548 -6859
rect -514 -6893 -508 -6859
rect -554 -6931 -508 -6893
rect -554 -6965 -548 -6931
rect -514 -6965 -508 -6931
rect -554 -7003 -508 -6965
rect -554 -7037 -548 -7003
rect -514 -7037 -508 -7003
rect -554 -7075 -508 -7037
rect -554 -7109 -548 -7075
rect -514 -7109 -508 -7075
rect -554 -7147 -508 -7109
rect -554 -7181 -548 -7147
rect -514 -7181 -508 -7147
rect -554 -7219 -508 -7181
rect -554 -7253 -548 -7219
rect -514 -7253 -508 -7219
rect -554 -7291 -508 -7253
rect -554 -7325 -548 -7291
rect -514 -7325 -508 -7291
rect -554 -7363 -508 -7325
rect -554 -7397 -548 -7363
rect -514 -7397 -508 -7363
rect -554 -7435 -508 -7397
rect -554 -7469 -548 -7435
rect -514 -7469 -508 -7435
rect -554 -7507 -508 -7469
rect -554 -7541 -548 -7507
rect -514 -7541 -508 -7507
rect -554 -7579 -508 -7541
rect -554 -7613 -548 -7579
rect -514 -7613 -508 -7579
rect -554 -7651 -508 -7613
rect -554 -7685 -548 -7651
rect -514 -7685 -508 -7651
rect -554 -7723 -508 -7685
rect -554 -7757 -548 -7723
rect -514 -7757 -508 -7723
rect -554 -7795 -508 -7757
rect -554 -7829 -548 -7795
rect -514 -7829 -508 -7795
rect -554 -7867 -508 -7829
rect -554 -7901 -548 -7867
rect -514 -7901 -508 -7867
rect -554 -7939 -508 -7901
rect -554 -7973 -548 -7939
rect -514 -7973 -508 -7939
rect -554 -8011 -508 -7973
rect -554 -8045 -548 -8011
rect -514 -8045 -508 -8011
rect -554 -8083 -508 -8045
rect -554 -8117 -548 -8083
rect -514 -8117 -508 -8083
rect -554 -8155 -508 -8117
rect -554 -8189 -548 -8155
rect -514 -8189 -508 -8155
rect -554 -8227 -508 -8189
rect -554 -8261 -548 -8227
rect -514 -8261 -508 -8227
rect -554 -8299 -508 -8261
rect -554 -8333 -548 -8299
rect -514 -8333 -508 -8299
rect -554 -8371 -508 -8333
rect -554 -8405 -548 -8371
rect -514 -8405 -508 -8371
rect -554 -8443 -508 -8405
rect -554 -8477 -548 -8443
rect -514 -8477 -508 -8443
rect -554 -8515 -508 -8477
rect -554 -8549 -548 -8515
rect -514 -8549 -508 -8515
rect -554 -8587 -508 -8549
rect -554 -8621 -548 -8587
rect -514 -8621 -508 -8587
rect -554 -8659 -508 -8621
rect -554 -8693 -548 -8659
rect -514 -8693 -508 -8659
rect -554 -8731 -508 -8693
rect -554 -8765 -548 -8731
rect -514 -8765 -508 -8731
rect -554 -8803 -508 -8765
rect -554 -8837 -548 -8803
rect -514 -8837 -508 -8803
rect -554 -8875 -508 -8837
rect -554 -8909 -548 -8875
rect -514 -8909 -508 -8875
rect -554 -8947 -508 -8909
rect -554 -8981 -548 -8947
rect -514 -8981 -508 -8947
rect -554 -9019 -508 -8981
rect -554 -9053 -548 -9019
rect -514 -9053 -508 -9019
rect -554 -9091 -508 -9053
rect -554 -9125 -548 -9091
rect -514 -9125 -508 -9091
rect -554 -9163 -508 -9125
rect -554 -9197 -548 -9163
rect -514 -9197 -508 -9163
rect -554 -9235 -508 -9197
rect -554 -9269 -548 -9235
rect -514 -9269 -508 -9235
rect -554 -9307 -508 -9269
rect -554 -9341 -548 -9307
rect -514 -9341 -508 -9307
rect -554 -9379 -508 -9341
rect -554 -9413 -548 -9379
rect -514 -9413 -508 -9379
rect -554 -9451 -508 -9413
rect -554 -9485 -548 -9451
rect -514 -9485 -508 -9451
rect -554 -9523 -508 -9485
rect -554 -9557 -548 -9523
rect -514 -9557 -508 -9523
rect -554 -9600 -508 -9557
rect -436 9557 -390 9600
rect -436 9523 -430 9557
rect -396 9523 -390 9557
rect -436 9485 -390 9523
rect -436 9451 -430 9485
rect -396 9451 -390 9485
rect -436 9413 -390 9451
rect -436 9379 -430 9413
rect -396 9379 -390 9413
rect -436 9341 -390 9379
rect -436 9307 -430 9341
rect -396 9307 -390 9341
rect -436 9269 -390 9307
rect -436 9235 -430 9269
rect -396 9235 -390 9269
rect -436 9197 -390 9235
rect -436 9163 -430 9197
rect -396 9163 -390 9197
rect -436 9125 -390 9163
rect -436 9091 -430 9125
rect -396 9091 -390 9125
rect -436 9053 -390 9091
rect -436 9019 -430 9053
rect -396 9019 -390 9053
rect -436 8981 -390 9019
rect -436 8947 -430 8981
rect -396 8947 -390 8981
rect -436 8909 -390 8947
rect -436 8875 -430 8909
rect -396 8875 -390 8909
rect -436 8837 -390 8875
rect -436 8803 -430 8837
rect -396 8803 -390 8837
rect -436 8765 -390 8803
rect -436 8731 -430 8765
rect -396 8731 -390 8765
rect -436 8693 -390 8731
rect -436 8659 -430 8693
rect -396 8659 -390 8693
rect -436 8621 -390 8659
rect -436 8587 -430 8621
rect -396 8587 -390 8621
rect -436 8549 -390 8587
rect -436 8515 -430 8549
rect -396 8515 -390 8549
rect -436 8477 -390 8515
rect -436 8443 -430 8477
rect -396 8443 -390 8477
rect -436 8405 -390 8443
rect -436 8371 -430 8405
rect -396 8371 -390 8405
rect -436 8333 -390 8371
rect -436 8299 -430 8333
rect -396 8299 -390 8333
rect -436 8261 -390 8299
rect -436 8227 -430 8261
rect -396 8227 -390 8261
rect -436 8189 -390 8227
rect -436 8155 -430 8189
rect -396 8155 -390 8189
rect -436 8117 -390 8155
rect -436 8083 -430 8117
rect -396 8083 -390 8117
rect -436 8045 -390 8083
rect -436 8011 -430 8045
rect -396 8011 -390 8045
rect -436 7973 -390 8011
rect -436 7939 -430 7973
rect -396 7939 -390 7973
rect -436 7901 -390 7939
rect -436 7867 -430 7901
rect -396 7867 -390 7901
rect -436 7829 -390 7867
rect -436 7795 -430 7829
rect -396 7795 -390 7829
rect -436 7757 -390 7795
rect -436 7723 -430 7757
rect -396 7723 -390 7757
rect -436 7685 -390 7723
rect -436 7651 -430 7685
rect -396 7651 -390 7685
rect -436 7613 -390 7651
rect -436 7579 -430 7613
rect -396 7579 -390 7613
rect -436 7541 -390 7579
rect -436 7507 -430 7541
rect -396 7507 -390 7541
rect -436 7469 -390 7507
rect -436 7435 -430 7469
rect -396 7435 -390 7469
rect -436 7397 -390 7435
rect -436 7363 -430 7397
rect -396 7363 -390 7397
rect -436 7325 -390 7363
rect -436 7291 -430 7325
rect -396 7291 -390 7325
rect -436 7253 -390 7291
rect -436 7219 -430 7253
rect -396 7219 -390 7253
rect -436 7181 -390 7219
rect -436 7147 -430 7181
rect -396 7147 -390 7181
rect -436 7109 -390 7147
rect -436 7075 -430 7109
rect -396 7075 -390 7109
rect -436 7037 -390 7075
rect -436 7003 -430 7037
rect -396 7003 -390 7037
rect -436 6965 -390 7003
rect -436 6931 -430 6965
rect -396 6931 -390 6965
rect -436 6893 -390 6931
rect -436 6859 -430 6893
rect -396 6859 -390 6893
rect -436 6821 -390 6859
rect -436 6787 -430 6821
rect -396 6787 -390 6821
rect -436 6749 -390 6787
rect -436 6715 -430 6749
rect -396 6715 -390 6749
rect -436 6677 -390 6715
rect -436 6643 -430 6677
rect -396 6643 -390 6677
rect -436 6605 -390 6643
rect -436 6571 -430 6605
rect -396 6571 -390 6605
rect -436 6533 -390 6571
rect -436 6499 -430 6533
rect -396 6499 -390 6533
rect -436 6461 -390 6499
rect -436 6427 -430 6461
rect -396 6427 -390 6461
rect -436 6389 -390 6427
rect -436 6355 -430 6389
rect -396 6355 -390 6389
rect -436 6317 -390 6355
rect -436 6283 -430 6317
rect -396 6283 -390 6317
rect -436 6245 -390 6283
rect -436 6211 -430 6245
rect -396 6211 -390 6245
rect -436 6173 -390 6211
rect -436 6139 -430 6173
rect -396 6139 -390 6173
rect -436 6101 -390 6139
rect -436 6067 -430 6101
rect -396 6067 -390 6101
rect -436 6029 -390 6067
rect -436 5995 -430 6029
rect -396 5995 -390 6029
rect -436 5957 -390 5995
rect -436 5923 -430 5957
rect -396 5923 -390 5957
rect -436 5885 -390 5923
rect -436 5851 -430 5885
rect -396 5851 -390 5885
rect -436 5813 -390 5851
rect -436 5779 -430 5813
rect -396 5779 -390 5813
rect -436 5741 -390 5779
rect -436 5707 -430 5741
rect -396 5707 -390 5741
rect -436 5669 -390 5707
rect -436 5635 -430 5669
rect -396 5635 -390 5669
rect -436 5597 -390 5635
rect -436 5563 -430 5597
rect -396 5563 -390 5597
rect -436 5525 -390 5563
rect -436 5491 -430 5525
rect -396 5491 -390 5525
rect -436 5453 -390 5491
rect -436 5419 -430 5453
rect -396 5419 -390 5453
rect -436 5381 -390 5419
rect -436 5347 -430 5381
rect -396 5347 -390 5381
rect -436 5309 -390 5347
rect -436 5275 -430 5309
rect -396 5275 -390 5309
rect -436 5237 -390 5275
rect -436 5203 -430 5237
rect -396 5203 -390 5237
rect -436 5165 -390 5203
rect -436 5131 -430 5165
rect -396 5131 -390 5165
rect -436 5093 -390 5131
rect -436 5059 -430 5093
rect -396 5059 -390 5093
rect -436 5021 -390 5059
rect -436 4987 -430 5021
rect -396 4987 -390 5021
rect -436 4949 -390 4987
rect -436 4915 -430 4949
rect -396 4915 -390 4949
rect -436 4877 -390 4915
rect -436 4843 -430 4877
rect -396 4843 -390 4877
rect -436 4805 -390 4843
rect -436 4771 -430 4805
rect -396 4771 -390 4805
rect -436 4733 -390 4771
rect -436 4699 -430 4733
rect -396 4699 -390 4733
rect -436 4661 -390 4699
rect -436 4627 -430 4661
rect -396 4627 -390 4661
rect -436 4589 -390 4627
rect -436 4555 -430 4589
rect -396 4555 -390 4589
rect -436 4517 -390 4555
rect -436 4483 -430 4517
rect -396 4483 -390 4517
rect -436 4445 -390 4483
rect -436 4411 -430 4445
rect -396 4411 -390 4445
rect -436 4373 -390 4411
rect -436 4339 -430 4373
rect -396 4339 -390 4373
rect -436 4301 -390 4339
rect -436 4267 -430 4301
rect -396 4267 -390 4301
rect -436 4229 -390 4267
rect -436 4195 -430 4229
rect -396 4195 -390 4229
rect -436 4157 -390 4195
rect -436 4123 -430 4157
rect -396 4123 -390 4157
rect -436 4085 -390 4123
rect -436 4051 -430 4085
rect -396 4051 -390 4085
rect -436 4013 -390 4051
rect -436 3979 -430 4013
rect -396 3979 -390 4013
rect -436 3941 -390 3979
rect -436 3907 -430 3941
rect -396 3907 -390 3941
rect -436 3869 -390 3907
rect -436 3835 -430 3869
rect -396 3835 -390 3869
rect -436 3797 -390 3835
rect -436 3763 -430 3797
rect -396 3763 -390 3797
rect -436 3725 -390 3763
rect -436 3691 -430 3725
rect -396 3691 -390 3725
rect -436 3653 -390 3691
rect -436 3619 -430 3653
rect -396 3619 -390 3653
rect -436 3581 -390 3619
rect -436 3547 -430 3581
rect -396 3547 -390 3581
rect -436 3509 -390 3547
rect -436 3475 -430 3509
rect -396 3475 -390 3509
rect -436 3437 -390 3475
rect -436 3403 -430 3437
rect -396 3403 -390 3437
rect -436 3365 -390 3403
rect -436 3331 -430 3365
rect -396 3331 -390 3365
rect -436 3293 -390 3331
rect -436 3259 -430 3293
rect -396 3259 -390 3293
rect -436 3221 -390 3259
rect -436 3187 -430 3221
rect -396 3187 -390 3221
rect -436 3149 -390 3187
rect -436 3115 -430 3149
rect -396 3115 -390 3149
rect -436 3077 -390 3115
rect -436 3043 -430 3077
rect -396 3043 -390 3077
rect -436 3005 -390 3043
rect -436 2971 -430 3005
rect -396 2971 -390 3005
rect -436 2933 -390 2971
rect -436 2899 -430 2933
rect -396 2899 -390 2933
rect -436 2861 -390 2899
rect -436 2827 -430 2861
rect -396 2827 -390 2861
rect -436 2789 -390 2827
rect -436 2755 -430 2789
rect -396 2755 -390 2789
rect -436 2717 -390 2755
rect -436 2683 -430 2717
rect -396 2683 -390 2717
rect -436 2645 -390 2683
rect -436 2611 -430 2645
rect -396 2611 -390 2645
rect -436 2573 -390 2611
rect -436 2539 -430 2573
rect -396 2539 -390 2573
rect -436 2501 -390 2539
rect -436 2467 -430 2501
rect -396 2467 -390 2501
rect -436 2429 -390 2467
rect -436 2395 -430 2429
rect -396 2395 -390 2429
rect -436 2357 -390 2395
rect -436 2323 -430 2357
rect -396 2323 -390 2357
rect -436 2285 -390 2323
rect -436 2251 -430 2285
rect -396 2251 -390 2285
rect -436 2213 -390 2251
rect -436 2179 -430 2213
rect -396 2179 -390 2213
rect -436 2141 -390 2179
rect -436 2107 -430 2141
rect -396 2107 -390 2141
rect -436 2069 -390 2107
rect -436 2035 -430 2069
rect -396 2035 -390 2069
rect -436 1997 -390 2035
rect -436 1963 -430 1997
rect -396 1963 -390 1997
rect -436 1925 -390 1963
rect -436 1891 -430 1925
rect -396 1891 -390 1925
rect -436 1853 -390 1891
rect -436 1819 -430 1853
rect -396 1819 -390 1853
rect -436 1781 -390 1819
rect -436 1747 -430 1781
rect -396 1747 -390 1781
rect -436 1709 -390 1747
rect -436 1675 -430 1709
rect -396 1675 -390 1709
rect -436 1637 -390 1675
rect -436 1603 -430 1637
rect -396 1603 -390 1637
rect -436 1565 -390 1603
rect -436 1531 -430 1565
rect -396 1531 -390 1565
rect -436 1493 -390 1531
rect -436 1459 -430 1493
rect -396 1459 -390 1493
rect -436 1421 -390 1459
rect -436 1387 -430 1421
rect -396 1387 -390 1421
rect -436 1349 -390 1387
rect -436 1315 -430 1349
rect -396 1315 -390 1349
rect -436 1277 -390 1315
rect -436 1243 -430 1277
rect -396 1243 -390 1277
rect -436 1205 -390 1243
rect -436 1171 -430 1205
rect -396 1171 -390 1205
rect -436 1133 -390 1171
rect -436 1099 -430 1133
rect -396 1099 -390 1133
rect -436 1061 -390 1099
rect -436 1027 -430 1061
rect -396 1027 -390 1061
rect -436 989 -390 1027
rect -436 955 -430 989
rect -396 955 -390 989
rect -436 917 -390 955
rect -436 883 -430 917
rect -396 883 -390 917
rect -436 845 -390 883
rect -436 811 -430 845
rect -396 811 -390 845
rect -436 773 -390 811
rect -436 739 -430 773
rect -396 739 -390 773
rect -436 701 -390 739
rect -436 667 -430 701
rect -396 667 -390 701
rect -436 629 -390 667
rect -436 595 -430 629
rect -396 595 -390 629
rect -436 557 -390 595
rect -436 523 -430 557
rect -396 523 -390 557
rect -436 485 -390 523
rect -436 451 -430 485
rect -396 451 -390 485
rect -436 413 -390 451
rect -436 379 -430 413
rect -396 379 -390 413
rect -436 341 -390 379
rect -436 307 -430 341
rect -396 307 -390 341
rect -436 269 -390 307
rect -436 235 -430 269
rect -396 235 -390 269
rect -436 197 -390 235
rect -436 163 -430 197
rect -396 163 -390 197
rect -436 125 -390 163
rect -436 91 -430 125
rect -396 91 -390 125
rect -436 53 -390 91
rect -436 19 -430 53
rect -396 19 -390 53
rect -436 -19 -390 19
rect -436 -53 -430 -19
rect -396 -53 -390 -19
rect -436 -91 -390 -53
rect -436 -125 -430 -91
rect -396 -125 -390 -91
rect -436 -163 -390 -125
rect -436 -197 -430 -163
rect -396 -197 -390 -163
rect -436 -235 -390 -197
rect -436 -269 -430 -235
rect -396 -269 -390 -235
rect -436 -307 -390 -269
rect -436 -341 -430 -307
rect -396 -341 -390 -307
rect -436 -379 -390 -341
rect -436 -413 -430 -379
rect -396 -413 -390 -379
rect -436 -451 -390 -413
rect -436 -485 -430 -451
rect -396 -485 -390 -451
rect -436 -523 -390 -485
rect -436 -557 -430 -523
rect -396 -557 -390 -523
rect -436 -595 -390 -557
rect -436 -629 -430 -595
rect -396 -629 -390 -595
rect -436 -667 -390 -629
rect -436 -701 -430 -667
rect -396 -701 -390 -667
rect -436 -739 -390 -701
rect -436 -773 -430 -739
rect -396 -773 -390 -739
rect -436 -811 -390 -773
rect -436 -845 -430 -811
rect -396 -845 -390 -811
rect -436 -883 -390 -845
rect -436 -917 -430 -883
rect -396 -917 -390 -883
rect -436 -955 -390 -917
rect -436 -989 -430 -955
rect -396 -989 -390 -955
rect -436 -1027 -390 -989
rect -436 -1061 -430 -1027
rect -396 -1061 -390 -1027
rect -436 -1099 -390 -1061
rect -436 -1133 -430 -1099
rect -396 -1133 -390 -1099
rect -436 -1171 -390 -1133
rect -436 -1205 -430 -1171
rect -396 -1205 -390 -1171
rect -436 -1243 -390 -1205
rect -436 -1277 -430 -1243
rect -396 -1277 -390 -1243
rect -436 -1315 -390 -1277
rect -436 -1349 -430 -1315
rect -396 -1349 -390 -1315
rect -436 -1387 -390 -1349
rect -436 -1421 -430 -1387
rect -396 -1421 -390 -1387
rect -436 -1459 -390 -1421
rect -436 -1493 -430 -1459
rect -396 -1493 -390 -1459
rect -436 -1531 -390 -1493
rect -436 -1565 -430 -1531
rect -396 -1565 -390 -1531
rect -436 -1603 -390 -1565
rect -436 -1637 -430 -1603
rect -396 -1637 -390 -1603
rect -436 -1675 -390 -1637
rect -436 -1709 -430 -1675
rect -396 -1709 -390 -1675
rect -436 -1747 -390 -1709
rect -436 -1781 -430 -1747
rect -396 -1781 -390 -1747
rect -436 -1819 -390 -1781
rect -436 -1853 -430 -1819
rect -396 -1853 -390 -1819
rect -436 -1891 -390 -1853
rect -436 -1925 -430 -1891
rect -396 -1925 -390 -1891
rect -436 -1963 -390 -1925
rect -436 -1997 -430 -1963
rect -396 -1997 -390 -1963
rect -436 -2035 -390 -1997
rect -436 -2069 -430 -2035
rect -396 -2069 -390 -2035
rect -436 -2107 -390 -2069
rect -436 -2141 -430 -2107
rect -396 -2141 -390 -2107
rect -436 -2179 -390 -2141
rect -436 -2213 -430 -2179
rect -396 -2213 -390 -2179
rect -436 -2251 -390 -2213
rect -436 -2285 -430 -2251
rect -396 -2285 -390 -2251
rect -436 -2323 -390 -2285
rect -436 -2357 -430 -2323
rect -396 -2357 -390 -2323
rect -436 -2395 -390 -2357
rect -436 -2429 -430 -2395
rect -396 -2429 -390 -2395
rect -436 -2467 -390 -2429
rect -436 -2501 -430 -2467
rect -396 -2501 -390 -2467
rect -436 -2539 -390 -2501
rect -436 -2573 -430 -2539
rect -396 -2573 -390 -2539
rect -436 -2611 -390 -2573
rect -436 -2645 -430 -2611
rect -396 -2645 -390 -2611
rect -436 -2683 -390 -2645
rect -436 -2717 -430 -2683
rect -396 -2717 -390 -2683
rect -436 -2755 -390 -2717
rect -436 -2789 -430 -2755
rect -396 -2789 -390 -2755
rect -436 -2827 -390 -2789
rect -436 -2861 -430 -2827
rect -396 -2861 -390 -2827
rect -436 -2899 -390 -2861
rect -436 -2933 -430 -2899
rect -396 -2933 -390 -2899
rect -436 -2971 -390 -2933
rect -436 -3005 -430 -2971
rect -396 -3005 -390 -2971
rect -436 -3043 -390 -3005
rect -436 -3077 -430 -3043
rect -396 -3077 -390 -3043
rect -436 -3115 -390 -3077
rect -436 -3149 -430 -3115
rect -396 -3149 -390 -3115
rect -436 -3187 -390 -3149
rect -436 -3221 -430 -3187
rect -396 -3221 -390 -3187
rect -436 -3259 -390 -3221
rect -436 -3293 -430 -3259
rect -396 -3293 -390 -3259
rect -436 -3331 -390 -3293
rect -436 -3365 -430 -3331
rect -396 -3365 -390 -3331
rect -436 -3403 -390 -3365
rect -436 -3437 -430 -3403
rect -396 -3437 -390 -3403
rect -436 -3475 -390 -3437
rect -436 -3509 -430 -3475
rect -396 -3509 -390 -3475
rect -436 -3547 -390 -3509
rect -436 -3581 -430 -3547
rect -396 -3581 -390 -3547
rect -436 -3619 -390 -3581
rect -436 -3653 -430 -3619
rect -396 -3653 -390 -3619
rect -436 -3691 -390 -3653
rect -436 -3725 -430 -3691
rect -396 -3725 -390 -3691
rect -436 -3763 -390 -3725
rect -436 -3797 -430 -3763
rect -396 -3797 -390 -3763
rect -436 -3835 -390 -3797
rect -436 -3869 -430 -3835
rect -396 -3869 -390 -3835
rect -436 -3907 -390 -3869
rect -436 -3941 -430 -3907
rect -396 -3941 -390 -3907
rect -436 -3979 -390 -3941
rect -436 -4013 -430 -3979
rect -396 -4013 -390 -3979
rect -436 -4051 -390 -4013
rect -436 -4085 -430 -4051
rect -396 -4085 -390 -4051
rect -436 -4123 -390 -4085
rect -436 -4157 -430 -4123
rect -396 -4157 -390 -4123
rect -436 -4195 -390 -4157
rect -436 -4229 -430 -4195
rect -396 -4229 -390 -4195
rect -436 -4267 -390 -4229
rect -436 -4301 -430 -4267
rect -396 -4301 -390 -4267
rect -436 -4339 -390 -4301
rect -436 -4373 -430 -4339
rect -396 -4373 -390 -4339
rect -436 -4411 -390 -4373
rect -436 -4445 -430 -4411
rect -396 -4445 -390 -4411
rect -436 -4483 -390 -4445
rect -436 -4517 -430 -4483
rect -396 -4517 -390 -4483
rect -436 -4555 -390 -4517
rect -436 -4589 -430 -4555
rect -396 -4589 -390 -4555
rect -436 -4627 -390 -4589
rect -436 -4661 -430 -4627
rect -396 -4661 -390 -4627
rect -436 -4699 -390 -4661
rect -436 -4733 -430 -4699
rect -396 -4733 -390 -4699
rect -436 -4771 -390 -4733
rect -436 -4805 -430 -4771
rect -396 -4805 -390 -4771
rect -436 -4843 -390 -4805
rect -436 -4877 -430 -4843
rect -396 -4877 -390 -4843
rect -436 -4915 -390 -4877
rect -436 -4949 -430 -4915
rect -396 -4949 -390 -4915
rect -436 -4987 -390 -4949
rect -436 -5021 -430 -4987
rect -396 -5021 -390 -4987
rect -436 -5059 -390 -5021
rect -436 -5093 -430 -5059
rect -396 -5093 -390 -5059
rect -436 -5131 -390 -5093
rect -436 -5165 -430 -5131
rect -396 -5165 -390 -5131
rect -436 -5203 -390 -5165
rect -436 -5237 -430 -5203
rect -396 -5237 -390 -5203
rect -436 -5275 -390 -5237
rect -436 -5309 -430 -5275
rect -396 -5309 -390 -5275
rect -436 -5347 -390 -5309
rect -436 -5381 -430 -5347
rect -396 -5381 -390 -5347
rect -436 -5419 -390 -5381
rect -436 -5453 -430 -5419
rect -396 -5453 -390 -5419
rect -436 -5491 -390 -5453
rect -436 -5525 -430 -5491
rect -396 -5525 -390 -5491
rect -436 -5563 -390 -5525
rect -436 -5597 -430 -5563
rect -396 -5597 -390 -5563
rect -436 -5635 -390 -5597
rect -436 -5669 -430 -5635
rect -396 -5669 -390 -5635
rect -436 -5707 -390 -5669
rect -436 -5741 -430 -5707
rect -396 -5741 -390 -5707
rect -436 -5779 -390 -5741
rect -436 -5813 -430 -5779
rect -396 -5813 -390 -5779
rect -436 -5851 -390 -5813
rect -436 -5885 -430 -5851
rect -396 -5885 -390 -5851
rect -436 -5923 -390 -5885
rect -436 -5957 -430 -5923
rect -396 -5957 -390 -5923
rect -436 -5995 -390 -5957
rect -436 -6029 -430 -5995
rect -396 -6029 -390 -5995
rect -436 -6067 -390 -6029
rect -436 -6101 -430 -6067
rect -396 -6101 -390 -6067
rect -436 -6139 -390 -6101
rect -436 -6173 -430 -6139
rect -396 -6173 -390 -6139
rect -436 -6211 -390 -6173
rect -436 -6245 -430 -6211
rect -396 -6245 -390 -6211
rect -436 -6283 -390 -6245
rect -436 -6317 -430 -6283
rect -396 -6317 -390 -6283
rect -436 -6355 -390 -6317
rect -436 -6389 -430 -6355
rect -396 -6389 -390 -6355
rect -436 -6427 -390 -6389
rect -436 -6461 -430 -6427
rect -396 -6461 -390 -6427
rect -436 -6499 -390 -6461
rect -436 -6533 -430 -6499
rect -396 -6533 -390 -6499
rect -436 -6571 -390 -6533
rect -436 -6605 -430 -6571
rect -396 -6605 -390 -6571
rect -436 -6643 -390 -6605
rect -436 -6677 -430 -6643
rect -396 -6677 -390 -6643
rect -436 -6715 -390 -6677
rect -436 -6749 -430 -6715
rect -396 -6749 -390 -6715
rect -436 -6787 -390 -6749
rect -436 -6821 -430 -6787
rect -396 -6821 -390 -6787
rect -436 -6859 -390 -6821
rect -436 -6893 -430 -6859
rect -396 -6893 -390 -6859
rect -436 -6931 -390 -6893
rect -436 -6965 -430 -6931
rect -396 -6965 -390 -6931
rect -436 -7003 -390 -6965
rect -436 -7037 -430 -7003
rect -396 -7037 -390 -7003
rect -436 -7075 -390 -7037
rect -436 -7109 -430 -7075
rect -396 -7109 -390 -7075
rect -436 -7147 -390 -7109
rect -436 -7181 -430 -7147
rect -396 -7181 -390 -7147
rect -436 -7219 -390 -7181
rect -436 -7253 -430 -7219
rect -396 -7253 -390 -7219
rect -436 -7291 -390 -7253
rect -436 -7325 -430 -7291
rect -396 -7325 -390 -7291
rect -436 -7363 -390 -7325
rect -436 -7397 -430 -7363
rect -396 -7397 -390 -7363
rect -436 -7435 -390 -7397
rect -436 -7469 -430 -7435
rect -396 -7469 -390 -7435
rect -436 -7507 -390 -7469
rect -436 -7541 -430 -7507
rect -396 -7541 -390 -7507
rect -436 -7579 -390 -7541
rect -436 -7613 -430 -7579
rect -396 -7613 -390 -7579
rect -436 -7651 -390 -7613
rect -436 -7685 -430 -7651
rect -396 -7685 -390 -7651
rect -436 -7723 -390 -7685
rect -436 -7757 -430 -7723
rect -396 -7757 -390 -7723
rect -436 -7795 -390 -7757
rect -436 -7829 -430 -7795
rect -396 -7829 -390 -7795
rect -436 -7867 -390 -7829
rect -436 -7901 -430 -7867
rect -396 -7901 -390 -7867
rect -436 -7939 -390 -7901
rect -436 -7973 -430 -7939
rect -396 -7973 -390 -7939
rect -436 -8011 -390 -7973
rect -436 -8045 -430 -8011
rect -396 -8045 -390 -8011
rect -436 -8083 -390 -8045
rect -436 -8117 -430 -8083
rect -396 -8117 -390 -8083
rect -436 -8155 -390 -8117
rect -436 -8189 -430 -8155
rect -396 -8189 -390 -8155
rect -436 -8227 -390 -8189
rect -436 -8261 -430 -8227
rect -396 -8261 -390 -8227
rect -436 -8299 -390 -8261
rect -436 -8333 -430 -8299
rect -396 -8333 -390 -8299
rect -436 -8371 -390 -8333
rect -436 -8405 -430 -8371
rect -396 -8405 -390 -8371
rect -436 -8443 -390 -8405
rect -436 -8477 -430 -8443
rect -396 -8477 -390 -8443
rect -436 -8515 -390 -8477
rect -436 -8549 -430 -8515
rect -396 -8549 -390 -8515
rect -436 -8587 -390 -8549
rect -436 -8621 -430 -8587
rect -396 -8621 -390 -8587
rect -436 -8659 -390 -8621
rect -436 -8693 -430 -8659
rect -396 -8693 -390 -8659
rect -436 -8731 -390 -8693
rect -436 -8765 -430 -8731
rect -396 -8765 -390 -8731
rect -436 -8803 -390 -8765
rect -436 -8837 -430 -8803
rect -396 -8837 -390 -8803
rect -436 -8875 -390 -8837
rect -436 -8909 -430 -8875
rect -396 -8909 -390 -8875
rect -436 -8947 -390 -8909
rect -436 -8981 -430 -8947
rect -396 -8981 -390 -8947
rect -436 -9019 -390 -8981
rect -436 -9053 -430 -9019
rect -396 -9053 -390 -9019
rect -436 -9091 -390 -9053
rect -436 -9125 -430 -9091
rect -396 -9125 -390 -9091
rect -436 -9163 -390 -9125
rect -436 -9197 -430 -9163
rect -396 -9197 -390 -9163
rect -436 -9235 -390 -9197
rect -436 -9269 -430 -9235
rect -396 -9269 -390 -9235
rect -436 -9307 -390 -9269
rect -436 -9341 -430 -9307
rect -396 -9341 -390 -9307
rect -436 -9379 -390 -9341
rect -436 -9413 -430 -9379
rect -396 -9413 -390 -9379
rect -436 -9451 -390 -9413
rect -436 -9485 -430 -9451
rect -396 -9485 -390 -9451
rect -436 -9523 -390 -9485
rect -436 -9557 -430 -9523
rect -396 -9557 -390 -9523
rect -436 -9600 -390 -9557
rect -318 9557 -272 9600
rect -318 9523 -312 9557
rect -278 9523 -272 9557
rect -318 9485 -272 9523
rect -318 9451 -312 9485
rect -278 9451 -272 9485
rect -318 9413 -272 9451
rect -318 9379 -312 9413
rect -278 9379 -272 9413
rect -318 9341 -272 9379
rect -318 9307 -312 9341
rect -278 9307 -272 9341
rect -318 9269 -272 9307
rect -318 9235 -312 9269
rect -278 9235 -272 9269
rect -318 9197 -272 9235
rect -318 9163 -312 9197
rect -278 9163 -272 9197
rect -318 9125 -272 9163
rect -318 9091 -312 9125
rect -278 9091 -272 9125
rect -318 9053 -272 9091
rect -318 9019 -312 9053
rect -278 9019 -272 9053
rect -318 8981 -272 9019
rect -318 8947 -312 8981
rect -278 8947 -272 8981
rect -318 8909 -272 8947
rect -318 8875 -312 8909
rect -278 8875 -272 8909
rect -318 8837 -272 8875
rect -318 8803 -312 8837
rect -278 8803 -272 8837
rect -318 8765 -272 8803
rect -318 8731 -312 8765
rect -278 8731 -272 8765
rect -318 8693 -272 8731
rect -318 8659 -312 8693
rect -278 8659 -272 8693
rect -318 8621 -272 8659
rect -318 8587 -312 8621
rect -278 8587 -272 8621
rect -318 8549 -272 8587
rect -318 8515 -312 8549
rect -278 8515 -272 8549
rect -318 8477 -272 8515
rect -318 8443 -312 8477
rect -278 8443 -272 8477
rect -318 8405 -272 8443
rect -318 8371 -312 8405
rect -278 8371 -272 8405
rect -318 8333 -272 8371
rect -318 8299 -312 8333
rect -278 8299 -272 8333
rect -318 8261 -272 8299
rect -318 8227 -312 8261
rect -278 8227 -272 8261
rect -318 8189 -272 8227
rect -318 8155 -312 8189
rect -278 8155 -272 8189
rect -318 8117 -272 8155
rect -318 8083 -312 8117
rect -278 8083 -272 8117
rect -318 8045 -272 8083
rect -318 8011 -312 8045
rect -278 8011 -272 8045
rect -318 7973 -272 8011
rect -318 7939 -312 7973
rect -278 7939 -272 7973
rect -318 7901 -272 7939
rect -318 7867 -312 7901
rect -278 7867 -272 7901
rect -318 7829 -272 7867
rect -318 7795 -312 7829
rect -278 7795 -272 7829
rect -318 7757 -272 7795
rect -318 7723 -312 7757
rect -278 7723 -272 7757
rect -318 7685 -272 7723
rect -318 7651 -312 7685
rect -278 7651 -272 7685
rect -318 7613 -272 7651
rect -318 7579 -312 7613
rect -278 7579 -272 7613
rect -318 7541 -272 7579
rect -318 7507 -312 7541
rect -278 7507 -272 7541
rect -318 7469 -272 7507
rect -318 7435 -312 7469
rect -278 7435 -272 7469
rect -318 7397 -272 7435
rect -318 7363 -312 7397
rect -278 7363 -272 7397
rect -318 7325 -272 7363
rect -318 7291 -312 7325
rect -278 7291 -272 7325
rect -318 7253 -272 7291
rect -318 7219 -312 7253
rect -278 7219 -272 7253
rect -318 7181 -272 7219
rect -318 7147 -312 7181
rect -278 7147 -272 7181
rect -318 7109 -272 7147
rect -318 7075 -312 7109
rect -278 7075 -272 7109
rect -318 7037 -272 7075
rect -318 7003 -312 7037
rect -278 7003 -272 7037
rect -318 6965 -272 7003
rect -318 6931 -312 6965
rect -278 6931 -272 6965
rect -318 6893 -272 6931
rect -318 6859 -312 6893
rect -278 6859 -272 6893
rect -318 6821 -272 6859
rect -318 6787 -312 6821
rect -278 6787 -272 6821
rect -318 6749 -272 6787
rect -318 6715 -312 6749
rect -278 6715 -272 6749
rect -318 6677 -272 6715
rect -318 6643 -312 6677
rect -278 6643 -272 6677
rect -318 6605 -272 6643
rect -318 6571 -312 6605
rect -278 6571 -272 6605
rect -318 6533 -272 6571
rect -318 6499 -312 6533
rect -278 6499 -272 6533
rect -318 6461 -272 6499
rect -318 6427 -312 6461
rect -278 6427 -272 6461
rect -318 6389 -272 6427
rect -318 6355 -312 6389
rect -278 6355 -272 6389
rect -318 6317 -272 6355
rect -318 6283 -312 6317
rect -278 6283 -272 6317
rect -318 6245 -272 6283
rect -318 6211 -312 6245
rect -278 6211 -272 6245
rect -318 6173 -272 6211
rect -318 6139 -312 6173
rect -278 6139 -272 6173
rect -318 6101 -272 6139
rect -318 6067 -312 6101
rect -278 6067 -272 6101
rect -318 6029 -272 6067
rect -318 5995 -312 6029
rect -278 5995 -272 6029
rect -318 5957 -272 5995
rect -318 5923 -312 5957
rect -278 5923 -272 5957
rect -318 5885 -272 5923
rect -318 5851 -312 5885
rect -278 5851 -272 5885
rect -318 5813 -272 5851
rect -318 5779 -312 5813
rect -278 5779 -272 5813
rect -318 5741 -272 5779
rect -318 5707 -312 5741
rect -278 5707 -272 5741
rect -318 5669 -272 5707
rect -318 5635 -312 5669
rect -278 5635 -272 5669
rect -318 5597 -272 5635
rect -318 5563 -312 5597
rect -278 5563 -272 5597
rect -318 5525 -272 5563
rect -318 5491 -312 5525
rect -278 5491 -272 5525
rect -318 5453 -272 5491
rect -318 5419 -312 5453
rect -278 5419 -272 5453
rect -318 5381 -272 5419
rect -318 5347 -312 5381
rect -278 5347 -272 5381
rect -318 5309 -272 5347
rect -318 5275 -312 5309
rect -278 5275 -272 5309
rect -318 5237 -272 5275
rect -318 5203 -312 5237
rect -278 5203 -272 5237
rect -318 5165 -272 5203
rect -318 5131 -312 5165
rect -278 5131 -272 5165
rect -318 5093 -272 5131
rect -318 5059 -312 5093
rect -278 5059 -272 5093
rect -318 5021 -272 5059
rect -318 4987 -312 5021
rect -278 4987 -272 5021
rect -318 4949 -272 4987
rect -318 4915 -312 4949
rect -278 4915 -272 4949
rect -318 4877 -272 4915
rect -318 4843 -312 4877
rect -278 4843 -272 4877
rect -318 4805 -272 4843
rect -318 4771 -312 4805
rect -278 4771 -272 4805
rect -318 4733 -272 4771
rect -318 4699 -312 4733
rect -278 4699 -272 4733
rect -318 4661 -272 4699
rect -318 4627 -312 4661
rect -278 4627 -272 4661
rect -318 4589 -272 4627
rect -318 4555 -312 4589
rect -278 4555 -272 4589
rect -318 4517 -272 4555
rect -318 4483 -312 4517
rect -278 4483 -272 4517
rect -318 4445 -272 4483
rect -318 4411 -312 4445
rect -278 4411 -272 4445
rect -318 4373 -272 4411
rect -318 4339 -312 4373
rect -278 4339 -272 4373
rect -318 4301 -272 4339
rect -318 4267 -312 4301
rect -278 4267 -272 4301
rect -318 4229 -272 4267
rect -318 4195 -312 4229
rect -278 4195 -272 4229
rect -318 4157 -272 4195
rect -318 4123 -312 4157
rect -278 4123 -272 4157
rect -318 4085 -272 4123
rect -318 4051 -312 4085
rect -278 4051 -272 4085
rect -318 4013 -272 4051
rect -318 3979 -312 4013
rect -278 3979 -272 4013
rect -318 3941 -272 3979
rect -318 3907 -312 3941
rect -278 3907 -272 3941
rect -318 3869 -272 3907
rect -318 3835 -312 3869
rect -278 3835 -272 3869
rect -318 3797 -272 3835
rect -318 3763 -312 3797
rect -278 3763 -272 3797
rect -318 3725 -272 3763
rect -318 3691 -312 3725
rect -278 3691 -272 3725
rect -318 3653 -272 3691
rect -318 3619 -312 3653
rect -278 3619 -272 3653
rect -318 3581 -272 3619
rect -318 3547 -312 3581
rect -278 3547 -272 3581
rect -318 3509 -272 3547
rect -318 3475 -312 3509
rect -278 3475 -272 3509
rect -318 3437 -272 3475
rect -318 3403 -312 3437
rect -278 3403 -272 3437
rect -318 3365 -272 3403
rect -318 3331 -312 3365
rect -278 3331 -272 3365
rect -318 3293 -272 3331
rect -318 3259 -312 3293
rect -278 3259 -272 3293
rect -318 3221 -272 3259
rect -318 3187 -312 3221
rect -278 3187 -272 3221
rect -318 3149 -272 3187
rect -318 3115 -312 3149
rect -278 3115 -272 3149
rect -318 3077 -272 3115
rect -318 3043 -312 3077
rect -278 3043 -272 3077
rect -318 3005 -272 3043
rect -318 2971 -312 3005
rect -278 2971 -272 3005
rect -318 2933 -272 2971
rect -318 2899 -312 2933
rect -278 2899 -272 2933
rect -318 2861 -272 2899
rect -318 2827 -312 2861
rect -278 2827 -272 2861
rect -318 2789 -272 2827
rect -318 2755 -312 2789
rect -278 2755 -272 2789
rect -318 2717 -272 2755
rect -318 2683 -312 2717
rect -278 2683 -272 2717
rect -318 2645 -272 2683
rect -318 2611 -312 2645
rect -278 2611 -272 2645
rect -318 2573 -272 2611
rect -318 2539 -312 2573
rect -278 2539 -272 2573
rect -318 2501 -272 2539
rect -318 2467 -312 2501
rect -278 2467 -272 2501
rect -318 2429 -272 2467
rect -318 2395 -312 2429
rect -278 2395 -272 2429
rect -318 2357 -272 2395
rect -318 2323 -312 2357
rect -278 2323 -272 2357
rect -318 2285 -272 2323
rect -318 2251 -312 2285
rect -278 2251 -272 2285
rect -318 2213 -272 2251
rect -318 2179 -312 2213
rect -278 2179 -272 2213
rect -318 2141 -272 2179
rect -318 2107 -312 2141
rect -278 2107 -272 2141
rect -318 2069 -272 2107
rect -318 2035 -312 2069
rect -278 2035 -272 2069
rect -318 1997 -272 2035
rect -318 1963 -312 1997
rect -278 1963 -272 1997
rect -318 1925 -272 1963
rect -318 1891 -312 1925
rect -278 1891 -272 1925
rect -318 1853 -272 1891
rect -318 1819 -312 1853
rect -278 1819 -272 1853
rect -318 1781 -272 1819
rect -318 1747 -312 1781
rect -278 1747 -272 1781
rect -318 1709 -272 1747
rect -318 1675 -312 1709
rect -278 1675 -272 1709
rect -318 1637 -272 1675
rect -318 1603 -312 1637
rect -278 1603 -272 1637
rect -318 1565 -272 1603
rect -318 1531 -312 1565
rect -278 1531 -272 1565
rect -318 1493 -272 1531
rect -318 1459 -312 1493
rect -278 1459 -272 1493
rect -318 1421 -272 1459
rect -318 1387 -312 1421
rect -278 1387 -272 1421
rect -318 1349 -272 1387
rect -318 1315 -312 1349
rect -278 1315 -272 1349
rect -318 1277 -272 1315
rect -318 1243 -312 1277
rect -278 1243 -272 1277
rect -318 1205 -272 1243
rect -318 1171 -312 1205
rect -278 1171 -272 1205
rect -318 1133 -272 1171
rect -318 1099 -312 1133
rect -278 1099 -272 1133
rect -318 1061 -272 1099
rect -318 1027 -312 1061
rect -278 1027 -272 1061
rect -318 989 -272 1027
rect -318 955 -312 989
rect -278 955 -272 989
rect -318 917 -272 955
rect -318 883 -312 917
rect -278 883 -272 917
rect -318 845 -272 883
rect -318 811 -312 845
rect -278 811 -272 845
rect -318 773 -272 811
rect -318 739 -312 773
rect -278 739 -272 773
rect -318 701 -272 739
rect -318 667 -312 701
rect -278 667 -272 701
rect -318 629 -272 667
rect -318 595 -312 629
rect -278 595 -272 629
rect -318 557 -272 595
rect -318 523 -312 557
rect -278 523 -272 557
rect -318 485 -272 523
rect -318 451 -312 485
rect -278 451 -272 485
rect -318 413 -272 451
rect -318 379 -312 413
rect -278 379 -272 413
rect -318 341 -272 379
rect -318 307 -312 341
rect -278 307 -272 341
rect -318 269 -272 307
rect -318 235 -312 269
rect -278 235 -272 269
rect -318 197 -272 235
rect -318 163 -312 197
rect -278 163 -272 197
rect -318 125 -272 163
rect -318 91 -312 125
rect -278 91 -272 125
rect -318 53 -272 91
rect -318 19 -312 53
rect -278 19 -272 53
rect -318 -19 -272 19
rect -318 -53 -312 -19
rect -278 -53 -272 -19
rect -318 -91 -272 -53
rect -318 -125 -312 -91
rect -278 -125 -272 -91
rect -318 -163 -272 -125
rect -318 -197 -312 -163
rect -278 -197 -272 -163
rect -318 -235 -272 -197
rect -318 -269 -312 -235
rect -278 -269 -272 -235
rect -318 -307 -272 -269
rect -318 -341 -312 -307
rect -278 -341 -272 -307
rect -318 -379 -272 -341
rect -318 -413 -312 -379
rect -278 -413 -272 -379
rect -318 -451 -272 -413
rect -318 -485 -312 -451
rect -278 -485 -272 -451
rect -318 -523 -272 -485
rect -318 -557 -312 -523
rect -278 -557 -272 -523
rect -318 -595 -272 -557
rect -318 -629 -312 -595
rect -278 -629 -272 -595
rect -318 -667 -272 -629
rect -318 -701 -312 -667
rect -278 -701 -272 -667
rect -318 -739 -272 -701
rect -318 -773 -312 -739
rect -278 -773 -272 -739
rect -318 -811 -272 -773
rect -318 -845 -312 -811
rect -278 -845 -272 -811
rect -318 -883 -272 -845
rect -318 -917 -312 -883
rect -278 -917 -272 -883
rect -318 -955 -272 -917
rect -318 -989 -312 -955
rect -278 -989 -272 -955
rect -318 -1027 -272 -989
rect -318 -1061 -312 -1027
rect -278 -1061 -272 -1027
rect -318 -1099 -272 -1061
rect -318 -1133 -312 -1099
rect -278 -1133 -272 -1099
rect -318 -1171 -272 -1133
rect -318 -1205 -312 -1171
rect -278 -1205 -272 -1171
rect -318 -1243 -272 -1205
rect -318 -1277 -312 -1243
rect -278 -1277 -272 -1243
rect -318 -1315 -272 -1277
rect -318 -1349 -312 -1315
rect -278 -1349 -272 -1315
rect -318 -1387 -272 -1349
rect -318 -1421 -312 -1387
rect -278 -1421 -272 -1387
rect -318 -1459 -272 -1421
rect -318 -1493 -312 -1459
rect -278 -1493 -272 -1459
rect -318 -1531 -272 -1493
rect -318 -1565 -312 -1531
rect -278 -1565 -272 -1531
rect -318 -1603 -272 -1565
rect -318 -1637 -312 -1603
rect -278 -1637 -272 -1603
rect -318 -1675 -272 -1637
rect -318 -1709 -312 -1675
rect -278 -1709 -272 -1675
rect -318 -1747 -272 -1709
rect -318 -1781 -312 -1747
rect -278 -1781 -272 -1747
rect -318 -1819 -272 -1781
rect -318 -1853 -312 -1819
rect -278 -1853 -272 -1819
rect -318 -1891 -272 -1853
rect -318 -1925 -312 -1891
rect -278 -1925 -272 -1891
rect -318 -1963 -272 -1925
rect -318 -1997 -312 -1963
rect -278 -1997 -272 -1963
rect -318 -2035 -272 -1997
rect -318 -2069 -312 -2035
rect -278 -2069 -272 -2035
rect -318 -2107 -272 -2069
rect -318 -2141 -312 -2107
rect -278 -2141 -272 -2107
rect -318 -2179 -272 -2141
rect -318 -2213 -312 -2179
rect -278 -2213 -272 -2179
rect -318 -2251 -272 -2213
rect -318 -2285 -312 -2251
rect -278 -2285 -272 -2251
rect -318 -2323 -272 -2285
rect -318 -2357 -312 -2323
rect -278 -2357 -272 -2323
rect -318 -2395 -272 -2357
rect -318 -2429 -312 -2395
rect -278 -2429 -272 -2395
rect -318 -2467 -272 -2429
rect -318 -2501 -312 -2467
rect -278 -2501 -272 -2467
rect -318 -2539 -272 -2501
rect -318 -2573 -312 -2539
rect -278 -2573 -272 -2539
rect -318 -2611 -272 -2573
rect -318 -2645 -312 -2611
rect -278 -2645 -272 -2611
rect -318 -2683 -272 -2645
rect -318 -2717 -312 -2683
rect -278 -2717 -272 -2683
rect -318 -2755 -272 -2717
rect -318 -2789 -312 -2755
rect -278 -2789 -272 -2755
rect -318 -2827 -272 -2789
rect -318 -2861 -312 -2827
rect -278 -2861 -272 -2827
rect -318 -2899 -272 -2861
rect -318 -2933 -312 -2899
rect -278 -2933 -272 -2899
rect -318 -2971 -272 -2933
rect -318 -3005 -312 -2971
rect -278 -3005 -272 -2971
rect -318 -3043 -272 -3005
rect -318 -3077 -312 -3043
rect -278 -3077 -272 -3043
rect -318 -3115 -272 -3077
rect -318 -3149 -312 -3115
rect -278 -3149 -272 -3115
rect -318 -3187 -272 -3149
rect -318 -3221 -312 -3187
rect -278 -3221 -272 -3187
rect -318 -3259 -272 -3221
rect -318 -3293 -312 -3259
rect -278 -3293 -272 -3259
rect -318 -3331 -272 -3293
rect -318 -3365 -312 -3331
rect -278 -3365 -272 -3331
rect -318 -3403 -272 -3365
rect -318 -3437 -312 -3403
rect -278 -3437 -272 -3403
rect -318 -3475 -272 -3437
rect -318 -3509 -312 -3475
rect -278 -3509 -272 -3475
rect -318 -3547 -272 -3509
rect -318 -3581 -312 -3547
rect -278 -3581 -272 -3547
rect -318 -3619 -272 -3581
rect -318 -3653 -312 -3619
rect -278 -3653 -272 -3619
rect -318 -3691 -272 -3653
rect -318 -3725 -312 -3691
rect -278 -3725 -272 -3691
rect -318 -3763 -272 -3725
rect -318 -3797 -312 -3763
rect -278 -3797 -272 -3763
rect -318 -3835 -272 -3797
rect -318 -3869 -312 -3835
rect -278 -3869 -272 -3835
rect -318 -3907 -272 -3869
rect -318 -3941 -312 -3907
rect -278 -3941 -272 -3907
rect -318 -3979 -272 -3941
rect -318 -4013 -312 -3979
rect -278 -4013 -272 -3979
rect -318 -4051 -272 -4013
rect -318 -4085 -312 -4051
rect -278 -4085 -272 -4051
rect -318 -4123 -272 -4085
rect -318 -4157 -312 -4123
rect -278 -4157 -272 -4123
rect -318 -4195 -272 -4157
rect -318 -4229 -312 -4195
rect -278 -4229 -272 -4195
rect -318 -4267 -272 -4229
rect -318 -4301 -312 -4267
rect -278 -4301 -272 -4267
rect -318 -4339 -272 -4301
rect -318 -4373 -312 -4339
rect -278 -4373 -272 -4339
rect -318 -4411 -272 -4373
rect -318 -4445 -312 -4411
rect -278 -4445 -272 -4411
rect -318 -4483 -272 -4445
rect -318 -4517 -312 -4483
rect -278 -4517 -272 -4483
rect -318 -4555 -272 -4517
rect -318 -4589 -312 -4555
rect -278 -4589 -272 -4555
rect -318 -4627 -272 -4589
rect -318 -4661 -312 -4627
rect -278 -4661 -272 -4627
rect -318 -4699 -272 -4661
rect -318 -4733 -312 -4699
rect -278 -4733 -272 -4699
rect -318 -4771 -272 -4733
rect -318 -4805 -312 -4771
rect -278 -4805 -272 -4771
rect -318 -4843 -272 -4805
rect -318 -4877 -312 -4843
rect -278 -4877 -272 -4843
rect -318 -4915 -272 -4877
rect -318 -4949 -312 -4915
rect -278 -4949 -272 -4915
rect -318 -4987 -272 -4949
rect -318 -5021 -312 -4987
rect -278 -5021 -272 -4987
rect -318 -5059 -272 -5021
rect -318 -5093 -312 -5059
rect -278 -5093 -272 -5059
rect -318 -5131 -272 -5093
rect -318 -5165 -312 -5131
rect -278 -5165 -272 -5131
rect -318 -5203 -272 -5165
rect -318 -5237 -312 -5203
rect -278 -5237 -272 -5203
rect -318 -5275 -272 -5237
rect -318 -5309 -312 -5275
rect -278 -5309 -272 -5275
rect -318 -5347 -272 -5309
rect -318 -5381 -312 -5347
rect -278 -5381 -272 -5347
rect -318 -5419 -272 -5381
rect -318 -5453 -312 -5419
rect -278 -5453 -272 -5419
rect -318 -5491 -272 -5453
rect -318 -5525 -312 -5491
rect -278 -5525 -272 -5491
rect -318 -5563 -272 -5525
rect -318 -5597 -312 -5563
rect -278 -5597 -272 -5563
rect -318 -5635 -272 -5597
rect -318 -5669 -312 -5635
rect -278 -5669 -272 -5635
rect -318 -5707 -272 -5669
rect -318 -5741 -312 -5707
rect -278 -5741 -272 -5707
rect -318 -5779 -272 -5741
rect -318 -5813 -312 -5779
rect -278 -5813 -272 -5779
rect -318 -5851 -272 -5813
rect -318 -5885 -312 -5851
rect -278 -5885 -272 -5851
rect -318 -5923 -272 -5885
rect -318 -5957 -312 -5923
rect -278 -5957 -272 -5923
rect -318 -5995 -272 -5957
rect -318 -6029 -312 -5995
rect -278 -6029 -272 -5995
rect -318 -6067 -272 -6029
rect -318 -6101 -312 -6067
rect -278 -6101 -272 -6067
rect -318 -6139 -272 -6101
rect -318 -6173 -312 -6139
rect -278 -6173 -272 -6139
rect -318 -6211 -272 -6173
rect -318 -6245 -312 -6211
rect -278 -6245 -272 -6211
rect -318 -6283 -272 -6245
rect -318 -6317 -312 -6283
rect -278 -6317 -272 -6283
rect -318 -6355 -272 -6317
rect -318 -6389 -312 -6355
rect -278 -6389 -272 -6355
rect -318 -6427 -272 -6389
rect -318 -6461 -312 -6427
rect -278 -6461 -272 -6427
rect -318 -6499 -272 -6461
rect -318 -6533 -312 -6499
rect -278 -6533 -272 -6499
rect -318 -6571 -272 -6533
rect -318 -6605 -312 -6571
rect -278 -6605 -272 -6571
rect -318 -6643 -272 -6605
rect -318 -6677 -312 -6643
rect -278 -6677 -272 -6643
rect -318 -6715 -272 -6677
rect -318 -6749 -312 -6715
rect -278 -6749 -272 -6715
rect -318 -6787 -272 -6749
rect -318 -6821 -312 -6787
rect -278 -6821 -272 -6787
rect -318 -6859 -272 -6821
rect -318 -6893 -312 -6859
rect -278 -6893 -272 -6859
rect -318 -6931 -272 -6893
rect -318 -6965 -312 -6931
rect -278 -6965 -272 -6931
rect -318 -7003 -272 -6965
rect -318 -7037 -312 -7003
rect -278 -7037 -272 -7003
rect -318 -7075 -272 -7037
rect -318 -7109 -312 -7075
rect -278 -7109 -272 -7075
rect -318 -7147 -272 -7109
rect -318 -7181 -312 -7147
rect -278 -7181 -272 -7147
rect -318 -7219 -272 -7181
rect -318 -7253 -312 -7219
rect -278 -7253 -272 -7219
rect -318 -7291 -272 -7253
rect -318 -7325 -312 -7291
rect -278 -7325 -272 -7291
rect -318 -7363 -272 -7325
rect -318 -7397 -312 -7363
rect -278 -7397 -272 -7363
rect -318 -7435 -272 -7397
rect -318 -7469 -312 -7435
rect -278 -7469 -272 -7435
rect -318 -7507 -272 -7469
rect -318 -7541 -312 -7507
rect -278 -7541 -272 -7507
rect -318 -7579 -272 -7541
rect -318 -7613 -312 -7579
rect -278 -7613 -272 -7579
rect -318 -7651 -272 -7613
rect -318 -7685 -312 -7651
rect -278 -7685 -272 -7651
rect -318 -7723 -272 -7685
rect -318 -7757 -312 -7723
rect -278 -7757 -272 -7723
rect -318 -7795 -272 -7757
rect -318 -7829 -312 -7795
rect -278 -7829 -272 -7795
rect -318 -7867 -272 -7829
rect -318 -7901 -312 -7867
rect -278 -7901 -272 -7867
rect -318 -7939 -272 -7901
rect -318 -7973 -312 -7939
rect -278 -7973 -272 -7939
rect -318 -8011 -272 -7973
rect -318 -8045 -312 -8011
rect -278 -8045 -272 -8011
rect -318 -8083 -272 -8045
rect -318 -8117 -312 -8083
rect -278 -8117 -272 -8083
rect -318 -8155 -272 -8117
rect -318 -8189 -312 -8155
rect -278 -8189 -272 -8155
rect -318 -8227 -272 -8189
rect -318 -8261 -312 -8227
rect -278 -8261 -272 -8227
rect -318 -8299 -272 -8261
rect -318 -8333 -312 -8299
rect -278 -8333 -272 -8299
rect -318 -8371 -272 -8333
rect -318 -8405 -312 -8371
rect -278 -8405 -272 -8371
rect -318 -8443 -272 -8405
rect -318 -8477 -312 -8443
rect -278 -8477 -272 -8443
rect -318 -8515 -272 -8477
rect -318 -8549 -312 -8515
rect -278 -8549 -272 -8515
rect -318 -8587 -272 -8549
rect -318 -8621 -312 -8587
rect -278 -8621 -272 -8587
rect -318 -8659 -272 -8621
rect -318 -8693 -312 -8659
rect -278 -8693 -272 -8659
rect -318 -8731 -272 -8693
rect -318 -8765 -312 -8731
rect -278 -8765 -272 -8731
rect -318 -8803 -272 -8765
rect -318 -8837 -312 -8803
rect -278 -8837 -272 -8803
rect -318 -8875 -272 -8837
rect -318 -8909 -312 -8875
rect -278 -8909 -272 -8875
rect -318 -8947 -272 -8909
rect -318 -8981 -312 -8947
rect -278 -8981 -272 -8947
rect -318 -9019 -272 -8981
rect -318 -9053 -312 -9019
rect -278 -9053 -272 -9019
rect -318 -9091 -272 -9053
rect -318 -9125 -312 -9091
rect -278 -9125 -272 -9091
rect -318 -9163 -272 -9125
rect -318 -9197 -312 -9163
rect -278 -9197 -272 -9163
rect -318 -9235 -272 -9197
rect -318 -9269 -312 -9235
rect -278 -9269 -272 -9235
rect -318 -9307 -272 -9269
rect -318 -9341 -312 -9307
rect -278 -9341 -272 -9307
rect -318 -9379 -272 -9341
rect -318 -9413 -312 -9379
rect -278 -9413 -272 -9379
rect -318 -9451 -272 -9413
rect -318 -9485 -312 -9451
rect -278 -9485 -272 -9451
rect -318 -9523 -272 -9485
rect -318 -9557 -312 -9523
rect -278 -9557 -272 -9523
rect -318 -9600 -272 -9557
rect -200 9557 -154 9600
rect -200 9523 -194 9557
rect -160 9523 -154 9557
rect -200 9485 -154 9523
rect -200 9451 -194 9485
rect -160 9451 -154 9485
rect -200 9413 -154 9451
rect -200 9379 -194 9413
rect -160 9379 -154 9413
rect -200 9341 -154 9379
rect -200 9307 -194 9341
rect -160 9307 -154 9341
rect -200 9269 -154 9307
rect -200 9235 -194 9269
rect -160 9235 -154 9269
rect -200 9197 -154 9235
rect -200 9163 -194 9197
rect -160 9163 -154 9197
rect -200 9125 -154 9163
rect -200 9091 -194 9125
rect -160 9091 -154 9125
rect -200 9053 -154 9091
rect -200 9019 -194 9053
rect -160 9019 -154 9053
rect -200 8981 -154 9019
rect -200 8947 -194 8981
rect -160 8947 -154 8981
rect -200 8909 -154 8947
rect -200 8875 -194 8909
rect -160 8875 -154 8909
rect -200 8837 -154 8875
rect -200 8803 -194 8837
rect -160 8803 -154 8837
rect -200 8765 -154 8803
rect -200 8731 -194 8765
rect -160 8731 -154 8765
rect -200 8693 -154 8731
rect -200 8659 -194 8693
rect -160 8659 -154 8693
rect -200 8621 -154 8659
rect -200 8587 -194 8621
rect -160 8587 -154 8621
rect -200 8549 -154 8587
rect -200 8515 -194 8549
rect -160 8515 -154 8549
rect -200 8477 -154 8515
rect -200 8443 -194 8477
rect -160 8443 -154 8477
rect -200 8405 -154 8443
rect -200 8371 -194 8405
rect -160 8371 -154 8405
rect -200 8333 -154 8371
rect -200 8299 -194 8333
rect -160 8299 -154 8333
rect -200 8261 -154 8299
rect -200 8227 -194 8261
rect -160 8227 -154 8261
rect -200 8189 -154 8227
rect -200 8155 -194 8189
rect -160 8155 -154 8189
rect -200 8117 -154 8155
rect -200 8083 -194 8117
rect -160 8083 -154 8117
rect -200 8045 -154 8083
rect -200 8011 -194 8045
rect -160 8011 -154 8045
rect -200 7973 -154 8011
rect -200 7939 -194 7973
rect -160 7939 -154 7973
rect -200 7901 -154 7939
rect -200 7867 -194 7901
rect -160 7867 -154 7901
rect -200 7829 -154 7867
rect -200 7795 -194 7829
rect -160 7795 -154 7829
rect -200 7757 -154 7795
rect -200 7723 -194 7757
rect -160 7723 -154 7757
rect -200 7685 -154 7723
rect -200 7651 -194 7685
rect -160 7651 -154 7685
rect -200 7613 -154 7651
rect -200 7579 -194 7613
rect -160 7579 -154 7613
rect -200 7541 -154 7579
rect -200 7507 -194 7541
rect -160 7507 -154 7541
rect -200 7469 -154 7507
rect -200 7435 -194 7469
rect -160 7435 -154 7469
rect -200 7397 -154 7435
rect -200 7363 -194 7397
rect -160 7363 -154 7397
rect -200 7325 -154 7363
rect -200 7291 -194 7325
rect -160 7291 -154 7325
rect -200 7253 -154 7291
rect -200 7219 -194 7253
rect -160 7219 -154 7253
rect -200 7181 -154 7219
rect -200 7147 -194 7181
rect -160 7147 -154 7181
rect -200 7109 -154 7147
rect -200 7075 -194 7109
rect -160 7075 -154 7109
rect -200 7037 -154 7075
rect -200 7003 -194 7037
rect -160 7003 -154 7037
rect -200 6965 -154 7003
rect -200 6931 -194 6965
rect -160 6931 -154 6965
rect -200 6893 -154 6931
rect -200 6859 -194 6893
rect -160 6859 -154 6893
rect -200 6821 -154 6859
rect -200 6787 -194 6821
rect -160 6787 -154 6821
rect -200 6749 -154 6787
rect -200 6715 -194 6749
rect -160 6715 -154 6749
rect -200 6677 -154 6715
rect -200 6643 -194 6677
rect -160 6643 -154 6677
rect -200 6605 -154 6643
rect -200 6571 -194 6605
rect -160 6571 -154 6605
rect -200 6533 -154 6571
rect -200 6499 -194 6533
rect -160 6499 -154 6533
rect -200 6461 -154 6499
rect -200 6427 -194 6461
rect -160 6427 -154 6461
rect -200 6389 -154 6427
rect -200 6355 -194 6389
rect -160 6355 -154 6389
rect -200 6317 -154 6355
rect -200 6283 -194 6317
rect -160 6283 -154 6317
rect -200 6245 -154 6283
rect -200 6211 -194 6245
rect -160 6211 -154 6245
rect -200 6173 -154 6211
rect -200 6139 -194 6173
rect -160 6139 -154 6173
rect -200 6101 -154 6139
rect -200 6067 -194 6101
rect -160 6067 -154 6101
rect -200 6029 -154 6067
rect -200 5995 -194 6029
rect -160 5995 -154 6029
rect -200 5957 -154 5995
rect -200 5923 -194 5957
rect -160 5923 -154 5957
rect -200 5885 -154 5923
rect -200 5851 -194 5885
rect -160 5851 -154 5885
rect -200 5813 -154 5851
rect -200 5779 -194 5813
rect -160 5779 -154 5813
rect -200 5741 -154 5779
rect -200 5707 -194 5741
rect -160 5707 -154 5741
rect -200 5669 -154 5707
rect -200 5635 -194 5669
rect -160 5635 -154 5669
rect -200 5597 -154 5635
rect -200 5563 -194 5597
rect -160 5563 -154 5597
rect -200 5525 -154 5563
rect -200 5491 -194 5525
rect -160 5491 -154 5525
rect -200 5453 -154 5491
rect -200 5419 -194 5453
rect -160 5419 -154 5453
rect -200 5381 -154 5419
rect -200 5347 -194 5381
rect -160 5347 -154 5381
rect -200 5309 -154 5347
rect -200 5275 -194 5309
rect -160 5275 -154 5309
rect -200 5237 -154 5275
rect -200 5203 -194 5237
rect -160 5203 -154 5237
rect -200 5165 -154 5203
rect -200 5131 -194 5165
rect -160 5131 -154 5165
rect -200 5093 -154 5131
rect -200 5059 -194 5093
rect -160 5059 -154 5093
rect -200 5021 -154 5059
rect -200 4987 -194 5021
rect -160 4987 -154 5021
rect -200 4949 -154 4987
rect -200 4915 -194 4949
rect -160 4915 -154 4949
rect -200 4877 -154 4915
rect -200 4843 -194 4877
rect -160 4843 -154 4877
rect -200 4805 -154 4843
rect -200 4771 -194 4805
rect -160 4771 -154 4805
rect -200 4733 -154 4771
rect -200 4699 -194 4733
rect -160 4699 -154 4733
rect -200 4661 -154 4699
rect -200 4627 -194 4661
rect -160 4627 -154 4661
rect -200 4589 -154 4627
rect -200 4555 -194 4589
rect -160 4555 -154 4589
rect -200 4517 -154 4555
rect -200 4483 -194 4517
rect -160 4483 -154 4517
rect -200 4445 -154 4483
rect -200 4411 -194 4445
rect -160 4411 -154 4445
rect -200 4373 -154 4411
rect -200 4339 -194 4373
rect -160 4339 -154 4373
rect -200 4301 -154 4339
rect -200 4267 -194 4301
rect -160 4267 -154 4301
rect -200 4229 -154 4267
rect -200 4195 -194 4229
rect -160 4195 -154 4229
rect -200 4157 -154 4195
rect -200 4123 -194 4157
rect -160 4123 -154 4157
rect -200 4085 -154 4123
rect -200 4051 -194 4085
rect -160 4051 -154 4085
rect -200 4013 -154 4051
rect -200 3979 -194 4013
rect -160 3979 -154 4013
rect -200 3941 -154 3979
rect -200 3907 -194 3941
rect -160 3907 -154 3941
rect -200 3869 -154 3907
rect -200 3835 -194 3869
rect -160 3835 -154 3869
rect -200 3797 -154 3835
rect -200 3763 -194 3797
rect -160 3763 -154 3797
rect -200 3725 -154 3763
rect -200 3691 -194 3725
rect -160 3691 -154 3725
rect -200 3653 -154 3691
rect -200 3619 -194 3653
rect -160 3619 -154 3653
rect -200 3581 -154 3619
rect -200 3547 -194 3581
rect -160 3547 -154 3581
rect -200 3509 -154 3547
rect -200 3475 -194 3509
rect -160 3475 -154 3509
rect -200 3437 -154 3475
rect -200 3403 -194 3437
rect -160 3403 -154 3437
rect -200 3365 -154 3403
rect -200 3331 -194 3365
rect -160 3331 -154 3365
rect -200 3293 -154 3331
rect -200 3259 -194 3293
rect -160 3259 -154 3293
rect -200 3221 -154 3259
rect -200 3187 -194 3221
rect -160 3187 -154 3221
rect -200 3149 -154 3187
rect -200 3115 -194 3149
rect -160 3115 -154 3149
rect -200 3077 -154 3115
rect -200 3043 -194 3077
rect -160 3043 -154 3077
rect -200 3005 -154 3043
rect -200 2971 -194 3005
rect -160 2971 -154 3005
rect -200 2933 -154 2971
rect -200 2899 -194 2933
rect -160 2899 -154 2933
rect -200 2861 -154 2899
rect -200 2827 -194 2861
rect -160 2827 -154 2861
rect -200 2789 -154 2827
rect -200 2755 -194 2789
rect -160 2755 -154 2789
rect -200 2717 -154 2755
rect -200 2683 -194 2717
rect -160 2683 -154 2717
rect -200 2645 -154 2683
rect -200 2611 -194 2645
rect -160 2611 -154 2645
rect -200 2573 -154 2611
rect -200 2539 -194 2573
rect -160 2539 -154 2573
rect -200 2501 -154 2539
rect -200 2467 -194 2501
rect -160 2467 -154 2501
rect -200 2429 -154 2467
rect -200 2395 -194 2429
rect -160 2395 -154 2429
rect -200 2357 -154 2395
rect -200 2323 -194 2357
rect -160 2323 -154 2357
rect -200 2285 -154 2323
rect -200 2251 -194 2285
rect -160 2251 -154 2285
rect -200 2213 -154 2251
rect -200 2179 -194 2213
rect -160 2179 -154 2213
rect -200 2141 -154 2179
rect -200 2107 -194 2141
rect -160 2107 -154 2141
rect -200 2069 -154 2107
rect -200 2035 -194 2069
rect -160 2035 -154 2069
rect -200 1997 -154 2035
rect -200 1963 -194 1997
rect -160 1963 -154 1997
rect -200 1925 -154 1963
rect -200 1891 -194 1925
rect -160 1891 -154 1925
rect -200 1853 -154 1891
rect -200 1819 -194 1853
rect -160 1819 -154 1853
rect -200 1781 -154 1819
rect -200 1747 -194 1781
rect -160 1747 -154 1781
rect -200 1709 -154 1747
rect -200 1675 -194 1709
rect -160 1675 -154 1709
rect -200 1637 -154 1675
rect -200 1603 -194 1637
rect -160 1603 -154 1637
rect -200 1565 -154 1603
rect -200 1531 -194 1565
rect -160 1531 -154 1565
rect -200 1493 -154 1531
rect -200 1459 -194 1493
rect -160 1459 -154 1493
rect -200 1421 -154 1459
rect -200 1387 -194 1421
rect -160 1387 -154 1421
rect -200 1349 -154 1387
rect -200 1315 -194 1349
rect -160 1315 -154 1349
rect -200 1277 -154 1315
rect -200 1243 -194 1277
rect -160 1243 -154 1277
rect -200 1205 -154 1243
rect -200 1171 -194 1205
rect -160 1171 -154 1205
rect -200 1133 -154 1171
rect -200 1099 -194 1133
rect -160 1099 -154 1133
rect -200 1061 -154 1099
rect -200 1027 -194 1061
rect -160 1027 -154 1061
rect -200 989 -154 1027
rect -200 955 -194 989
rect -160 955 -154 989
rect -200 917 -154 955
rect -200 883 -194 917
rect -160 883 -154 917
rect -200 845 -154 883
rect -200 811 -194 845
rect -160 811 -154 845
rect -200 773 -154 811
rect -200 739 -194 773
rect -160 739 -154 773
rect -200 701 -154 739
rect -200 667 -194 701
rect -160 667 -154 701
rect -200 629 -154 667
rect -200 595 -194 629
rect -160 595 -154 629
rect -200 557 -154 595
rect -200 523 -194 557
rect -160 523 -154 557
rect -200 485 -154 523
rect -200 451 -194 485
rect -160 451 -154 485
rect -200 413 -154 451
rect -200 379 -194 413
rect -160 379 -154 413
rect -200 341 -154 379
rect -200 307 -194 341
rect -160 307 -154 341
rect -200 269 -154 307
rect -200 235 -194 269
rect -160 235 -154 269
rect -200 197 -154 235
rect -200 163 -194 197
rect -160 163 -154 197
rect -200 125 -154 163
rect -200 91 -194 125
rect -160 91 -154 125
rect -200 53 -154 91
rect -200 19 -194 53
rect -160 19 -154 53
rect -200 -19 -154 19
rect -200 -53 -194 -19
rect -160 -53 -154 -19
rect -200 -91 -154 -53
rect -200 -125 -194 -91
rect -160 -125 -154 -91
rect -200 -163 -154 -125
rect -200 -197 -194 -163
rect -160 -197 -154 -163
rect -200 -235 -154 -197
rect -200 -269 -194 -235
rect -160 -269 -154 -235
rect -200 -307 -154 -269
rect -200 -341 -194 -307
rect -160 -341 -154 -307
rect -200 -379 -154 -341
rect -200 -413 -194 -379
rect -160 -413 -154 -379
rect -200 -451 -154 -413
rect -200 -485 -194 -451
rect -160 -485 -154 -451
rect -200 -523 -154 -485
rect -200 -557 -194 -523
rect -160 -557 -154 -523
rect -200 -595 -154 -557
rect -200 -629 -194 -595
rect -160 -629 -154 -595
rect -200 -667 -154 -629
rect -200 -701 -194 -667
rect -160 -701 -154 -667
rect -200 -739 -154 -701
rect -200 -773 -194 -739
rect -160 -773 -154 -739
rect -200 -811 -154 -773
rect -200 -845 -194 -811
rect -160 -845 -154 -811
rect -200 -883 -154 -845
rect -200 -917 -194 -883
rect -160 -917 -154 -883
rect -200 -955 -154 -917
rect -200 -989 -194 -955
rect -160 -989 -154 -955
rect -200 -1027 -154 -989
rect -200 -1061 -194 -1027
rect -160 -1061 -154 -1027
rect -200 -1099 -154 -1061
rect -200 -1133 -194 -1099
rect -160 -1133 -154 -1099
rect -200 -1171 -154 -1133
rect -200 -1205 -194 -1171
rect -160 -1205 -154 -1171
rect -200 -1243 -154 -1205
rect -200 -1277 -194 -1243
rect -160 -1277 -154 -1243
rect -200 -1315 -154 -1277
rect -200 -1349 -194 -1315
rect -160 -1349 -154 -1315
rect -200 -1387 -154 -1349
rect -200 -1421 -194 -1387
rect -160 -1421 -154 -1387
rect -200 -1459 -154 -1421
rect -200 -1493 -194 -1459
rect -160 -1493 -154 -1459
rect -200 -1531 -154 -1493
rect -200 -1565 -194 -1531
rect -160 -1565 -154 -1531
rect -200 -1603 -154 -1565
rect -200 -1637 -194 -1603
rect -160 -1637 -154 -1603
rect -200 -1675 -154 -1637
rect -200 -1709 -194 -1675
rect -160 -1709 -154 -1675
rect -200 -1747 -154 -1709
rect -200 -1781 -194 -1747
rect -160 -1781 -154 -1747
rect -200 -1819 -154 -1781
rect -200 -1853 -194 -1819
rect -160 -1853 -154 -1819
rect -200 -1891 -154 -1853
rect -200 -1925 -194 -1891
rect -160 -1925 -154 -1891
rect -200 -1963 -154 -1925
rect -200 -1997 -194 -1963
rect -160 -1997 -154 -1963
rect -200 -2035 -154 -1997
rect -200 -2069 -194 -2035
rect -160 -2069 -154 -2035
rect -200 -2107 -154 -2069
rect -200 -2141 -194 -2107
rect -160 -2141 -154 -2107
rect -200 -2179 -154 -2141
rect -200 -2213 -194 -2179
rect -160 -2213 -154 -2179
rect -200 -2251 -154 -2213
rect -200 -2285 -194 -2251
rect -160 -2285 -154 -2251
rect -200 -2323 -154 -2285
rect -200 -2357 -194 -2323
rect -160 -2357 -154 -2323
rect -200 -2395 -154 -2357
rect -200 -2429 -194 -2395
rect -160 -2429 -154 -2395
rect -200 -2467 -154 -2429
rect -200 -2501 -194 -2467
rect -160 -2501 -154 -2467
rect -200 -2539 -154 -2501
rect -200 -2573 -194 -2539
rect -160 -2573 -154 -2539
rect -200 -2611 -154 -2573
rect -200 -2645 -194 -2611
rect -160 -2645 -154 -2611
rect -200 -2683 -154 -2645
rect -200 -2717 -194 -2683
rect -160 -2717 -154 -2683
rect -200 -2755 -154 -2717
rect -200 -2789 -194 -2755
rect -160 -2789 -154 -2755
rect -200 -2827 -154 -2789
rect -200 -2861 -194 -2827
rect -160 -2861 -154 -2827
rect -200 -2899 -154 -2861
rect -200 -2933 -194 -2899
rect -160 -2933 -154 -2899
rect -200 -2971 -154 -2933
rect -200 -3005 -194 -2971
rect -160 -3005 -154 -2971
rect -200 -3043 -154 -3005
rect -200 -3077 -194 -3043
rect -160 -3077 -154 -3043
rect -200 -3115 -154 -3077
rect -200 -3149 -194 -3115
rect -160 -3149 -154 -3115
rect -200 -3187 -154 -3149
rect -200 -3221 -194 -3187
rect -160 -3221 -154 -3187
rect -200 -3259 -154 -3221
rect -200 -3293 -194 -3259
rect -160 -3293 -154 -3259
rect -200 -3331 -154 -3293
rect -200 -3365 -194 -3331
rect -160 -3365 -154 -3331
rect -200 -3403 -154 -3365
rect -200 -3437 -194 -3403
rect -160 -3437 -154 -3403
rect -200 -3475 -154 -3437
rect -200 -3509 -194 -3475
rect -160 -3509 -154 -3475
rect -200 -3547 -154 -3509
rect -200 -3581 -194 -3547
rect -160 -3581 -154 -3547
rect -200 -3619 -154 -3581
rect -200 -3653 -194 -3619
rect -160 -3653 -154 -3619
rect -200 -3691 -154 -3653
rect -200 -3725 -194 -3691
rect -160 -3725 -154 -3691
rect -200 -3763 -154 -3725
rect -200 -3797 -194 -3763
rect -160 -3797 -154 -3763
rect -200 -3835 -154 -3797
rect -200 -3869 -194 -3835
rect -160 -3869 -154 -3835
rect -200 -3907 -154 -3869
rect -200 -3941 -194 -3907
rect -160 -3941 -154 -3907
rect -200 -3979 -154 -3941
rect -200 -4013 -194 -3979
rect -160 -4013 -154 -3979
rect -200 -4051 -154 -4013
rect -200 -4085 -194 -4051
rect -160 -4085 -154 -4051
rect -200 -4123 -154 -4085
rect -200 -4157 -194 -4123
rect -160 -4157 -154 -4123
rect -200 -4195 -154 -4157
rect -200 -4229 -194 -4195
rect -160 -4229 -154 -4195
rect -200 -4267 -154 -4229
rect -200 -4301 -194 -4267
rect -160 -4301 -154 -4267
rect -200 -4339 -154 -4301
rect -200 -4373 -194 -4339
rect -160 -4373 -154 -4339
rect -200 -4411 -154 -4373
rect -200 -4445 -194 -4411
rect -160 -4445 -154 -4411
rect -200 -4483 -154 -4445
rect -200 -4517 -194 -4483
rect -160 -4517 -154 -4483
rect -200 -4555 -154 -4517
rect -200 -4589 -194 -4555
rect -160 -4589 -154 -4555
rect -200 -4627 -154 -4589
rect -200 -4661 -194 -4627
rect -160 -4661 -154 -4627
rect -200 -4699 -154 -4661
rect -200 -4733 -194 -4699
rect -160 -4733 -154 -4699
rect -200 -4771 -154 -4733
rect -200 -4805 -194 -4771
rect -160 -4805 -154 -4771
rect -200 -4843 -154 -4805
rect -200 -4877 -194 -4843
rect -160 -4877 -154 -4843
rect -200 -4915 -154 -4877
rect -200 -4949 -194 -4915
rect -160 -4949 -154 -4915
rect -200 -4987 -154 -4949
rect -200 -5021 -194 -4987
rect -160 -5021 -154 -4987
rect -200 -5059 -154 -5021
rect -200 -5093 -194 -5059
rect -160 -5093 -154 -5059
rect -200 -5131 -154 -5093
rect -200 -5165 -194 -5131
rect -160 -5165 -154 -5131
rect -200 -5203 -154 -5165
rect -200 -5237 -194 -5203
rect -160 -5237 -154 -5203
rect -200 -5275 -154 -5237
rect -200 -5309 -194 -5275
rect -160 -5309 -154 -5275
rect -200 -5347 -154 -5309
rect -200 -5381 -194 -5347
rect -160 -5381 -154 -5347
rect -200 -5419 -154 -5381
rect -200 -5453 -194 -5419
rect -160 -5453 -154 -5419
rect -200 -5491 -154 -5453
rect -200 -5525 -194 -5491
rect -160 -5525 -154 -5491
rect -200 -5563 -154 -5525
rect -200 -5597 -194 -5563
rect -160 -5597 -154 -5563
rect -200 -5635 -154 -5597
rect -200 -5669 -194 -5635
rect -160 -5669 -154 -5635
rect -200 -5707 -154 -5669
rect -200 -5741 -194 -5707
rect -160 -5741 -154 -5707
rect -200 -5779 -154 -5741
rect -200 -5813 -194 -5779
rect -160 -5813 -154 -5779
rect -200 -5851 -154 -5813
rect -200 -5885 -194 -5851
rect -160 -5885 -154 -5851
rect -200 -5923 -154 -5885
rect -200 -5957 -194 -5923
rect -160 -5957 -154 -5923
rect -200 -5995 -154 -5957
rect -200 -6029 -194 -5995
rect -160 -6029 -154 -5995
rect -200 -6067 -154 -6029
rect -200 -6101 -194 -6067
rect -160 -6101 -154 -6067
rect -200 -6139 -154 -6101
rect -200 -6173 -194 -6139
rect -160 -6173 -154 -6139
rect -200 -6211 -154 -6173
rect -200 -6245 -194 -6211
rect -160 -6245 -154 -6211
rect -200 -6283 -154 -6245
rect -200 -6317 -194 -6283
rect -160 -6317 -154 -6283
rect -200 -6355 -154 -6317
rect -200 -6389 -194 -6355
rect -160 -6389 -154 -6355
rect -200 -6427 -154 -6389
rect -200 -6461 -194 -6427
rect -160 -6461 -154 -6427
rect -200 -6499 -154 -6461
rect -200 -6533 -194 -6499
rect -160 -6533 -154 -6499
rect -200 -6571 -154 -6533
rect -200 -6605 -194 -6571
rect -160 -6605 -154 -6571
rect -200 -6643 -154 -6605
rect -200 -6677 -194 -6643
rect -160 -6677 -154 -6643
rect -200 -6715 -154 -6677
rect -200 -6749 -194 -6715
rect -160 -6749 -154 -6715
rect -200 -6787 -154 -6749
rect -200 -6821 -194 -6787
rect -160 -6821 -154 -6787
rect -200 -6859 -154 -6821
rect -200 -6893 -194 -6859
rect -160 -6893 -154 -6859
rect -200 -6931 -154 -6893
rect -200 -6965 -194 -6931
rect -160 -6965 -154 -6931
rect -200 -7003 -154 -6965
rect -200 -7037 -194 -7003
rect -160 -7037 -154 -7003
rect -200 -7075 -154 -7037
rect -200 -7109 -194 -7075
rect -160 -7109 -154 -7075
rect -200 -7147 -154 -7109
rect -200 -7181 -194 -7147
rect -160 -7181 -154 -7147
rect -200 -7219 -154 -7181
rect -200 -7253 -194 -7219
rect -160 -7253 -154 -7219
rect -200 -7291 -154 -7253
rect -200 -7325 -194 -7291
rect -160 -7325 -154 -7291
rect -200 -7363 -154 -7325
rect -200 -7397 -194 -7363
rect -160 -7397 -154 -7363
rect -200 -7435 -154 -7397
rect -200 -7469 -194 -7435
rect -160 -7469 -154 -7435
rect -200 -7507 -154 -7469
rect -200 -7541 -194 -7507
rect -160 -7541 -154 -7507
rect -200 -7579 -154 -7541
rect -200 -7613 -194 -7579
rect -160 -7613 -154 -7579
rect -200 -7651 -154 -7613
rect -200 -7685 -194 -7651
rect -160 -7685 -154 -7651
rect -200 -7723 -154 -7685
rect -200 -7757 -194 -7723
rect -160 -7757 -154 -7723
rect -200 -7795 -154 -7757
rect -200 -7829 -194 -7795
rect -160 -7829 -154 -7795
rect -200 -7867 -154 -7829
rect -200 -7901 -194 -7867
rect -160 -7901 -154 -7867
rect -200 -7939 -154 -7901
rect -200 -7973 -194 -7939
rect -160 -7973 -154 -7939
rect -200 -8011 -154 -7973
rect -200 -8045 -194 -8011
rect -160 -8045 -154 -8011
rect -200 -8083 -154 -8045
rect -200 -8117 -194 -8083
rect -160 -8117 -154 -8083
rect -200 -8155 -154 -8117
rect -200 -8189 -194 -8155
rect -160 -8189 -154 -8155
rect -200 -8227 -154 -8189
rect -200 -8261 -194 -8227
rect -160 -8261 -154 -8227
rect -200 -8299 -154 -8261
rect -200 -8333 -194 -8299
rect -160 -8333 -154 -8299
rect -200 -8371 -154 -8333
rect -200 -8405 -194 -8371
rect -160 -8405 -154 -8371
rect -200 -8443 -154 -8405
rect -200 -8477 -194 -8443
rect -160 -8477 -154 -8443
rect -200 -8515 -154 -8477
rect -200 -8549 -194 -8515
rect -160 -8549 -154 -8515
rect -200 -8587 -154 -8549
rect -200 -8621 -194 -8587
rect -160 -8621 -154 -8587
rect -200 -8659 -154 -8621
rect -200 -8693 -194 -8659
rect -160 -8693 -154 -8659
rect -200 -8731 -154 -8693
rect -200 -8765 -194 -8731
rect -160 -8765 -154 -8731
rect -200 -8803 -154 -8765
rect -200 -8837 -194 -8803
rect -160 -8837 -154 -8803
rect -200 -8875 -154 -8837
rect -200 -8909 -194 -8875
rect -160 -8909 -154 -8875
rect -200 -8947 -154 -8909
rect -200 -8981 -194 -8947
rect -160 -8981 -154 -8947
rect -200 -9019 -154 -8981
rect -200 -9053 -194 -9019
rect -160 -9053 -154 -9019
rect -200 -9091 -154 -9053
rect -200 -9125 -194 -9091
rect -160 -9125 -154 -9091
rect -200 -9163 -154 -9125
rect -200 -9197 -194 -9163
rect -160 -9197 -154 -9163
rect -200 -9235 -154 -9197
rect -200 -9269 -194 -9235
rect -160 -9269 -154 -9235
rect -200 -9307 -154 -9269
rect -200 -9341 -194 -9307
rect -160 -9341 -154 -9307
rect -200 -9379 -154 -9341
rect -200 -9413 -194 -9379
rect -160 -9413 -154 -9379
rect -200 -9451 -154 -9413
rect -200 -9485 -194 -9451
rect -160 -9485 -154 -9451
rect -200 -9523 -154 -9485
rect -200 -9557 -194 -9523
rect -160 -9557 -154 -9523
rect -200 -9600 -154 -9557
rect -82 9557 -36 9600
rect -82 9523 -76 9557
rect -42 9523 -36 9557
rect -82 9485 -36 9523
rect -82 9451 -76 9485
rect -42 9451 -36 9485
rect -82 9413 -36 9451
rect -82 9379 -76 9413
rect -42 9379 -36 9413
rect -82 9341 -36 9379
rect -82 9307 -76 9341
rect -42 9307 -36 9341
rect -82 9269 -36 9307
rect -82 9235 -76 9269
rect -42 9235 -36 9269
rect -82 9197 -36 9235
rect -82 9163 -76 9197
rect -42 9163 -36 9197
rect -82 9125 -36 9163
rect -82 9091 -76 9125
rect -42 9091 -36 9125
rect -82 9053 -36 9091
rect -82 9019 -76 9053
rect -42 9019 -36 9053
rect -82 8981 -36 9019
rect -82 8947 -76 8981
rect -42 8947 -36 8981
rect -82 8909 -36 8947
rect -82 8875 -76 8909
rect -42 8875 -36 8909
rect -82 8837 -36 8875
rect -82 8803 -76 8837
rect -42 8803 -36 8837
rect -82 8765 -36 8803
rect -82 8731 -76 8765
rect -42 8731 -36 8765
rect -82 8693 -36 8731
rect -82 8659 -76 8693
rect -42 8659 -36 8693
rect -82 8621 -36 8659
rect -82 8587 -76 8621
rect -42 8587 -36 8621
rect -82 8549 -36 8587
rect -82 8515 -76 8549
rect -42 8515 -36 8549
rect -82 8477 -36 8515
rect -82 8443 -76 8477
rect -42 8443 -36 8477
rect -82 8405 -36 8443
rect -82 8371 -76 8405
rect -42 8371 -36 8405
rect -82 8333 -36 8371
rect -82 8299 -76 8333
rect -42 8299 -36 8333
rect -82 8261 -36 8299
rect -82 8227 -76 8261
rect -42 8227 -36 8261
rect -82 8189 -36 8227
rect -82 8155 -76 8189
rect -42 8155 -36 8189
rect -82 8117 -36 8155
rect -82 8083 -76 8117
rect -42 8083 -36 8117
rect -82 8045 -36 8083
rect -82 8011 -76 8045
rect -42 8011 -36 8045
rect -82 7973 -36 8011
rect -82 7939 -76 7973
rect -42 7939 -36 7973
rect -82 7901 -36 7939
rect -82 7867 -76 7901
rect -42 7867 -36 7901
rect -82 7829 -36 7867
rect -82 7795 -76 7829
rect -42 7795 -36 7829
rect -82 7757 -36 7795
rect -82 7723 -76 7757
rect -42 7723 -36 7757
rect -82 7685 -36 7723
rect -82 7651 -76 7685
rect -42 7651 -36 7685
rect -82 7613 -36 7651
rect -82 7579 -76 7613
rect -42 7579 -36 7613
rect -82 7541 -36 7579
rect -82 7507 -76 7541
rect -42 7507 -36 7541
rect -82 7469 -36 7507
rect -82 7435 -76 7469
rect -42 7435 -36 7469
rect -82 7397 -36 7435
rect -82 7363 -76 7397
rect -42 7363 -36 7397
rect -82 7325 -36 7363
rect -82 7291 -76 7325
rect -42 7291 -36 7325
rect -82 7253 -36 7291
rect -82 7219 -76 7253
rect -42 7219 -36 7253
rect -82 7181 -36 7219
rect -82 7147 -76 7181
rect -42 7147 -36 7181
rect -82 7109 -36 7147
rect -82 7075 -76 7109
rect -42 7075 -36 7109
rect -82 7037 -36 7075
rect -82 7003 -76 7037
rect -42 7003 -36 7037
rect -82 6965 -36 7003
rect -82 6931 -76 6965
rect -42 6931 -36 6965
rect -82 6893 -36 6931
rect -82 6859 -76 6893
rect -42 6859 -36 6893
rect -82 6821 -36 6859
rect -82 6787 -76 6821
rect -42 6787 -36 6821
rect -82 6749 -36 6787
rect -82 6715 -76 6749
rect -42 6715 -36 6749
rect -82 6677 -36 6715
rect -82 6643 -76 6677
rect -42 6643 -36 6677
rect -82 6605 -36 6643
rect -82 6571 -76 6605
rect -42 6571 -36 6605
rect -82 6533 -36 6571
rect -82 6499 -76 6533
rect -42 6499 -36 6533
rect -82 6461 -36 6499
rect -82 6427 -76 6461
rect -42 6427 -36 6461
rect -82 6389 -36 6427
rect -82 6355 -76 6389
rect -42 6355 -36 6389
rect -82 6317 -36 6355
rect -82 6283 -76 6317
rect -42 6283 -36 6317
rect -82 6245 -36 6283
rect -82 6211 -76 6245
rect -42 6211 -36 6245
rect -82 6173 -36 6211
rect -82 6139 -76 6173
rect -42 6139 -36 6173
rect -82 6101 -36 6139
rect -82 6067 -76 6101
rect -42 6067 -36 6101
rect -82 6029 -36 6067
rect -82 5995 -76 6029
rect -42 5995 -36 6029
rect -82 5957 -36 5995
rect -82 5923 -76 5957
rect -42 5923 -36 5957
rect -82 5885 -36 5923
rect -82 5851 -76 5885
rect -42 5851 -36 5885
rect -82 5813 -36 5851
rect -82 5779 -76 5813
rect -42 5779 -36 5813
rect -82 5741 -36 5779
rect -82 5707 -76 5741
rect -42 5707 -36 5741
rect -82 5669 -36 5707
rect -82 5635 -76 5669
rect -42 5635 -36 5669
rect -82 5597 -36 5635
rect -82 5563 -76 5597
rect -42 5563 -36 5597
rect -82 5525 -36 5563
rect -82 5491 -76 5525
rect -42 5491 -36 5525
rect -82 5453 -36 5491
rect -82 5419 -76 5453
rect -42 5419 -36 5453
rect -82 5381 -36 5419
rect -82 5347 -76 5381
rect -42 5347 -36 5381
rect -82 5309 -36 5347
rect -82 5275 -76 5309
rect -42 5275 -36 5309
rect -82 5237 -36 5275
rect -82 5203 -76 5237
rect -42 5203 -36 5237
rect -82 5165 -36 5203
rect -82 5131 -76 5165
rect -42 5131 -36 5165
rect -82 5093 -36 5131
rect -82 5059 -76 5093
rect -42 5059 -36 5093
rect -82 5021 -36 5059
rect -82 4987 -76 5021
rect -42 4987 -36 5021
rect -82 4949 -36 4987
rect -82 4915 -76 4949
rect -42 4915 -36 4949
rect -82 4877 -36 4915
rect -82 4843 -76 4877
rect -42 4843 -36 4877
rect -82 4805 -36 4843
rect -82 4771 -76 4805
rect -42 4771 -36 4805
rect -82 4733 -36 4771
rect -82 4699 -76 4733
rect -42 4699 -36 4733
rect -82 4661 -36 4699
rect -82 4627 -76 4661
rect -42 4627 -36 4661
rect -82 4589 -36 4627
rect -82 4555 -76 4589
rect -42 4555 -36 4589
rect -82 4517 -36 4555
rect -82 4483 -76 4517
rect -42 4483 -36 4517
rect -82 4445 -36 4483
rect -82 4411 -76 4445
rect -42 4411 -36 4445
rect -82 4373 -36 4411
rect -82 4339 -76 4373
rect -42 4339 -36 4373
rect -82 4301 -36 4339
rect -82 4267 -76 4301
rect -42 4267 -36 4301
rect -82 4229 -36 4267
rect -82 4195 -76 4229
rect -42 4195 -36 4229
rect -82 4157 -36 4195
rect -82 4123 -76 4157
rect -42 4123 -36 4157
rect -82 4085 -36 4123
rect -82 4051 -76 4085
rect -42 4051 -36 4085
rect -82 4013 -36 4051
rect -82 3979 -76 4013
rect -42 3979 -36 4013
rect -82 3941 -36 3979
rect -82 3907 -76 3941
rect -42 3907 -36 3941
rect -82 3869 -36 3907
rect -82 3835 -76 3869
rect -42 3835 -36 3869
rect -82 3797 -36 3835
rect -82 3763 -76 3797
rect -42 3763 -36 3797
rect -82 3725 -36 3763
rect -82 3691 -76 3725
rect -42 3691 -36 3725
rect -82 3653 -36 3691
rect -82 3619 -76 3653
rect -42 3619 -36 3653
rect -82 3581 -36 3619
rect -82 3547 -76 3581
rect -42 3547 -36 3581
rect -82 3509 -36 3547
rect -82 3475 -76 3509
rect -42 3475 -36 3509
rect -82 3437 -36 3475
rect -82 3403 -76 3437
rect -42 3403 -36 3437
rect -82 3365 -36 3403
rect -82 3331 -76 3365
rect -42 3331 -36 3365
rect -82 3293 -36 3331
rect -82 3259 -76 3293
rect -42 3259 -36 3293
rect -82 3221 -36 3259
rect -82 3187 -76 3221
rect -42 3187 -36 3221
rect -82 3149 -36 3187
rect -82 3115 -76 3149
rect -42 3115 -36 3149
rect -82 3077 -36 3115
rect -82 3043 -76 3077
rect -42 3043 -36 3077
rect -82 3005 -36 3043
rect -82 2971 -76 3005
rect -42 2971 -36 3005
rect -82 2933 -36 2971
rect -82 2899 -76 2933
rect -42 2899 -36 2933
rect -82 2861 -36 2899
rect -82 2827 -76 2861
rect -42 2827 -36 2861
rect -82 2789 -36 2827
rect -82 2755 -76 2789
rect -42 2755 -36 2789
rect -82 2717 -36 2755
rect -82 2683 -76 2717
rect -42 2683 -36 2717
rect -82 2645 -36 2683
rect -82 2611 -76 2645
rect -42 2611 -36 2645
rect -82 2573 -36 2611
rect -82 2539 -76 2573
rect -42 2539 -36 2573
rect -82 2501 -36 2539
rect -82 2467 -76 2501
rect -42 2467 -36 2501
rect -82 2429 -36 2467
rect -82 2395 -76 2429
rect -42 2395 -36 2429
rect -82 2357 -36 2395
rect -82 2323 -76 2357
rect -42 2323 -36 2357
rect -82 2285 -36 2323
rect -82 2251 -76 2285
rect -42 2251 -36 2285
rect -82 2213 -36 2251
rect -82 2179 -76 2213
rect -42 2179 -36 2213
rect -82 2141 -36 2179
rect -82 2107 -76 2141
rect -42 2107 -36 2141
rect -82 2069 -36 2107
rect -82 2035 -76 2069
rect -42 2035 -36 2069
rect -82 1997 -36 2035
rect -82 1963 -76 1997
rect -42 1963 -36 1997
rect -82 1925 -36 1963
rect -82 1891 -76 1925
rect -42 1891 -36 1925
rect -82 1853 -36 1891
rect -82 1819 -76 1853
rect -42 1819 -36 1853
rect -82 1781 -36 1819
rect -82 1747 -76 1781
rect -42 1747 -36 1781
rect -82 1709 -36 1747
rect -82 1675 -76 1709
rect -42 1675 -36 1709
rect -82 1637 -36 1675
rect -82 1603 -76 1637
rect -42 1603 -36 1637
rect -82 1565 -36 1603
rect -82 1531 -76 1565
rect -42 1531 -36 1565
rect -82 1493 -36 1531
rect -82 1459 -76 1493
rect -42 1459 -36 1493
rect -82 1421 -36 1459
rect -82 1387 -76 1421
rect -42 1387 -36 1421
rect -82 1349 -36 1387
rect -82 1315 -76 1349
rect -42 1315 -36 1349
rect -82 1277 -36 1315
rect -82 1243 -76 1277
rect -42 1243 -36 1277
rect -82 1205 -36 1243
rect -82 1171 -76 1205
rect -42 1171 -36 1205
rect -82 1133 -36 1171
rect -82 1099 -76 1133
rect -42 1099 -36 1133
rect -82 1061 -36 1099
rect -82 1027 -76 1061
rect -42 1027 -36 1061
rect -82 989 -36 1027
rect -82 955 -76 989
rect -42 955 -36 989
rect -82 917 -36 955
rect -82 883 -76 917
rect -42 883 -36 917
rect -82 845 -36 883
rect -82 811 -76 845
rect -42 811 -36 845
rect -82 773 -36 811
rect -82 739 -76 773
rect -42 739 -36 773
rect -82 701 -36 739
rect -82 667 -76 701
rect -42 667 -36 701
rect -82 629 -36 667
rect -82 595 -76 629
rect -42 595 -36 629
rect -82 557 -36 595
rect -82 523 -76 557
rect -42 523 -36 557
rect -82 485 -36 523
rect -82 451 -76 485
rect -42 451 -36 485
rect -82 413 -36 451
rect -82 379 -76 413
rect -42 379 -36 413
rect -82 341 -36 379
rect -82 307 -76 341
rect -42 307 -36 341
rect -82 269 -36 307
rect -82 235 -76 269
rect -42 235 -36 269
rect -82 197 -36 235
rect -82 163 -76 197
rect -42 163 -36 197
rect -82 125 -36 163
rect -82 91 -76 125
rect -42 91 -36 125
rect -82 53 -36 91
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -91 -36 -53
rect -82 -125 -76 -91
rect -42 -125 -36 -91
rect -82 -163 -36 -125
rect -82 -197 -76 -163
rect -42 -197 -36 -163
rect -82 -235 -36 -197
rect -82 -269 -76 -235
rect -42 -269 -36 -235
rect -82 -307 -36 -269
rect -82 -341 -76 -307
rect -42 -341 -36 -307
rect -82 -379 -36 -341
rect -82 -413 -76 -379
rect -42 -413 -36 -379
rect -82 -451 -36 -413
rect -82 -485 -76 -451
rect -42 -485 -36 -451
rect -82 -523 -36 -485
rect -82 -557 -76 -523
rect -42 -557 -36 -523
rect -82 -595 -36 -557
rect -82 -629 -76 -595
rect -42 -629 -36 -595
rect -82 -667 -36 -629
rect -82 -701 -76 -667
rect -42 -701 -36 -667
rect -82 -739 -36 -701
rect -82 -773 -76 -739
rect -42 -773 -36 -739
rect -82 -811 -36 -773
rect -82 -845 -76 -811
rect -42 -845 -36 -811
rect -82 -883 -36 -845
rect -82 -917 -76 -883
rect -42 -917 -36 -883
rect -82 -955 -36 -917
rect -82 -989 -76 -955
rect -42 -989 -36 -955
rect -82 -1027 -36 -989
rect -82 -1061 -76 -1027
rect -42 -1061 -36 -1027
rect -82 -1099 -36 -1061
rect -82 -1133 -76 -1099
rect -42 -1133 -36 -1099
rect -82 -1171 -36 -1133
rect -82 -1205 -76 -1171
rect -42 -1205 -36 -1171
rect -82 -1243 -36 -1205
rect -82 -1277 -76 -1243
rect -42 -1277 -36 -1243
rect -82 -1315 -36 -1277
rect -82 -1349 -76 -1315
rect -42 -1349 -36 -1315
rect -82 -1387 -36 -1349
rect -82 -1421 -76 -1387
rect -42 -1421 -36 -1387
rect -82 -1459 -36 -1421
rect -82 -1493 -76 -1459
rect -42 -1493 -36 -1459
rect -82 -1531 -36 -1493
rect -82 -1565 -76 -1531
rect -42 -1565 -36 -1531
rect -82 -1603 -36 -1565
rect -82 -1637 -76 -1603
rect -42 -1637 -36 -1603
rect -82 -1675 -36 -1637
rect -82 -1709 -76 -1675
rect -42 -1709 -36 -1675
rect -82 -1747 -36 -1709
rect -82 -1781 -76 -1747
rect -42 -1781 -36 -1747
rect -82 -1819 -36 -1781
rect -82 -1853 -76 -1819
rect -42 -1853 -36 -1819
rect -82 -1891 -36 -1853
rect -82 -1925 -76 -1891
rect -42 -1925 -36 -1891
rect -82 -1963 -36 -1925
rect -82 -1997 -76 -1963
rect -42 -1997 -36 -1963
rect -82 -2035 -36 -1997
rect -82 -2069 -76 -2035
rect -42 -2069 -36 -2035
rect -82 -2107 -36 -2069
rect -82 -2141 -76 -2107
rect -42 -2141 -36 -2107
rect -82 -2179 -36 -2141
rect -82 -2213 -76 -2179
rect -42 -2213 -36 -2179
rect -82 -2251 -36 -2213
rect -82 -2285 -76 -2251
rect -42 -2285 -36 -2251
rect -82 -2323 -36 -2285
rect -82 -2357 -76 -2323
rect -42 -2357 -36 -2323
rect -82 -2395 -36 -2357
rect -82 -2429 -76 -2395
rect -42 -2429 -36 -2395
rect -82 -2467 -36 -2429
rect -82 -2501 -76 -2467
rect -42 -2501 -36 -2467
rect -82 -2539 -36 -2501
rect -82 -2573 -76 -2539
rect -42 -2573 -36 -2539
rect -82 -2611 -36 -2573
rect -82 -2645 -76 -2611
rect -42 -2645 -36 -2611
rect -82 -2683 -36 -2645
rect -82 -2717 -76 -2683
rect -42 -2717 -36 -2683
rect -82 -2755 -36 -2717
rect -82 -2789 -76 -2755
rect -42 -2789 -36 -2755
rect -82 -2827 -36 -2789
rect -82 -2861 -76 -2827
rect -42 -2861 -36 -2827
rect -82 -2899 -36 -2861
rect -82 -2933 -76 -2899
rect -42 -2933 -36 -2899
rect -82 -2971 -36 -2933
rect -82 -3005 -76 -2971
rect -42 -3005 -36 -2971
rect -82 -3043 -36 -3005
rect -82 -3077 -76 -3043
rect -42 -3077 -36 -3043
rect -82 -3115 -36 -3077
rect -82 -3149 -76 -3115
rect -42 -3149 -36 -3115
rect -82 -3187 -36 -3149
rect -82 -3221 -76 -3187
rect -42 -3221 -36 -3187
rect -82 -3259 -36 -3221
rect -82 -3293 -76 -3259
rect -42 -3293 -36 -3259
rect -82 -3331 -36 -3293
rect -82 -3365 -76 -3331
rect -42 -3365 -36 -3331
rect -82 -3403 -36 -3365
rect -82 -3437 -76 -3403
rect -42 -3437 -36 -3403
rect -82 -3475 -36 -3437
rect -82 -3509 -76 -3475
rect -42 -3509 -36 -3475
rect -82 -3547 -36 -3509
rect -82 -3581 -76 -3547
rect -42 -3581 -36 -3547
rect -82 -3619 -36 -3581
rect -82 -3653 -76 -3619
rect -42 -3653 -36 -3619
rect -82 -3691 -36 -3653
rect -82 -3725 -76 -3691
rect -42 -3725 -36 -3691
rect -82 -3763 -36 -3725
rect -82 -3797 -76 -3763
rect -42 -3797 -36 -3763
rect -82 -3835 -36 -3797
rect -82 -3869 -76 -3835
rect -42 -3869 -36 -3835
rect -82 -3907 -36 -3869
rect -82 -3941 -76 -3907
rect -42 -3941 -36 -3907
rect -82 -3979 -36 -3941
rect -82 -4013 -76 -3979
rect -42 -4013 -36 -3979
rect -82 -4051 -36 -4013
rect -82 -4085 -76 -4051
rect -42 -4085 -36 -4051
rect -82 -4123 -36 -4085
rect -82 -4157 -76 -4123
rect -42 -4157 -36 -4123
rect -82 -4195 -36 -4157
rect -82 -4229 -76 -4195
rect -42 -4229 -36 -4195
rect -82 -4267 -36 -4229
rect -82 -4301 -76 -4267
rect -42 -4301 -36 -4267
rect -82 -4339 -36 -4301
rect -82 -4373 -76 -4339
rect -42 -4373 -36 -4339
rect -82 -4411 -36 -4373
rect -82 -4445 -76 -4411
rect -42 -4445 -36 -4411
rect -82 -4483 -36 -4445
rect -82 -4517 -76 -4483
rect -42 -4517 -36 -4483
rect -82 -4555 -36 -4517
rect -82 -4589 -76 -4555
rect -42 -4589 -36 -4555
rect -82 -4627 -36 -4589
rect -82 -4661 -76 -4627
rect -42 -4661 -36 -4627
rect -82 -4699 -36 -4661
rect -82 -4733 -76 -4699
rect -42 -4733 -36 -4699
rect -82 -4771 -36 -4733
rect -82 -4805 -76 -4771
rect -42 -4805 -36 -4771
rect -82 -4843 -36 -4805
rect -82 -4877 -76 -4843
rect -42 -4877 -36 -4843
rect -82 -4915 -36 -4877
rect -82 -4949 -76 -4915
rect -42 -4949 -36 -4915
rect -82 -4987 -36 -4949
rect -82 -5021 -76 -4987
rect -42 -5021 -36 -4987
rect -82 -5059 -36 -5021
rect -82 -5093 -76 -5059
rect -42 -5093 -36 -5059
rect -82 -5131 -36 -5093
rect -82 -5165 -76 -5131
rect -42 -5165 -36 -5131
rect -82 -5203 -36 -5165
rect -82 -5237 -76 -5203
rect -42 -5237 -36 -5203
rect -82 -5275 -36 -5237
rect -82 -5309 -76 -5275
rect -42 -5309 -36 -5275
rect -82 -5347 -36 -5309
rect -82 -5381 -76 -5347
rect -42 -5381 -36 -5347
rect -82 -5419 -36 -5381
rect -82 -5453 -76 -5419
rect -42 -5453 -36 -5419
rect -82 -5491 -36 -5453
rect -82 -5525 -76 -5491
rect -42 -5525 -36 -5491
rect -82 -5563 -36 -5525
rect -82 -5597 -76 -5563
rect -42 -5597 -36 -5563
rect -82 -5635 -36 -5597
rect -82 -5669 -76 -5635
rect -42 -5669 -36 -5635
rect -82 -5707 -36 -5669
rect -82 -5741 -76 -5707
rect -42 -5741 -36 -5707
rect -82 -5779 -36 -5741
rect -82 -5813 -76 -5779
rect -42 -5813 -36 -5779
rect -82 -5851 -36 -5813
rect -82 -5885 -76 -5851
rect -42 -5885 -36 -5851
rect -82 -5923 -36 -5885
rect -82 -5957 -76 -5923
rect -42 -5957 -36 -5923
rect -82 -5995 -36 -5957
rect -82 -6029 -76 -5995
rect -42 -6029 -36 -5995
rect -82 -6067 -36 -6029
rect -82 -6101 -76 -6067
rect -42 -6101 -36 -6067
rect -82 -6139 -36 -6101
rect -82 -6173 -76 -6139
rect -42 -6173 -36 -6139
rect -82 -6211 -36 -6173
rect -82 -6245 -76 -6211
rect -42 -6245 -36 -6211
rect -82 -6283 -36 -6245
rect -82 -6317 -76 -6283
rect -42 -6317 -36 -6283
rect -82 -6355 -36 -6317
rect -82 -6389 -76 -6355
rect -42 -6389 -36 -6355
rect -82 -6427 -36 -6389
rect -82 -6461 -76 -6427
rect -42 -6461 -36 -6427
rect -82 -6499 -36 -6461
rect -82 -6533 -76 -6499
rect -42 -6533 -36 -6499
rect -82 -6571 -36 -6533
rect -82 -6605 -76 -6571
rect -42 -6605 -36 -6571
rect -82 -6643 -36 -6605
rect -82 -6677 -76 -6643
rect -42 -6677 -36 -6643
rect -82 -6715 -36 -6677
rect -82 -6749 -76 -6715
rect -42 -6749 -36 -6715
rect -82 -6787 -36 -6749
rect -82 -6821 -76 -6787
rect -42 -6821 -36 -6787
rect -82 -6859 -36 -6821
rect -82 -6893 -76 -6859
rect -42 -6893 -36 -6859
rect -82 -6931 -36 -6893
rect -82 -6965 -76 -6931
rect -42 -6965 -36 -6931
rect -82 -7003 -36 -6965
rect -82 -7037 -76 -7003
rect -42 -7037 -36 -7003
rect -82 -7075 -36 -7037
rect -82 -7109 -76 -7075
rect -42 -7109 -36 -7075
rect -82 -7147 -36 -7109
rect -82 -7181 -76 -7147
rect -42 -7181 -36 -7147
rect -82 -7219 -36 -7181
rect -82 -7253 -76 -7219
rect -42 -7253 -36 -7219
rect -82 -7291 -36 -7253
rect -82 -7325 -76 -7291
rect -42 -7325 -36 -7291
rect -82 -7363 -36 -7325
rect -82 -7397 -76 -7363
rect -42 -7397 -36 -7363
rect -82 -7435 -36 -7397
rect -82 -7469 -76 -7435
rect -42 -7469 -36 -7435
rect -82 -7507 -36 -7469
rect -82 -7541 -76 -7507
rect -42 -7541 -36 -7507
rect -82 -7579 -36 -7541
rect -82 -7613 -76 -7579
rect -42 -7613 -36 -7579
rect -82 -7651 -36 -7613
rect -82 -7685 -76 -7651
rect -42 -7685 -36 -7651
rect -82 -7723 -36 -7685
rect -82 -7757 -76 -7723
rect -42 -7757 -36 -7723
rect -82 -7795 -36 -7757
rect -82 -7829 -76 -7795
rect -42 -7829 -36 -7795
rect -82 -7867 -36 -7829
rect -82 -7901 -76 -7867
rect -42 -7901 -36 -7867
rect -82 -7939 -36 -7901
rect -82 -7973 -76 -7939
rect -42 -7973 -36 -7939
rect -82 -8011 -36 -7973
rect -82 -8045 -76 -8011
rect -42 -8045 -36 -8011
rect -82 -8083 -36 -8045
rect -82 -8117 -76 -8083
rect -42 -8117 -36 -8083
rect -82 -8155 -36 -8117
rect -82 -8189 -76 -8155
rect -42 -8189 -36 -8155
rect -82 -8227 -36 -8189
rect -82 -8261 -76 -8227
rect -42 -8261 -36 -8227
rect -82 -8299 -36 -8261
rect -82 -8333 -76 -8299
rect -42 -8333 -36 -8299
rect -82 -8371 -36 -8333
rect -82 -8405 -76 -8371
rect -42 -8405 -36 -8371
rect -82 -8443 -36 -8405
rect -82 -8477 -76 -8443
rect -42 -8477 -36 -8443
rect -82 -8515 -36 -8477
rect -82 -8549 -76 -8515
rect -42 -8549 -36 -8515
rect -82 -8587 -36 -8549
rect -82 -8621 -76 -8587
rect -42 -8621 -36 -8587
rect -82 -8659 -36 -8621
rect -82 -8693 -76 -8659
rect -42 -8693 -36 -8659
rect -82 -8731 -36 -8693
rect -82 -8765 -76 -8731
rect -42 -8765 -36 -8731
rect -82 -8803 -36 -8765
rect -82 -8837 -76 -8803
rect -42 -8837 -36 -8803
rect -82 -8875 -36 -8837
rect -82 -8909 -76 -8875
rect -42 -8909 -36 -8875
rect -82 -8947 -36 -8909
rect -82 -8981 -76 -8947
rect -42 -8981 -36 -8947
rect -82 -9019 -36 -8981
rect -82 -9053 -76 -9019
rect -42 -9053 -36 -9019
rect -82 -9091 -36 -9053
rect -82 -9125 -76 -9091
rect -42 -9125 -36 -9091
rect -82 -9163 -36 -9125
rect -82 -9197 -76 -9163
rect -42 -9197 -36 -9163
rect -82 -9235 -36 -9197
rect -82 -9269 -76 -9235
rect -42 -9269 -36 -9235
rect -82 -9307 -36 -9269
rect -82 -9341 -76 -9307
rect -42 -9341 -36 -9307
rect -82 -9379 -36 -9341
rect -82 -9413 -76 -9379
rect -42 -9413 -36 -9379
rect -82 -9451 -36 -9413
rect -82 -9485 -76 -9451
rect -42 -9485 -36 -9451
rect -82 -9523 -36 -9485
rect -82 -9557 -76 -9523
rect -42 -9557 -36 -9523
rect -82 -9600 -36 -9557
rect 36 9557 82 9600
rect 36 9523 42 9557
rect 76 9523 82 9557
rect 36 9485 82 9523
rect 36 9451 42 9485
rect 76 9451 82 9485
rect 36 9413 82 9451
rect 36 9379 42 9413
rect 76 9379 82 9413
rect 36 9341 82 9379
rect 36 9307 42 9341
rect 76 9307 82 9341
rect 36 9269 82 9307
rect 36 9235 42 9269
rect 76 9235 82 9269
rect 36 9197 82 9235
rect 36 9163 42 9197
rect 76 9163 82 9197
rect 36 9125 82 9163
rect 36 9091 42 9125
rect 76 9091 82 9125
rect 36 9053 82 9091
rect 36 9019 42 9053
rect 76 9019 82 9053
rect 36 8981 82 9019
rect 36 8947 42 8981
rect 76 8947 82 8981
rect 36 8909 82 8947
rect 36 8875 42 8909
rect 76 8875 82 8909
rect 36 8837 82 8875
rect 36 8803 42 8837
rect 76 8803 82 8837
rect 36 8765 82 8803
rect 36 8731 42 8765
rect 76 8731 82 8765
rect 36 8693 82 8731
rect 36 8659 42 8693
rect 76 8659 82 8693
rect 36 8621 82 8659
rect 36 8587 42 8621
rect 76 8587 82 8621
rect 36 8549 82 8587
rect 36 8515 42 8549
rect 76 8515 82 8549
rect 36 8477 82 8515
rect 36 8443 42 8477
rect 76 8443 82 8477
rect 36 8405 82 8443
rect 36 8371 42 8405
rect 76 8371 82 8405
rect 36 8333 82 8371
rect 36 8299 42 8333
rect 76 8299 82 8333
rect 36 8261 82 8299
rect 36 8227 42 8261
rect 76 8227 82 8261
rect 36 8189 82 8227
rect 36 8155 42 8189
rect 76 8155 82 8189
rect 36 8117 82 8155
rect 36 8083 42 8117
rect 76 8083 82 8117
rect 36 8045 82 8083
rect 36 8011 42 8045
rect 76 8011 82 8045
rect 36 7973 82 8011
rect 36 7939 42 7973
rect 76 7939 82 7973
rect 36 7901 82 7939
rect 36 7867 42 7901
rect 76 7867 82 7901
rect 36 7829 82 7867
rect 36 7795 42 7829
rect 76 7795 82 7829
rect 36 7757 82 7795
rect 36 7723 42 7757
rect 76 7723 82 7757
rect 36 7685 82 7723
rect 36 7651 42 7685
rect 76 7651 82 7685
rect 36 7613 82 7651
rect 36 7579 42 7613
rect 76 7579 82 7613
rect 36 7541 82 7579
rect 36 7507 42 7541
rect 76 7507 82 7541
rect 36 7469 82 7507
rect 36 7435 42 7469
rect 76 7435 82 7469
rect 36 7397 82 7435
rect 36 7363 42 7397
rect 76 7363 82 7397
rect 36 7325 82 7363
rect 36 7291 42 7325
rect 76 7291 82 7325
rect 36 7253 82 7291
rect 36 7219 42 7253
rect 76 7219 82 7253
rect 36 7181 82 7219
rect 36 7147 42 7181
rect 76 7147 82 7181
rect 36 7109 82 7147
rect 36 7075 42 7109
rect 76 7075 82 7109
rect 36 7037 82 7075
rect 36 7003 42 7037
rect 76 7003 82 7037
rect 36 6965 82 7003
rect 36 6931 42 6965
rect 76 6931 82 6965
rect 36 6893 82 6931
rect 36 6859 42 6893
rect 76 6859 82 6893
rect 36 6821 82 6859
rect 36 6787 42 6821
rect 76 6787 82 6821
rect 36 6749 82 6787
rect 36 6715 42 6749
rect 76 6715 82 6749
rect 36 6677 82 6715
rect 36 6643 42 6677
rect 76 6643 82 6677
rect 36 6605 82 6643
rect 36 6571 42 6605
rect 76 6571 82 6605
rect 36 6533 82 6571
rect 36 6499 42 6533
rect 76 6499 82 6533
rect 36 6461 82 6499
rect 36 6427 42 6461
rect 76 6427 82 6461
rect 36 6389 82 6427
rect 36 6355 42 6389
rect 76 6355 82 6389
rect 36 6317 82 6355
rect 36 6283 42 6317
rect 76 6283 82 6317
rect 36 6245 82 6283
rect 36 6211 42 6245
rect 76 6211 82 6245
rect 36 6173 82 6211
rect 36 6139 42 6173
rect 76 6139 82 6173
rect 36 6101 82 6139
rect 36 6067 42 6101
rect 76 6067 82 6101
rect 36 6029 82 6067
rect 36 5995 42 6029
rect 76 5995 82 6029
rect 36 5957 82 5995
rect 36 5923 42 5957
rect 76 5923 82 5957
rect 36 5885 82 5923
rect 36 5851 42 5885
rect 76 5851 82 5885
rect 36 5813 82 5851
rect 36 5779 42 5813
rect 76 5779 82 5813
rect 36 5741 82 5779
rect 36 5707 42 5741
rect 76 5707 82 5741
rect 36 5669 82 5707
rect 36 5635 42 5669
rect 76 5635 82 5669
rect 36 5597 82 5635
rect 36 5563 42 5597
rect 76 5563 82 5597
rect 36 5525 82 5563
rect 36 5491 42 5525
rect 76 5491 82 5525
rect 36 5453 82 5491
rect 36 5419 42 5453
rect 76 5419 82 5453
rect 36 5381 82 5419
rect 36 5347 42 5381
rect 76 5347 82 5381
rect 36 5309 82 5347
rect 36 5275 42 5309
rect 76 5275 82 5309
rect 36 5237 82 5275
rect 36 5203 42 5237
rect 76 5203 82 5237
rect 36 5165 82 5203
rect 36 5131 42 5165
rect 76 5131 82 5165
rect 36 5093 82 5131
rect 36 5059 42 5093
rect 76 5059 82 5093
rect 36 5021 82 5059
rect 36 4987 42 5021
rect 76 4987 82 5021
rect 36 4949 82 4987
rect 36 4915 42 4949
rect 76 4915 82 4949
rect 36 4877 82 4915
rect 36 4843 42 4877
rect 76 4843 82 4877
rect 36 4805 82 4843
rect 36 4771 42 4805
rect 76 4771 82 4805
rect 36 4733 82 4771
rect 36 4699 42 4733
rect 76 4699 82 4733
rect 36 4661 82 4699
rect 36 4627 42 4661
rect 76 4627 82 4661
rect 36 4589 82 4627
rect 36 4555 42 4589
rect 76 4555 82 4589
rect 36 4517 82 4555
rect 36 4483 42 4517
rect 76 4483 82 4517
rect 36 4445 82 4483
rect 36 4411 42 4445
rect 76 4411 82 4445
rect 36 4373 82 4411
rect 36 4339 42 4373
rect 76 4339 82 4373
rect 36 4301 82 4339
rect 36 4267 42 4301
rect 76 4267 82 4301
rect 36 4229 82 4267
rect 36 4195 42 4229
rect 76 4195 82 4229
rect 36 4157 82 4195
rect 36 4123 42 4157
rect 76 4123 82 4157
rect 36 4085 82 4123
rect 36 4051 42 4085
rect 76 4051 82 4085
rect 36 4013 82 4051
rect 36 3979 42 4013
rect 76 3979 82 4013
rect 36 3941 82 3979
rect 36 3907 42 3941
rect 76 3907 82 3941
rect 36 3869 82 3907
rect 36 3835 42 3869
rect 76 3835 82 3869
rect 36 3797 82 3835
rect 36 3763 42 3797
rect 76 3763 82 3797
rect 36 3725 82 3763
rect 36 3691 42 3725
rect 76 3691 82 3725
rect 36 3653 82 3691
rect 36 3619 42 3653
rect 76 3619 82 3653
rect 36 3581 82 3619
rect 36 3547 42 3581
rect 76 3547 82 3581
rect 36 3509 82 3547
rect 36 3475 42 3509
rect 76 3475 82 3509
rect 36 3437 82 3475
rect 36 3403 42 3437
rect 76 3403 82 3437
rect 36 3365 82 3403
rect 36 3331 42 3365
rect 76 3331 82 3365
rect 36 3293 82 3331
rect 36 3259 42 3293
rect 76 3259 82 3293
rect 36 3221 82 3259
rect 36 3187 42 3221
rect 76 3187 82 3221
rect 36 3149 82 3187
rect 36 3115 42 3149
rect 76 3115 82 3149
rect 36 3077 82 3115
rect 36 3043 42 3077
rect 76 3043 82 3077
rect 36 3005 82 3043
rect 36 2971 42 3005
rect 76 2971 82 3005
rect 36 2933 82 2971
rect 36 2899 42 2933
rect 76 2899 82 2933
rect 36 2861 82 2899
rect 36 2827 42 2861
rect 76 2827 82 2861
rect 36 2789 82 2827
rect 36 2755 42 2789
rect 76 2755 82 2789
rect 36 2717 82 2755
rect 36 2683 42 2717
rect 76 2683 82 2717
rect 36 2645 82 2683
rect 36 2611 42 2645
rect 76 2611 82 2645
rect 36 2573 82 2611
rect 36 2539 42 2573
rect 76 2539 82 2573
rect 36 2501 82 2539
rect 36 2467 42 2501
rect 76 2467 82 2501
rect 36 2429 82 2467
rect 36 2395 42 2429
rect 76 2395 82 2429
rect 36 2357 82 2395
rect 36 2323 42 2357
rect 76 2323 82 2357
rect 36 2285 82 2323
rect 36 2251 42 2285
rect 76 2251 82 2285
rect 36 2213 82 2251
rect 36 2179 42 2213
rect 76 2179 82 2213
rect 36 2141 82 2179
rect 36 2107 42 2141
rect 76 2107 82 2141
rect 36 2069 82 2107
rect 36 2035 42 2069
rect 76 2035 82 2069
rect 36 1997 82 2035
rect 36 1963 42 1997
rect 76 1963 82 1997
rect 36 1925 82 1963
rect 36 1891 42 1925
rect 76 1891 82 1925
rect 36 1853 82 1891
rect 36 1819 42 1853
rect 76 1819 82 1853
rect 36 1781 82 1819
rect 36 1747 42 1781
rect 76 1747 82 1781
rect 36 1709 82 1747
rect 36 1675 42 1709
rect 76 1675 82 1709
rect 36 1637 82 1675
rect 36 1603 42 1637
rect 76 1603 82 1637
rect 36 1565 82 1603
rect 36 1531 42 1565
rect 76 1531 82 1565
rect 36 1493 82 1531
rect 36 1459 42 1493
rect 76 1459 82 1493
rect 36 1421 82 1459
rect 36 1387 42 1421
rect 76 1387 82 1421
rect 36 1349 82 1387
rect 36 1315 42 1349
rect 76 1315 82 1349
rect 36 1277 82 1315
rect 36 1243 42 1277
rect 76 1243 82 1277
rect 36 1205 82 1243
rect 36 1171 42 1205
rect 76 1171 82 1205
rect 36 1133 82 1171
rect 36 1099 42 1133
rect 76 1099 82 1133
rect 36 1061 82 1099
rect 36 1027 42 1061
rect 76 1027 82 1061
rect 36 989 82 1027
rect 36 955 42 989
rect 76 955 82 989
rect 36 917 82 955
rect 36 883 42 917
rect 76 883 82 917
rect 36 845 82 883
rect 36 811 42 845
rect 76 811 82 845
rect 36 773 82 811
rect 36 739 42 773
rect 76 739 82 773
rect 36 701 82 739
rect 36 667 42 701
rect 76 667 82 701
rect 36 629 82 667
rect 36 595 42 629
rect 76 595 82 629
rect 36 557 82 595
rect 36 523 42 557
rect 76 523 82 557
rect 36 485 82 523
rect 36 451 42 485
rect 76 451 82 485
rect 36 413 82 451
rect 36 379 42 413
rect 76 379 82 413
rect 36 341 82 379
rect 36 307 42 341
rect 76 307 82 341
rect 36 269 82 307
rect 36 235 42 269
rect 76 235 82 269
rect 36 197 82 235
rect 36 163 42 197
rect 76 163 82 197
rect 36 125 82 163
rect 36 91 42 125
rect 76 91 82 125
rect 36 53 82 91
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -91 82 -53
rect 36 -125 42 -91
rect 76 -125 82 -91
rect 36 -163 82 -125
rect 36 -197 42 -163
rect 76 -197 82 -163
rect 36 -235 82 -197
rect 36 -269 42 -235
rect 76 -269 82 -235
rect 36 -307 82 -269
rect 36 -341 42 -307
rect 76 -341 82 -307
rect 36 -379 82 -341
rect 36 -413 42 -379
rect 76 -413 82 -379
rect 36 -451 82 -413
rect 36 -485 42 -451
rect 76 -485 82 -451
rect 36 -523 82 -485
rect 36 -557 42 -523
rect 76 -557 82 -523
rect 36 -595 82 -557
rect 36 -629 42 -595
rect 76 -629 82 -595
rect 36 -667 82 -629
rect 36 -701 42 -667
rect 76 -701 82 -667
rect 36 -739 82 -701
rect 36 -773 42 -739
rect 76 -773 82 -739
rect 36 -811 82 -773
rect 36 -845 42 -811
rect 76 -845 82 -811
rect 36 -883 82 -845
rect 36 -917 42 -883
rect 76 -917 82 -883
rect 36 -955 82 -917
rect 36 -989 42 -955
rect 76 -989 82 -955
rect 36 -1027 82 -989
rect 36 -1061 42 -1027
rect 76 -1061 82 -1027
rect 36 -1099 82 -1061
rect 36 -1133 42 -1099
rect 76 -1133 82 -1099
rect 36 -1171 82 -1133
rect 36 -1205 42 -1171
rect 76 -1205 82 -1171
rect 36 -1243 82 -1205
rect 36 -1277 42 -1243
rect 76 -1277 82 -1243
rect 36 -1315 82 -1277
rect 36 -1349 42 -1315
rect 76 -1349 82 -1315
rect 36 -1387 82 -1349
rect 36 -1421 42 -1387
rect 76 -1421 82 -1387
rect 36 -1459 82 -1421
rect 36 -1493 42 -1459
rect 76 -1493 82 -1459
rect 36 -1531 82 -1493
rect 36 -1565 42 -1531
rect 76 -1565 82 -1531
rect 36 -1603 82 -1565
rect 36 -1637 42 -1603
rect 76 -1637 82 -1603
rect 36 -1675 82 -1637
rect 36 -1709 42 -1675
rect 76 -1709 82 -1675
rect 36 -1747 82 -1709
rect 36 -1781 42 -1747
rect 76 -1781 82 -1747
rect 36 -1819 82 -1781
rect 36 -1853 42 -1819
rect 76 -1853 82 -1819
rect 36 -1891 82 -1853
rect 36 -1925 42 -1891
rect 76 -1925 82 -1891
rect 36 -1963 82 -1925
rect 36 -1997 42 -1963
rect 76 -1997 82 -1963
rect 36 -2035 82 -1997
rect 36 -2069 42 -2035
rect 76 -2069 82 -2035
rect 36 -2107 82 -2069
rect 36 -2141 42 -2107
rect 76 -2141 82 -2107
rect 36 -2179 82 -2141
rect 36 -2213 42 -2179
rect 76 -2213 82 -2179
rect 36 -2251 82 -2213
rect 36 -2285 42 -2251
rect 76 -2285 82 -2251
rect 36 -2323 82 -2285
rect 36 -2357 42 -2323
rect 76 -2357 82 -2323
rect 36 -2395 82 -2357
rect 36 -2429 42 -2395
rect 76 -2429 82 -2395
rect 36 -2467 82 -2429
rect 36 -2501 42 -2467
rect 76 -2501 82 -2467
rect 36 -2539 82 -2501
rect 36 -2573 42 -2539
rect 76 -2573 82 -2539
rect 36 -2611 82 -2573
rect 36 -2645 42 -2611
rect 76 -2645 82 -2611
rect 36 -2683 82 -2645
rect 36 -2717 42 -2683
rect 76 -2717 82 -2683
rect 36 -2755 82 -2717
rect 36 -2789 42 -2755
rect 76 -2789 82 -2755
rect 36 -2827 82 -2789
rect 36 -2861 42 -2827
rect 76 -2861 82 -2827
rect 36 -2899 82 -2861
rect 36 -2933 42 -2899
rect 76 -2933 82 -2899
rect 36 -2971 82 -2933
rect 36 -3005 42 -2971
rect 76 -3005 82 -2971
rect 36 -3043 82 -3005
rect 36 -3077 42 -3043
rect 76 -3077 82 -3043
rect 36 -3115 82 -3077
rect 36 -3149 42 -3115
rect 76 -3149 82 -3115
rect 36 -3187 82 -3149
rect 36 -3221 42 -3187
rect 76 -3221 82 -3187
rect 36 -3259 82 -3221
rect 36 -3293 42 -3259
rect 76 -3293 82 -3259
rect 36 -3331 82 -3293
rect 36 -3365 42 -3331
rect 76 -3365 82 -3331
rect 36 -3403 82 -3365
rect 36 -3437 42 -3403
rect 76 -3437 82 -3403
rect 36 -3475 82 -3437
rect 36 -3509 42 -3475
rect 76 -3509 82 -3475
rect 36 -3547 82 -3509
rect 36 -3581 42 -3547
rect 76 -3581 82 -3547
rect 36 -3619 82 -3581
rect 36 -3653 42 -3619
rect 76 -3653 82 -3619
rect 36 -3691 82 -3653
rect 36 -3725 42 -3691
rect 76 -3725 82 -3691
rect 36 -3763 82 -3725
rect 36 -3797 42 -3763
rect 76 -3797 82 -3763
rect 36 -3835 82 -3797
rect 36 -3869 42 -3835
rect 76 -3869 82 -3835
rect 36 -3907 82 -3869
rect 36 -3941 42 -3907
rect 76 -3941 82 -3907
rect 36 -3979 82 -3941
rect 36 -4013 42 -3979
rect 76 -4013 82 -3979
rect 36 -4051 82 -4013
rect 36 -4085 42 -4051
rect 76 -4085 82 -4051
rect 36 -4123 82 -4085
rect 36 -4157 42 -4123
rect 76 -4157 82 -4123
rect 36 -4195 82 -4157
rect 36 -4229 42 -4195
rect 76 -4229 82 -4195
rect 36 -4267 82 -4229
rect 36 -4301 42 -4267
rect 76 -4301 82 -4267
rect 36 -4339 82 -4301
rect 36 -4373 42 -4339
rect 76 -4373 82 -4339
rect 36 -4411 82 -4373
rect 36 -4445 42 -4411
rect 76 -4445 82 -4411
rect 36 -4483 82 -4445
rect 36 -4517 42 -4483
rect 76 -4517 82 -4483
rect 36 -4555 82 -4517
rect 36 -4589 42 -4555
rect 76 -4589 82 -4555
rect 36 -4627 82 -4589
rect 36 -4661 42 -4627
rect 76 -4661 82 -4627
rect 36 -4699 82 -4661
rect 36 -4733 42 -4699
rect 76 -4733 82 -4699
rect 36 -4771 82 -4733
rect 36 -4805 42 -4771
rect 76 -4805 82 -4771
rect 36 -4843 82 -4805
rect 36 -4877 42 -4843
rect 76 -4877 82 -4843
rect 36 -4915 82 -4877
rect 36 -4949 42 -4915
rect 76 -4949 82 -4915
rect 36 -4987 82 -4949
rect 36 -5021 42 -4987
rect 76 -5021 82 -4987
rect 36 -5059 82 -5021
rect 36 -5093 42 -5059
rect 76 -5093 82 -5059
rect 36 -5131 82 -5093
rect 36 -5165 42 -5131
rect 76 -5165 82 -5131
rect 36 -5203 82 -5165
rect 36 -5237 42 -5203
rect 76 -5237 82 -5203
rect 36 -5275 82 -5237
rect 36 -5309 42 -5275
rect 76 -5309 82 -5275
rect 36 -5347 82 -5309
rect 36 -5381 42 -5347
rect 76 -5381 82 -5347
rect 36 -5419 82 -5381
rect 36 -5453 42 -5419
rect 76 -5453 82 -5419
rect 36 -5491 82 -5453
rect 36 -5525 42 -5491
rect 76 -5525 82 -5491
rect 36 -5563 82 -5525
rect 36 -5597 42 -5563
rect 76 -5597 82 -5563
rect 36 -5635 82 -5597
rect 36 -5669 42 -5635
rect 76 -5669 82 -5635
rect 36 -5707 82 -5669
rect 36 -5741 42 -5707
rect 76 -5741 82 -5707
rect 36 -5779 82 -5741
rect 36 -5813 42 -5779
rect 76 -5813 82 -5779
rect 36 -5851 82 -5813
rect 36 -5885 42 -5851
rect 76 -5885 82 -5851
rect 36 -5923 82 -5885
rect 36 -5957 42 -5923
rect 76 -5957 82 -5923
rect 36 -5995 82 -5957
rect 36 -6029 42 -5995
rect 76 -6029 82 -5995
rect 36 -6067 82 -6029
rect 36 -6101 42 -6067
rect 76 -6101 82 -6067
rect 36 -6139 82 -6101
rect 36 -6173 42 -6139
rect 76 -6173 82 -6139
rect 36 -6211 82 -6173
rect 36 -6245 42 -6211
rect 76 -6245 82 -6211
rect 36 -6283 82 -6245
rect 36 -6317 42 -6283
rect 76 -6317 82 -6283
rect 36 -6355 82 -6317
rect 36 -6389 42 -6355
rect 76 -6389 82 -6355
rect 36 -6427 82 -6389
rect 36 -6461 42 -6427
rect 76 -6461 82 -6427
rect 36 -6499 82 -6461
rect 36 -6533 42 -6499
rect 76 -6533 82 -6499
rect 36 -6571 82 -6533
rect 36 -6605 42 -6571
rect 76 -6605 82 -6571
rect 36 -6643 82 -6605
rect 36 -6677 42 -6643
rect 76 -6677 82 -6643
rect 36 -6715 82 -6677
rect 36 -6749 42 -6715
rect 76 -6749 82 -6715
rect 36 -6787 82 -6749
rect 36 -6821 42 -6787
rect 76 -6821 82 -6787
rect 36 -6859 82 -6821
rect 36 -6893 42 -6859
rect 76 -6893 82 -6859
rect 36 -6931 82 -6893
rect 36 -6965 42 -6931
rect 76 -6965 82 -6931
rect 36 -7003 82 -6965
rect 36 -7037 42 -7003
rect 76 -7037 82 -7003
rect 36 -7075 82 -7037
rect 36 -7109 42 -7075
rect 76 -7109 82 -7075
rect 36 -7147 82 -7109
rect 36 -7181 42 -7147
rect 76 -7181 82 -7147
rect 36 -7219 82 -7181
rect 36 -7253 42 -7219
rect 76 -7253 82 -7219
rect 36 -7291 82 -7253
rect 36 -7325 42 -7291
rect 76 -7325 82 -7291
rect 36 -7363 82 -7325
rect 36 -7397 42 -7363
rect 76 -7397 82 -7363
rect 36 -7435 82 -7397
rect 36 -7469 42 -7435
rect 76 -7469 82 -7435
rect 36 -7507 82 -7469
rect 36 -7541 42 -7507
rect 76 -7541 82 -7507
rect 36 -7579 82 -7541
rect 36 -7613 42 -7579
rect 76 -7613 82 -7579
rect 36 -7651 82 -7613
rect 36 -7685 42 -7651
rect 76 -7685 82 -7651
rect 36 -7723 82 -7685
rect 36 -7757 42 -7723
rect 76 -7757 82 -7723
rect 36 -7795 82 -7757
rect 36 -7829 42 -7795
rect 76 -7829 82 -7795
rect 36 -7867 82 -7829
rect 36 -7901 42 -7867
rect 76 -7901 82 -7867
rect 36 -7939 82 -7901
rect 36 -7973 42 -7939
rect 76 -7973 82 -7939
rect 36 -8011 82 -7973
rect 36 -8045 42 -8011
rect 76 -8045 82 -8011
rect 36 -8083 82 -8045
rect 36 -8117 42 -8083
rect 76 -8117 82 -8083
rect 36 -8155 82 -8117
rect 36 -8189 42 -8155
rect 76 -8189 82 -8155
rect 36 -8227 82 -8189
rect 36 -8261 42 -8227
rect 76 -8261 82 -8227
rect 36 -8299 82 -8261
rect 36 -8333 42 -8299
rect 76 -8333 82 -8299
rect 36 -8371 82 -8333
rect 36 -8405 42 -8371
rect 76 -8405 82 -8371
rect 36 -8443 82 -8405
rect 36 -8477 42 -8443
rect 76 -8477 82 -8443
rect 36 -8515 82 -8477
rect 36 -8549 42 -8515
rect 76 -8549 82 -8515
rect 36 -8587 82 -8549
rect 36 -8621 42 -8587
rect 76 -8621 82 -8587
rect 36 -8659 82 -8621
rect 36 -8693 42 -8659
rect 76 -8693 82 -8659
rect 36 -8731 82 -8693
rect 36 -8765 42 -8731
rect 76 -8765 82 -8731
rect 36 -8803 82 -8765
rect 36 -8837 42 -8803
rect 76 -8837 82 -8803
rect 36 -8875 82 -8837
rect 36 -8909 42 -8875
rect 76 -8909 82 -8875
rect 36 -8947 82 -8909
rect 36 -8981 42 -8947
rect 76 -8981 82 -8947
rect 36 -9019 82 -8981
rect 36 -9053 42 -9019
rect 76 -9053 82 -9019
rect 36 -9091 82 -9053
rect 36 -9125 42 -9091
rect 76 -9125 82 -9091
rect 36 -9163 82 -9125
rect 36 -9197 42 -9163
rect 76 -9197 82 -9163
rect 36 -9235 82 -9197
rect 36 -9269 42 -9235
rect 76 -9269 82 -9235
rect 36 -9307 82 -9269
rect 36 -9341 42 -9307
rect 76 -9341 82 -9307
rect 36 -9379 82 -9341
rect 36 -9413 42 -9379
rect 76 -9413 82 -9379
rect 36 -9451 82 -9413
rect 36 -9485 42 -9451
rect 76 -9485 82 -9451
rect 36 -9523 82 -9485
rect 36 -9557 42 -9523
rect 76 -9557 82 -9523
rect 36 -9600 82 -9557
rect 154 9557 200 9600
rect 154 9523 160 9557
rect 194 9523 200 9557
rect 154 9485 200 9523
rect 154 9451 160 9485
rect 194 9451 200 9485
rect 154 9413 200 9451
rect 154 9379 160 9413
rect 194 9379 200 9413
rect 154 9341 200 9379
rect 154 9307 160 9341
rect 194 9307 200 9341
rect 154 9269 200 9307
rect 154 9235 160 9269
rect 194 9235 200 9269
rect 154 9197 200 9235
rect 154 9163 160 9197
rect 194 9163 200 9197
rect 154 9125 200 9163
rect 154 9091 160 9125
rect 194 9091 200 9125
rect 154 9053 200 9091
rect 154 9019 160 9053
rect 194 9019 200 9053
rect 154 8981 200 9019
rect 154 8947 160 8981
rect 194 8947 200 8981
rect 154 8909 200 8947
rect 154 8875 160 8909
rect 194 8875 200 8909
rect 154 8837 200 8875
rect 154 8803 160 8837
rect 194 8803 200 8837
rect 154 8765 200 8803
rect 154 8731 160 8765
rect 194 8731 200 8765
rect 154 8693 200 8731
rect 154 8659 160 8693
rect 194 8659 200 8693
rect 154 8621 200 8659
rect 154 8587 160 8621
rect 194 8587 200 8621
rect 154 8549 200 8587
rect 154 8515 160 8549
rect 194 8515 200 8549
rect 154 8477 200 8515
rect 154 8443 160 8477
rect 194 8443 200 8477
rect 154 8405 200 8443
rect 154 8371 160 8405
rect 194 8371 200 8405
rect 154 8333 200 8371
rect 154 8299 160 8333
rect 194 8299 200 8333
rect 154 8261 200 8299
rect 154 8227 160 8261
rect 194 8227 200 8261
rect 154 8189 200 8227
rect 154 8155 160 8189
rect 194 8155 200 8189
rect 154 8117 200 8155
rect 154 8083 160 8117
rect 194 8083 200 8117
rect 154 8045 200 8083
rect 154 8011 160 8045
rect 194 8011 200 8045
rect 154 7973 200 8011
rect 154 7939 160 7973
rect 194 7939 200 7973
rect 154 7901 200 7939
rect 154 7867 160 7901
rect 194 7867 200 7901
rect 154 7829 200 7867
rect 154 7795 160 7829
rect 194 7795 200 7829
rect 154 7757 200 7795
rect 154 7723 160 7757
rect 194 7723 200 7757
rect 154 7685 200 7723
rect 154 7651 160 7685
rect 194 7651 200 7685
rect 154 7613 200 7651
rect 154 7579 160 7613
rect 194 7579 200 7613
rect 154 7541 200 7579
rect 154 7507 160 7541
rect 194 7507 200 7541
rect 154 7469 200 7507
rect 154 7435 160 7469
rect 194 7435 200 7469
rect 154 7397 200 7435
rect 154 7363 160 7397
rect 194 7363 200 7397
rect 154 7325 200 7363
rect 154 7291 160 7325
rect 194 7291 200 7325
rect 154 7253 200 7291
rect 154 7219 160 7253
rect 194 7219 200 7253
rect 154 7181 200 7219
rect 154 7147 160 7181
rect 194 7147 200 7181
rect 154 7109 200 7147
rect 154 7075 160 7109
rect 194 7075 200 7109
rect 154 7037 200 7075
rect 154 7003 160 7037
rect 194 7003 200 7037
rect 154 6965 200 7003
rect 154 6931 160 6965
rect 194 6931 200 6965
rect 154 6893 200 6931
rect 154 6859 160 6893
rect 194 6859 200 6893
rect 154 6821 200 6859
rect 154 6787 160 6821
rect 194 6787 200 6821
rect 154 6749 200 6787
rect 154 6715 160 6749
rect 194 6715 200 6749
rect 154 6677 200 6715
rect 154 6643 160 6677
rect 194 6643 200 6677
rect 154 6605 200 6643
rect 154 6571 160 6605
rect 194 6571 200 6605
rect 154 6533 200 6571
rect 154 6499 160 6533
rect 194 6499 200 6533
rect 154 6461 200 6499
rect 154 6427 160 6461
rect 194 6427 200 6461
rect 154 6389 200 6427
rect 154 6355 160 6389
rect 194 6355 200 6389
rect 154 6317 200 6355
rect 154 6283 160 6317
rect 194 6283 200 6317
rect 154 6245 200 6283
rect 154 6211 160 6245
rect 194 6211 200 6245
rect 154 6173 200 6211
rect 154 6139 160 6173
rect 194 6139 200 6173
rect 154 6101 200 6139
rect 154 6067 160 6101
rect 194 6067 200 6101
rect 154 6029 200 6067
rect 154 5995 160 6029
rect 194 5995 200 6029
rect 154 5957 200 5995
rect 154 5923 160 5957
rect 194 5923 200 5957
rect 154 5885 200 5923
rect 154 5851 160 5885
rect 194 5851 200 5885
rect 154 5813 200 5851
rect 154 5779 160 5813
rect 194 5779 200 5813
rect 154 5741 200 5779
rect 154 5707 160 5741
rect 194 5707 200 5741
rect 154 5669 200 5707
rect 154 5635 160 5669
rect 194 5635 200 5669
rect 154 5597 200 5635
rect 154 5563 160 5597
rect 194 5563 200 5597
rect 154 5525 200 5563
rect 154 5491 160 5525
rect 194 5491 200 5525
rect 154 5453 200 5491
rect 154 5419 160 5453
rect 194 5419 200 5453
rect 154 5381 200 5419
rect 154 5347 160 5381
rect 194 5347 200 5381
rect 154 5309 200 5347
rect 154 5275 160 5309
rect 194 5275 200 5309
rect 154 5237 200 5275
rect 154 5203 160 5237
rect 194 5203 200 5237
rect 154 5165 200 5203
rect 154 5131 160 5165
rect 194 5131 200 5165
rect 154 5093 200 5131
rect 154 5059 160 5093
rect 194 5059 200 5093
rect 154 5021 200 5059
rect 154 4987 160 5021
rect 194 4987 200 5021
rect 154 4949 200 4987
rect 154 4915 160 4949
rect 194 4915 200 4949
rect 154 4877 200 4915
rect 154 4843 160 4877
rect 194 4843 200 4877
rect 154 4805 200 4843
rect 154 4771 160 4805
rect 194 4771 200 4805
rect 154 4733 200 4771
rect 154 4699 160 4733
rect 194 4699 200 4733
rect 154 4661 200 4699
rect 154 4627 160 4661
rect 194 4627 200 4661
rect 154 4589 200 4627
rect 154 4555 160 4589
rect 194 4555 200 4589
rect 154 4517 200 4555
rect 154 4483 160 4517
rect 194 4483 200 4517
rect 154 4445 200 4483
rect 154 4411 160 4445
rect 194 4411 200 4445
rect 154 4373 200 4411
rect 154 4339 160 4373
rect 194 4339 200 4373
rect 154 4301 200 4339
rect 154 4267 160 4301
rect 194 4267 200 4301
rect 154 4229 200 4267
rect 154 4195 160 4229
rect 194 4195 200 4229
rect 154 4157 200 4195
rect 154 4123 160 4157
rect 194 4123 200 4157
rect 154 4085 200 4123
rect 154 4051 160 4085
rect 194 4051 200 4085
rect 154 4013 200 4051
rect 154 3979 160 4013
rect 194 3979 200 4013
rect 154 3941 200 3979
rect 154 3907 160 3941
rect 194 3907 200 3941
rect 154 3869 200 3907
rect 154 3835 160 3869
rect 194 3835 200 3869
rect 154 3797 200 3835
rect 154 3763 160 3797
rect 194 3763 200 3797
rect 154 3725 200 3763
rect 154 3691 160 3725
rect 194 3691 200 3725
rect 154 3653 200 3691
rect 154 3619 160 3653
rect 194 3619 200 3653
rect 154 3581 200 3619
rect 154 3547 160 3581
rect 194 3547 200 3581
rect 154 3509 200 3547
rect 154 3475 160 3509
rect 194 3475 200 3509
rect 154 3437 200 3475
rect 154 3403 160 3437
rect 194 3403 200 3437
rect 154 3365 200 3403
rect 154 3331 160 3365
rect 194 3331 200 3365
rect 154 3293 200 3331
rect 154 3259 160 3293
rect 194 3259 200 3293
rect 154 3221 200 3259
rect 154 3187 160 3221
rect 194 3187 200 3221
rect 154 3149 200 3187
rect 154 3115 160 3149
rect 194 3115 200 3149
rect 154 3077 200 3115
rect 154 3043 160 3077
rect 194 3043 200 3077
rect 154 3005 200 3043
rect 154 2971 160 3005
rect 194 2971 200 3005
rect 154 2933 200 2971
rect 154 2899 160 2933
rect 194 2899 200 2933
rect 154 2861 200 2899
rect 154 2827 160 2861
rect 194 2827 200 2861
rect 154 2789 200 2827
rect 154 2755 160 2789
rect 194 2755 200 2789
rect 154 2717 200 2755
rect 154 2683 160 2717
rect 194 2683 200 2717
rect 154 2645 200 2683
rect 154 2611 160 2645
rect 194 2611 200 2645
rect 154 2573 200 2611
rect 154 2539 160 2573
rect 194 2539 200 2573
rect 154 2501 200 2539
rect 154 2467 160 2501
rect 194 2467 200 2501
rect 154 2429 200 2467
rect 154 2395 160 2429
rect 194 2395 200 2429
rect 154 2357 200 2395
rect 154 2323 160 2357
rect 194 2323 200 2357
rect 154 2285 200 2323
rect 154 2251 160 2285
rect 194 2251 200 2285
rect 154 2213 200 2251
rect 154 2179 160 2213
rect 194 2179 200 2213
rect 154 2141 200 2179
rect 154 2107 160 2141
rect 194 2107 200 2141
rect 154 2069 200 2107
rect 154 2035 160 2069
rect 194 2035 200 2069
rect 154 1997 200 2035
rect 154 1963 160 1997
rect 194 1963 200 1997
rect 154 1925 200 1963
rect 154 1891 160 1925
rect 194 1891 200 1925
rect 154 1853 200 1891
rect 154 1819 160 1853
rect 194 1819 200 1853
rect 154 1781 200 1819
rect 154 1747 160 1781
rect 194 1747 200 1781
rect 154 1709 200 1747
rect 154 1675 160 1709
rect 194 1675 200 1709
rect 154 1637 200 1675
rect 154 1603 160 1637
rect 194 1603 200 1637
rect 154 1565 200 1603
rect 154 1531 160 1565
rect 194 1531 200 1565
rect 154 1493 200 1531
rect 154 1459 160 1493
rect 194 1459 200 1493
rect 154 1421 200 1459
rect 154 1387 160 1421
rect 194 1387 200 1421
rect 154 1349 200 1387
rect 154 1315 160 1349
rect 194 1315 200 1349
rect 154 1277 200 1315
rect 154 1243 160 1277
rect 194 1243 200 1277
rect 154 1205 200 1243
rect 154 1171 160 1205
rect 194 1171 200 1205
rect 154 1133 200 1171
rect 154 1099 160 1133
rect 194 1099 200 1133
rect 154 1061 200 1099
rect 154 1027 160 1061
rect 194 1027 200 1061
rect 154 989 200 1027
rect 154 955 160 989
rect 194 955 200 989
rect 154 917 200 955
rect 154 883 160 917
rect 194 883 200 917
rect 154 845 200 883
rect 154 811 160 845
rect 194 811 200 845
rect 154 773 200 811
rect 154 739 160 773
rect 194 739 200 773
rect 154 701 200 739
rect 154 667 160 701
rect 194 667 200 701
rect 154 629 200 667
rect 154 595 160 629
rect 194 595 200 629
rect 154 557 200 595
rect 154 523 160 557
rect 194 523 200 557
rect 154 485 200 523
rect 154 451 160 485
rect 194 451 200 485
rect 154 413 200 451
rect 154 379 160 413
rect 194 379 200 413
rect 154 341 200 379
rect 154 307 160 341
rect 194 307 200 341
rect 154 269 200 307
rect 154 235 160 269
rect 194 235 200 269
rect 154 197 200 235
rect 154 163 160 197
rect 194 163 200 197
rect 154 125 200 163
rect 154 91 160 125
rect 194 91 200 125
rect 154 53 200 91
rect 154 19 160 53
rect 194 19 200 53
rect 154 -19 200 19
rect 154 -53 160 -19
rect 194 -53 200 -19
rect 154 -91 200 -53
rect 154 -125 160 -91
rect 194 -125 200 -91
rect 154 -163 200 -125
rect 154 -197 160 -163
rect 194 -197 200 -163
rect 154 -235 200 -197
rect 154 -269 160 -235
rect 194 -269 200 -235
rect 154 -307 200 -269
rect 154 -341 160 -307
rect 194 -341 200 -307
rect 154 -379 200 -341
rect 154 -413 160 -379
rect 194 -413 200 -379
rect 154 -451 200 -413
rect 154 -485 160 -451
rect 194 -485 200 -451
rect 154 -523 200 -485
rect 154 -557 160 -523
rect 194 -557 200 -523
rect 154 -595 200 -557
rect 154 -629 160 -595
rect 194 -629 200 -595
rect 154 -667 200 -629
rect 154 -701 160 -667
rect 194 -701 200 -667
rect 154 -739 200 -701
rect 154 -773 160 -739
rect 194 -773 200 -739
rect 154 -811 200 -773
rect 154 -845 160 -811
rect 194 -845 200 -811
rect 154 -883 200 -845
rect 154 -917 160 -883
rect 194 -917 200 -883
rect 154 -955 200 -917
rect 154 -989 160 -955
rect 194 -989 200 -955
rect 154 -1027 200 -989
rect 154 -1061 160 -1027
rect 194 -1061 200 -1027
rect 154 -1099 200 -1061
rect 154 -1133 160 -1099
rect 194 -1133 200 -1099
rect 154 -1171 200 -1133
rect 154 -1205 160 -1171
rect 194 -1205 200 -1171
rect 154 -1243 200 -1205
rect 154 -1277 160 -1243
rect 194 -1277 200 -1243
rect 154 -1315 200 -1277
rect 154 -1349 160 -1315
rect 194 -1349 200 -1315
rect 154 -1387 200 -1349
rect 154 -1421 160 -1387
rect 194 -1421 200 -1387
rect 154 -1459 200 -1421
rect 154 -1493 160 -1459
rect 194 -1493 200 -1459
rect 154 -1531 200 -1493
rect 154 -1565 160 -1531
rect 194 -1565 200 -1531
rect 154 -1603 200 -1565
rect 154 -1637 160 -1603
rect 194 -1637 200 -1603
rect 154 -1675 200 -1637
rect 154 -1709 160 -1675
rect 194 -1709 200 -1675
rect 154 -1747 200 -1709
rect 154 -1781 160 -1747
rect 194 -1781 200 -1747
rect 154 -1819 200 -1781
rect 154 -1853 160 -1819
rect 194 -1853 200 -1819
rect 154 -1891 200 -1853
rect 154 -1925 160 -1891
rect 194 -1925 200 -1891
rect 154 -1963 200 -1925
rect 154 -1997 160 -1963
rect 194 -1997 200 -1963
rect 154 -2035 200 -1997
rect 154 -2069 160 -2035
rect 194 -2069 200 -2035
rect 154 -2107 200 -2069
rect 154 -2141 160 -2107
rect 194 -2141 200 -2107
rect 154 -2179 200 -2141
rect 154 -2213 160 -2179
rect 194 -2213 200 -2179
rect 154 -2251 200 -2213
rect 154 -2285 160 -2251
rect 194 -2285 200 -2251
rect 154 -2323 200 -2285
rect 154 -2357 160 -2323
rect 194 -2357 200 -2323
rect 154 -2395 200 -2357
rect 154 -2429 160 -2395
rect 194 -2429 200 -2395
rect 154 -2467 200 -2429
rect 154 -2501 160 -2467
rect 194 -2501 200 -2467
rect 154 -2539 200 -2501
rect 154 -2573 160 -2539
rect 194 -2573 200 -2539
rect 154 -2611 200 -2573
rect 154 -2645 160 -2611
rect 194 -2645 200 -2611
rect 154 -2683 200 -2645
rect 154 -2717 160 -2683
rect 194 -2717 200 -2683
rect 154 -2755 200 -2717
rect 154 -2789 160 -2755
rect 194 -2789 200 -2755
rect 154 -2827 200 -2789
rect 154 -2861 160 -2827
rect 194 -2861 200 -2827
rect 154 -2899 200 -2861
rect 154 -2933 160 -2899
rect 194 -2933 200 -2899
rect 154 -2971 200 -2933
rect 154 -3005 160 -2971
rect 194 -3005 200 -2971
rect 154 -3043 200 -3005
rect 154 -3077 160 -3043
rect 194 -3077 200 -3043
rect 154 -3115 200 -3077
rect 154 -3149 160 -3115
rect 194 -3149 200 -3115
rect 154 -3187 200 -3149
rect 154 -3221 160 -3187
rect 194 -3221 200 -3187
rect 154 -3259 200 -3221
rect 154 -3293 160 -3259
rect 194 -3293 200 -3259
rect 154 -3331 200 -3293
rect 154 -3365 160 -3331
rect 194 -3365 200 -3331
rect 154 -3403 200 -3365
rect 154 -3437 160 -3403
rect 194 -3437 200 -3403
rect 154 -3475 200 -3437
rect 154 -3509 160 -3475
rect 194 -3509 200 -3475
rect 154 -3547 200 -3509
rect 154 -3581 160 -3547
rect 194 -3581 200 -3547
rect 154 -3619 200 -3581
rect 154 -3653 160 -3619
rect 194 -3653 200 -3619
rect 154 -3691 200 -3653
rect 154 -3725 160 -3691
rect 194 -3725 200 -3691
rect 154 -3763 200 -3725
rect 154 -3797 160 -3763
rect 194 -3797 200 -3763
rect 154 -3835 200 -3797
rect 154 -3869 160 -3835
rect 194 -3869 200 -3835
rect 154 -3907 200 -3869
rect 154 -3941 160 -3907
rect 194 -3941 200 -3907
rect 154 -3979 200 -3941
rect 154 -4013 160 -3979
rect 194 -4013 200 -3979
rect 154 -4051 200 -4013
rect 154 -4085 160 -4051
rect 194 -4085 200 -4051
rect 154 -4123 200 -4085
rect 154 -4157 160 -4123
rect 194 -4157 200 -4123
rect 154 -4195 200 -4157
rect 154 -4229 160 -4195
rect 194 -4229 200 -4195
rect 154 -4267 200 -4229
rect 154 -4301 160 -4267
rect 194 -4301 200 -4267
rect 154 -4339 200 -4301
rect 154 -4373 160 -4339
rect 194 -4373 200 -4339
rect 154 -4411 200 -4373
rect 154 -4445 160 -4411
rect 194 -4445 200 -4411
rect 154 -4483 200 -4445
rect 154 -4517 160 -4483
rect 194 -4517 200 -4483
rect 154 -4555 200 -4517
rect 154 -4589 160 -4555
rect 194 -4589 200 -4555
rect 154 -4627 200 -4589
rect 154 -4661 160 -4627
rect 194 -4661 200 -4627
rect 154 -4699 200 -4661
rect 154 -4733 160 -4699
rect 194 -4733 200 -4699
rect 154 -4771 200 -4733
rect 154 -4805 160 -4771
rect 194 -4805 200 -4771
rect 154 -4843 200 -4805
rect 154 -4877 160 -4843
rect 194 -4877 200 -4843
rect 154 -4915 200 -4877
rect 154 -4949 160 -4915
rect 194 -4949 200 -4915
rect 154 -4987 200 -4949
rect 154 -5021 160 -4987
rect 194 -5021 200 -4987
rect 154 -5059 200 -5021
rect 154 -5093 160 -5059
rect 194 -5093 200 -5059
rect 154 -5131 200 -5093
rect 154 -5165 160 -5131
rect 194 -5165 200 -5131
rect 154 -5203 200 -5165
rect 154 -5237 160 -5203
rect 194 -5237 200 -5203
rect 154 -5275 200 -5237
rect 154 -5309 160 -5275
rect 194 -5309 200 -5275
rect 154 -5347 200 -5309
rect 154 -5381 160 -5347
rect 194 -5381 200 -5347
rect 154 -5419 200 -5381
rect 154 -5453 160 -5419
rect 194 -5453 200 -5419
rect 154 -5491 200 -5453
rect 154 -5525 160 -5491
rect 194 -5525 200 -5491
rect 154 -5563 200 -5525
rect 154 -5597 160 -5563
rect 194 -5597 200 -5563
rect 154 -5635 200 -5597
rect 154 -5669 160 -5635
rect 194 -5669 200 -5635
rect 154 -5707 200 -5669
rect 154 -5741 160 -5707
rect 194 -5741 200 -5707
rect 154 -5779 200 -5741
rect 154 -5813 160 -5779
rect 194 -5813 200 -5779
rect 154 -5851 200 -5813
rect 154 -5885 160 -5851
rect 194 -5885 200 -5851
rect 154 -5923 200 -5885
rect 154 -5957 160 -5923
rect 194 -5957 200 -5923
rect 154 -5995 200 -5957
rect 154 -6029 160 -5995
rect 194 -6029 200 -5995
rect 154 -6067 200 -6029
rect 154 -6101 160 -6067
rect 194 -6101 200 -6067
rect 154 -6139 200 -6101
rect 154 -6173 160 -6139
rect 194 -6173 200 -6139
rect 154 -6211 200 -6173
rect 154 -6245 160 -6211
rect 194 -6245 200 -6211
rect 154 -6283 200 -6245
rect 154 -6317 160 -6283
rect 194 -6317 200 -6283
rect 154 -6355 200 -6317
rect 154 -6389 160 -6355
rect 194 -6389 200 -6355
rect 154 -6427 200 -6389
rect 154 -6461 160 -6427
rect 194 -6461 200 -6427
rect 154 -6499 200 -6461
rect 154 -6533 160 -6499
rect 194 -6533 200 -6499
rect 154 -6571 200 -6533
rect 154 -6605 160 -6571
rect 194 -6605 200 -6571
rect 154 -6643 200 -6605
rect 154 -6677 160 -6643
rect 194 -6677 200 -6643
rect 154 -6715 200 -6677
rect 154 -6749 160 -6715
rect 194 -6749 200 -6715
rect 154 -6787 200 -6749
rect 154 -6821 160 -6787
rect 194 -6821 200 -6787
rect 154 -6859 200 -6821
rect 154 -6893 160 -6859
rect 194 -6893 200 -6859
rect 154 -6931 200 -6893
rect 154 -6965 160 -6931
rect 194 -6965 200 -6931
rect 154 -7003 200 -6965
rect 154 -7037 160 -7003
rect 194 -7037 200 -7003
rect 154 -7075 200 -7037
rect 154 -7109 160 -7075
rect 194 -7109 200 -7075
rect 154 -7147 200 -7109
rect 154 -7181 160 -7147
rect 194 -7181 200 -7147
rect 154 -7219 200 -7181
rect 154 -7253 160 -7219
rect 194 -7253 200 -7219
rect 154 -7291 200 -7253
rect 154 -7325 160 -7291
rect 194 -7325 200 -7291
rect 154 -7363 200 -7325
rect 154 -7397 160 -7363
rect 194 -7397 200 -7363
rect 154 -7435 200 -7397
rect 154 -7469 160 -7435
rect 194 -7469 200 -7435
rect 154 -7507 200 -7469
rect 154 -7541 160 -7507
rect 194 -7541 200 -7507
rect 154 -7579 200 -7541
rect 154 -7613 160 -7579
rect 194 -7613 200 -7579
rect 154 -7651 200 -7613
rect 154 -7685 160 -7651
rect 194 -7685 200 -7651
rect 154 -7723 200 -7685
rect 154 -7757 160 -7723
rect 194 -7757 200 -7723
rect 154 -7795 200 -7757
rect 154 -7829 160 -7795
rect 194 -7829 200 -7795
rect 154 -7867 200 -7829
rect 154 -7901 160 -7867
rect 194 -7901 200 -7867
rect 154 -7939 200 -7901
rect 154 -7973 160 -7939
rect 194 -7973 200 -7939
rect 154 -8011 200 -7973
rect 154 -8045 160 -8011
rect 194 -8045 200 -8011
rect 154 -8083 200 -8045
rect 154 -8117 160 -8083
rect 194 -8117 200 -8083
rect 154 -8155 200 -8117
rect 154 -8189 160 -8155
rect 194 -8189 200 -8155
rect 154 -8227 200 -8189
rect 154 -8261 160 -8227
rect 194 -8261 200 -8227
rect 154 -8299 200 -8261
rect 154 -8333 160 -8299
rect 194 -8333 200 -8299
rect 154 -8371 200 -8333
rect 154 -8405 160 -8371
rect 194 -8405 200 -8371
rect 154 -8443 200 -8405
rect 154 -8477 160 -8443
rect 194 -8477 200 -8443
rect 154 -8515 200 -8477
rect 154 -8549 160 -8515
rect 194 -8549 200 -8515
rect 154 -8587 200 -8549
rect 154 -8621 160 -8587
rect 194 -8621 200 -8587
rect 154 -8659 200 -8621
rect 154 -8693 160 -8659
rect 194 -8693 200 -8659
rect 154 -8731 200 -8693
rect 154 -8765 160 -8731
rect 194 -8765 200 -8731
rect 154 -8803 200 -8765
rect 154 -8837 160 -8803
rect 194 -8837 200 -8803
rect 154 -8875 200 -8837
rect 154 -8909 160 -8875
rect 194 -8909 200 -8875
rect 154 -8947 200 -8909
rect 154 -8981 160 -8947
rect 194 -8981 200 -8947
rect 154 -9019 200 -8981
rect 154 -9053 160 -9019
rect 194 -9053 200 -9019
rect 154 -9091 200 -9053
rect 154 -9125 160 -9091
rect 194 -9125 200 -9091
rect 154 -9163 200 -9125
rect 154 -9197 160 -9163
rect 194 -9197 200 -9163
rect 154 -9235 200 -9197
rect 154 -9269 160 -9235
rect 194 -9269 200 -9235
rect 154 -9307 200 -9269
rect 154 -9341 160 -9307
rect 194 -9341 200 -9307
rect 154 -9379 200 -9341
rect 154 -9413 160 -9379
rect 194 -9413 200 -9379
rect 154 -9451 200 -9413
rect 154 -9485 160 -9451
rect 194 -9485 200 -9451
rect 154 -9523 200 -9485
rect 154 -9557 160 -9523
rect 194 -9557 200 -9523
rect 154 -9600 200 -9557
rect 272 9557 318 9600
rect 272 9523 278 9557
rect 312 9523 318 9557
rect 272 9485 318 9523
rect 272 9451 278 9485
rect 312 9451 318 9485
rect 272 9413 318 9451
rect 272 9379 278 9413
rect 312 9379 318 9413
rect 272 9341 318 9379
rect 272 9307 278 9341
rect 312 9307 318 9341
rect 272 9269 318 9307
rect 272 9235 278 9269
rect 312 9235 318 9269
rect 272 9197 318 9235
rect 272 9163 278 9197
rect 312 9163 318 9197
rect 272 9125 318 9163
rect 272 9091 278 9125
rect 312 9091 318 9125
rect 272 9053 318 9091
rect 272 9019 278 9053
rect 312 9019 318 9053
rect 272 8981 318 9019
rect 272 8947 278 8981
rect 312 8947 318 8981
rect 272 8909 318 8947
rect 272 8875 278 8909
rect 312 8875 318 8909
rect 272 8837 318 8875
rect 272 8803 278 8837
rect 312 8803 318 8837
rect 272 8765 318 8803
rect 272 8731 278 8765
rect 312 8731 318 8765
rect 272 8693 318 8731
rect 272 8659 278 8693
rect 312 8659 318 8693
rect 272 8621 318 8659
rect 272 8587 278 8621
rect 312 8587 318 8621
rect 272 8549 318 8587
rect 272 8515 278 8549
rect 312 8515 318 8549
rect 272 8477 318 8515
rect 272 8443 278 8477
rect 312 8443 318 8477
rect 272 8405 318 8443
rect 272 8371 278 8405
rect 312 8371 318 8405
rect 272 8333 318 8371
rect 272 8299 278 8333
rect 312 8299 318 8333
rect 272 8261 318 8299
rect 272 8227 278 8261
rect 312 8227 318 8261
rect 272 8189 318 8227
rect 272 8155 278 8189
rect 312 8155 318 8189
rect 272 8117 318 8155
rect 272 8083 278 8117
rect 312 8083 318 8117
rect 272 8045 318 8083
rect 272 8011 278 8045
rect 312 8011 318 8045
rect 272 7973 318 8011
rect 272 7939 278 7973
rect 312 7939 318 7973
rect 272 7901 318 7939
rect 272 7867 278 7901
rect 312 7867 318 7901
rect 272 7829 318 7867
rect 272 7795 278 7829
rect 312 7795 318 7829
rect 272 7757 318 7795
rect 272 7723 278 7757
rect 312 7723 318 7757
rect 272 7685 318 7723
rect 272 7651 278 7685
rect 312 7651 318 7685
rect 272 7613 318 7651
rect 272 7579 278 7613
rect 312 7579 318 7613
rect 272 7541 318 7579
rect 272 7507 278 7541
rect 312 7507 318 7541
rect 272 7469 318 7507
rect 272 7435 278 7469
rect 312 7435 318 7469
rect 272 7397 318 7435
rect 272 7363 278 7397
rect 312 7363 318 7397
rect 272 7325 318 7363
rect 272 7291 278 7325
rect 312 7291 318 7325
rect 272 7253 318 7291
rect 272 7219 278 7253
rect 312 7219 318 7253
rect 272 7181 318 7219
rect 272 7147 278 7181
rect 312 7147 318 7181
rect 272 7109 318 7147
rect 272 7075 278 7109
rect 312 7075 318 7109
rect 272 7037 318 7075
rect 272 7003 278 7037
rect 312 7003 318 7037
rect 272 6965 318 7003
rect 272 6931 278 6965
rect 312 6931 318 6965
rect 272 6893 318 6931
rect 272 6859 278 6893
rect 312 6859 318 6893
rect 272 6821 318 6859
rect 272 6787 278 6821
rect 312 6787 318 6821
rect 272 6749 318 6787
rect 272 6715 278 6749
rect 312 6715 318 6749
rect 272 6677 318 6715
rect 272 6643 278 6677
rect 312 6643 318 6677
rect 272 6605 318 6643
rect 272 6571 278 6605
rect 312 6571 318 6605
rect 272 6533 318 6571
rect 272 6499 278 6533
rect 312 6499 318 6533
rect 272 6461 318 6499
rect 272 6427 278 6461
rect 312 6427 318 6461
rect 272 6389 318 6427
rect 272 6355 278 6389
rect 312 6355 318 6389
rect 272 6317 318 6355
rect 272 6283 278 6317
rect 312 6283 318 6317
rect 272 6245 318 6283
rect 272 6211 278 6245
rect 312 6211 318 6245
rect 272 6173 318 6211
rect 272 6139 278 6173
rect 312 6139 318 6173
rect 272 6101 318 6139
rect 272 6067 278 6101
rect 312 6067 318 6101
rect 272 6029 318 6067
rect 272 5995 278 6029
rect 312 5995 318 6029
rect 272 5957 318 5995
rect 272 5923 278 5957
rect 312 5923 318 5957
rect 272 5885 318 5923
rect 272 5851 278 5885
rect 312 5851 318 5885
rect 272 5813 318 5851
rect 272 5779 278 5813
rect 312 5779 318 5813
rect 272 5741 318 5779
rect 272 5707 278 5741
rect 312 5707 318 5741
rect 272 5669 318 5707
rect 272 5635 278 5669
rect 312 5635 318 5669
rect 272 5597 318 5635
rect 272 5563 278 5597
rect 312 5563 318 5597
rect 272 5525 318 5563
rect 272 5491 278 5525
rect 312 5491 318 5525
rect 272 5453 318 5491
rect 272 5419 278 5453
rect 312 5419 318 5453
rect 272 5381 318 5419
rect 272 5347 278 5381
rect 312 5347 318 5381
rect 272 5309 318 5347
rect 272 5275 278 5309
rect 312 5275 318 5309
rect 272 5237 318 5275
rect 272 5203 278 5237
rect 312 5203 318 5237
rect 272 5165 318 5203
rect 272 5131 278 5165
rect 312 5131 318 5165
rect 272 5093 318 5131
rect 272 5059 278 5093
rect 312 5059 318 5093
rect 272 5021 318 5059
rect 272 4987 278 5021
rect 312 4987 318 5021
rect 272 4949 318 4987
rect 272 4915 278 4949
rect 312 4915 318 4949
rect 272 4877 318 4915
rect 272 4843 278 4877
rect 312 4843 318 4877
rect 272 4805 318 4843
rect 272 4771 278 4805
rect 312 4771 318 4805
rect 272 4733 318 4771
rect 272 4699 278 4733
rect 312 4699 318 4733
rect 272 4661 318 4699
rect 272 4627 278 4661
rect 312 4627 318 4661
rect 272 4589 318 4627
rect 272 4555 278 4589
rect 312 4555 318 4589
rect 272 4517 318 4555
rect 272 4483 278 4517
rect 312 4483 318 4517
rect 272 4445 318 4483
rect 272 4411 278 4445
rect 312 4411 318 4445
rect 272 4373 318 4411
rect 272 4339 278 4373
rect 312 4339 318 4373
rect 272 4301 318 4339
rect 272 4267 278 4301
rect 312 4267 318 4301
rect 272 4229 318 4267
rect 272 4195 278 4229
rect 312 4195 318 4229
rect 272 4157 318 4195
rect 272 4123 278 4157
rect 312 4123 318 4157
rect 272 4085 318 4123
rect 272 4051 278 4085
rect 312 4051 318 4085
rect 272 4013 318 4051
rect 272 3979 278 4013
rect 312 3979 318 4013
rect 272 3941 318 3979
rect 272 3907 278 3941
rect 312 3907 318 3941
rect 272 3869 318 3907
rect 272 3835 278 3869
rect 312 3835 318 3869
rect 272 3797 318 3835
rect 272 3763 278 3797
rect 312 3763 318 3797
rect 272 3725 318 3763
rect 272 3691 278 3725
rect 312 3691 318 3725
rect 272 3653 318 3691
rect 272 3619 278 3653
rect 312 3619 318 3653
rect 272 3581 318 3619
rect 272 3547 278 3581
rect 312 3547 318 3581
rect 272 3509 318 3547
rect 272 3475 278 3509
rect 312 3475 318 3509
rect 272 3437 318 3475
rect 272 3403 278 3437
rect 312 3403 318 3437
rect 272 3365 318 3403
rect 272 3331 278 3365
rect 312 3331 318 3365
rect 272 3293 318 3331
rect 272 3259 278 3293
rect 312 3259 318 3293
rect 272 3221 318 3259
rect 272 3187 278 3221
rect 312 3187 318 3221
rect 272 3149 318 3187
rect 272 3115 278 3149
rect 312 3115 318 3149
rect 272 3077 318 3115
rect 272 3043 278 3077
rect 312 3043 318 3077
rect 272 3005 318 3043
rect 272 2971 278 3005
rect 312 2971 318 3005
rect 272 2933 318 2971
rect 272 2899 278 2933
rect 312 2899 318 2933
rect 272 2861 318 2899
rect 272 2827 278 2861
rect 312 2827 318 2861
rect 272 2789 318 2827
rect 272 2755 278 2789
rect 312 2755 318 2789
rect 272 2717 318 2755
rect 272 2683 278 2717
rect 312 2683 318 2717
rect 272 2645 318 2683
rect 272 2611 278 2645
rect 312 2611 318 2645
rect 272 2573 318 2611
rect 272 2539 278 2573
rect 312 2539 318 2573
rect 272 2501 318 2539
rect 272 2467 278 2501
rect 312 2467 318 2501
rect 272 2429 318 2467
rect 272 2395 278 2429
rect 312 2395 318 2429
rect 272 2357 318 2395
rect 272 2323 278 2357
rect 312 2323 318 2357
rect 272 2285 318 2323
rect 272 2251 278 2285
rect 312 2251 318 2285
rect 272 2213 318 2251
rect 272 2179 278 2213
rect 312 2179 318 2213
rect 272 2141 318 2179
rect 272 2107 278 2141
rect 312 2107 318 2141
rect 272 2069 318 2107
rect 272 2035 278 2069
rect 312 2035 318 2069
rect 272 1997 318 2035
rect 272 1963 278 1997
rect 312 1963 318 1997
rect 272 1925 318 1963
rect 272 1891 278 1925
rect 312 1891 318 1925
rect 272 1853 318 1891
rect 272 1819 278 1853
rect 312 1819 318 1853
rect 272 1781 318 1819
rect 272 1747 278 1781
rect 312 1747 318 1781
rect 272 1709 318 1747
rect 272 1675 278 1709
rect 312 1675 318 1709
rect 272 1637 318 1675
rect 272 1603 278 1637
rect 312 1603 318 1637
rect 272 1565 318 1603
rect 272 1531 278 1565
rect 312 1531 318 1565
rect 272 1493 318 1531
rect 272 1459 278 1493
rect 312 1459 318 1493
rect 272 1421 318 1459
rect 272 1387 278 1421
rect 312 1387 318 1421
rect 272 1349 318 1387
rect 272 1315 278 1349
rect 312 1315 318 1349
rect 272 1277 318 1315
rect 272 1243 278 1277
rect 312 1243 318 1277
rect 272 1205 318 1243
rect 272 1171 278 1205
rect 312 1171 318 1205
rect 272 1133 318 1171
rect 272 1099 278 1133
rect 312 1099 318 1133
rect 272 1061 318 1099
rect 272 1027 278 1061
rect 312 1027 318 1061
rect 272 989 318 1027
rect 272 955 278 989
rect 312 955 318 989
rect 272 917 318 955
rect 272 883 278 917
rect 312 883 318 917
rect 272 845 318 883
rect 272 811 278 845
rect 312 811 318 845
rect 272 773 318 811
rect 272 739 278 773
rect 312 739 318 773
rect 272 701 318 739
rect 272 667 278 701
rect 312 667 318 701
rect 272 629 318 667
rect 272 595 278 629
rect 312 595 318 629
rect 272 557 318 595
rect 272 523 278 557
rect 312 523 318 557
rect 272 485 318 523
rect 272 451 278 485
rect 312 451 318 485
rect 272 413 318 451
rect 272 379 278 413
rect 312 379 318 413
rect 272 341 318 379
rect 272 307 278 341
rect 312 307 318 341
rect 272 269 318 307
rect 272 235 278 269
rect 312 235 318 269
rect 272 197 318 235
rect 272 163 278 197
rect 312 163 318 197
rect 272 125 318 163
rect 272 91 278 125
rect 312 91 318 125
rect 272 53 318 91
rect 272 19 278 53
rect 312 19 318 53
rect 272 -19 318 19
rect 272 -53 278 -19
rect 312 -53 318 -19
rect 272 -91 318 -53
rect 272 -125 278 -91
rect 312 -125 318 -91
rect 272 -163 318 -125
rect 272 -197 278 -163
rect 312 -197 318 -163
rect 272 -235 318 -197
rect 272 -269 278 -235
rect 312 -269 318 -235
rect 272 -307 318 -269
rect 272 -341 278 -307
rect 312 -341 318 -307
rect 272 -379 318 -341
rect 272 -413 278 -379
rect 312 -413 318 -379
rect 272 -451 318 -413
rect 272 -485 278 -451
rect 312 -485 318 -451
rect 272 -523 318 -485
rect 272 -557 278 -523
rect 312 -557 318 -523
rect 272 -595 318 -557
rect 272 -629 278 -595
rect 312 -629 318 -595
rect 272 -667 318 -629
rect 272 -701 278 -667
rect 312 -701 318 -667
rect 272 -739 318 -701
rect 272 -773 278 -739
rect 312 -773 318 -739
rect 272 -811 318 -773
rect 272 -845 278 -811
rect 312 -845 318 -811
rect 272 -883 318 -845
rect 272 -917 278 -883
rect 312 -917 318 -883
rect 272 -955 318 -917
rect 272 -989 278 -955
rect 312 -989 318 -955
rect 272 -1027 318 -989
rect 272 -1061 278 -1027
rect 312 -1061 318 -1027
rect 272 -1099 318 -1061
rect 272 -1133 278 -1099
rect 312 -1133 318 -1099
rect 272 -1171 318 -1133
rect 272 -1205 278 -1171
rect 312 -1205 318 -1171
rect 272 -1243 318 -1205
rect 272 -1277 278 -1243
rect 312 -1277 318 -1243
rect 272 -1315 318 -1277
rect 272 -1349 278 -1315
rect 312 -1349 318 -1315
rect 272 -1387 318 -1349
rect 272 -1421 278 -1387
rect 312 -1421 318 -1387
rect 272 -1459 318 -1421
rect 272 -1493 278 -1459
rect 312 -1493 318 -1459
rect 272 -1531 318 -1493
rect 272 -1565 278 -1531
rect 312 -1565 318 -1531
rect 272 -1603 318 -1565
rect 272 -1637 278 -1603
rect 312 -1637 318 -1603
rect 272 -1675 318 -1637
rect 272 -1709 278 -1675
rect 312 -1709 318 -1675
rect 272 -1747 318 -1709
rect 272 -1781 278 -1747
rect 312 -1781 318 -1747
rect 272 -1819 318 -1781
rect 272 -1853 278 -1819
rect 312 -1853 318 -1819
rect 272 -1891 318 -1853
rect 272 -1925 278 -1891
rect 312 -1925 318 -1891
rect 272 -1963 318 -1925
rect 272 -1997 278 -1963
rect 312 -1997 318 -1963
rect 272 -2035 318 -1997
rect 272 -2069 278 -2035
rect 312 -2069 318 -2035
rect 272 -2107 318 -2069
rect 272 -2141 278 -2107
rect 312 -2141 318 -2107
rect 272 -2179 318 -2141
rect 272 -2213 278 -2179
rect 312 -2213 318 -2179
rect 272 -2251 318 -2213
rect 272 -2285 278 -2251
rect 312 -2285 318 -2251
rect 272 -2323 318 -2285
rect 272 -2357 278 -2323
rect 312 -2357 318 -2323
rect 272 -2395 318 -2357
rect 272 -2429 278 -2395
rect 312 -2429 318 -2395
rect 272 -2467 318 -2429
rect 272 -2501 278 -2467
rect 312 -2501 318 -2467
rect 272 -2539 318 -2501
rect 272 -2573 278 -2539
rect 312 -2573 318 -2539
rect 272 -2611 318 -2573
rect 272 -2645 278 -2611
rect 312 -2645 318 -2611
rect 272 -2683 318 -2645
rect 272 -2717 278 -2683
rect 312 -2717 318 -2683
rect 272 -2755 318 -2717
rect 272 -2789 278 -2755
rect 312 -2789 318 -2755
rect 272 -2827 318 -2789
rect 272 -2861 278 -2827
rect 312 -2861 318 -2827
rect 272 -2899 318 -2861
rect 272 -2933 278 -2899
rect 312 -2933 318 -2899
rect 272 -2971 318 -2933
rect 272 -3005 278 -2971
rect 312 -3005 318 -2971
rect 272 -3043 318 -3005
rect 272 -3077 278 -3043
rect 312 -3077 318 -3043
rect 272 -3115 318 -3077
rect 272 -3149 278 -3115
rect 312 -3149 318 -3115
rect 272 -3187 318 -3149
rect 272 -3221 278 -3187
rect 312 -3221 318 -3187
rect 272 -3259 318 -3221
rect 272 -3293 278 -3259
rect 312 -3293 318 -3259
rect 272 -3331 318 -3293
rect 272 -3365 278 -3331
rect 312 -3365 318 -3331
rect 272 -3403 318 -3365
rect 272 -3437 278 -3403
rect 312 -3437 318 -3403
rect 272 -3475 318 -3437
rect 272 -3509 278 -3475
rect 312 -3509 318 -3475
rect 272 -3547 318 -3509
rect 272 -3581 278 -3547
rect 312 -3581 318 -3547
rect 272 -3619 318 -3581
rect 272 -3653 278 -3619
rect 312 -3653 318 -3619
rect 272 -3691 318 -3653
rect 272 -3725 278 -3691
rect 312 -3725 318 -3691
rect 272 -3763 318 -3725
rect 272 -3797 278 -3763
rect 312 -3797 318 -3763
rect 272 -3835 318 -3797
rect 272 -3869 278 -3835
rect 312 -3869 318 -3835
rect 272 -3907 318 -3869
rect 272 -3941 278 -3907
rect 312 -3941 318 -3907
rect 272 -3979 318 -3941
rect 272 -4013 278 -3979
rect 312 -4013 318 -3979
rect 272 -4051 318 -4013
rect 272 -4085 278 -4051
rect 312 -4085 318 -4051
rect 272 -4123 318 -4085
rect 272 -4157 278 -4123
rect 312 -4157 318 -4123
rect 272 -4195 318 -4157
rect 272 -4229 278 -4195
rect 312 -4229 318 -4195
rect 272 -4267 318 -4229
rect 272 -4301 278 -4267
rect 312 -4301 318 -4267
rect 272 -4339 318 -4301
rect 272 -4373 278 -4339
rect 312 -4373 318 -4339
rect 272 -4411 318 -4373
rect 272 -4445 278 -4411
rect 312 -4445 318 -4411
rect 272 -4483 318 -4445
rect 272 -4517 278 -4483
rect 312 -4517 318 -4483
rect 272 -4555 318 -4517
rect 272 -4589 278 -4555
rect 312 -4589 318 -4555
rect 272 -4627 318 -4589
rect 272 -4661 278 -4627
rect 312 -4661 318 -4627
rect 272 -4699 318 -4661
rect 272 -4733 278 -4699
rect 312 -4733 318 -4699
rect 272 -4771 318 -4733
rect 272 -4805 278 -4771
rect 312 -4805 318 -4771
rect 272 -4843 318 -4805
rect 272 -4877 278 -4843
rect 312 -4877 318 -4843
rect 272 -4915 318 -4877
rect 272 -4949 278 -4915
rect 312 -4949 318 -4915
rect 272 -4987 318 -4949
rect 272 -5021 278 -4987
rect 312 -5021 318 -4987
rect 272 -5059 318 -5021
rect 272 -5093 278 -5059
rect 312 -5093 318 -5059
rect 272 -5131 318 -5093
rect 272 -5165 278 -5131
rect 312 -5165 318 -5131
rect 272 -5203 318 -5165
rect 272 -5237 278 -5203
rect 312 -5237 318 -5203
rect 272 -5275 318 -5237
rect 272 -5309 278 -5275
rect 312 -5309 318 -5275
rect 272 -5347 318 -5309
rect 272 -5381 278 -5347
rect 312 -5381 318 -5347
rect 272 -5419 318 -5381
rect 272 -5453 278 -5419
rect 312 -5453 318 -5419
rect 272 -5491 318 -5453
rect 272 -5525 278 -5491
rect 312 -5525 318 -5491
rect 272 -5563 318 -5525
rect 272 -5597 278 -5563
rect 312 -5597 318 -5563
rect 272 -5635 318 -5597
rect 272 -5669 278 -5635
rect 312 -5669 318 -5635
rect 272 -5707 318 -5669
rect 272 -5741 278 -5707
rect 312 -5741 318 -5707
rect 272 -5779 318 -5741
rect 272 -5813 278 -5779
rect 312 -5813 318 -5779
rect 272 -5851 318 -5813
rect 272 -5885 278 -5851
rect 312 -5885 318 -5851
rect 272 -5923 318 -5885
rect 272 -5957 278 -5923
rect 312 -5957 318 -5923
rect 272 -5995 318 -5957
rect 272 -6029 278 -5995
rect 312 -6029 318 -5995
rect 272 -6067 318 -6029
rect 272 -6101 278 -6067
rect 312 -6101 318 -6067
rect 272 -6139 318 -6101
rect 272 -6173 278 -6139
rect 312 -6173 318 -6139
rect 272 -6211 318 -6173
rect 272 -6245 278 -6211
rect 312 -6245 318 -6211
rect 272 -6283 318 -6245
rect 272 -6317 278 -6283
rect 312 -6317 318 -6283
rect 272 -6355 318 -6317
rect 272 -6389 278 -6355
rect 312 -6389 318 -6355
rect 272 -6427 318 -6389
rect 272 -6461 278 -6427
rect 312 -6461 318 -6427
rect 272 -6499 318 -6461
rect 272 -6533 278 -6499
rect 312 -6533 318 -6499
rect 272 -6571 318 -6533
rect 272 -6605 278 -6571
rect 312 -6605 318 -6571
rect 272 -6643 318 -6605
rect 272 -6677 278 -6643
rect 312 -6677 318 -6643
rect 272 -6715 318 -6677
rect 272 -6749 278 -6715
rect 312 -6749 318 -6715
rect 272 -6787 318 -6749
rect 272 -6821 278 -6787
rect 312 -6821 318 -6787
rect 272 -6859 318 -6821
rect 272 -6893 278 -6859
rect 312 -6893 318 -6859
rect 272 -6931 318 -6893
rect 272 -6965 278 -6931
rect 312 -6965 318 -6931
rect 272 -7003 318 -6965
rect 272 -7037 278 -7003
rect 312 -7037 318 -7003
rect 272 -7075 318 -7037
rect 272 -7109 278 -7075
rect 312 -7109 318 -7075
rect 272 -7147 318 -7109
rect 272 -7181 278 -7147
rect 312 -7181 318 -7147
rect 272 -7219 318 -7181
rect 272 -7253 278 -7219
rect 312 -7253 318 -7219
rect 272 -7291 318 -7253
rect 272 -7325 278 -7291
rect 312 -7325 318 -7291
rect 272 -7363 318 -7325
rect 272 -7397 278 -7363
rect 312 -7397 318 -7363
rect 272 -7435 318 -7397
rect 272 -7469 278 -7435
rect 312 -7469 318 -7435
rect 272 -7507 318 -7469
rect 272 -7541 278 -7507
rect 312 -7541 318 -7507
rect 272 -7579 318 -7541
rect 272 -7613 278 -7579
rect 312 -7613 318 -7579
rect 272 -7651 318 -7613
rect 272 -7685 278 -7651
rect 312 -7685 318 -7651
rect 272 -7723 318 -7685
rect 272 -7757 278 -7723
rect 312 -7757 318 -7723
rect 272 -7795 318 -7757
rect 272 -7829 278 -7795
rect 312 -7829 318 -7795
rect 272 -7867 318 -7829
rect 272 -7901 278 -7867
rect 312 -7901 318 -7867
rect 272 -7939 318 -7901
rect 272 -7973 278 -7939
rect 312 -7973 318 -7939
rect 272 -8011 318 -7973
rect 272 -8045 278 -8011
rect 312 -8045 318 -8011
rect 272 -8083 318 -8045
rect 272 -8117 278 -8083
rect 312 -8117 318 -8083
rect 272 -8155 318 -8117
rect 272 -8189 278 -8155
rect 312 -8189 318 -8155
rect 272 -8227 318 -8189
rect 272 -8261 278 -8227
rect 312 -8261 318 -8227
rect 272 -8299 318 -8261
rect 272 -8333 278 -8299
rect 312 -8333 318 -8299
rect 272 -8371 318 -8333
rect 272 -8405 278 -8371
rect 312 -8405 318 -8371
rect 272 -8443 318 -8405
rect 272 -8477 278 -8443
rect 312 -8477 318 -8443
rect 272 -8515 318 -8477
rect 272 -8549 278 -8515
rect 312 -8549 318 -8515
rect 272 -8587 318 -8549
rect 272 -8621 278 -8587
rect 312 -8621 318 -8587
rect 272 -8659 318 -8621
rect 272 -8693 278 -8659
rect 312 -8693 318 -8659
rect 272 -8731 318 -8693
rect 272 -8765 278 -8731
rect 312 -8765 318 -8731
rect 272 -8803 318 -8765
rect 272 -8837 278 -8803
rect 312 -8837 318 -8803
rect 272 -8875 318 -8837
rect 272 -8909 278 -8875
rect 312 -8909 318 -8875
rect 272 -8947 318 -8909
rect 272 -8981 278 -8947
rect 312 -8981 318 -8947
rect 272 -9019 318 -8981
rect 272 -9053 278 -9019
rect 312 -9053 318 -9019
rect 272 -9091 318 -9053
rect 272 -9125 278 -9091
rect 312 -9125 318 -9091
rect 272 -9163 318 -9125
rect 272 -9197 278 -9163
rect 312 -9197 318 -9163
rect 272 -9235 318 -9197
rect 272 -9269 278 -9235
rect 312 -9269 318 -9235
rect 272 -9307 318 -9269
rect 272 -9341 278 -9307
rect 312 -9341 318 -9307
rect 272 -9379 318 -9341
rect 272 -9413 278 -9379
rect 312 -9413 318 -9379
rect 272 -9451 318 -9413
rect 272 -9485 278 -9451
rect 312 -9485 318 -9451
rect 272 -9523 318 -9485
rect 272 -9557 278 -9523
rect 312 -9557 318 -9523
rect 272 -9600 318 -9557
rect 390 9557 436 9600
rect 390 9523 396 9557
rect 430 9523 436 9557
rect 390 9485 436 9523
rect 390 9451 396 9485
rect 430 9451 436 9485
rect 390 9413 436 9451
rect 390 9379 396 9413
rect 430 9379 436 9413
rect 390 9341 436 9379
rect 390 9307 396 9341
rect 430 9307 436 9341
rect 390 9269 436 9307
rect 390 9235 396 9269
rect 430 9235 436 9269
rect 390 9197 436 9235
rect 390 9163 396 9197
rect 430 9163 436 9197
rect 390 9125 436 9163
rect 390 9091 396 9125
rect 430 9091 436 9125
rect 390 9053 436 9091
rect 390 9019 396 9053
rect 430 9019 436 9053
rect 390 8981 436 9019
rect 390 8947 396 8981
rect 430 8947 436 8981
rect 390 8909 436 8947
rect 390 8875 396 8909
rect 430 8875 436 8909
rect 390 8837 436 8875
rect 390 8803 396 8837
rect 430 8803 436 8837
rect 390 8765 436 8803
rect 390 8731 396 8765
rect 430 8731 436 8765
rect 390 8693 436 8731
rect 390 8659 396 8693
rect 430 8659 436 8693
rect 390 8621 436 8659
rect 390 8587 396 8621
rect 430 8587 436 8621
rect 390 8549 436 8587
rect 390 8515 396 8549
rect 430 8515 436 8549
rect 390 8477 436 8515
rect 390 8443 396 8477
rect 430 8443 436 8477
rect 390 8405 436 8443
rect 390 8371 396 8405
rect 430 8371 436 8405
rect 390 8333 436 8371
rect 390 8299 396 8333
rect 430 8299 436 8333
rect 390 8261 436 8299
rect 390 8227 396 8261
rect 430 8227 436 8261
rect 390 8189 436 8227
rect 390 8155 396 8189
rect 430 8155 436 8189
rect 390 8117 436 8155
rect 390 8083 396 8117
rect 430 8083 436 8117
rect 390 8045 436 8083
rect 390 8011 396 8045
rect 430 8011 436 8045
rect 390 7973 436 8011
rect 390 7939 396 7973
rect 430 7939 436 7973
rect 390 7901 436 7939
rect 390 7867 396 7901
rect 430 7867 436 7901
rect 390 7829 436 7867
rect 390 7795 396 7829
rect 430 7795 436 7829
rect 390 7757 436 7795
rect 390 7723 396 7757
rect 430 7723 436 7757
rect 390 7685 436 7723
rect 390 7651 396 7685
rect 430 7651 436 7685
rect 390 7613 436 7651
rect 390 7579 396 7613
rect 430 7579 436 7613
rect 390 7541 436 7579
rect 390 7507 396 7541
rect 430 7507 436 7541
rect 390 7469 436 7507
rect 390 7435 396 7469
rect 430 7435 436 7469
rect 390 7397 436 7435
rect 390 7363 396 7397
rect 430 7363 436 7397
rect 390 7325 436 7363
rect 390 7291 396 7325
rect 430 7291 436 7325
rect 390 7253 436 7291
rect 390 7219 396 7253
rect 430 7219 436 7253
rect 390 7181 436 7219
rect 390 7147 396 7181
rect 430 7147 436 7181
rect 390 7109 436 7147
rect 390 7075 396 7109
rect 430 7075 436 7109
rect 390 7037 436 7075
rect 390 7003 396 7037
rect 430 7003 436 7037
rect 390 6965 436 7003
rect 390 6931 396 6965
rect 430 6931 436 6965
rect 390 6893 436 6931
rect 390 6859 396 6893
rect 430 6859 436 6893
rect 390 6821 436 6859
rect 390 6787 396 6821
rect 430 6787 436 6821
rect 390 6749 436 6787
rect 390 6715 396 6749
rect 430 6715 436 6749
rect 390 6677 436 6715
rect 390 6643 396 6677
rect 430 6643 436 6677
rect 390 6605 436 6643
rect 390 6571 396 6605
rect 430 6571 436 6605
rect 390 6533 436 6571
rect 390 6499 396 6533
rect 430 6499 436 6533
rect 390 6461 436 6499
rect 390 6427 396 6461
rect 430 6427 436 6461
rect 390 6389 436 6427
rect 390 6355 396 6389
rect 430 6355 436 6389
rect 390 6317 436 6355
rect 390 6283 396 6317
rect 430 6283 436 6317
rect 390 6245 436 6283
rect 390 6211 396 6245
rect 430 6211 436 6245
rect 390 6173 436 6211
rect 390 6139 396 6173
rect 430 6139 436 6173
rect 390 6101 436 6139
rect 390 6067 396 6101
rect 430 6067 436 6101
rect 390 6029 436 6067
rect 390 5995 396 6029
rect 430 5995 436 6029
rect 390 5957 436 5995
rect 390 5923 396 5957
rect 430 5923 436 5957
rect 390 5885 436 5923
rect 390 5851 396 5885
rect 430 5851 436 5885
rect 390 5813 436 5851
rect 390 5779 396 5813
rect 430 5779 436 5813
rect 390 5741 436 5779
rect 390 5707 396 5741
rect 430 5707 436 5741
rect 390 5669 436 5707
rect 390 5635 396 5669
rect 430 5635 436 5669
rect 390 5597 436 5635
rect 390 5563 396 5597
rect 430 5563 436 5597
rect 390 5525 436 5563
rect 390 5491 396 5525
rect 430 5491 436 5525
rect 390 5453 436 5491
rect 390 5419 396 5453
rect 430 5419 436 5453
rect 390 5381 436 5419
rect 390 5347 396 5381
rect 430 5347 436 5381
rect 390 5309 436 5347
rect 390 5275 396 5309
rect 430 5275 436 5309
rect 390 5237 436 5275
rect 390 5203 396 5237
rect 430 5203 436 5237
rect 390 5165 436 5203
rect 390 5131 396 5165
rect 430 5131 436 5165
rect 390 5093 436 5131
rect 390 5059 396 5093
rect 430 5059 436 5093
rect 390 5021 436 5059
rect 390 4987 396 5021
rect 430 4987 436 5021
rect 390 4949 436 4987
rect 390 4915 396 4949
rect 430 4915 436 4949
rect 390 4877 436 4915
rect 390 4843 396 4877
rect 430 4843 436 4877
rect 390 4805 436 4843
rect 390 4771 396 4805
rect 430 4771 436 4805
rect 390 4733 436 4771
rect 390 4699 396 4733
rect 430 4699 436 4733
rect 390 4661 436 4699
rect 390 4627 396 4661
rect 430 4627 436 4661
rect 390 4589 436 4627
rect 390 4555 396 4589
rect 430 4555 436 4589
rect 390 4517 436 4555
rect 390 4483 396 4517
rect 430 4483 436 4517
rect 390 4445 436 4483
rect 390 4411 396 4445
rect 430 4411 436 4445
rect 390 4373 436 4411
rect 390 4339 396 4373
rect 430 4339 436 4373
rect 390 4301 436 4339
rect 390 4267 396 4301
rect 430 4267 436 4301
rect 390 4229 436 4267
rect 390 4195 396 4229
rect 430 4195 436 4229
rect 390 4157 436 4195
rect 390 4123 396 4157
rect 430 4123 436 4157
rect 390 4085 436 4123
rect 390 4051 396 4085
rect 430 4051 436 4085
rect 390 4013 436 4051
rect 390 3979 396 4013
rect 430 3979 436 4013
rect 390 3941 436 3979
rect 390 3907 396 3941
rect 430 3907 436 3941
rect 390 3869 436 3907
rect 390 3835 396 3869
rect 430 3835 436 3869
rect 390 3797 436 3835
rect 390 3763 396 3797
rect 430 3763 436 3797
rect 390 3725 436 3763
rect 390 3691 396 3725
rect 430 3691 436 3725
rect 390 3653 436 3691
rect 390 3619 396 3653
rect 430 3619 436 3653
rect 390 3581 436 3619
rect 390 3547 396 3581
rect 430 3547 436 3581
rect 390 3509 436 3547
rect 390 3475 396 3509
rect 430 3475 436 3509
rect 390 3437 436 3475
rect 390 3403 396 3437
rect 430 3403 436 3437
rect 390 3365 436 3403
rect 390 3331 396 3365
rect 430 3331 436 3365
rect 390 3293 436 3331
rect 390 3259 396 3293
rect 430 3259 436 3293
rect 390 3221 436 3259
rect 390 3187 396 3221
rect 430 3187 436 3221
rect 390 3149 436 3187
rect 390 3115 396 3149
rect 430 3115 436 3149
rect 390 3077 436 3115
rect 390 3043 396 3077
rect 430 3043 436 3077
rect 390 3005 436 3043
rect 390 2971 396 3005
rect 430 2971 436 3005
rect 390 2933 436 2971
rect 390 2899 396 2933
rect 430 2899 436 2933
rect 390 2861 436 2899
rect 390 2827 396 2861
rect 430 2827 436 2861
rect 390 2789 436 2827
rect 390 2755 396 2789
rect 430 2755 436 2789
rect 390 2717 436 2755
rect 390 2683 396 2717
rect 430 2683 436 2717
rect 390 2645 436 2683
rect 390 2611 396 2645
rect 430 2611 436 2645
rect 390 2573 436 2611
rect 390 2539 396 2573
rect 430 2539 436 2573
rect 390 2501 436 2539
rect 390 2467 396 2501
rect 430 2467 436 2501
rect 390 2429 436 2467
rect 390 2395 396 2429
rect 430 2395 436 2429
rect 390 2357 436 2395
rect 390 2323 396 2357
rect 430 2323 436 2357
rect 390 2285 436 2323
rect 390 2251 396 2285
rect 430 2251 436 2285
rect 390 2213 436 2251
rect 390 2179 396 2213
rect 430 2179 436 2213
rect 390 2141 436 2179
rect 390 2107 396 2141
rect 430 2107 436 2141
rect 390 2069 436 2107
rect 390 2035 396 2069
rect 430 2035 436 2069
rect 390 1997 436 2035
rect 390 1963 396 1997
rect 430 1963 436 1997
rect 390 1925 436 1963
rect 390 1891 396 1925
rect 430 1891 436 1925
rect 390 1853 436 1891
rect 390 1819 396 1853
rect 430 1819 436 1853
rect 390 1781 436 1819
rect 390 1747 396 1781
rect 430 1747 436 1781
rect 390 1709 436 1747
rect 390 1675 396 1709
rect 430 1675 436 1709
rect 390 1637 436 1675
rect 390 1603 396 1637
rect 430 1603 436 1637
rect 390 1565 436 1603
rect 390 1531 396 1565
rect 430 1531 436 1565
rect 390 1493 436 1531
rect 390 1459 396 1493
rect 430 1459 436 1493
rect 390 1421 436 1459
rect 390 1387 396 1421
rect 430 1387 436 1421
rect 390 1349 436 1387
rect 390 1315 396 1349
rect 430 1315 436 1349
rect 390 1277 436 1315
rect 390 1243 396 1277
rect 430 1243 436 1277
rect 390 1205 436 1243
rect 390 1171 396 1205
rect 430 1171 436 1205
rect 390 1133 436 1171
rect 390 1099 396 1133
rect 430 1099 436 1133
rect 390 1061 436 1099
rect 390 1027 396 1061
rect 430 1027 436 1061
rect 390 989 436 1027
rect 390 955 396 989
rect 430 955 436 989
rect 390 917 436 955
rect 390 883 396 917
rect 430 883 436 917
rect 390 845 436 883
rect 390 811 396 845
rect 430 811 436 845
rect 390 773 436 811
rect 390 739 396 773
rect 430 739 436 773
rect 390 701 436 739
rect 390 667 396 701
rect 430 667 436 701
rect 390 629 436 667
rect 390 595 396 629
rect 430 595 436 629
rect 390 557 436 595
rect 390 523 396 557
rect 430 523 436 557
rect 390 485 436 523
rect 390 451 396 485
rect 430 451 436 485
rect 390 413 436 451
rect 390 379 396 413
rect 430 379 436 413
rect 390 341 436 379
rect 390 307 396 341
rect 430 307 436 341
rect 390 269 436 307
rect 390 235 396 269
rect 430 235 436 269
rect 390 197 436 235
rect 390 163 396 197
rect 430 163 436 197
rect 390 125 436 163
rect 390 91 396 125
rect 430 91 436 125
rect 390 53 436 91
rect 390 19 396 53
rect 430 19 436 53
rect 390 -19 436 19
rect 390 -53 396 -19
rect 430 -53 436 -19
rect 390 -91 436 -53
rect 390 -125 396 -91
rect 430 -125 436 -91
rect 390 -163 436 -125
rect 390 -197 396 -163
rect 430 -197 436 -163
rect 390 -235 436 -197
rect 390 -269 396 -235
rect 430 -269 436 -235
rect 390 -307 436 -269
rect 390 -341 396 -307
rect 430 -341 436 -307
rect 390 -379 436 -341
rect 390 -413 396 -379
rect 430 -413 436 -379
rect 390 -451 436 -413
rect 390 -485 396 -451
rect 430 -485 436 -451
rect 390 -523 436 -485
rect 390 -557 396 -523
rect 430 -557 436 -523
rect 390 -595 436 -557
rect 390 -629 396 -595
rect 430 -629 436 -595
rect 390 -667 436 -629
rect 390 -701 396 -667
rect 430 -701 436 -667
rect 390 -739 436 -701
rect 390 -773 396 -739
rect 430 -773 436 -739
rect 390 -811 436 -773
rect 390 -845 396 -811
rect 430 -845 436 -811
rect 390 -883 436 -845
rect 390 -917 396 -883
rect 430 -917 436 -883
rect 390 -955 436 -917
rect 390 -989 396 -955
rect 430 -989 436 -955
rect 390 -1027 436 -989
rect 390 -1061 396 -1027
rect 430 -1061 436 -1027
rect 390 -1099 436 -1061
rect 390 -1133 396 -1099
rect 430 -1133 436 -1099
rect 390 -1171 436 -1133
rect 390 -1205 396 -1171
rect 430 -1205 436 -1171
rect 390 -1243 436 -1205
rect 390 -1277 396 -1243
rect 430 -1277 436 -1243
rect 390 -1315 436 -1277
rect 390 -1349 396 -1315
rect 430 -1349 436 -1315
rect 390 -1387 436 -1349
rect 390 -1421 396 -1387
rect 430 -1421 436 -1387
rect 390 -1459 436 -1421
rect 390 -1493 396 -1459
rect 430 -1493 436 -1459
rect 390 -1531 436 -1493
rect 390 -1565 396 -1531
rect 430 -1565 436 -1531
rect 390 -1603 436 -1565
rect 390 -1637 396 -1603
rect 430 -1637 436 -1603
rect 390 -1675 436 -1637
rect 390 -1709 396 -1675
rect 430 -1709 436 -1675
rect 390 -1747 436 -1709
rect 390 -1781 396 -1747
rect 430 -1781 436 -1747
rect 390 -1819 436 -1781
rect 390 -1853 396 -1819
rect 430 -1853 436 -1819
rect 390 -1891 436 -1853
rect 390 -1925 396 -1891
rect 430 -1925 436 -1891
rect 390 -1963 436 -1925
rect 390 -1997 396 -1963
rect 430 -1997 436 -1963
rect 390 -2035 436 -1997
rect 390 -2069 396 -2035
rect 430 -2069 436 -2035
rect 390 -2107 436 -2069
rect 390 -2141 396 -2107
rect 430 -2141 436 -2107
rect 390 -2179 436 -2141
rect 390 -2213 396 -2179
rect 430 -2213 436 -2179
rect 390 -2251 436 -2213
rect 390 -2285 396 -2251
rect 430 -2285 436 -2251
rect 390 -2323 436 -2285
rect 390 -2357 396 -2323
rect 430 -2357 436 -2323
rect 390 -2395 436 -2357
rect 390 -2429 396 -2395
rect 430 -2429 436 -2395
rect 390 -2467 436 -2429
rect 390 -2501 396 -2467
rect 430 -2501 436 -2467
rect 390 -2539 436 -2501
rect 390 -2573 396 -2539
rect 430 -2573 436 -2539
rect 390 -2611 436 -2573
rect 390 -2645 396 -2611
rect 430 -2645 436 -2611
rect 390 -2683 436 -2645
rect 390 -2717 396 -2683
rect 430 -2717 436 -2683
rect 390 -2755 436 -2717
rect 390 -2789 396 -2755
rect 430 -2789 436 -2755
rect 390 -2827 436 -2789
rect 390 -2861 396 -2827
rect 430 -2861 436 -2827
rect 390 -2899 436 -2861
rect 390 -2933 396 -2899
rect 430 -2933 436 -2899
rect 390 -2971 436 -2933
rect 390 -3005 396 -2971
rect 430 -3005 436 -2971
rect 390 -3043 436 -3005
rect 390 -3077 396 -3043
rect 430 -3077 436 -3043
rect 390 -3115 436 -3077
rect 390 -3149 396 -3115
rect 430 -3149 436 -3115
rect 390 -3187 436 -3149
rect 390 -3221 396 -3187
rect 430 -3221 436 -3187
rect 390 -3259 436 -3221
rect 390 -3293 396 -3259
rect 430 -3293 436 -3259
rect 390 -3331 436 -3293
rect 390 -3365 396 -3331
rect 430 -3365 436 -3331
rect 390 -3403 436 -3365
rect 390 -3437 396 -3403
rect 430 -3437 436 -3403
rect 390 -3475 436 -3437
rect 390 -3509 396 -3475
rect 430 -3509 436 -3475
rect 390 -3547 436 -3509
rect 390 -3581 396 -3547
rect 430 -3581 436 -3547
rect 390 -3619 436 -3581
rect 390 -3653 396 -3619
rect 430 -3653 436 -3619
rect 390 -3691 436 -3653
rect 390 -3725 396 -3691
rect 430 -3725 436 -3691
rect 390 -3763 436 -3725
rect 390 -3797 396 -3763
rect 430 -3797 436 -3763
rect 390 -3835 436 -3797
rect 390 -3869 396 -3835
rect 430 -3869 436 -3835
rect 390 -3907 436 -3869
rect 390 -3941 396 -3907
rect 430 -3941 436 -3907
rect 390 -3979 436 -3941
rect 390 -4013 396 -3979
rect 430 -4013 436 -3979
rect 390 -4051 436 -4013
rect 390 -4085 396 -4051
rect 430 -4085 436 -4051
rect 390 -4123 436 -4085
rect 390 -4157 396 -4123
rect 430 -4157 436 -4123
rect 390 -4195 436 -4157
rect 390 -4229 396 -4195
rect 430 -4229 436 -4195
rect 390 -4267 436 -4229
rect 390 -4301 396 -4267
rect 430 -4301 436 -4267
rect 390 -4339 436 -4301
rect 390 -4373 396 -4339
rect 430 -4373 436 -4339
rect 390 -4411 436 -4373
rect 390 -4445 396 -4411
rect 430 -4445 436 -4411
rect 390 -4483 436 -4445
rect 390 -4517 396 -4483
rect 430 -4517 436 -4483
rect 390 -4555 436 -4517
rect 390 -4589 396 -4555
rect 430 -4589 436 -4555
rect 390 -4627 436 -4589
rect 390 -4661 396 -4627
rect 430 -4661 436 -4627
rect 390 -4699 436 -4661
rect 390 -4733 396 -4699
rect 430 -4733 436 -4699
rect 390 -4771 436 -4733
rect 390 -4805 396 -4771
rect 430 -4805 436 -4771
rect 390 -4843 436 -4805
rect 390 -4877 396 -4843
rect 430 -4877 436 -4843
rect 390 -4915 436 -4877
rect 390 -4949 396 -4915
rect 430 -4949 436 -4915
rect 390 -4987 436 -4949
rect 390 -5021 396 -4987
rect 430 -5021 436 -4987
rect 390 -5059 436 -5021
rect 390 -5093 396 -5059
rect 430 -5093 436 -5059
rect 390 -5131 436 -5093
rect 390 -5165 396 -5131
rect 430 -5165 436 -5131
rect 390 -5203 436 -5165
rect 390 -5237 396 -5203
rect 430 -5237 436 -5203
rect 390 -5275 436 -5237
rect 390 -5309 396 -5275
rect 430 -5309 436 -5275
rect 390 -5347 436 -5309
rect 390 -5381 396 -5347
rect 430 -5381 436 -5347
rect 390 -5419 436 -5381
rect 390 -5453 396 -5419
rect 430 -5453 436 -5419
rect 390 -5491 436 -5453
rect 390 -5525 396 -5491
rect 430 -5525 436 -5491
rect 390 -5563 436 -5525
rect 390 -5597 396 -5563
rect 430 -5597 436 -5563
rect 390 -5635 436 -5597
rect 390 -5669 396 -5635
rect 430 -5669 436 -5635
rect 390 -5707 436 -5669
rect 390 -5741 396 -5707
rect 430 -5741 436 -5707
rect 390 -5779 436 -5741
rect 390 -5813 396 -5779
rect 430 -5813 436 -5779
rect 390 -5851 436 -5813
rect 390 -5885 396 -5851
rect 430 -5885 436 -5851
rect 390 -5923 436 -5885
rect 390 -5957 396 -5923
rect 430 -5957 436 -5923
rect 390 -5995 436 -5957
rect 390 -6029 396 -5995
rect 430 -6029 436 -5995
rect 390 -6067 436 -6029
rect 390 -6101 396 -6067
rect 430 -6101 436 -6067
rect 390 -6139 436 -6101
rect 390 -6173 396 -6139
rect 430 -6173 436 -6139
rect 390 -6211 436 -6173
rect 390 -6245 396 -6211
rect 430 -6245 436 -6211
rect 390 -6283 436 -6245
rect 390 -6317 396 -6283
rect 430 -6317 436 -6283
rect 390 -6355 436 -6317
rect 390 -6389 396 -6355
rect 430 -6389 436 -6355
rect 390 -6427 436 -6389
rect 390 -6461 396 -6427
rect 430 -6461 436 -6427
rect 390 -6499 436 -6461
rect 390 -6533 396 -6499
rect 430 -6533 436 -6499
rect 390 -6571 436 -6533
rect 390 -6605 396 -6571
rect 430 -6605 436 -6571
rect 390 -6643 436 -6605
rect 390 -6677 396 -6643
rect 430 -6677 436 -6643
rect 390 -6715 436 -6677
rect 390 -6749 396 -6715
rect 430 -6749 436 -6715
rect 390 -6787 436 -6749
rect 390 -6821 396 -6787
rect 430 -6821 436 -6787
rect 390 -6859 436 -6821
rect 390 -6893 396 -6859
rect 430 -6893 436 -6859
rect 390 -6931 436 -6893
rect 390 -6965 396 -6931
rect 430 -6965 436 -6931
rect 390 -7003 436 -6965
rect 390 -7037 396 -7003
rect 430 -7037 436 -7003
rect 390 -7075 436 -7037
rect 390 -7109 396 -7075
rect 430 -7109 436 -7075
rect 390 -7147 436 -7109
rect 390 -7181 396 -7147
rect 430 -7181 436 -7147
rect 390 -7219 436 -7181
rect 390 -7253 396 -7219
rect 430 -7253 436 -7219
rect 390 -7291 436 -7253
rect 390 -7325 396 -7291
rect 430 -7325 436 -7291
rect 390 -7363 436 -7325
rect 390 -7397 396 -7363
rect 430 -7397 436 -7363
rect 390 -7435 436 -7397
rect 390 -7469 396 -7435
rect 430 -7469 436 -7435
rect 390 -7507 436 -7469
rect 390 -7541 396 -7507
rect 430 -7541 436 -7507
rect 390 -7579 436 -7541
rect 390 -7613 396 -7579
rect 430 -7613 436 -7579
rect 390 -7651 436 -7613
rect 390 -7685 396 -7651
rect 430 -7685 436 -7651
rect 390 -7723 436 -7685
rect 390 -7757 396 -7723
rect 430 -7757 436 -7723
rect 390 -7795 436 -7757
rect 390 -7829 396 -7795
rect 430 -7829 436 -7795
rect 390 -7867 436 -7829
rect 390 -7901 396 -7867
rect 430 -7901 436 -7867
rect 390 -7939 436 -7901
rect 390 -7973 396 -7939
rect 430 -7973 436 -7939
rect 390 -8011 436 -7973
rect 390 -8045 396 -8011
rect 430 -8045 436 -8011
rect 390 -8083 436 -8045
rect 390 -8117 396 -8083
rect 430 -8117 436 -8083
rect 390 -8155 436 -8117
rect 390 -8189 396 -8155
rect 430 -8189 436 -8155
rect 390 -8227 436 -8189
rect 390 -8261 396 -8227
rect 430 -8261 436 -8227
rect 390 -8299 436 -8261
rect 390 -8333 396 -8299
rect 430 -8333 436 -8299
rect 390 -8371 436 -8333
rect 390 -8405 396 -8371
rect 430 -8405 436 -8371
rect 390 -8443 436 -8405
rect 390 -8477 396 -8443
rect 430 -8477 436 -8443
rect 390 -8515 436 -8477
rect 390 -8549 396 -8515
rect 430 -8549 436 -8515
rect 390 -8587 436 -8549
rect 390 -8621 396 -8587
rect 430 -8621 436 -8587
rect 390 -8659 436 -8621
rect 390 -8693 396 -8659
rect 430 -8693 436 -8659
rect 390 -8731 436 -8693
rect 390 -8765 396 -8731
rect 430 -8765 436 -8731
rect 390 -8803 436 -8765
rect 390 -8837 396 -8803
rect 430 -8837 436 -8803
rect 390 -8875 436 -8837
rect 390 -8909 396 -8875
rect 430 -8909 436 -8875
rect 390 -8947 436 -8909
rect 390 -8981 396 -8947
rect 430 -8981 436 -8947
rect 390 -9019 436 -8981
rect 390 -9053 396 -9019
rect 430 -9053 436 -9019
rect 390 -9091 436 -9053
rect 390 -9125 396 -9091
rect 430 -9125 436 -9091
rect 390 -9163 436 -9125
rect 390 -9197 396 -9163
rect 430 -9197 436 -9163
rect 390 -9235 436 -9197
rect 390 -9269 396 -9235
rect 430 -9269 436 -9235
rect 390 -9307 436 -9269
rect 390 -9341 396 -9307
rect 430 -9341 436 -9307
rect 390 -9379 436 -9341
rect 390 -9413 396 -9379
rect 430 -9413 436 -9379
rect 390 -9451 436 -9413
rect 390 -9485 396 -9451
rect 430 -9485 436 -9451
rect 390 -9523 436 -9485
rect 390 -9557 396 -9523
rect 430 -9557 436 -9523
rect 390 -9600 436 -9557
rect 508 9557 554 9600
rect 508 9523 514 9557
rect 548 9523 554 9557
rect 508 9485 554 9523
rect 508 9451 514 9485
rect 548 9451 554 9485
rect 508 9413 554 9451
rect 508 9379 514 9413
rect 548 9379 554 9413
rect 508 9341 554 9379
rect 508 9307 514 9341
rect 548 9307 554 9341
rect 508 9269 554 9307
rect 508 9235 514 9269
rect 548 9235 554 9269
rect 508 9197 554 9235
rect 508 9163 514 9197
rect 548 9163 554 9197
rect 508 9125 554 9163
rect 508 9091 514 9125
rect 548 9091 554 9125
rect 508 9053 554 9091
rect 508 9019 514 9053
rect 548 9019 554 9053
rect 508 8981 554 9019
rect 508 8947 514 8981
rect 548 8947 554 8981
rect 508 8909 554 8947
rect 508 8875 514 8909
rect 548 8875 554 8909
rect 508 8837 554 8875
rect 508 8803 514 8837
rect 548 8803 554 8837
rect 508 8765 554 8803
rect 508 8731 514 8765
rect 548 8731 554 8765
rect 508 8693 554 8731
rect 508 8659 514 8693
rect 548 8659 554 8693
rect 508 8621 554 8659
rect 508 8587 514 8621
rect 548 8587 554 8621
rect 508 8549 554 8587
rect 508 8515 514 8549
rect 548 8515 554 8549
rect 508 8477 554 8515
rect 508 8443 514 8477
rect 548 8443 554 8477
rect 508 8405 554 8443
rect 508 8371 514 8405
rect 548 8371 554 8405
rect 508 8333 554 8371
rect 508 8299 514 8333
rect 548 8299 554 8333
rect 508 8261 554 8299
rect 508 8227 514 8261
rect 548 8227 554 8261
rect 508 8189 554 8227
rect 508 8155 514 8189
rect 548 8155 554 8189
rect 508 8117 554 8155
rect 508 8083 514 8117
rect 548 8083 554 8117
rect 508 8045 554 8083
rect 508 8011 514 8045
rect 548 8011 554 8045
rect 508 7973 554 8011
rect 508 7939 514 7973
rect 548 7939 554 7973
rect 508 7901 554 7939
rect 508 7867 514 7901
rect 548 7867 554 7901
rect 508 7829 554 7867
rect 508 7795 514 7829
rect 548 7795 554 7829
rect 508 7757 554 7795
rect 508 7723 514 7757
rect 548 7723 554 7757
rect 508 7685 554 7723
rect 508 7651 514 7685
rect 548 7651 554 7685
rect 508 7613 554 7651
rect 508 7579 514 7613
rect 548 7579 554 7613
rect 508 7541 554 7579
rect 508 7507 514 7541
rect 548 7507 554 7541
rect 508 7469 554 7507
rect 508 7435 514 7469
rect 548 7435 554 7469
rect 508 7397 554 7435
rect 508 7363 514 7397
rect 548 7363 554 7397
rect 508 7325 554 7363
rect 508 7291 514 7325
rect 548 7291 554 7325
rect 508 7253 554 7291
rect 508 7219 514 7253
rect 548 7219 554 7253
rect 508 7181 554 7219
rect 508 7147 514 7181
rect 548 7147 554 7181
rect 508 7109 554 7147
rect 508 7075 514 7109
rect 548 7075 554 7109
rect 508 7037 554 7075
rect 508 7003 514 7037
rect 548 7003 554 7037
rect 508 6965 554 7003
rect 508 6931 514 6965
rect 548 6931 554 6965
rect 508 6893 554 6931
rect 508 6859 514 6893
rect 548 6859 554 6893
rect 508 6821 554 6859
rect 508 6787 514 6821
rect 548 6787 554 6821
rect 508 6749 554 6787
rect 508 6715 514 6749
rect 548 6715 554 6749
rect 508 6677 554 6715
rect 508 6643 514 6677
rect 548 6643 554 6677
rect 508 6605 554 6643
rect 508 6571 514 6605
rect 548 6571 554 6605
rect 508 6533 554 6571
rect 508 6499 514 6533
rect 548 6499 554 6533
rect 508 6461 554 6499
rect 508 6427 514 6461
rect 548 6427 554 6461
rect 508 6389 554 6427
rect 508 6355 514 6389
rect 548 6355 554 6389
rect 508 6317 554 6355
rect 508 6283 514 6317
rect 548 6283 554 6317
rect 508 6245 554 6283
rect 508 6211 514 6245
rect 548 6211 554 6245
rect 508 6173 554 6211
rect 508 6139 514 6173
rect 548 6139 554 6173
rect 508 6101 554 6139
rect 508 6067 514 6101
rect 548 6067 554 6101
rect 508 6029 554 6067
rect 508 5995 514 6029
rect 548 5995 554 6029
rect 508 5957 554 5995
rect 508 5923 514 5957
rect 548 5923 554 5957
rect 508 5885 554 5923
rect 508 5851 514 5885
rect 548 5851 554 5885
rect 508 5813 554 5851
rect 508 5779 514 5813
rect 548 5779 554 5813
rect 508 5741 554 5779
rect 508 5707 514 5741
rect 548 5707 554 5741
rect 508 5669 554 5707
rect 508 5635 514 5669
rect 548 5635 554 5669
rect 508 5597 554 5635
rect 508 5563 514 5597
rect 548 5563 554 5597
rect 508 5525 554 5563
rect 508 5491 514 5525
rect 548 5491 554 5525
rect 508 5453 554 5491
rect 508 5419 514 5453
rect 548 5419 554 5453
rect 508 5381 554 5419
rect 508 5347 514 5381
rect 548 5347 554 5381
rect 508 5309 554 5347
rect 508 5275 514 5309
rect 548 5275 554 5309
rect 508 5237 554 5275
rect 508 5203 514 5237
rect 548 5203 554 5237
rect 508 5165 554 5203
rect 508 5131 514 5165
rect 548 5131 554 5165
rect 508 5093 554 5131
rect 508 5059 514 5093
rect 548 5059 554 5093
rect 508 5021 554 5059
rect 508 4987 514 5021
rect 548 4987 554 5021
rect 508 4949 554 4987
rect 508 4915 514 4949
rect 548 4915 554 4949
rect 508 4877 554 4915
rect 508 4843 514 4877
rect 548 4843 554 4877
rect 508 4805 554 4843
rect 508 4771 514 4805
rect 548 4771 554 4805
rect 508 4733 554 4771
rect 508 4699 514 4733
rect 548 4699 554 4733
rect 508 4661 554 4699
rect 508 4627 514 4661
rect 548 4627 554 4661
rect 508 4589 554 4627
rect 508 4555 514 4589
rect 548 4555 554 4589
rect 508 4517 554 4555
rect 508 4483 514 4517
rect 548 4483 554 4517
rect 508 4445 554 4483
rect 508 4411 514 4445
rect 548 4411 554 4445
rect 508 4373 554 4411
rect 508 4339 514 4373
rect 548 4339 554 4373
rect 508 4301 554 4339
rect 508 4267 514 4301
rect 548 4267 554 4301
rect 508 4229 554 4267
rect 508 4195 514 4229
rect 548 4195 554 4229
rect 508 4157 554 4195
rect 508 4123 514 4157
rect 548 4123 554 4157
rect 508 4085 554 4123
rect 508 4051 514 4085
rect 548 4051 554 4085
rect 508 4013 554 4051
rect 508 3979 514 4013
rect 548 3979 554 4013
rect 508 3941 554 3979
rect 508 3907 514 3941
rect 548 3907 554 3941
rect 508 3869 554 3907
rect 508 3835 514 3869
rect 548 3835 554 3869
rect 508 3797 554 3835
rect 508 3763 514 3797
rect 548 3763 554 3797
rect 508 3725 554 3763
rect 508 3691 514 3725
rect 548 3691 554 3725
rect 508 3653 554 3691
rect 508 3619 514 3653
rect 548 3619 554 3653
rect 508 3581 554 3619
rect 508 3547 514 3581
rect 548 3547 554 3581
rect 508 3509 554 3547
rect 508 3475 514 3509
rect 548 3475 554 3509
rect 508 3437 554 3475
rect 508 3403 514 3437
rect 548 3403 554 3437
rect 508 3365 554 3403
rect 508 3331 514 3365
rect 548 3331 554 3365
rect 508 3293 554 3331
rect 508 3259 514 3293
rect 548 3259 554 3293
rect 508 3221 554 3259
rect 508 3187 514 3221
rect 548 3187 554 3221
rect 508 3149 554 3187
rect 508 3115 514 3149
rect 548 3115 554 3149
rect 508 3077 554 3115
rect 508 3043 514 3077
rect 548 3043 554 3077
rect 508 3005 554 3043
rect 508 2971 514 3005
rect 548 2971 554 3005
rect 508 2933 554 2971
rect 508 2899 514 2933
rect 548 2899 554 2933
rect 508 2861 554 2899
rect 508 2827 514 2861
rect 548 2827 554 2861
rect 508 2789 554 2827
rect 508 2755 514 2789
rect 548 2755 554 2789
rect 508 2717 554 2755
rect 508 2683 514 2717
rect 548 2683 554 2717
rect 508 2645 554 2683
rect 508 2611 514 2645
rect 548 2611 554 2645
rect 508 2573 554 2611
rect 508 2539 514 2573
rect 548 2539 554 2573
rect 508 2501 554 2539
rect 508 2467 514 2501
rect 548 2467 554 2501
rect 508 2429 554 2467
rect 508 2395 514 2429
rect 548 2395 554 2429
rect 508 2357 554 2395
rect 508 2323 514 2357
rect 548 2323 554 2357
rect 508 2285 554 2323
rect 508 2251 514 2285
rect 548 2251 554 2285
rect 508 2213 554 2251
rect 508 2179 514 2213
rect 548 2179 554 2213
rect 508 2141 554 2179
rect 508 2107 514 2141
rect 548 2107 554 2141
rect 508 2069 554 2107
rect 508 2035 514 2069
rect 548 2035 554 2069
rect 508 1997 554 2035
rect 508 1963 514 1997
rect 548 1963 554 1997
rect 508 1925 554 1963
rect 508 1891 514 1925
rect 548 1891 554 1925
rect 508 1853 554 1891
rect 508 1819 514 1853
rect 548 1819 554 1853
rect 508 1781 554 1819
rect 508 1747 514 1781
rect 548 1747 554 1781
rect 508 1709 554 1747
rect 508 1675 514 1709
rect 548 1675 554 1709
rect 508 1637 554 1675
rect 508 1603 514 1637
rect 548 1603 554 1637
rect 508 1565 554 1603
rect 508 1531 514 1565
rect 548 1531 554 1565
rect 508 1493 554 1531
rect 508 1459 514 1493
rect 548 1459 554 1493
rect 508 1421 554 1459
rect 508 1387 514 1421
rect 548 1387 554 1421
rect 508 1349 554 1387
rect 508 1315 514 1349
rect 548 1315 554 1349
rect 508 1277 554 1315
rect 508 1243 514 1277
rect 548 1243 554 1277
rect 508 1205 554 1243
rect 508 1171 514 1205
rect 548 1171 554 1205
rect 508 1133 554 1171
rect 508 1099 514 1133
rect 548 1099 554 1133
rect 508 1061 554 1099
rect 508 1027 514 1061
rect 548 1027 554 1061
rect 508 989 554 1027
rect 508 955 514 989
rect 548 955 554 989
rect 508 917 554 955
rect 508 883 514 917
rect 548 883 554 917
rect 508 845 554 883
rect 508 811 514 845
rect 548 811 554 845
rect 508 773 554 811
rect 508 739 514 773
rect 548 739 554 773
rect 508 701 554 739
rect 508 667 514 701
rect 548 667 554 701
rect 508 629 554 667
rect 508 595 514 629
rect 548 595 554 629
rect 508 557 554 595
rect 508 523 514 557
rect 548 523 554 557
rect 508 485 554 523
rect 508 451 514 485
rect 548 451 554 485
rect 508 413 554 451
rect 508 379 514 413
rect 548 379 554 413
rect 508 341 554 379
rect 508 307 514 341
rect 548 307 554 341
rect 508 269 554 307
rect 508 235 514 269
rect 548 235 554 269
rect 508 197 554 235
rect 508 163 514 197
rect 548 163 554 197
rect 508 125 554 163
rect 508 91 514 125
rect 548 91 554 125
rect 508 53 554 91
rect 508 19 514 53
rect 548 19 554 53
rect 508 -19 554 19
rect 508 -53 514 -19
rect 548 -53 554 -19
rect 508 -91 554 -53
rect 508 -125 514 -91
rect 548 -125 554 -91
rect 508 -163 554 -125
rect 508 -197 514 -163
rect 548 -197 554 -163
rect 508 -235 554 -197
rect 508 -269 514 -235
rect 548 -269 554 -235
rect 508 -307 554 -269
rect 508 -341 514 -307
rect 548 -341 554 -307
rect 508 -379 554 -341
rect 508 -413 514 -379
rect 548 -413 554 -379
rect 508 -451 554 -413
rect 508 -485 514 -451
rect 548 -485 554 -451
rect 508 -523 554 -485
rect 508 -557 514 -523
rect 548 -557 554 -523
rect 508 -595 554 -557
rect 508 -629 514 -595
rect 548 -629 554 -595
rect 508 -667 554 -629
rect 508 -701 514 -667
rect 548 -701 554 -667
rect 508 -739 554 -701
rect 508 -773 514 -739
rect 548 -773 554 -739
rect 508 -811 554 -773
rect 508 -845 514 -811
rect 548 -845 554 -811
rect 508 -883 554 -845
rect 508 -917 514 -883
rect 548 -917 554 -883
rect 508 -955 554 -917
rect 508 -989 514 -955
rect 548 -989 554 -955
rect 508 -1027 554 -989
rect 508 -1061 514 -1027
rect 548 -1061 554 -1027
rect 508 -1099 554 -1061
rect 508 -1133 514 -1099
rect 548 -1133 554 -1099
rect 508 -1171 554 -1133
rect 508 -1205 514 -1171
rect 548 -1205 554 -1171
rect 508 -1243 554 -1205
rect 508 -1277 514 -1243
rect 548 -1277 554 -1243
rect 508 -1315 554 -1277
rect 508 -1349 514 -1315
rect 548 -1349 554 -1315
rect 508 -1387 554 -1349
rect 508 -1421 514 -1387
rect 548 -1421 554 -1387
rect 508 -1459 554 -1421
rect 508 -1493 514 -1459
rect 548 -1493 554 -1459
rect 508 -1531 554 -1493
rect 508 -1565 514 -1531
rect 548 -1565 554 -1531
rect 508 -1603 554 -1565
rect 508 -1637 514 -1603
rect 548 -1637 554 -1603
rect 508 -1675 554 -1637
rect 508 -1709 514 -1675
rect 548 -1709 554 -1675
rect 508 -1747 554 -1709
rect 508 -1781 514 -1747
rect 548 -1781 554 -1747
rect 508 -1819 554 -1781
rect 508 -1853 514 -1819
rect 548 -1853 554 -1819
rect 508 -1891 554 -1853
rect 508 -1925 514 -1891
rect 548 -1925 554 -1891
rect 508 -1963 554 -1925
rect 508 -1997 514 -1963
rect 548 -1997 554 -1963
rect 508 -2035 554 -1997
rect 508 -2069 514 -2035
rect 548 -2069 554 -2035
rect 508 -2107 554 -2069
rect 508 -2141 514 -2107
rect 548 -2141 554 -2107
rect 508 -2179 554 -2141
rect 508 -2213 514 -2179
rect 548 -2213 554 -2179
rect 508 -2251 554 -2213
rect 508 -2285 514 -2251
rect 548 -2285 554 -2251
rect 508 -2323 554 -2285
rect 508 -2357 514 -2323
rect 548 -2357 554 -2323
rect 508 -2395 554 -2357
rect 508 -2429 514 -2395
rect 548 -2429 554 -2395
rect 508 -2467 554 -2429
rect 508 -2501 514 -2467
rect 548 -2501 554 -2467
rect 508 -2539 554 -2501
rect 508 -2573 514 -2539
rect 548 -2573 554 -2539
rect 508 -2611 554 -2573
rect 508 -2645 514 -2611
rect 548 -2645 554 -2611
rect 508 -2683 554 -2645
rect 508 -2717 514 -2683
rect 548 -2717 554 -2683
rect 508 -2755 554 -2717
rect 508 -2789 514 -2755
rect 548 -2789 554 -2755
rect 508 -2827 554 -2789
rect 508 -2861 514 -2827
rect 548 -2861 554 -2827
rect 508 -2899 554 -2861
rect 508 -2933 514 -2899
rect 548 -2933 554 -2899
rect 508 -2971 554 -2933
rect 508 -3005 514 -2971
rect 548 -3005 554 -2971
rect 508 -3043 554 -3005
rect 508 -3077 514 -3043
rect 548 -3077 554 -3043
rect 508 -3115 554 -3077
rect 508 -3149 514 -3115
rect 548 -3149 554 -3115
rect 508 -3187 554 -3149
rect 508 -3221 514 -3187
rect 548 -3221 554 -3187
rect 508 -3259 554 -3221
rect 508 -3293 514 -3259
rect 548 -3293 554 -3259
rect 508 -3331 554 -3293
rect 508 -3365 514 -3331
rect 548 -3365 554 -3331
rect 508 -3403 554 -3365
rect 508 -3437 514 -3403
rect 548 -3437 554 -3403
rect 508 -3475 554 -3437
rect 508 -3509 514 -3475
rect 548 -3509 554 -3475
rect 508 -3547 554 -3509
rect 508 -3581 514 -3547
rect 548 -3581 554 -3547
rect 508 -3619 554 -3581
rect 508 -3653 514 -3619
rect 548 -3653 554 -3619
rect 508 -3691 554 -3653
rect 508 -3725 514 -3691
rect 548 -3725 554 -3691
rect 508 -3763 554 -3725
rect 508 -3797 514 -3763
rect 548 -3797 554 -3763
rect 508 -3835 554 -3797
rect 508 -3869 514 -3835
rect 548 -3869 554 -3835
rect 508 -3907 554 -3869
rect 508 -3941 514 -3907
rect 548 -3941 554 -3907
rect 508 -3979 554 -3941
rect 508 -4013 514 -3979
rect 548 -4013 554 -3979
rect 508 -4051 554 -4013
rect 508 -4085 514 -4051
rect 548 -4085 554 -4051
rect 508 -4123 554 -4085
rect 508 -4157 514 -4123
rect 548 -4157 554 -4123
rect 508 -4195 554 -4157
rect 508 -4229 514 -4195
rect 548 -4229 554 -4195
rect 508 -4267 554 -4229
rect 508 -4301 514 -4267
rect 548 -4301 554 -4267
rect 508 -4339 554 -4301
rect 508 -4373 514 -4339
rect 548 -4373 554 -4339
rect 508 -4411 554 -4373
rect 508 -4445 514 -4411
rect 548 -4445 554 -4411
rect 508 -4483 554 -4445
rect 508 -4517 514 -4483
rect 548 -4517 554 -4483
rect 508 -4555 554 -4517
rect 508 -4589 514 -4555
rect 548 -4589 554 -4555
rect 508 -4627 554 -4589
rect 508 -4661 514 -4627
rect 548 -4661 554 -4627
rect 508 -4699 554 -4661
rect 508 -4733 514 -4699
rect 548 -4733 554 -4699
rect 508 -4771 554 -4733
rect 508 -4805 514 -4771
rect 548 -4805 554 -4771
rect 508 -4843 554 -4805
rect 508 -4877 514 -4843
rect 548 -4877 554 -4843
rect 508 -4915 554 -4877
rect 508 -4949 514 -4915
rect 548 -4949 554 -4915
rect 508 -4987 554 -4949
rect 508 -5021 514 -4987
rect 548 -5021 554 -4987
rect 508 -5059 554 -5021
rect 508 -5093 514 -5059
rect 548 -5093 554 -5059
rect 508 -5131 554 -5093
rect 508 -5165 514 -5131
rect 548 -5165 554 -5131
rect 508 -5203 554 -5165
rect 508 -5237 514 -5203
rect 548 -5237 554 -5203
rect 508 -5275 554 -5237
rect 508 -5309 514 -5275
rect 548 -5309 554 -5275
rect 508 -5347 554 -5309
rect 508 -5381 514 -5347
rect 548 -5381 554 -5347
rect 508 -5419 554 -5381
rect 508 -5453 514 -5419
rect 548 -5453 554 -5419
rect 508 -5491 554 -5453
rect 508 -5525 514 -5491
rect 548 -5525 554 -5491
rect 508 -5563 554 -5525
rect 508 -5597 514 -5563
rect 548 -5597 554 -5563
rect 508 -5635 554 -5597
rect 508 -5669 514 -5635
rect 548 -5669 554 -5635
rect 508 -5707 554 -5669
rect 508 -5741 514 -5707
rect 548 -5741 554 -5707
rect 508 -5779 554 -5741
rect 508 -5813 514 -5779
rect 548 -5813 554 -5779
rect 508 -5851 554 -5813
rect 508 -5885 514 -5851
rect 548 -5885 554 -5851
rect 508 -5923 554 -5885
rect 508 -5957 514 -5923
rect 548 -5957 554 -5923
rect 508 -5995 554 -5957
rect 508 -6029 514 -5995
rect 548 -6029 554 -5995
rect 508 -6067 554 -6029
rect 508 -6101 514 -6067
rect 548 -6101 554 -6067
rect 508 -6139 554 -6101
rect 508 -6173 514 -6139
rect 548 -6173 554 -6139
rect 508 -6211 554 -6173
rect 508 -6245 514 -6211
rect 548 -6245 554 -6211
rect 508 -6283 554 -6245
rect 508 -6317 514 -6283
rect 548 -6317 554 -6283
rect 508 -6355 554 -6317
rect 508 -6389 514 -6355
rect 548 -6389 554 -6355
rect 508 -6427 554 -6389
rect 508 -6461 514 -6427
rect 548 -6461 554 -6427
rect 508 -6499 554 -6461
rect 508 -6533 514 -6499
rect 548 -6533 554 -6499
rect 508 -6571 554 -6533
rect 508 -6605 514 -6571
rect 548 -6605 554 -6571
rect 508 -6643 554 -6605
rect 508 -6677 514 -6643
rect 548 -6677 554 -6643
rect 508 -6715 554 -6677
rect 508 -6749 514 -6715
rect 548 -6749 554 -6715
rect 508 -6787 554 -6749
rect 508 -6821 514 -6787
rect 548 -6821 554 -6787
rect 508 -6859 554 -6821
rect 508 -6893 514 -6859
rect 548 -6893 554 -6859
rect 508 -6931 554 -6893
rect 508 -6965 514 -6931
rect 548 -6965 554 -6931
rect 508 -7003 554 -6965
rect 508 -7037 514 -7003
rect 548 -7037 554 -7003
rect 508 -7075 554 -7037
rect 508 -7109 514 -7075
rect 548 -7109 554 -7075
rect 508 -7147 554 -7109
rect 508 -7181 514 -7147
rect 548 -7181 554 -7147
rect 508 -7219 554 -7181
rect 508 -7253 514 -7219
rect 548 -7253 554 -7219
rect 508 -7291 554 -7253
rect 508 -7325 514 -7291
rect 548 -7325 554 -7291
rect 508 -7363 554 -7325
rect 508 -7397 514 -7363
rect 548 -7397 554 -7363
rect 508 -7435 554 -7397
rect 508 -7469 514 -7435
rect 548 -7469 554 -7435
rect 508 -7507 554 -7469
rect 508 -7541 514 -7507
rect 548 -7541 554 -7507
rect 508 -7579 554 -7541
rect 508 -7613 514 -7579
rect 548 -7613 554 -7579
rect 508 -7651 554 -7613
rect 508 -7685 514 -7651
rect 548 -7685 554 -7651
rect 508 -7723 554 -7685
rect 508 -7757 514 -7723
rect 548 -7757 554 -7723
rect 508 -7795 554 -7757
rect 508 -7829 514 -7795
rect 548 -7829 554 -7795
rect 508 -7867 554 -7829
rect 508 -7901 514 -7867
rect 548 -7901 554 -7867
rect 508 -7939 554 -7901
rect 508 -7973 514 -7939
rect 548 -7973 554 -7939
rect 508 -8011 554 -7973
rect 508 -8045 514 -8011
rect 548 -8045 554 -8011
rect 508 -8083 554 -8045
rect 508 -8117 514 -8083
rect 548 -8117 554 -8083
rect 508 -8155 554 -8117
rect 508 -8189 514 -8155
rect 548 -8189 554 -8155
rect 508 -8227 554 -8189
rect 508 -8261 514 -8227
rect 548 -8261 554 -8227
rect 508 -8299 554 -8261
rect 508 -8333 514 -8299
rect 548 -8333 554 -8299
rect 508 -8371 554 -8333
rect 508 -8405 514 -8371
rect 548 -8405 554 -8371
rect 508 -8443 554 -8405
rect 508 -8477 514 -8443
rect 548 -8477 554 -8443
rect 508 -8515 554 -8477
rect 508 -8549 514 -8515
rect 548 -8549 554 -8515
rect 508 -8587 554 -8549
rect 508 -8621 514 -8587
rect 548 -8621 554 -8587
rect 508 -8659 554 -8621
rect 508 -8693 514 -8659
rect 548 -8693 554 -8659
rect 508 -8731 554 -8693
rect 508 -8765 514 -8731
rect 548 -8765 554 -8731
rect 508 -8803 554 -8765
rect 508 -8837 514 -8803
rect 548 -8837 554 -8803
rect 508 -8875 554 -8837
rect 508 -8909 514 -8875
rect 548 -8909 554 -8875
rect 508 -8947 554 -8909
rect 508 -8981 514 -8947
rect 548 -8981 554 -8947
rect 508 -9019 554 -8981
rect 508 -9053 514 -9019
rect 548 -9053 554 -9019
rect 508 -9091 554 -9053
rect 508 -9125 514 -9091
rect 548 -9125 554 -9091
rect 508 -9163 554 -9125
rect 508 -9197 514 -9163
rect 548 -9197 554 -9163
rect 508 -9235 554 -9197
rect 508 -9269 514 -9235
rect 548 -9269 554 -9235
rect 508 -9307 554 -9269
rect 508 -9341 514 -9307
rect 548 -9341 554 -9307
rect 508 -9379 554 -9341
rect 508 -9413 514 -9379
rect 548 -9413 554 -9379
rect 508 -9451 554 -9413
rect 508 -9485 514 -9451
rect 548 -9485 554 -9451
rect 508 -9523 554 -9485
rect 508 -9557 514 -9523
rect 548 -9557 554 -9523
rect 508 -9600 554 -9557
rect 626 9557 672 9600
rect 626 9523 632 9557
rect 666 9523 672 9557
rect 626 9485 672 9523
rect 626 9451 632 9485
rect 666 9451 672 9485
rect 626 9413 672 9451
rect 626 9379 632 9413
rect 666 9379 672 9413
rect 626 9341 672 9379
rect 626 9307 632 9341
rect 666 9307 672 9341
rect 626 9269 672 9307
rect 626 9235 632 9269
rect 666 9235 672 9269
rect 626 9197 672 9235
rect 626 9163 632 9197
rect 666 9163 672 9197
rect 626 9125 672 9163
rect 626 9091 632 9125
rect 666 9091 672 9125
rect 626 9053 672 9091
rect 626 9019 632 9053
rect 666 9019 672 9053
rect 626 8981 672 9019
rect 626 8947 632 8981
rect 666 8947 672 8981
rect 626 8909 672 8947
rect 626 8875 632 8909
rect 666 8875 672 8909
rect 626 8837 672 8875
rect 626 8803 632 8837
rect 666 8803 672 8837
rect 626 8765 672 8803
rect 626 8731 632 8765
rect 666 8731 672 8765
rect 626 8693 672 8731
rect 626 8659 632 8693
rect 666 8659 672 8693
rect 626 8621 672 8659
rect 626 8587 632 8621
rect 666 8587 672 8621
rect 626 8549 672 8587
rect 626 8515 632 8549
rect 666 8515 672 8549
rect 626 8477 672 8515
rect 626 8443 632 8477
rect 666 8443 672 8477
rect 626 8405 672 8443
rect 626 8371 632 8405
rect 666 8371 672 8405
rect 626 8333 672 8371
rect 626 8299 632 8333
rect 666 8299 672 8333
rect 626 8261 672 8299
rect 626 8227 632 8261
rect 666 8227 672 8261
rect 626 8189 672 8227
rect 626 8155 632 8189
rect 666 8155 672 8189
rect 626 8117 672 8155
rect 626 8083 632 8117
rect 666 8083 672 8117
rect 626 8045 672 8083
rect 626 8011 632 8045
rect 666 8011 672 8045
rect 626 7973 672 8011
rect 626 7939 632 7973
rect 666 7939 672 7973
rect 626 7901 672 7939
rect 626 7867 632 7901
rect 666 7867 672 7901
rect 626 7829 672 7867
rect 626 7795 632 7829
rect 666 7795 672 7829
rect 626 7757 672 7795
rect 626 7723 632 7757
rect 666 7723 672 7757
rect 626 7685 672 7723
rect 626 7651 632 7685
rect 666 7651 672 7685
rect 626 7613 672 7651
rect 626 7579 632 7613
rect 666 7579 672 7613
rect 626 7541 672 7579
rect 626 7507 632 7541
rect 666 7507 672 7541
rect 626 7469 672 7507
rect 626 7435 632 7469
rect 666 7435 672 7469
rect 626 7397 672 7435
rect 626 7363 632 7397
rect 666 7363 672 7397
rect 626 7325 672 7363
rect 626 7291 632 7325
rect 666 7291 672 7325
rect 626 7253 672 7291
rect 626 7219 632 7253
rect 666 7219 672 7253
rect 626 7181 672 7219
rect 626 7147 632 7181
rect 666 7147 672 7181
rect 626 7109 672 7147
rect 626 7075 632 7109
rect 666 7075 672 7109
rect 626 7037 672 7075
rect 626 7003 632 7037
rect 666 7003 672 7037
rect 626 6965 672 7003
rect 626 6931 632 6965
rect 666 6931 672 6965
rect 626 6893 672 6931
rect 626 6859 632 6893
rect 666 6859 672 6893
rect 626 6821 672 6859
rect 626 6787 632 6821
rect 666 6787 672 6821
rect 626 6749 672 6787
rect 626 6715 632 6749
rect 666 6715 672 6749
rect 626 6677 672 6715
rect 626 6643 632 6677
rect 666 6643 672 6677
rect 626 6605 672 6643
rect 626 6571 632 6605
rect 666 6571 672 6605
rect 626 6533 672 6571
rect 626 6499 632 6533
rect 666 6499 672 6533
rect 626 6461 672 6499
rect 626 6427 632 6461
rect 666 6427 672 6461
rect 626 6389 672 6427
rect 626 6355 632 6389
rect 666 6355 672 6389
rect 626 6317 672 6355
rect 626 6283 632 6317
rect 666 6283 672 6317
rect 626 6245 672 6283
rect 626 6211 632 6245
rect 666 6211 672 6245
rect 626 6173 672 6211
rect 626 6139 632 6173
rect 666 6139 672 6173
rect 626 6101 672 6139
rect 626 6067 632 6101
rect 666 6067 672 6101
rect 626 6029 672 6067
rect 626 5995 632 6029
rect 666 5995 672 6029
rect 626 5957 672 5995
rect 626 5923 632 5957
rect 666 5923 672 5957
rect 626 5885 672 5923
rect 626 5851 632 5885
rect 666 5851 672 5885
rect 626 5813 672 5851
rect 626 5779 632 5813
rect 666 5779 672 5813
rect 626 5741 672 5779
rect 626 5707 632 5741
rect 666 5707 672 5741
rect 626 5669 672 5707
rect 626 5635 632 5669
rect 666 5635 672 5669
rect 626 5597 672 5635
rect 626 5563 632 5597
rect 666 5563 672 5597
rect 626 5525 672 5563
rect 626 5491 632 5525
rect 666 5491 672 5525
rect 626 5453 672 5491
rect 626 5419 632 5453
rect 666 5419 672 5453
rect 626 5381 672 5419
rect 626 5347 632 5381
rect 666 5347 672 5381
rect 626 5309 672 5347
rect 626 5275 632 5309
rect 666 5275 672 5309
rect 626 5237 672 5275
rect 626 5203 632 5237
rect 666 5203 672 5237
rect 626 5165 672 5203
rect 626 5131 632 5165
rect 666 5131 672 5165
rect 626 5093 672 5131
rect 626 5059 632 5093
rect 666 5059 672 5093
rect 626 5021 672 5059
rect 626 4987 632 5021
rect 666 4987 672 5021
rect 626 4949 672 4987
rect 626 4915 632 4949
rect 666 4915 672 4949
rect 626 4877 672 4915
rect 626 4843 632 4877
rect 666 4843 672 4877
rect 626 4805 672 4843
rect 626 4771 632 4805
rect 666 4771 672 4805
rect 626 4733 672 4771
rect 626 4699 632 4733
rect 666 4699 672 4733
rect 626 4661 672 4699
rect 626 4627 632 4661
rect 666 4627 672 4661
rect 626 4589 672 4627
rect 626 4555 632 4589
rect 666 4555 672 4589
rect 626 4517 672 4555
rect 626 4483 632 4517
rect 666 4483 672 4517
rect 626 4445 672 4483
rect 626 4411 632 4445
rect 666 4411 672 4445
rect 626 4373 672 4411
rect 626 4339 632 4373
rect 666 4339 672 4373
rect 626 4301 672 4339
rect 626 4267 632 4301
rect 666 4267 672 4301
rect 626 4229 672 4267
rect 626 4195 632 4229
rect 666 4195 672 4229
rect 626 4157 672 4195
rect 626 4123 632 4157
rect 666 4123 672 4157
rect 626 4085 672 4123
rect 626 4051 632 4085
rect 666 4051 672 4085
rect 626 4013 672 4051
rect 626 3979 632 4013
rect 666 3979 672 4013
rect 626 3941 672 3979
rect 626 3907 632 3941
rect 666 3907 672 3941
rect 626 3869 672 3907
rect 626 3835 632 3869
rect 666 3835 672 3869
rect 626 3797 672 3835
rect 626 3763 632 3797
rect 666 3763 672 3797
rect 626 3725 672 3763
rect 626 3691 632 3725
rect 666 3691 672 3725
rect 626 3653 672 3691
rect 626 3619 632 3653
rect 666 3619 672 3653
rect 626 3581 672 3619
rect 626 3547 632 3581
rect 666 3547 672 3581
rect 626 3509 672 3547
rect 626 3475 632 3509
rect 666 3475 672 3509
rect 626 3437 672 3475
rect 626 3403 632 3437
rect 666 3403 672 3437
rect 626 3365 672 3403
rect 626 3331 632 3365
rect 666 3331 672 3365
rect 626 3293 672 3331
rect 626 3259 632 3293
rect 666 3259 672 3293
rect 626 3221 672 3259
rect 626 3187 632 3221
rect 666 3187 672 3221
rect 626 3149 672 3187
rect 626 3115 632 3149
rect 666 3115 672 3149
rect 626 3077 672 3115
rect 626 3043 632 3077
rect 666 3043 672 3077
rect 626 3005 672 3043
rect 626 2971 632 3005
rect 666 2971 672 3005
rect 626 2933 672 2971
rect 626 2899 632 2933
rect 666 2899 672 2933
rect 626 2861 672 2899
rect 626 2827 632 2861
rect 666 2827 672 2861
rect 626 2789 672 2827
rect 626 2755 632 2789
rect 666 2755 672 2789
rect 626 2717 672 2755
rect 626 2683 632 2717
rect 666 2683 672 2717
rect 626 2645 672 2683
rect 626 2611 632 2645
rect 666 2611 672 2645
rect 626 2573 672 2611
rect 626 2539 632 2573
rect 666 2539 672 2573
rect 626 2501 672 2539
rect 626 2467 632 2501
rect 666 2467 672 2501
rect 626 2429 672 2467
rect 626 2395 632 2429
rect 666 2395 672 2429
rect 626 2357 672 2395
rect 626 2323 632 2357
rect 666 2323 672 2357
rect 626 2285 672 2323
rect 626 2251 632 2285
rect 666 2251 672 2285
rect 626 2213 672 2251
rect 626 2179 632 2213
rect 666 2179 672 2213
rect 626 2141 672 2179
rect 626 2107 632 2141
rect 666 2107 672 2141
rect 626 2069 672 2107
rect 626 2035 632 2069
rect 666 2035 672 2069
rect 626 1997 672 2035
rect 626 1963 632 1997
rect 666 1963 672 1997
rect 626 1925 672 1963
rect 626 1891 632 1925
rect 666 1891 672 1925
rect 626 1853 672 1891
rect 626 1819 632 1853
rect 666 1819 672 1853
rect 626 1781 672 1819
rect 626 1747 632 1781
rect 666 1747 672 1781
rect 626 1709 672 1747
rect 626 1675 632 1709
rect 666 1675 672 1709
rect 626 1637 672 1675
rect 626 1603 632 1637
rect 666 1603 672 1637
rect 626 1565 672 1603
rect 626 1531 632 1565
rect 666 1531 672 1565
rect 626 1493 672 1531
rect 626 1459 632 1493
rect 666 1459 672 1493
rect 626 1421 672 1459
rect 626 1387 632 1421
rect 666 1387 672 1421
rect 626 1349 672 1387
rect 626 1315 632 1349
rect 666 1315 672 1349
rect 626 1277 672 1315
rect 626 1243 632 1277
rect 666 1243 672 1277
rect 626 1205 672 1243
rect 626 1171 632 1205
rect 666 1171 672 1205
rect 626 1133 672 1171
rect 626 1099 632 1133
rect 666 1099 672 1133
rect 626 1061 672 1099
rect 626 1027 632 1061
rect 666 1027 672 1061
rect 626 989 672 1027
rect 626 955 632 989
rect 666 955 672 989
rect 626 917 672 955
rect 626 883 632 917
rect 666 883 672 917
rect 626 845 672 883
rect 626 811 632 845
rect 666 811 672 845
rect 626 773 672 811
rect 626 739 632 773
rect 666 739 672 773
rect 626 701 672 739
rect 626 667 632 701
rect 666 667 672 701
rect 626 629 672 667
rect 626 595 632 629
rect 666 595 672 629
rect 626 557 672 595
rect 626 523 632 557
rect 666 523 672 557
rect 626 485 672 523
rect 626 451 632 485
rect 666 451 672 485
rect 626 413 672 451
rect 626 379 632 413
rect 666 379 672 413
rect 626 341 672 379
rect 626 307 632 341
rect 666 307 672 341
rect 626 269 672 307
rect 626 235 632 269
rect 666 235 672 269
rect 626 197 672 235
rect 626 163 632 197
rect 666 163 672 197
rect 626 125 672 163
rect 626 91 632 125
rect 666 91 672 125
rect 626 53 672 91
rect 626 19 632 53
rect 666 19 672 53
rect 626 -19 672 19
rect 626 -53 632 -19
rect 666 -53 672 -19
rect 626 -91 672 -53
rect 626 -125 632 -91
rect 666 -125 672 -91
rect 626 -163 672 -125
rect 626 -197 632 -163
rect 666 -197 672 -163
rect 626 -235 672 -197
rect 626 -269 632 -235
rect 666 -269 672 -235
rect 626 -307 672 -269
rect 626 -341 632 -307
rect 666 -341 672 -307
rect 626 -379 672 -341
rect 626 -413 632 -379
rect 666 -413 672 -379
rect 626 -451 672 -413
rect 626 -485 632 -451
rect 666 -485 672 -451
rect 626 -523 672 -485
rect 626 -557 632 -523
rect 666 -557 672 -523
rect 626 -595 672 -557
rect 626 -629 632 -595
rect 666 -629 672 -595
rect 626 -667 672 -629
rect 626 -701 632 -667
rect 666 -701 672 -667
rect 626 -739 672 -701
rect 626 -773 632 -739
rect 666 -773 672 -739
rect 626 -811 672 -773
rect 626 -845 632 -811
rect 666 -845 672 -811
rect 626 -883 672 -845
rect 626 -917 632 -883
rect 666 -917 672 -883
rect 626 -955 672 -917
rect 626 -989 632 -955
rect 666 -989 672 -955
rect 626 -1027 672 -989
rect 626 -1061 632 -1027
rect 666 -1061 672 -1027
rect 626 -1099 672 -1061
rect 626 -1133 632 -1099
rect 666 -1133 672 -1099
rect 626 -1171 672 -1133
rect 626 -1205 632 -1171
rect 666 -1205 672 -1171
rect 626 -1243 672 -1205
rect 626 -1277 632 -1243
rect 666 -1277 672 -1243
rect 626 -1315 672 -1277
rect 626 -1349 632 -1315
rect 666 -1349 672 -1315
rect 626 -1387 672 -1349
rect 626 -1421 632 -1387
rect 666 -1421 672 -1387
rect 626 -1459 672 -1421
rect 626 -1493 632 -1459
rect 666 -1493 672 -1459
rect 626 -1531 672 -1493
rect 626 -1565 632 -1531
rect 666 -1565 672 -1531
rect 626 -1603 672 -1565
rect 626 -1637 632 -1603
rect 666 -1637 672 -1603
rect 626 -1675 672 -1637
rect 626 -1709 632 -1675
rect 666 -1709 672 -1675
rect 626 -1747 672 -1709
rect 626 -1781 632 -1747
rect 666 -1781 672 -1747
rect 626 -1819 672 -1781
rect 626 -1853 632 -1819
rect 666 -1853 672 -1819
rect 626 -1891 672 -1853
rect 626 -1925 632 -1891
rect 666 -1925 672 -1891
rect 626 -1963 672 -1925
rect 626 -1997 632 -1963
rect 666 -1997 672 -1963
rect 626 -2035 672 -1997
rect 626 -2069 632 -2035
rect 666 -2069 672 -2035
rect 626 -2107 672 -2069
rect 626 -2141 632 -2107
rect 666 -2141 672 -2107
rect 626 -2179 672 -2141
rect 626 -2213 632 -2179
rect 666 -2213 672 -2179
rect 626 -2251 672 -2213
rect 626 -2285 632 -2251
rect 666 -2285 672 -2251
rect 626 -2323 672 -2285
rect 626 -2357 632 -2323
rect 666 -2357 672 -2323
rect 626 -2395 672 -2357
rect 626 -2429 632 -2395
rect 666 -2429 672 -2395
rect 626 -2467 672 -2429
rect 626 -2501 632 -2467
rect 666 -2501 672 -2467
rect 626 -2539 672 -2501
rect 626 -2573 632 -2539
rect 666 -2573 672 -2539
rect 626 -2611 672 -2573
rect 626 -2645 632 -2611
rect 666 -2645 672 -2611
rect 626 -2683 672 -2645
rect 626 -2717 632 -2683
rect 666 -2717 672 -2683
rect 626 -2755 672 -2717
rect 626 -2789 632 -2755
rect 666 -2789 672 -2755
rect 626 -2827 672 -2789
rect 626 -2861 632 -2827
rect 666 -2861 672 -2827
rect 626 -2899 672 -2861
rect 626 -2933 632 -2899
rect 666 -2933 672 -2899
rect 626 -2971 672 -2933
rect 626 -3005 632 -2971
rect 666 -3005 672 -2971
rect 626 -3043 672 -3005
rect 626 -3077 632 -3043
rect 666 -3077 672 -3043
rect 626 -3115 672 -3077
rect 626 -3149 632 -3115
rect 666 -3149 672 -3115
rect 626 -3187 672 -3149
rect 626 -3221 632 -3187
rect 666 -3221 672 -3187
rect 626 -3259 672 -3221
rect 626 -3293 632 -3259
rect 666 -3293 672 -3259
rect 626 -3331 672 -3293
rect 626 -3365 632 -3331
rect 666 -3365 672 -3331
rect 626 -3403 672 -3365
rect 626 -3437 632 -3403
rect 666 -3437 672 -3403
rect 626 -3475 672 -3437
rect 626 -3509 632 -3475
rect 666 -3509 672 -3475
rect 626 -3547 672 -3509
rect 626 -3581 632 -3547
rect 666 -3581 672 -3547
rect 626 -3619 672 -3581
rect 626 -3653 632 -3619
rect 666 -3653 672 -3619
rect 626 -3691 672 -3653
rect 626 -3725 632 -3691
rect 666 -3725 672 -3691
rect 626 -3763 672 -3725
rect 626 -3797 632 -3763
rect 666 -3797 672 -3763
rect 626 -3835 672 -3797
rect 626 -3869 632 -3835
rect 666 -3869 672 -3835
rect 626 -3907 672 -3869
rect 626 -3941 632 -3907
rect 666 -3941 672 -3907
rect 626 -3979 672 -3941
rect 626 -4013 632 -3979
rect 666 -4013 672 -3979
rect 626 -4051 672 -4013
rect 626 -4085 632 -4051
rect 666 -4085 672 -4051
rect 626 -4123 672 -4085
rect 626 -4157 632 -4123
rect 666 -4157 672 -4123
rect 626 -4195 672 -4157
rect 626 -4229 632 -4195
rect 666 -4229 672 -4195
rect 626 -4267 672 -4229
rect 626 -4301 632 -4267
rect 666 -4301 672 -4267
rect 626 -4339 672 -4301
rect 626 -4373 632 -4339
rect 666 -4373 672 -4339
rect 626 -4411 672 -4373
rect 626 -4445 632 -4411
rect 666 -4445 672 -4411
rect 626 -4483 672 -4445
rect 626 -4517 632 -4483
rect 666 -4517 672 -4483
rect 626 -4555 672 -4517
rect 626 -4589 632 -4555
rect 666 -4589 672 -4555
rect 626 -4627 672 -4589
rect 626 -4661 632 -4627
rect 666 -4661 672 -4627
rect 626 -4699 672 -4661
rect 626 -4733 632 -4699
rect 666 -4733 672 -4699
rect 626 -4771 672 -4733
rect 626 -4805 632 -4771
rect 666 -4805 672 -4771
rect 626 -4843 672 -4805
rect 626 -4877 632 -4843
rect 666 -4877 672 -4843
rect 626 -4915 672 -4877
rect 626 -4949 632 -4915
rect 666 -4949 672 -4915
rect 626 -4987 672 -4949
rect 626 -5021 632 -4987
rect 666 -5021 672 -4987
rect 626 -5059 672 -5021
rect 626 -5093 632 -5059
rect 666 -5093 672 -5059
rect 626 -5131 672 -5093
rect 626 -5165 632 -5131
rect 666 -5165 672 -5131
rect 626 -5203 672 -5165
rect 626 -5237 632 -5203
rect 666 -5237 672 -5203
rect 626 -5275 672 -5237
rect 626 -5309 632 -5275
rect 666 -5309 672 -5275
rect 626 -5347 672 -5309
rect 626 -5381 632 -5347
rect 666 -5381 672 -5347
rect 626 -5419 672 -5381
rect 626 -5453 632 -5419
rect 666 -5453 672 -5419
rect 626 -5491 672 -5453
rect 626 -5525 632 -5491
rect 666 -5525 672 -5491
rect 626 -5563 672 -5525
rect 626 -5597 632 -5563
rect 666 -5597 672 -5563
rect 626 -5635 672 -5597
rect 626 -5669 632 -5635
rect 666 -5669 672 -5635
rect 626 -5707 672 -5669
rect 626 -5741 632 -5707
rect 666 -5741 672 -5707
rect 626 -5779 672 -5741
rect 626 -5813 632 -5779
rect 666 -5813 672 -5779
rect 626 -5851 672 -5813
rect 626 -5885 632 -5851
rect 666 -5885 672 -5851
rect 626 -5923 672 -5885
rect 626 -5957 632 -5923
rect 666 -5957 672 -5923
rect 626 -5995 672 -5957
rect 626 -6029 632 -5995
rect 666 -6029 672 -5995
rect 626 -6067 672 -6029
rect 626 -6101 632 -6067
rect 666 -6101 672 -6067
rect 626 -6139 672 -6101
rect 626 -6173 632 -6139
rect 666 -6173 672 -6139
rect 626 -6211 672 -6173
rect 626 -6245 632 -6211
rect 666 -6245 672 -6211
rect 626 -6283 672 -6245
rect 626 -6317 632 -6283
rect 666 -6317 672 -6283
rect 626 -6355 672 -6317
rect 626 -6389 632 -6355
rect 666 -6389 672 -6355
rect 626 -6427 672 -6389
rect 626 -6461 632 -6427
rect 666 -6461 672 -6427
rect 626 -6499 672 -6461
rect 626 -6533 632 -6499
rect 666 -6533 672 -6499
rect 626 -6571 672 -6533
rect 626 -6605 632 -6571
rect 666 -6605 672 -6571
rect 626 -6643 672 -6605
rect 626 -6677 632 -6643
rect 666 -6677 672 -6643
rect 626 -6715 672 -6677
rect 626 -6749 632 -6715
rect 666 -6749 672 -6715
rect 626 -6787 672 -6749
rect 626 -6821 632 -6787
rect 666 -6821 672 -6787
rect 626 -6859 672 -6821
rect 626 -6893 632 -6859
rect 666 -6893 672 -6859
rect 626 -6931 672 -6893
rect 626 -6965 632 -6931
rect 666 -6965 672 -6931
rect 626 -7003 672 -6965
rect 626 -7037 632 -7003
rect 666 -7037 672 -7003
rect 626 -7075 672 -7037
rect 626 -7109 632 -7075
rect 666 -7109 672 -7075
rect 626 -7147 672 -7109
rect 626 -7181 632 -7147
rect 666 -7181 672 -7147
rect 626 -7219 672 -7181
rect 626 -7253 632 -7219
rect 666 -7253 672 -7219
rect 626 -7291 672 -7253
rect 626 -7325 632 -7291
rect 666 -7325 672 -7291
rect 626 -7363 672 -7325
rect 626 -7397 632 -7363
rect 666 -7397 672 -7363
rect 626 -7435 672 -7397
rect 626 -7469 632 -7435
rect 666 -7469 672 -7435
rect 626 -7507 672 -7469
rect 626 -7541 632 -7507
rect 666 -7541 672 -7507
rect 626 -7579 672 -7541
rect 626 -7613 632 -7579
rect 666 -7613 672 -7579
rect 626 -7651 672 -7613
rect 626 -7685 632 -7651
rect 666 -7685 672 -7651
rect 626 -7723 672 -7685
rect 626 -7757 632 -7723
rect 666 -7757 672 -7723
rect 626 -7795 672 -7757
rect 626 -7829 632 -7795
rect 666 -7829 672 -7795
rect 626 -7867 672 -7829
rect 626 -7901 632 -7867
rect 666 -7901 672 -7867
rect 626 -7939 672 -7901
rect 626 -7973 632 -7939
rect 666 -7973 672 -7939
rect 626 -8011 672 -7973
rect 626 -8045 632 -8011
rect 666 -8045 672 -8011
rect 626 -8083 672 -8045
rect 626 -8117 632 -8083
rect 666 -8117 672 -8083
rect 626 -8155 672 -8117
rect 626 -8189 632 -8155
rect 666 -8189 672 -8155
rect 626 -8227 672 -8189
rect 626 -8261 632 -8227
rect 666 -8261 672 -8227
rect 626 -8299 672 -8261
rect 626 -8333 632 -8299
rect 666 -8333 672 -8299
rect 626 -8371 672 -8333
rect 626 -8405 632 -8371
rect 666 -8405 672 -8371
rect 626 -8443 672 -8405
rect 626 -8477 632 -8443
rect 666 -8477 672 -8443
rect 626 -8515 672 -8477
rect 626 -8549 632 -8515
rect 666 -8549 672 -8515
rect 626 -8587 672 -8549
rect 626 -8621 632 -8587
rect 666 -8621 672 -8587
rect 626 -8659 672 -8621
rect 626 -8693 632 -8659
rect 666 -8693 672 -8659
rect 626 -8731 672 -8693
rect 626 -8765 632 -8731
rect 666 -8765 672 -8731
rect 626 -8803 672 -8765
rect 626 -8837 632 -8803
rect 666 -8837 672 -8803
rect 626 -8875 672 -8837
rect 626 -8909 632 -8875
rect 666 -8909 672 -8875
rect 626 -8947 672 -8909
rect 626 -8981 632 -8947
rect 666 -8981 672 -8947
rect 626 -9019 672 -8981
rect 626 -9053 632 -9019
rect 666 -9053 672 -9019
rect 626 -9091 672 -9053
rect 626 -9125 632 -9091
rect 666 -9125 672 -9091
rect 626 -9163 672 -9125
rect 626 -9197 632 -9163
rect 666 -9197 672 -9163
rect 626 -9235 672 -9197
rect 626 -9269 632 -9235
rect 666 -9269 672 -9235
rect 626 -9307 672 -9269
rect 626 -9341 632 -9307
rect 666 -9341 672 -9307
rect 626 -9379 672 -9341
rect 626 -9413 632 -9379
rect 666 -9413 672 -9379
rect 626 -9451 672 -9413
rect 626 -9485 632 -9451
rect 666 -9485 672 -9451
rect 626 -9523 672 -9485
rect 626 -9557 632 -9523
rect 666 -9557 672 -9523
rect 626 -9600 672 -9557
rect 744 9557 790 9600
rect 744 9523 750 9557
rect 784 9523 790 9557
rect 744 9485 790 9523
rect 744 9451 750 9485
rect 784 9451 790 9485
rect 744 9413 790 9451
rect 744 9379 750 9413
rect 784 9379 790 9413
rect 744 9341 790 9379
rect 744 9307 750 9341
rect 784 9307 790 9341
rect 744 9269 790 9307
rect 744 9235 750 9269
rect 784 9235 790 9269
rect 744 9197 790 9235
rect 744 9163 750 9197
rect 784 9163 790 9197
rect 744 9125 790 9163
rect 744 9091 750 9125
rect 784 9091 790 9125
rect 744 9053 790 9091
rect 744 9019 750 9053
rect 784 9019 790 9053
rect 744 8981 790 9019
rect 744 8947 750 8981
rect 784 8947 790 8981
rect 744 8909 790 8947
rect 744 8875 750 8909
rect 784 8875 790 8909
rect 744 8837 790 8875
rect 744 8803 750 8837
rect 784 8803 790 8837
rect 744 8765 790 8803
rect 744 8731 750 8765
rect 784 8731 790 8765
rect 744 8693 790 8731
rect 744 8659 750 8693
rect 784 8659 790 8693
rect 744 8621 790 8659
rect 744 8587 750 8621
rect 784 8587 790 8621
rect 744 8549 790 8587
rect 744 8515 750 8549
rect 784 8515 790 8549
rect 744 8477 790 8515
rect 744 8443 750 8477
rect 784 8443 790 8477
rect 744 8405 790 8443
rect 744 8371 750 8405
rect 784 8371 790 8405
rect 744 8333 790 8371
rect 744 8299 750 8333
rect 784 8299 790 8333
rect 744 8261 790 8299
rect 744 8227 750 8261
rect 784 8227 790 8261
rect 744 8189 790 8227
rect 744 8155 750 8189
rect 784 8155 790 8189
rect 744 8117 790 8155
rect 744 8083 750 8117
rect 784 8083 790 8117
rect 744 8045 790 8083
rect 744 8011 750 8045
rect 784 8011 790 8045
rect 744 7973 790 8011
rect 744 7939 750 7973
rect 784 7939 790 7973
rect 744 7901 790 7939
rect 744 7867 750 7901
rect 784 7867 790 7901
rect 744 7829 790 7867
rect 744 7795 750 7829
rect 784 7795 790 7829
rect 744 7757 790 7795
rect 744 7723 750 7757
rect 784 7723 790 7757
rect 744 7685 790 7723
rect 744 7651 750 7685
rect 784 7651 790 7685
rect 744 7613 790 7651
rect 744 7579 750 7613
rect 784 7579 790 7613
rect 744 7541 790 7579
rect 744 7507 750 7541
rect 784 7507 790 7541
rect 744 7469 790 7507
rect 744 7435 750 7469
rect 784 7435 790 7469
rect 744 7397 790 7435
rect 744 7363 750 7397
rect 784 7363 790 7397
rect 744 7325 790 7363
rect 744 7291 750 7325
rect 784 7291 790 7325
rect 744 7253 790 7291
rect 744 7219 750 7253
rect 784 7219 790 7253
rect 744 7181 790 7219
rect 744 7147 750 7181
rect 784 7147 790 7181
rect 744 7109 790 7147
rect 744 7075 750 7109
rect 784 7075 790 7109
rect 744 7037 790 7075
rect 744 7003 750 7037
rect 784 7003 790 7037
rect 744 6965 790 7003
rect 744 6931 750 6965
rect 784 6931 790 6965
rect 744 6893 790 6931
rect 744 6859 750 6893
rect 784 6859 790 6893
rect 744 6821 790 6859
rect 744 6787 750 6821
rect 784 6787 790 6821
rect 744 6749 790 6787
rect 744 6715 750 6749
rect 784 6715 790 6749
rect 744 6677 790 6715
rect 744 6643 750 6677
rect 784 6643 790 6677
rect 744 6605 790 6643
rect 744 6571 750 6605
rect 784 6571 790 6605
rect 744 6533 790 6571
rect 744 6499 750 6533
rect 784 6499 790 6533
rect 744 6461 790 6499
rect 744 6427 750 6461
rect 784 6427 790 6461
rect 744 6389 790 6427
rect 744 6355 750 6389
rect 784 6355 790 6389
rect 744 6317 790 6355
rect 744 6283 750 6317
rect 784 6283 790 6317
rect 744 6245 790 6283
rect 744 6211 750 6245
rect 784 6211 790 6245
rect 744 6173 790 6211
rect 744 6139 750 6173
rect 784 6139 790 6173
rect 744 6101 790 6139
rect 744 6067 750 6101
rect 784 6067 790 6101
rect 744 6029 790 6067
rect 744 5995 750 6029
rect 784 5995 790 6029
rect 744 5957 790 5995
rect 744 5923 750 5957
rect 784 5923 790 5957
rect 744 5885 790 5923
rect 744 5851 750 5885
rect 784 5851 790 5885
rect 744 5813 790 5851
rect 744 5779 750 5813
rect 784 5779 790 5813
rect 744 5741 790 5779
rect 744 5707 750 5741
rect 784 5707 790 5741
rect 744 5669 790 5707
rect 744 5635 750 5669
rect 784 5635 790 5669
rect 744 5597 790 5635
rect 744 5563 750 5597
rect 784 5563 790 5597
rect 744 5525 790 5563
rect 744 5491 750 5525
rect 784 5491 790 5525
rect 744 5453 790 5491
rect 744 5419 750 5453
rect 784 5419 790 5453
rect 744 5381 790 5419
rect 744 5347 750 5381
rect 784 5347 790 5381
rect 744 5309 790 5347
rect 744 5275 750 5309
rect 784 5275 790 5309
rect 744 5237 790 5275
rect 744 5203 750 5237
rect 784 5203 790 5237
rect 744 5165 790 5203
rect 744 5131 750 5165
rect 784 5131 790 5165
rect 744 5093 790 5131
rect 744 5059 750 5093
rect 784 5059 790 5093
rect 744 5021 790 5059
rect 744 4987 750 5021
rect 784 4987 790 5021
rect 744 4949 790 4987
rect 744 4915 750 4949
rect 784 4915 790 4949
rect 744 4877 790 4915
rect 744 4843 750 4877
rect 784 4843 790 4877
rect 744 4805 790 4843
rect 744 4771 750 4805
rect 784 4771 790 4805
rect 744 4733 790 4771
rect 744 4699 750 4733
rect 784 4699 790 4733
rect 744 4661 790 4699
rect 744 4627 750 4661
rect 784 4627 790 4661
rect 744 4589 790 4627
rect 744 4555 750 4589
rect 784 4555 790 4589
rect 744 4517 790 4555
rect 744 4483 750 4517
rect 784 4483 790 4517
rect 744 4445 790 4483
rect 744 4411 750 4445
rect 784 4411 790 4445
rect 744 4373 790 4411
rect 744 4339 750 4373
rect 784 4339 790 4373
rect 744 4301 790 4339
rect 744 4267 750 4301
rect 784 4267 790 4301
rect 744 4229 790 4267
rect 744 4195 750 4229
rect 784 4195 790 4229
rect 744 4157 790 4195
rect 744 4123 750 4157
rect 784 4123 790 4157
rect 744 4085 790 4123
rect 744 4051 750 4085
rect 784 4051 790 4085
rect 744 4013 790 4051
rect 744 3979 750 4013
rect 784 3979 790 4013
rect 744 3941 790 3979
rect 744 3907 750 3941
rect 784 3907 790 3941
rect 744 3869 790 3907
rect 744 3835 750 3869
rect 784 3835 790 3869
rect 744 3797 790 3835
rect 744 3763 750 3797
rect 784 3763 790 3797
rect 744 3725 790 3763
rect 744 3691 750 3725
rect 784 3691 790 3725
rect 744 3653 790 3691
rect 744 3619 750 3653
rect 784 3619 790 3653
rect 744 3581 790 3619
rect 744 3547 750 3581
rect 784 3547 790 3581
rect 744 3509 790 3547
rect 744 3475 750 3509
rect 784 3475 790 3509
rect 744 3437 790 3475
rect 744 3403 750 3437
rect 784 3403 790 3437
rect 744 3365 790 3403
rect 744 3331 750 3365
rect 784 3331 790 3365
rect 744 3293 790 3331
rect 744 3259 750 3293
rect 784 3259 790 3293
rect 744 3221 790 3259
rect 744 3187 750 3221
rect 784 3187 790 3221
rect 744 3149 790 3187
rect 744 3115 750 3149
rect 784 3115 790 3149
rect 744 3077 790 3115
rect 744 3043 750 3077
rect 784 3043 790 3077
rect 744 3005 790 3043
rect 744 2971 750 3005
rect 784 2971 790 3005
rect 744 2933 790 2971
rect 744 2899 750 2933
rect 784 2899 790 2933
rect 744 2861 790 2899
rect 744 2827 750 2861
rect 784 2827 790 2861
rect 744 2789 790 2827
rect 744 2755 750 2789
rect 784 2755 790 2789
rect 744 2717 790 2755
rect 744 2683 750 2717
rect 784 2683 790 2717
rect 744 2645 790 2683
rect 744 2611 750 2645
rect 784 2611 790 2645
rect 744 2573 790 2611
rect 744 2539 750 2573
rect 784 2539 790 2573
rect 744 2501 790 2539
rect 744 2467 750 2501
rect 784 2467 790 2501
rect 744 2429 790 2467
rect 744 2395 750 2429
rect 784 2395 790 2429
rect 744 2357 790 2395
rect 744 2323 750 2357
rect 784 2323 790 2357
rect 744 2285 790 2323
rect 744 2251 750 2285
rect 784 2251 790 2285
rect 744 2213 790 2251
rect 744 2179 750 2213
rect 784 2179 790 2213
rect 744 2141 790 2179
rect 744 2107 750 2141
rect 784 2107 790 2141
rect 744 2069 790 2107
rect 744 2035 750 2069
rect 784 2035 790 2069
rect 744 1997 790 2035
rect 744 1963 750 1997
rect 784 1963 790 1997
rect 744 1925 790 1963
rect 744 1891 750 1925
rect 784 1891 790 1925
rect 744 1853 790 1891
rect 744 1819 750 1853
rect 784 1819 790 1853
rect 744 1781 790 1819
rect 744 1747 750 1781
rect 784 1747 790 1781
rect 744 1709 790 1747
rect 744 1675 750 1709
rect 784 1675 790 1709
rect 744 1637 790 1675
rect 744 1603 750 1637
rect 784 1603 790 1637
rect 744 1565 790 1603
rect 744 1531 750 1565
rect 784 1531 790 1565
rect 744 1493 790 1531
rect 744 1459 750 1493
rect 784 1459 790 1493
rect 744 1421 790 1459
rect 744 1387 750 1421
rect 784 1387 790 1421
rect 744 1349 790 1387
rect 744 1315 750 1349
rect 784 1315 790 1349
rect 744 1277 790 1315
rect 744 1243 750 1277
rect 784 1243 790 1277
rect 744 1205 790 1243
rect 744 1171 750 1205
rect 784 1171 790 1205
rect 744 1133 790 1171
rect 744 1099 750 1133
rect 784 1099 790 1133
rect 744 1061 790 1099
rect 744 1027 750 1061
rect 784 1027 790 1061
rect 744 989 790 1027
rect 744 955 750 989
rect 784 955 790 989
rect 744 917 790 955
rect 744 883 750 917
rect 784 883 790 917
rect 744 845 790 883
rect 744 811 750 845
rect 784 811 790 845
rect 744 773 790 811
rect 744 739 750 773
rect 784 739 790 773
rect 744 701 790 739
rect 744 667 750 701
rect 784 667 790 701
rect 744 629 790 667
rect 744 595 750 629
rect 784 595 790 629
rect 744 557 790 595
rect 744 523 750 557
rect 784 523 790 557
rect 744 485 790 523
rect 744 451 750 485
rect 784 451 790 485
rect 744 413 790 451
rect 744 379 750 413
rect 784 379 790 413
rect 744 341 790 379
rect 744 307 750 341
rect 784 307 790 341
rect 744 269 790 307
rect 744 235 750 269
rect 784 235 790 269
rect 744 197 790 235
rect 744 163 750 197
rect 784 163 790 197
rect 744 125 790 163
rect 744 91 750 125
rect 784 91 790 125
rect 744 53 790 91
rect 744 19 750 53
rect 784 19 790 53
rect 744 -19 790 19
rect 744 -53 750 -19
rect 784 -53 790 -19
rect 744 -91 790 -53
rect 744 -125 750 -91
rect 784 -125 790 -91
rect 744 -163 790 -125
rect 744 -197 750 -163
rect 784 -197 790 -163
rect 744 -235 790 -197
rect 744 -269 750 -235
rect 784 -269 790 -235
rect 744 -307 790 -269
rect 744 -341 750 -307
rect 784 -341 790 -307
rect 744 -379 790 -341
rect 744 -413 750 -379
rect 784 -413 790 -379
rect 744 -451 790 -413
rect 744 -485 750 -451
rect 784 -485 790 -451
rect 744 -523 790 -485
rect 744 -557 750 -523
rect 784 -557 790 -523
rect 744 -595 790 -557
rect 744 -629 750 -595
rect 784 -629 790 -595
rect 744 -667 790 -629
rect 744 -701 750 -667
rect 784 -701 790 -667
rect 744 -739 790 -701
rect 744 -773 750 -739
rect 784 -773 790 -739
rect 744 -811 790 -773
rect 744 -845 750 -811
rect 784 -845 790 -811
rect 744 -883 790 -845
rect 744 -917 750 -883
rect 784 -917 790 -883
rect 744 -955 790 -917
rect 744 -989 750 -955
rect 784 -989 790 -955
rect 744 -1027 790 -989
rect 744 -1061 750 -1027
rect 784 -1061 790 -1027
rect 744 -1099 790 -1061
rect 744 -1133 750 -1099
rect 784 -1133 790 -1099
rect 744 -1171 790 -1133
rect 744 -1205 750 -1171
rect 784 -1205 790 -1171
rect 744 -1243 790 -1205
rect 744 -1277 750 -1243
rect 784 -1277 790 -1243
rect 744 -1315 790 -1277
rect 744 -1349 750 -1315
rect 784 -1349 790 -1315
rect 744 -1387 790 -1349
rect 744 -1421 750 -1387
rect 784 -1421 790 -1387
rect 744 -1459 790 -1421
rect 744 -1493 750 -1459
rect 784 -1493 790 -1459
rect 744 -1531 790 -1493
rect 744 -1565 750 -1531
rect 784 -1565 790 -1531
rect 744 -1603 790 -1565
rect 744 -1637 750 -1603
rect 784 -1637 790 -1603
rect 744 -1675 790 -1637
rect 744 -1709 750 -1675
rect 784 -1709 790 -1675
rect 744 -1747 790 -1709
rect 744 -1781 750 -1747
rect 784 -1781 790 -1747
rect 744 -1819 790 -1781
rect 744 -1853 750 -1819
rect 784 -1853 790 -1819
rect 744 -1891 790 -1853
rect 744 -1925 750 -1891
rect 784 -1925 790 -1891
rect 744 -1963 790 -1925
rect 744 -1997 750 -1963
rect 784 -1997 790 -1963
rect 744 -2035 790 -1997
rect 744 -2069 750 -2035
rect 784 -2069 790 -2035
rect 744 -2107 790 -2069
rect 744 -2141 750 -2107
rect 784 -2141 790 -2107
rect 744 -2179 790 -2141
rect 744 -2213 750 -2179
rect 784 -2213 790 -2179
rect 744 -2251 790 -2213
rect 744 -2285 750 -2251
rect 784 -2285 790 -2251
rect 744 -2323 790 -2285
rect 744 -2357 750 -2323
rect 784 -2357 790 -2323
rect 744 -2395 790 -2357
rect 744 -2429 750 -2395
rect 784 -2429 790 -2395
rect 744 -2467 790 -2429
rect 744 -2501 750 -2467
rect 784 -2501 790 -2467
rect 744 -2539 790 -2501
rect 744 -2573 750 -2539
rect 784 -2573 790 -2539
rect 744 -2611 790 -2573
rect 744 -2645 750 -2611
rect 784 -2645 790 -2611
rect 744 -2683 790 -2645
rect 744 -2717 750 -2683
rect 784 -2717 790 -2683
rect 744 -2755 790 -2717
rect 744 -2789 750 -2755
rect 784 -2789 790 -2755
rect 744 -2827 790 -2789
rect 744 -2861 750 -2827
rect 784 -2861 790 -2827
rect 744 -2899 790 -2861
rect 744 -2933 750 -2899
rect 784 -2933 790 -2899
rect 744 -2971 790 -2933
rect 744 -3005 750 -2971
rect 784 -3005 790 -2971
rect 744 -3043 790 -3005
rect 744 -3077 750 -3043
rect 784 -3077 790 -3043
rect 744 -3115 790 -3077
rect 744 -3149 750 -3115
rect 784 -3149 790 -3115
rect 744 -3187 790 -3149
rect 744 -3221 750 -3187
rect 784 -3221 790 -3187
rect 744 -3259 790 -3221
rect 744 -3293 750 -3259
rect 784 -3293 790 -3259
rect 744 -3331 790 -3293
rect 744 -3365 750 -3331
rect 784 -3365 790 -3331
rect 744 -3403 790 -3365
rect 744 -3437 750 -3403
rect 784 -3437 790 -3403
rect 744 -3475 790 -3437
rect 744 -3509 750 -3475
rect 784 -3509 790 -3475
rect 744 -3547 790 -3509
rect 744 -3581 750 -3547
rect 784 -3581 790 -3547
rect 744 -3619 790 -3581
rect 744 -3653 750 -3619
rect 784 -3653 790 -3619
rect 744 -3691 790 -3653
rect 744 -3725 750 -3691
rect 784 -3725 790 -3691
rect 744 -3763 790 -3725
rect 744 -3797 750 -3763
rect 784 -3797 790 -3763
rect 744 -3835 790 -3797
rect 744 -3869 750 -3835
rect 784 -3869 790 -3835
rect 744 -3907 790 -3869
rect 744 -3941 750 -3907
rect 784 -3941 790 -3907
rect 744 -3979 790 -3941
rect 744 -4013 750 -3979
rect 784 -4013 790 -3979
rect 744 -4051 790 -4013
rect 744 -4085 750 -4051
rect 784 -4085 790 -4051
rect 744 -4123 790 -4085
rect 744 -4157 750 -4123
rect 784 -4157 790 -4123
rect 744 -4195 790 -4157
rect 744 -4229 750 -4195
rect 784 -4229 790 -4195
rect 744 -4267 790 -4229
rect 744 -4301 750 -4267
rect 784 -4301 790 -4267
rect 744 -4339 790 -4301
rect 744 -4373 750 -4339
rect 784 -4373 790 -4339
rect 744 -4411 790 -4373
rect 744 -4445 750 -4411
rect 784 -4445 790 -4411
rect 744 -4483 790 -4445
rect 744 -4517 750 -4483
rect 784 -4517 790 -4483
rect 744 -4555 790 -4517
rect 744 -4589 750 -4555
rect 784 -4589 790 -4555
rect 744 -4627 790 -4589
rect 744 -4661 750 -4627
rect 784 -4661 790 -4627
rect 744 -4699 790 -4661
rect 744 -4733 750 -4699
rect 784 -4733 790 -4699
rect 744 -4771 790 -4733
rect 744 -4805 750 -4771
rect 784 -4805 790 -4771
rect 744 -4843 790 -4805
rect 744 -4877 750 -4843
rect 784 -4877 790 -4843
rect 744 -4915 790 -4877
rect 744 -4949 750 -4915
rect 784 -4949 790 -4915
rect 744 -4987 790 -4949
rect 744 -5021 750 -4987
rect 784 -5021 790 -4987
rect 744 -5059 790 -5021
rect 744 -5093 750 -5059
rect 784 -5093 790 -5059
rect 744 -5131 790 -5093
rect 744 -5165 750 -5131
rect 784 -5165 790 -5131
rect 744 -5203 790 -5165
rect 744 -5237 750 -5203
rect 784 -5237 790 -5203
rect 744 -5275 790 -5237
rect 744 -5309 750 -5275
rect 784 -5309 790 -5275
rect 744 -5347 790 -5309
rect 744 -5381 750 -5347
rect 784 -5381 790 -5347
rect 744 -5419 790 -5381
rect 744 -5453 750 -5419
rect 784 -5453 790 -5419
rect 744 -5491 790 -5453
rect 744 -5525 750 -5491
rect 784 -5525 790 -5491
rect 744 -5563 790 -5525
rect 744 -5597 750 -5563
rect 784 -5597 790 -5563
rect 744 -5635 790 -5597
rect 744 -5669 750 -5635
rect 784 -5669 790 -5635
rect 744 -5707 790 -5669
rect 744 -5741 750 -5707
rect 784 -5741 790 -5707
rect 744 -5779 790 -5741
rect 744 -5813 750 -5779
rect 784 -5813 790 -5779
rect 744 -5851 790 -5813
rect 744 -5885 750 -5851
rect 784 -5885 790 -5851
rect 744 -5923 790 -5885
rect 744 -5957 750 -5923
rect 784 -5957 790 -5923
rect 744 -5995 790 -5957
rect 744 -6029 750 -5995
rect 784 -6029 790 -5995
rect 744 -6067 790 -6029
rect 744 -6101 750 -6067
rect 784 -6101 790 -6067
rect 744 -6139 790 -6101
rect 744 -6173 750 -6139
rect 784 -6173 790 -6139
rect 744 -6211 790 -6173
rect 744 -6245 750 -6211
rect 784 -6245 790 -6211
rect 744 -6283 790 -6245
rect 744 -6317 750 -6283
rect 784 -6317 790 -6283
rect 744 -6355 790 -6317
rect 744 -6389 750 -6355
rect 784 -6389 790 -6355
rect 744 -6427 790 -6389
rect 744 -6461 750 -6427
rect 784 -6461 790 -6427
rect 744 -6499 790 -6461
rect 744 -6533 750 -6499
rect 784 -6533 790 -6499
rect 744 -6571 790 -6533
rect 744 -6605 750 -6571
rect 784 -6605 790 -6571
rect 744 -6643 790 -6605
rect 744 -6677 750 -6643
rect 784 -6677 790 -6643
rect 744 -6715 790 -6677
rect 744 -6749 750 -6715
rect 784 -6749 790 -6715
rect 744 -6787 790 -6749
rect 744 -6821 750 -6787
rect 784 -6821 790 -6787
rect 744 -6859 790 -6821
rect 744 -6893 750 -6859
rect 784 -6893 790 -6859
rect 744 -6931 790 -6893
rect 744 -6965 750 -6931
rect 784 -6965 790 -6931
rect 744 -7003 790 -6965
rect 744 -7037 750 -7003
rect 784 -7037 790 -7003
rect 744 -7075 790 -7037
rect 744 -7109 750 -7075
rect 784 -7109 790 -7075
rect 744 -7147 790 -7109
rect 744 -7181 750 -7147
rect 784 -7181 790 -7147
rect 744 -7219 790 -7181
rect 744 -7253 750 -7219
rect 784 -7253 790 -7219
rect 744 -7291 790 -7253
rect 744 -7325 750 -7291
rect 784 -7325 790 -7291
rect 744 -7363 790 -7325
rect 744 -7397 750 -7363
rect 784 -7397 790 -7363
rect 744 -7435 790 -7397
rect 744 -7469 750 -7435
rect 784 -7469 790 -7435
rect 744 -7507 790 -7469
rect 744 -7541 750 -7507
rect 784 -7541 790 -7507
rect 744 -7579 790 -7541
rect 744 -7613 750 -7579
rect 784 -7613 790 -7579
rect 744 -7651 790 -7613
rect 744 -7685 750 -7651
rect 784 -7685 790 -7651
rect 744 -7723 790 -7685
rect 744 -7757 750 -7723
rect 784 -7757 790 -7723
rect 744 -7795 790 -7757
rect 744 -7829 750 -7795
rect 784 -7829 790 -7795
rect 744 -7867 790 -7829
rect 744 -7901 750 -7867
rect 784 -7901 790 -7867
rect 744 -7939 790 -7901
rect 744 -7973 750 -7939
rect 784 -7973 790 -7939
rect 744 -8011 790 -7973
rect 744 -8045 750 -8011
rect 784 -8045 790 -8011
rect 744 -8083 790 -8045
rect 744 -8117 750 -8083
rect 784 -8117 790 -8083
rect 744 -8155 790 -8117
rect 744 -8189 750 -8155
rect 784 -8189 790 -8155
rect 744 -8227 790 -8189
rect 744 -8261 750 -8227
rect 784 -8261 790 -8227
rect 744 -8299 790 -8261
rect 744 -8333 750 -8299
rect 784 -8333 790 -8299
rect 744 -8371 790 -8333
rect 744 -8405 750 -8371
rect 784 -8405 790 -8371
rect 744 -8443 790 -8405
rect 744 -8477 750 -8443
rect 784 -8477 790 -8443
rect 744 -8515 790 -8477
rect 744 -8549 750 -8515
rect 784 -8549 790 -8515
rect 744 -8587 790 -8549
rect 744 -8621 750 -8587
rect 784 -8621 790 -8587
rect 744 -8659 790 -8621
rect 744 -8693 750 -8659
rect 784 -8693 790 -8659
rect 744 -8731 790 -8693
rect 744 -8765 750 -8731
rect 784 -8765 790 -8731
rect 744 -8803 790 -8765
rect 744 -8837 750 -8803
rect 784 -8837 790 -8803
rect 744 -8875 790 -8837
rect 744 -8909 750 -8875
rect 784 -8909 790 -8875
rect 744 -8947 790 -8909
rect 744 -8981 750 -8947
rect 784 -8981 790 -8947
rect 744 -9019 790 -8981
rect 744 -9053 750 -9019
rect 784 -9053 790 -9019
rect 744 -9091 790 -9053
rect 744 -9125 750 -9091
rect 784 -9125 790 -9091
rect 744 -9163 790 -9125
rect 744 -9197 750 -9163
rect 784 -9197 790 -9163
rect 744 -9235 790 -9197
rect 744 -9269 750 -9235
rect 784 -9269 790 -9235
rect 744 -9307 790 -9269
rect 744 -9341 750 -9307
rect 784 -9341 790 -9307
rect 744 -9379 790 -9341
rect 744 -9413 750 -9379
rect 784 -9413 790 -9379
rect 744 -9451 790 -9413
rect 744 -9485 750 -9451
rect 784 -9485 790 -9451
rect 744 -9523 790 -9485
rect 744 -9557 750 -9523
rect 784 -9557 790 -9523
rect 744 -9600 790 -9557
rect 862 9557 908 9600
rect 862 9523 868 9557
rect 902 9523 908 9557
rect 862 9485 908 9523
rect 862 9451 868 9485
rect 902 9451 908 9485
rect 862 9413 908 9451
rect 862 9379 868 9413
rect 902 9379 908 9413
rect 862 9341 908 9379
rect 862 9307 868 9341
rect 902 9307 908 9341
rect 862 9269 908 9307
rect 862 9235 868 9269
rect 902 9235 908 9269
rect 862 9197 908 9235
rect 862 9163 868 9197
rect 902 9163 908 9197
rect 862 9125 908 9163
rect 862 9091 868 9125
rect 902 9091 908 9125
rect 862 9053 908 9091
rect 862 9019 868 9053
rect 902 9019 908 9053
rect 862 8981 908 9019
rect 862 8947 868 8981
rect 902 8947 908 8981
rect 862 8909 908 8947
rect 862 8875 868 8909
rect 902 8875 908 8909
rect 862 8837 908 8875
rect 862 8803 868 8837
rect 902 8803 908 8837
rect 862 8765 908 8803
rect 862 8731 868 8765
rect 902 8731 908 8765
rect 862 8693 908 8731
rect 862 8659 868 8693
rect 902 8659 908 8693
rect 862 8621 908 8659
rect 862 8587 868 8621
rect 902 8587 908 8621
rect 862 8549 908 8587
rect 862 8515 868 8549
rect 902 8515 908 8549
rect 862 8477 908 8515
rect 862 8443 868 8477
rect 902 8443 908 8477
rect 862 8405 908 8443
rect 862 8371 868 8405
rect 902 8371 908 8405
rect 862 8333 908 8371
rect 862 8299 868 8333
rect 902 8299 908 8333
rect 862 8261 908 8299
rect 862 8227 868 8261
rect 902 8227 908 8261
rect 862 8189 908 8227
rect 862 8155 868 8189
rect 902 8155 908 8189
rect 862 8117 908 8155
rect 862 8083 868 8117
rect 902 8083 908 8117
rect 862 8045 908 8083
rect 862 8011 868 8045
rect 902 8011 908 8045
rect 862 7973 908 8011
rect 862 7939 868 7973
rect 902 7939 908 7973
rect 862 7901 908 7939
rect 862 7867 868 7901
rect 902 7867 908 7901
rect 862 7829 908 7867
rect 862 7795 868 7829
rect 902 7795 908 7829
rect 862 7757 908 7795
rect 862 7723 868 7757
rect 902 7723 908 7757
rect 862 7685 908 7723
rect 862 7651 868 7685
rect 902 7651 908 7685
rect 862 7613 908 7651
rect 862 7579 868 7613
rect 902 7579 908 7613
rect 862 7541 908 7579
rect 862 7507 868 7541
rect 902 7507 908 7541
rect 862 7469 908 7507
rect 862 7435 868 7469
rect 902 7435 908 7469
rect 862 7397 908 7435
rect 862 7363 868 7397
rect 902 7363 908 7397
rect 862 7325 908 7363
rect 862 7291 868 7325
rect 902 7291 908 7325
rect 862 7253 908 7291
rect 862 7219 868 7253
rect 902 7219 908 7253
rect 862 7181 908 7219
rect 862 7147 868 7181
rect 902 7147 908 7181
rect 862 7109 908 7147
rect 862 7075 868 7109
rect 902 7075 908 7109
rect 862 7037 908 7075
rect 862 7003 868 7037
rect 902 7003 908 7037
rect 862 6965 908 7003
rect 862 6931 868 6965
rect 902 6931 908 6965
rect 862 6893 908 6931
rect 862 6859 868 6893
rect 902 6859 908 6893
rect 862 6821 908 6859
rect 862 6787 868 6821
rect 902 6787 908 6821
rect 862 6749 908 6787
rect 862 6715 868 6749
rect 902 6715 908 6749
rect 862 6677 908 6715
rect 862 6643 868 6677
rect 902 6643 908 6677
rect 862 6605 908 6643
rect 862 6571 868 6605
rect 902 6571 908 6605
rect 862 6533 908 6571
rect 862 6499 868 6533
rect 902 6499 908 6533
rect 862 6461 908 6499
rect 862 6427 868 6461
rect 902 6427 908 6461
rect 862 6389 908 6427
rect 862 6355 868 6389
rect 902 6355 908 6389
rect 862 6317 908 6355
rect 862 6283 868 6317
rect 902 6283 908 6317
rect 862 6245 908 6283
rect 862 6211 868 6245
rect 902 6211 908 6245
rect 862 6173 908 6211
rect 862 6139 868 6173
rect 902 6139 908 6173
rect 862 6101 908 6139
rect 862 6067 868 6101
rect 902 6067 908 6101
rect 862 6029 908 6067
rect 862 5995 868 6029
rect 902 5995 908 6029
rect 862 5957 908 5995
rect 862 5923 868 5957
rect 902 5923 908 5957
rect 862 5885 908 5923
rect 862 5851 868 5885
rect 902 5851 908 5885
rect 862 5813 908 5851
rect 862 5779 868 5813
rect 902 5779 908 5813
rect 862 5741 908 5779
rect 862 5707 868 5741
rect 902 5707 908 5741
rect 862 5669 908 5707
rect 862 5635 868 5669
rect 902 5635 908 5669
rect 862 5597 908 5635
rect 862 5563 868 5597
rect 902 5563 908 5597
rect 862 5525 908 5563
rect 862 5491 868 5525
rect 902 5491 908 5525
rect 862 5453 908 5491
rect 862 5419 868 5453
rect 902 5419 908 5453
rect 862 5381 908 5419
rect 862 5347 868 5381
rect 902 5347 908 5381
rect 862 5309 908 5347
rect 862 5275 868 5309
rect 902 5275 908 5309
rect 862 5237 908 5275
rect 862 5203 868 5237
rect 902 5203 908 5237
rect 862 5165 908 5203
rect 862 5131 868 5165
rect 902 5131 908 5165
rect 862 5093 908 5131
rect 862 5059 868 5093
rect 902 5059 908 5093
rect 862 5021 908 5059
rect 862 4987 868 5021
rect 902 4987 908 5021
rect 862 4949 908 4987
rect 862 4915 868 4949
rect 902 4915 908 4949
rect 862 4877 908 4915
rect 862 4843 868 4877
rect 902 4843 908 4877
rect 862 4805 908 4843
rect 862 4771 868 4805
rect 902 4771 908 4805
rect 862 4733 908 4771
rect 862 4699 868 4733
rect 902 4699 908 4733
rect 862 4661 908 4699
rect 862 4627 868 4661
rect 902 4627 908 4661
rect 862 4589 908 4627
rect 862 4555 868 4589
rect 902 4555 908 4589
rect 862 4517 908 4555
rect 862 4483 868 4517
rect 902 4483 908 4517
rect 862 4445 908 4483
rect 862 4411 868 4445
rect 902 4411 908 4445
rect 862 4373 908 4411
rect 862 4339 868 4373
rect 902 4339 908 4373
rect 862 4301 908 4339
rect 862 4267 868 4301
rect 902 4267 908 4301
rect 862 4229 908 4267
rect 862 4195 868 4229
rect 902 4195 908 4229
rect 862 4157 908 4195
rect 862 4123 868 4157
rect 902 4123 908 4157
rect 862 4085 908 4123
rect 862 4051 868 4085
rect 902 4051 908 4085
rect 862 4013 908 4051
rect 862 3979 868 4013
rect 902 3979 908 4013
rect 862 3941 908 3979
rect 862 3907 868 3941
rect 902 3907 908 3941
rect 862 3869 908 3907
rect 862 3835 868 3869
rect 902 3835 908 3869
rect 862 3797 908 3835
rect 862 3763 868 3797
rect 902 3763 908 3797
rect 862 3725 908 3763
rect 862 3691 868 3725
rect 902 3691 908 3725
rect 862 3653 908 3691
rect 862 3619 868 3653
rect 902 3619 908 3653
rect 862 3581 908 3619
rect 862 3547 868 3581
rect 902 3547 908 3581
rect 862 3509 908 3547
rect 862 3475 868 3509
rect 902 3475 908 3509
rect 862 3437 908 3475
rect 862 3403 868 3437
rect 902 3403 908 3437
rect 862 3365 908 3403
rect 862 3331 868 3365
rect 902 3331 908 3365
rect 862 3293 908 3331
rect 862 3259 868 3293
rect 902 3259 908 3293
rect 862 3221 908 3259
rect 862 3187 868 3221
rect 902 3187 908 3221
rect 862 3149 908 3187
rect 862 3115 868 3149
rect 902 3115 908 3149
rect 862 3077 908 3115
rect 862 3043 868 3077
rect 902 3043 908 3077
rect 862 3005 908 3043
rect 862 2971 868 3005
rect 902 2971 908 3005
rect 862 2933 908 2971
rect 862 2899 868 2933
rect 902 2899 908 2933
rect 862 2861 908 2899
rect 862 2827 868 2861
rect 902 2827 908 2861
rect 862 2789 908 2827
rect 862 2755 868 2789
rect 902 2755 908 2789
rect 862 2717 908 2755
rect 862 2683 868 2717
rect 902 2683 908 2717
rect 862 2645 908 2683
rect 862 2611 868 2645
rect 902 2611 908 2645
rect 862 2573 908 2611
rect 862 2539 868 2573
rect 902 2539 908 2573
rect 862 2501 908 2539
rect 862 2467 868 2501
rect 902 2467 908 2501
rect 862 2429 908 2467
rect 862 2395 868 2429
rect 902 2395 908 2429
rect 862 2357 908 2395
rect 862 2323 868 2357
rect 902 2323 908 2357
rect 862 2285 908 2323
rect 862 2251 868 2285
rect 902 2251 908 2285
rect 862 2213 908 2251
rect 862 2179 868 2213
rect 902 2179 908 2213
rect 862 2141 908 2179
rect 862 2107 868 2141
rect 902 2107 908 2141
rect 862 2069 908 2107
rect 862 2035 868 2069
rect 902 2035 908 2069
rect 862 1997 908 2035
rect 862 1963 868 1997
rect 902 1963 908 1997
rect 862 1925 908 1963
rect 862 1891 868 1925
rect 902 1891 908 1925
rect 862 1853 908 1891
rect 862 1819 868 1853
rect 902 1819 908 1853
rect 862 1781 908 1819
rect 862 1747 868 1781
rect 902 1747 908 1781
rect 862 1709 908 1747
rect 862 1675 868 1709
rect 902 1675 908 1709
rect 862 1637 908 1675
rect 862 1603 868 1637
rect 902 1603 908 1637
rect 862 1565 908 1603
rect 862 1531 868 1565
rect 902 1531 908 1565
rect 862 1493 908 1531
rect 862 1459 868 1493
rect 902 1459 908 1493
rect 862 1421 908 1459
rect 862 1387 868 1421
rect 902 1387 908 1421
rect 862 1349 908 1387
rect 862 1315 868 1349
rect 902 1315 908 1349
rect 862 1277 908 1315
rect 862 1243 868 1277
rect 902 1243 908 1277
rect 862 1205 908 1243
rect 862 1171 868 1205
rect 902 1171 908 1205
rect 862 1133 908 1171
rect 862 1099 868 1133
rect 902 1099 908 1133
rect 862 1061 908 1099
rect 862 1027 868 1061
rect 902 1027 908 1061
rect 862 989 908 1027
rect 862 955 868 989
rect 902 955 908 989
rect 862 917 908 955
rect 862 883 868 917
rect 902 883 908 917
rect 862 845 908 883
rect 862 811 868 845
rect 902 811 908 845
rect 862 773 908 811
rect 862 739 868 773
rect 902 739 908 773
rect 862 701 908 739
rect 862 667 868 701
rect 902 667 908 701
rect 862 629 908 667
rect 862 595 868 629
rect 902 595 908 629
rect 862 557 908 595
rect 862 523 868 557
rect 902 523 908 557
rect 862 485 908 523
rect 862 451 868 485
rect 902 451 908 485
rect 862 413 908 451
rect 862 379 868 413
rect 902 379 908 413
rect 862 341 908 379
rect 862 307 868 341
rect 902 307 908 341
rect 862 269 908 307
rect 862 235 868 269
rect 902 235 908 269
rect 862 197 908 235
rect 862 163 868 197
rect 902 163 908 197
rect 862 125 908 163
rect 862 91 868 125
rect 902 91 908 125
rect 862 53 908 91
rect 862 19 868 53
rect 902 19 908 53
rect 862 -19 908 19
rect 862 -53 868 -19
rect 902 -53 908 -19
rect 862 -91 908 -53
rect 862 -125 868 -91
rect 902 -125 908 -91
rect 862 -163 908 -125
rect 862 -197 868 -163
rect 902 -197 908 -163
rect 862 -235 908 -197
rect 862 -269 868 -235
rect 902 -269 908 -235
rect 862 -307 908 -269
rect 862 -341 868 -307
rect 902 -341 908 -307
rect 862 -379 908 -341
rect 862 -413 868 -379
rect 902 -413 908 -379
rect 862 -451 908 -413
rect 862 -485 868 -451
rect 902 -485 908 -451
rect 862 -523 908 -485
rect 862 -557 868 -523
rect 902 -557 908 -523
rect 862 -595 908 -557
rect 862 -629 868 -595
rect 902 -629 908 -595
rect 862 -667 908 -629
rect 862 -701 868 -667
rect 902 -701 908 -667
rect 862 -739 908 -701
rect 862 -773 868 -739
rect 902 -773 908 -739
rect 862 -811 908 -773
rect 862 -845 868 -811
rect 902 -845 908 -811
rect 862 -883 908 -845
rect 862 -917 868 -883
rect 902 -917 908 -883
rect 862 -955 908 -917
rect 862 -989 868 -955
rect 902 -989 908 -955
rect 862 -1027 908 -989
rect 862 -1061 868 -1027
rect 902 -1061 908 -1027
rect 862 -1099 908 -1061
rect 862 -1133 868 -1099
rect 902 -1133 908 -1099
rect 862 -1171 908 -1133
rect 862 -1205 868 -1171
rect 902 -1205 908 -1171
rect 862 -1243 908 -1205
rect 862 -1277 868 -1243
rect 902 -1277 908 -1243
rect 862 -1315 908 -1277
rect 862 -1349 868 -1315
rect 902 -1349 908 -1315
rect 862 -1387 908 -1349
rect 862 -1421 868 -1387
rect 902 -1421 908 -1387
rect 862 -1459 908 -1421
rect 862 -1493 868 -1459
rect 902 -1493 908 -1459
rect 862 -1531 908 -1493
rect 862 -1565 868 -1531
rect 902 -1565 908 -1531
rect 862 -1603 908 -1565
rect 862 -1637 868 -1603
rect 902 -1637 908 -1603
rect 862 -1675 908 -1637
rect 862 -1709 868 -1675
rect 902 -1709 908 -1675
rect 862 -1747 908 -1709
rect 862 -1781 868 -1747
rect 902 -1781 908 -1747
rect 862 -1819 908 -1781
rect 862 -1853 868 -1819
rect 902 -1853 908 -1819
rect 862 -1891 908 -1853
rect 862 -1925 868 -1891
rect 902 -1925 908 -1891
rect 862 -1963 908 -1925
rect 862 -1997 868 -1963
rect 902 -1997 908 -1963
rect 862 -2035 908 -1997
rect 862 -2069 868 -2035
rect 902 -2069 908 -2035
rect 862 -2107 908 -2069
rect 862 -2141 868 -2107
rect 902 -2141 908 -2107
rect 862 -2179 908 -2141
rect 862 -2213 868 -2179
rect 902 -2213 908 -2179
rect 862 -2251 908 -2213
rect 862 -2285 868 -2251
rect 902 -2285 908 -2251
rect 862 -2323 908 -2285
rect 862 -2357 868 -2323
rect 902 -2357 908 -2323
rect 862 -2395 908 -2357
rect 862 -2429 868 -2395
rect 902 -2429 908 -2395
rect 862 -2467 908 -2429
rect 862 -2501 868 -2467
rect 902 -2501 908 -2467
rect 862 -2539 908 -2501
rect 862 -2573 868 -2539
rect 902 -2573 908 -2539
rect 862 -2611 908 -2573
rect 862 -2645 868 -2611
rect 902 -2645 908 -2611
rect 862 -2683 908 -2645
rect 862 -2717 868 -2683
rect 902 -2717 908 -2683
rect 862 -2755 908 -2717
rect 862 -2789 868 -2755
rect 902 -2789 908 -2755
rect 862 -2827 908 -2789
rect 862 -2861 868 -2827
rect 902 -2861 908 -2827
rect 862 -2899 908 -2861
rect 862 -2933 868 -2899
rect 902 -2933 908 -2899
rect 862 -2971 908 -2933
rect 862 -3005 868 -2971
rect 902 -3005 908 -2971
rect 862 -3043 908 -3005
rect 862 -3077 868 -3043
rect 902 -3077 908 -3043
rect 862 -3115 908 -3077
rect 862 -3149 868 -3115
rect 902 -3149 908 -3115
rect 862 -3187 908 -3149
rect 862 -3221 868 -3187
rect 902 -3221 908 -3187
rect 862 -3259 908 -3221
rect 862 -3293 868 -3259
rect 902 -3293 908 -3259
rect 862 -3331 908 -3293
rect 862 -3365 868 -3331
rect 902 -3365 908 -3331
rect 862 -3403 908 -3365
rect 862 -3437 868 -3403
rect 902 -3437 908 -3403
rect 862 -3475 908 -3437
rect 862 -3509 868 -3475
rect 902 -3509 908 -3475
rect 862 -3547 908 -3509
rect 862 -3581 868 -3547
rect 902 -3581 908 -3547
rect 862 -3619 908 -3581
rect 862 -3653 868 -3619
rect 902 -3653 908 -3619
rect 862 -3691 908 -3653
rect 862 -3725 868 -3691
rect 902 -3725 908 -3691
rect 862 -3763 908 -3725
rect 862 -3797 868 -3763
rect 902 -3797 908 -3763
rect 862 -3835 908 -3797
rect 862 -3869 868 -3835
rect 902 -3869 908 -3835
rect 862 -3907 908 -3869
rect 862 -3941 868 -3907
rect 902 -3941 908 -3907
rect 862 -3979 908 -3941
rect 862 -4013 868 -3979
rect 902 -4013 908 -3979
rect 862 -4051 908 -4013
rect 862 -4085 868 -4051
rect 902 -4085 908 -4051
rect 862 -4123 908 -4085
rect 862 -4157 868 -4123
rect 902 -4157 908 -4123
rect 862 -4195 908 -4157
rect 862 -4229 868 -4195
rect 902 -4229 908 -4195
rect 862 -4267 908 -4229
rect 862 -4301 868 -4267
rect 902 -4301 908 -4267
rect 862 -4339 908 -4301
rect 862 -4373 868 -4339
rect 902 -4373 908 -4339
rect 862 -4411 908 -4373
rect 862 -4445 868 -4411
rect 902 -4445 908 -4411
rect 862 -4483 908 -4445
rect 862 -4517 868 -4483
rect 902 -4517 908 -4483
rect 862 -4555 908 -4517
rect 862 -4589 868 -4555
rect 902 -4589 908 -4555
rect 862 -4627 908 -4589
rect 862 -4661 868 -4627
rect 902 -4661 908 -4627
rect 862 -4699 908 -4661
rect 862 -4733 868 -4699
rect 902 -4733 908 -4699
rect 862 -4771 908 -4733
rect 862 -4805 868 -4771
rect 902 -4805 908 -4771
rect 862 -4843 908 -4805
rect 862 -4877 868 -4843
rect 902 -4877 908 -4843
rect 862 -4915 908 -4877
rect 862 -4949 868 -4915
rect 902 -4949 908 -4915
rect 862 -4987 908 -4949
rect 862 -5021 868 -4987
rect 902 -5021 908 -4987
rect 862 -5059 908 -5021
rect 862 -5093 868 -5059
rect 902 -5093 908 -5059
rect 862 -5131 908 -5093
rect 862 -5165 868 -5131
rect 902 -5165 908 -5131
rect 862 -5203 908 -5165
rect 862 -5237 868 -5203
rect 902 -5237 908 -5203
rect 862 -5275 908 -5237
rect 862 -5309 868 -5275
rect 902 -5309 908 -5275
rect 862 -5347 908 -5309
rect 862 -5381 868 -5347
rect 902 -5381 908 -5347
rect 862 -5419 908 -5381
rect 862 -5453 868 -5419
rect 902 -5453 908 -5419
rect 862 -5491 908 -5453
rect 862 -5525 868 -5491
rect 902 -5525 908 -5491
rect 862 -5563 908 -5525
rect 862 -5597 868 -5563
rect 902 -5597 908 -5563
rect 862 -5635 908 -5597
rect 862 -5669 868 -5635
rect 902 -5669 908 -5635
rect 862 -5707 908 -5669
rect 862 -5741 868 -5707
rect 902 -5741 908 -5707
rect 862 -5779 908 -5741
rect 862 -5813 868 -5779
rect 902 -5813 908 -5779
rect 862 -5851 908 -5813
rect 862 -5885 868 -5851
rect 902 -5885 908 -5851
rect 862 -5923 908 -5885
rect 862 -5957 868 -5923
rect 902 -5957 908 -5923
rect 862 -5995 908 -5957
rect 862 -6029 868 -5995
rect 902 -6029 908 -5995
rect 862 -6067 908 -6029
rect 862 -6101 868 -6067
rect 902 -6101 908 -6067
rect 862 -6139 908 -6101
rect 862 -6173 868 -6139
rect 902 -6173 908 -6139
rect 862 -6211 908 -6173
rect 862 -6245 868 -6211
rect 902 -6245 908 -6211
rect 862 -6283 908 -6245
rect 862 -6317 868 -6283
rect 902 -6317 908 -6283
rect 862 -6355 908 -6317
rect 862 -6389 868 -6355
rect 902 -6389 908 -6355
rect 862 -6427 908 -6389
rect 862 -6461 868 -6427
rect 902 -6461 908 -6427
rect 862 -6499 908 -6461
rect 862 -6533 868 -6499
rect 902 -6533 908 -6499
rect 862 -6571 908 -6533
rect 862 -6605 868 -6571
rect 902 -6605 908 -6571
rect 862 -6643 908 -6605
rect 862 -6677 868 -6643
rect 902 -6677 908 -6643
rect 862 -6715 908 -6677
rect 862 -6749 868 -6715
rect 902 -6749 908 -6715
rect 862 -6787 908 -6749
rect 862 -6821 868 -6787
rect 902 -6821 908 -6787
rect 862 -6859 908 -6821
rect 862 -6893 868 -6859
rect 902 -6893 908 -6859
rect 862 -6931 908 -6893
rect 862 -6965 868 -6931
rect 902 -6965 908 -6931
rect 862 -7003 908 -6965
rect 862 -7037 868 -7003
rect 902 -7037 908 -7003
rect 862 -7075 908 -7037
rect 862 -7109 868 -7075
rect 902 -7109 908 -7075
rect 862 -7147 908 -7109
rect 862 -7181 868 -7147
rect 902 -7181 908 -7147
rect 862 -7219 908 -7181
rect 862 -7253 868 -7219
rect 902 -7253 908 -7219
rect 862 -7291 908 -7253
rect 862 -7325 868 -7291
rect 902 -7325 908 -7291
rect 862 -7363 908 -7325
rect 862 -7397 868 -7363
rect 902 -7397 908 -7363
rect 862 -7435 908 -7397
rect 862 -7469 868 -7435
rect 902 -7469 908 -7435
rect 862 -7507 908 -7469
rect 862 -7541 868 -7507
rect 902 -7541 908 -7507
rect 862 -7579 908 -7541
rect 862 -7613 868 -7579
rect 902 -7613 908 -7579
rect 862 -7651 908 -7613
rect 862 -7685 868 -7651
rect 902 -7685 908 -7651
rect 862 -7723 908 -7685
rect 862 -7757 868 -7723
rect 902 -7757 908 -7723
rect 862 -7795 908 -7757
rect 862 -7829 868 -7795
rect 902 -7829 908 -7795
rect 862 -7867 908 -7829
rect 862 -7901 868 -7867
rect 902 -7901 908 -7867
rect 862 -7939 908 -7901
rect 862 -7973 868 -7939
rect 902 -7973 908 -7939
rect 862 -8011 908 -7973
rect 862 -8045 868 -8011
rect 902 -8045 908 -8011
rect 862 -8083 908 -8045
rect 862 -8117 868 -8083
rect 902 -8117 908 -8083
rect 862 -8155 908 -8117
rect 862 -8189 868 -8155
rect 902 -8189 908 -8155
rect 862 -8227 908 -8189
rect 862 -8261 868 -8227
rect 902 -8261 908 -8227
rect 862 -8299 908 -8261
rect 862 -8333 868 -8299
rect 902 -8333 908 -8299
rect 862 -8371 908 -8333
rect 862 -8405 868 -8371
rect 902 -8405 908 -8371
rect 862 -8443 908 -8405
rect 862 -8477 868 -8443
rect 902 -8477 908 -8443
rect 862 -8515 908 -8477
rect 862 -8549 868 -8515
rect 902 -8549 908 -8515
rect 862 -8587 908 -8549
rect 862 -8621 868 -8587
rect 902 -8621 908 -8587
rect 862 -8659 908 -8621
rect 862 -8693 868 -8659
rect 902 -8693 908 -8659
rect 862 -8731 908 -8693
rect 862 -8765 868 -8731
rect 902 -8765 908 -8731
rect 862 -8803 908 -8765
rect 862 -8837 868 -8803
rect 902 -8837 908 -8803
rect 862 -8875 908 -8837
rect 862 -8909 868 -8875
rect 902 -8909 908 -8875
rect 862 -8947 908 -8909
rect 862 -8981 868 -8947
rect 902 -8981 908 -8947
rect 862 -9019 908 -8981
rect 862 -9053 868 -9019
rect 902 -9053 908 -9019
rect 862 -9091 908 -9053
rect 862 -9125 868 -9091
rect 902 -9125 908 -9091
rect 862 -9163 908 -9125
rect 862 -9197 868 -9163
rect 902 -9197 908 -9163
rect 862 -9235 908 -9197
rect 862 -9269 868 -9235
rect 902 -9269 908 -9235
rect 862 -9307 908 -9269
rect 862 -9341 868 -9307
rect 902 -9341 908 -9307
rect 862 -9379 908 -9341
rect 862 -9413 868 -9379
rect 902 -9413 908 -9379
rect 862 -9451 908 -9413
rect 862 -9485 868 -9451
rect 902 -9485 908 -9451
rect 862 -9523 908 -9485
rect 862 -9557 868 -9523
rect 902 -9557 908 -9523
rect 862 -9600 908 -9557
rect 980 9557 1026 9600
rect 980 9523 986 9557
rect 1020 9523 1026 9557
rect 980 9485 1026 9523
rect 980 9451 986 9485
rect 1020 9451 1026 9485
rect 980 9413 1026 9451
rect 980 9379 986 9413
rect 1020 9379 1026 9413
rect 980 9341 1026 9379
rect 980 9307 986 9341
rect 1020 9307 1026 9341
rect 980 9269 1026 9307
rect 980 9235 986 9269
rect 1020 9235 1026 9269
rect 980 9197 1026 9235
rect 980 9163 986 9197
rect 1020 9163 1026 9197
rect 980 9125 1026 9163
rect 980 9091 986 9125
rect 1020 9091 1026 9125
rect 980 9053 1026 9091
rect 980 9019 986 9053
rect 1020 9019 1026 9053
rect 980 8981 1026 9019
rect 980 8947 986 8981
rect 1020 8947 1026 8981
rect 980 8909 1026 8947
rect 980 8875 986 8909
rect 1020 8875 1026 8909
rect 980 8837 1026 8875
rect 980 8803 986 8837
rect 1020 8803 1026 8837
rect 980 8765 1026 8803
rect 980 8731 986 8765
rect 1020 8731 1026 8765
rect 980 8693 1026 8731
rect 980 8659 986 8693
rect 1020 8659 1026 8693
rect 980 8621 1026 8659
rect 980 8587 986 8621
rect 1020 8587 1026 8621
rect 980 8549 1026 8587
rect 980 8515 986 8549
rect 1020 8515 1026 8549
rect 980 8477 1026 8515
rect 980 8443 986 8477
rect 1020 8443 1026 8477
rect 980 8405 1026 8443
rect 980 8371 986 8405
rect 1020 8371 1026 8405
rect 980 8333 1026 8371
rect 980 8299 986 8333
rect 1020 8299 1026 8333
rect 980 8261 1026 8299
rect 980 8227 986 8261
rect 1020 8227 1026 8261
rect 980 8189 1026 8227
rect 980 8155 986 8189
rect 1020 8155 1026 8189
rect 980 8117 1026 8155
rect 980 8083 986 8117
rect 1020 8083 1026 8117
rect 980 8045 1026 8083
rect 980 8011 986 8045
rect 1020 8011 1026 8045
rect 980 7973 1026 8011
rect 980 7939 986 7973
rect 1020 7939 1026 7973
rect 980 7901 1026 7939
rect 980 7867 986 7901
rect 1020 7867 1026 7901
rect 980 7829 1026 7867
rect 980 7795 986 7829
rect 1020 7795 1026 7829
rect 980 7757 1026 7795
rect 980 7723 986 7757
rect 1020 7723 1026 7757
rect 980 7685 1026 7723
rect 980 7651 986 7685
rect 1020 7651 1026 7685
rect 980 7613 1026 7651
rect 980 7579 986 7613
rect 1020 7579 1026 7613
rect 980 7541 1026 7579
rect 980 7507 986 7541
rect 1020 7507 1026 7541
rect 980 7469 1026 7507
rect 980 7435 986 7469
rect 1020 7435 1026 7469
rect 980 7397 1026 7435
rect 980 7363 986 7397
rect 1020 7363 1026 7397
rect 980 7325 1026 7363
rect 980 7291 986 7325
rect 1020 7291 1026 7325
rect 980 7253 1026 7291
rect 980 7219 986 7253
rect 1020 7219 1026 7253
rect 980 7181 1026 7219
rect 980 7147 986 7181
rect 1020 7147 1026 7181
rect 980 7109 1026 7147
rect 980 7075 986 7109
rect 1020 7075 1026 7109
rect 980 7037 1026 7075
rect 980 7003 986 7037
rect 1020 7003 1026 7037
rect 980 6965 1026 7003
rect 980 6931 986 6965
rect 1020 6931 1026 6965
rect 980 6893 1026 6931
rect 980 6859 986 6893
rect 1020 6859 1026 6893
rect 980 6821 1026 6859
rect 980 6787 986 6821
rect 1020 6787 1026 6821
rect 980 6749 1026 6787
rect 980 6715 986 6749
rect 1020 6715 1026 6749
rect 980 6677 1026 6715
rect 980 6643 986 6677
rect 1020 6643 1026 6677
rect 980 6605 1026 6643
rect 980 6571 986 6605
rect 1020 6571 1026 6605
rect 980 6533 1026 6571
rect 980 6499 986 6533
rect 1020 6499 1026 6533
rect 980 6461 1026 6499
rect 980 6427 986 6461
rect 1020 6427 1026 6461
rect 980 6389 1026 6427
rect 980 6355 986 6389
rect 1020 6355 1026 6389
rect 980 6317 1026 6355
rect 980 6283 986 6317
rect 1020 6283 1026 6317
rect 980 6245 1026 6283
rect 980 6211 986 6245
rect 1020 6211 1026 6245
rect 980 6173 1026 6211
rect 980 6139 986 6173
rect 1020 6139 1026 6173
rect 980 6101 1026 6139
rect 980 6067 986 6101
rect 1020 6067 1026 6101
rect 980 6029 1026 6067
rect 980 5995 986 6029
rect 1020 5995 1026 6029
rect 980 5957 1026 5995
rect 980 5923 986 5957
rect 1020 5923 1026 5957
rect 980 5885 1026 5923
rect 980 5851 986 5885
rect 1020 5851 1026 5885
rect 980 5813 1026 5851
rect 980 5779 986 5813
rect 1020 5779 1026 5813
rect 980 5741 1026 5779
rect 980 5707 986 5741
rect 1020 5707 1026 5741
rect 980 5669 1026 5707
rect 980 5635 986 5669
rect 1020 5635 1026 5669
rect 980 5597 1026 5635
rect 980 5563 986 5597
rect 1020 5563 1026 5597
rect 980 5525 1026 5563
rect 980 5491 986 5525
rect 1020 5491 1026 5525
rect 980 5453 1026 5491
rect 980 5419 986 5453
rect 1020 5419 1026 5453
rect 980 5381 1026 5419
rect 980 5347 986 5381
rect 1020 5347 1026 5381
rect 980 5309 1026 5347
rect 980 5275 986 5309
rect 1020 5275 1026 5309
rect 980 5237 1026 5275
rect 980 5203 986 5237
rect 1020 5203 1026 5237
rect 980 5165 1026 5203
rect 980 5131 986 5165
rect 1020 5131 1026 5165
rect 980 5093 1026 5131
rect 980 5059 986 5093
rect 1020 5059 1026 5093
rect 980 5021 1026 5059
rect 980 4987 986 5021
rect 1020 4987 1026 5021
rect 980 4949 1026 4987
rect 980 4915 986 4949
rect 1020 4915 1026 4949
rect 980 4877 1026 4915
rect 980 4843 986 4877
rect 1020 4843 1026 4877
rect 980 4805 1026 4843
rect 980 4771 986 4805
rect 1020 4771 1026 4805
rect 980 4733 1026 4771
rect 980 4699 986 4733
rect 1020 4699 1026 4733
rect 980 4661 1026 4699
rect 980 4627 986 4661
rect 1020 4627 1026 4661
rect 980 4589 1026 4627
rect 980 4555 986 4589
rect 1020 4555 1026 4589
rect 980 4517 1026 4555
rect 980 4483 986 4517
rect 1020 4483 1026 4517
rect 980 4445 1026 4483
rect 980 4411 986 4445
rect 1020 4411 1026 4445
rect 980 4373 1026 4411
rect 980 4339 986 4373
rect 1020 4339 1026 4373
rect 980 4301 1026 4339
rect 980 4267 986 4301
rect 1020 4267 1026 4301
rect 980 4229 1026 4267
rect 980 4195 986 4229
rect 1020 4195 1026 4229
rect 980 4157 1026 4195
rect 980 4123 986 4157
rect 1020 4123 1026 4157
rect 980 4085 1026 4123
rect 980 4051 986 4085
rect 1020 4051 1026 4085
rect 980 4013 1026 4051
rect 980 3979 986 4013
rect 1020 3979 1026 4013
rect 980 3941 1026 3979
rect 980 3907 986 3941
rect 1020 3907 1026 3941
rect 980 3869 1026 3907
rect 980 3835 986 3869
rect 1020 3835 1026 3869
rect 980 3797 1026 3835
rect 980 3763 986 3797
rect 1020 3763 1026 3797
rect 980 3725 1026 3763
rect 980 3691 986 3725
rect 1020 3691 1026 3725
rect 980 3653 1026 3691
rect 980 3619 986 3653
rect 1020 3619 1026 3653
rect 980 3581 1026 3619
rect 980 3547 986 3581
rect 1020 3547 1026 3581
rect 980 3509 1026 3547
rect 980 3475 986 3509
rect 1020 3475 1026 3509
rect 980 3437 1026 3475
rect 980 3403 986 3437
rect 1020 3403 1026 3437
rect 980 3365 1026 3403
rect 980 3331 986 3365
rect 1020 3331 1026 3365
rect 980 3293 1026 3331
rect 980 3259 986 3293
rect 1020 3259 1026 3293
rect 980 3221 1026 3259
rect 980 3187 986 3221
rect 1020 3187 1026 3221
rect 980 3149 1026 3187
rect 980 3115 986 3149
rect 1020 3115 1026 3149
rect 980 3077 1026 3115
rect 980 3043 986 3077
rect 1020 3043 1026 3077
rect 980 3005 1026 3043
rect 980 2971 986 3005
rect 1020 2971 1026 3005
rect 980 2933 1026 2971
rect 980 2899 986 2933
rect 1020 2899 1026 2933
rect 980 2861 1026 2899
rect 980 2827 986 2861
rect 1020 2827 1026 2861
rect 980 2789 1026 2827
rect 980 2755 986 2789
rect 1020 2755 1026 2789
rect 980 2717 1026 2755
rect 980 2683 986 2717
rect 1020 2683 1026 2717
rect 980 2645 1026 2683
rect 980 2611 986 2645
rect 1020 2611 1026 2645
rect 980 2573 1026 2611
rect 980 2539 986 2573
rect 1020 2539 1026 2573
rect 980 2501 1026 2539
rect 980 2467 986 2501
rect 1020 2467 1026 2501
rect 980 2429 1026 2467
rect 980 2395 986 2429
rect 1020 2395 1026 2429
rect 980 2357 1026 2395
rect 980 2323 986 2357
rect 1020 2323 1026 2357
rect 980 2285 1026 2323
rect 980 2251 986 2285
rect 1020 2251 1026 2285
rect 980 2213 1026 2251
rect 980 2179 986 2213
rect 1020 2179 1026 2213
rect 980 2141 1026 2179
rect 980 2107 986 2141
rect 1020 2107 1026 2141
rect 980 2069 1026 2107
rect 980 2035 986 2069
rect 1020 2035 1026 2069
rect 980 1997 1026 2035
rect 980 1963 986 1997
rect 1020 1963 1026 1997
rect 980 1925 1026 1963
rect 980 1891 986 1925
rect 1020 1891 1026 1925
rect 980 1853 1026 1891
rect 980 1819 986 1853
rect 1020 1819 1026 1853
rect 980 1781 1026 1819
rect 980 1747 986 1781
rect 1020 1747 1026 1781
rect 980 1709 1026 1747
rect 980 1675 986 1709
rect 1020 1675 1026 1709
rect 980 1637 1026 1675
rect 980 1603 986 1637
rect 1020 1603 1026 1637
rect 980 1565 1026 1603
rect 980 1531 986 1565
rect 1020 1531 1026 1565
rect 980 1493 1026 1531
rect 980 1459 986 1493
rect 1020 1459 1026 1493
rect 980 1421 1026 1459
rect 980 1387 986 1421
rect 1020 1387 1026 1421
rect 980 1349 1026 1387
rect 980 1315 986 1349
rect 1020 1315 1026 1349
rect 980 1277 1026 1315
rect 980 1243 986 1277
rect 1020 1243 1026 1277
rect 980 1205 1026 1243
rect 980 1171 986 1205
rect 1020 1171 1026 1205
rect 980 1133 1026 1171
rect 980 1099 986 1133
rect 1020 1099 1026 1133
rect 980 1061 1026 1099
rect 980 1027 986 1061
rect 1020 1027 1026 1061
rect 980 989 1026 1027
rect 980 955 986 989
rect 1020 955 1026 989
rect 980 917 1026 955
rect 980 883 986 917
rect 1020 883 1026 917
rect 980 845 1026 883
rect 980 811 986 845
rect 1020 811 1026 845
rect 980 773 1026 811
rect 980 739 986 773
rect 1020 739 1026 773
rect 980 701 1026 739
rect 980 667 986 701
rect 1020 667 1026 701
rect 980 629 1026 667
rect 980 595 986 629
rect 1020 595 1026 629
rect 980 557 1026 595
rect 980 523 986 557
rect 1020 523 1026 557
rect 980 485 1026 523
rect 980 451 986 485
rect 1020 451 1026 485
rect 980 413 1026 451
rect 980 379 986 413
rect 1020 379 1026 413
rect 980 341 1026 379
rect 980 307 986 341
rect 1020 307 1026 341
rect 980 269 1026 307
rect 980 235 986 269
rect 1020 235 1026 269
rect 980 197 1026 235
rect 980 163 986 197
rect 1020 163 1026 197
rect 980 125 1026 163
rect 980 91 986 125
rect 1020 91 1026 125
rect 980 53 1026 91
rect 980 19 986 53
rect 1020 19 1026 53
rect 980 -19 1026 19
rect 980 -53 986 -19
rect 1020 -53 1026 -19
rect 980 -91 1026 -53
rect 980 -125 986 -91
rect 1020 -125 1026 -91
rect 980 -163 1026 -125
rect 980 -197 986 -163
rect 1020 -197 1026 -163
rect 980 -235 1026 -197
rect 980 -269 986 -235
rect 1020 -269 1026 -235
rect 980 -307 1026 -269
rect 980 -341 986 -307
rect 1020 -341 1026 -307
rect 980 -379 1026 -341
rect 980 -413 986 -379
rect 1020 -413 1026 -379
rect 980 -451 1026 -413
rect 980 -485 986 -451
rect 1020 -485 1026 -451
rect 980 -523 1026 -485
rect 980 -557 986 -523
rect 1020 -557 1026 -523
rect 980 -595 1026 -557
rect 980 -629 986 -595
rect 1020 -629 1026 -595
rect 980 -667 1026 -629
rect 980 -701 986 -667
rect 1020 -701 1026 -667
rect 980 -739 1026 -701
rect 980 -773 986 -739
rect 1020 -773 1026 -739
rect 980 -811 1026 -773
rect 980 -845 986 -811
rect 1020 -845 1026 -811
rect 980 -883 1026 -845
rect 980 -917 986 -883
rect 1020 -917 1026 -883
rect 980 -955 1026 -917
rect 980 -989 986 -955
rect 1020 -989 1026 -955
rect 980 -1027 1026 -989
rect 980 -1061 986 -1027
rect 1020 -1061 1026 -1027
rect 980 -1099 1026 -1061
rect 980 -1133 986 -1099
rect 1020 -1133 1026 -1099
rect 980 -1171 1026 -1133
rect 980 -1205 986 -1171
rect 1020 -1205 1026 -1171
rect 980 -1243 1026 -1205
rect 980 -1277 986 -1243
rect 1020 -1277 1026 -1243
rect 980 -1315 1026 -1277
rect 980 -1349 986 -1315
rect 1020 -1349 1026 -1315
rect 980 -1387 1026 -1349
rect 980 -1421 986 -1387
rect 1020 -1421 1026 -1387
rect 980 -1459 1026 -1421
rect 980 -1493 986 -1459
rect 1020 -1493 1026 -1459
rect 980 -1531 1026 -1493
rect 980 -1565 986 -1531
rect 1020 -1565 1026 -1531
rect 980 -1603 1026 -1565
rect 980 -1637 986 -1603
rect 1020 -1637 1026 -1603
rect 980 -1675 1026 -1637
rect 980 -1709 986 -1675
rect 1020 -1709 1026 -1675
rect 980 -1747 1026 -1709
rect 980 -1781 986 -1747
rect 1020 -1781 1026 -1747
rect 980 -1819 1026 -1781
rect 980 -1853 986 -1819
rect 1020 -1853 1026 -1819
rect 980 -1891 1026 -1853
rect 980 -1925 986 -1891
rect 1020 -1925 1026 -1891
rect 980 -1963 1026 -1925
rect 980 -1997 986 -1963
rect 1020 -1997 1026 -1963
rect 980 -2035 1026 -1997
rect 980 -2069 986 -2035
rect 1020 -2069 1026 -2035
rect 980 -2107 1026 -2069
rect 980 -2141 986 -2107
rect 1020 -2141 1026 -2107
rect 980 -2179 1026 -2141
rect 980 -2213 986 -2179
rect 1020 -2213 1026 -2179
rect 980 -2251 1026 -2213
rect 980 -2285 986 -2251
rect 1020 -2285 1026 -2251
rect 980 -2323 1026 -2285
rect 980 -2357 986 -2323
rect 1020 -2357 1026 -2323
rect 980 -2395 1026 -2357
rect 980 -2429 986 -2395
rect 1020 -2429 1026 -2395
rect 980 -2467 1026 -2429
rect 980 -2501 986 -2467
rect 1020 -2501 1026 -2467
rect 980 -2539 1026 -2501
rect 980 -2573 986 -2539
rect 1020 -2573 1026 -2539
rect 980 -2611 1026 -2573
rect 980 -2645 986 -2611
rect 1020 -2645 1026 -2611
rect 980 -2683 1026 -2645
rect 980 -2717 986 -2683
rect 1020 -2717 1026 -2683
rect 980 -2755 1026 -2717
rect 980 -2789 986 -2755
rect 1020 -2789 1026 -2755
rect 980 -2827 1026 -2789
rect 980 -2861 986 -2827
rect 1020 -2861 1026 -2827
rect 980 -2899 1026 -2861
rect 980 -2933 986 -2899
rect 1020 -2933 1026 -2899
rect 980 -2971 1026 -2933
rect 980 -3005 986 -2971
rect 1020 -3005 1026 -2971
rect 980 -3043 1026 -3005
rect 980 -3077 986 -3043
rect 1020 -3077 1026 -3043
rect 980 -3115 1026 -3077
rect 980 -3149 986 -3115
rect 1020 -3149 1026 -3115
rect 980 -3187 1026 -3149
rect 980 -3221 986 -3187
rect 1020 -3221 1026 -3187
rect 980 -3259 1026 -3221
rect 980 -3293 986 -3259
rect 1020 -3293 1026 -3259
rect 980 -3331 1026 -3293
rect 980 -3365 986 -3331
rect 1020 -3365 1026 -3331
rect 980 -3403 1026 -3365
rect 980 -3437 986 -3403
rect 1020 -3437 1026 -3403
rect 980 -3475 1026 -3437
rect 980 -3509 986 -3475
rect 1020 -3509 1026 -3475
rect 980 -3547 1026 -3509
rect 980 -3581 986 -3547
rect 1020 -3581 1026 -3547
rect 980 -3619 1026 -3581
rect 980 -3653 986 -3619
rect 1020 -3653 1026 -3619
rect 980 -3691 1026 -3653
rect 980 -3725 986 -3691
rect 1020 -3725 1026 -3691
rect 980 -3763 1026 -3725
rect 980 -3797 986 -3763
rect 1020 -3797 1026 -3763
rect 980 -3835 1026 -3797
rect 980 -3869 986 -3835
rect 1020 -3869 1026 -3835
rect 980 -3907 1026 -3869
rect 980 -3941 986 -3907
rect 1020 -3941 1026 -3907
rect 980 -3979 1026 -3941
rect 980 -4013 986 -3979
rect 1020 -4013 1026 -3979
rect 980 -4051 1026 -4013
rect 980 -4085 986 -4051
rect 1020 -4085 1026 -4051
rect 980 -4123 1026 -4085
rect 980 -4157 986 -4123
rect 1020 -4157 1026 -4123
rect 980 -4195 1026 -4157
rect 980 -4229 986 -4195
rect 1020 -4229 1026 -4195
rect 980 -4267 1026 -4229
rect 980 -4301 986 -4267
rect 1020 -4301 1026 -4267
rect 980 -4339 1026 -4301
rect 980 -4373 986 -4339
rect 1020 -4373 1026 -4339
rect 980 -4411 1026 -4373
rect 980 -4445 986 -4411
rect 1020 -4445 1026 -4411
rect 980 -4483 1026 -4445
rect 980 -4517 986 -4483
rect 1020 -4517 1026 -4483
rect 980 -4555 1026 -4517
rect 980 -4589 986 -4555
rect 1020 -4589 1026 -4555
rect 980 -4627 1026 -4589
rect 980 -4661 986 -4627
rect 1020 -4661 1026 -4627
rect 980 -4699 1026 -4661
rect 980 -4733 986 -4699
rect 1020 -4733 1026 -4699
rect 980 -4771 1026 -4733
rect 980 -4805 986 -4771
rect 1020 -4805 1026 -4771
rect 980 -4843 1026 -4805
rect 980 -4877 986 -4843
rect 1020 -4877 1026 -4843
rect 980 -4915 1026 -4877
rect 980 -4949 986 -4915
rect 1020 -4949 1026 -4915
rect 980 -4987 1026 -4949
rect 980 -5021 986 -4987
rect 1020 -5021 1026 -4987
rect 980 -5059 1026 -5021
rect 980 -5093 986 -5059
rect 1020 -5093 1026 -5059
rect 980 -5131 1026 -5093
rect 980 -5165 986 -5131
rect 1020 -5165 1026 -5131
rect 980 -5203 1026 -5165
rect 980 -5237 986 -5203
rect 1020 -5237 1026 -5203
rect 980 -5275 1026 -5237
rect 980 -5309 986 -5275
rect 1020 -5309 1026 -5275
rect 980 -5347 1026 -5309
rect 980 -5381 986 -5347
rect 1020 -5381 1026 -5347
rect 980 -5419 1026 -5381
rect 980 -5453 986 -5419
rect 1020 -5453 1026 -5419
rect 980 -5491 1026 -5453
rect 980 -5525 986 -5491
rect 1020 -5525 1026 -5491
rect 980 -5563 1026 -5525
rect 980 -5597 986 -5563
rect 1020 -5597 1026 -5563
rect 980 -5635 1026 -5597
rect 980 -5669 986 -5635
rect 1020 -5669 1026 -5635
rect 980 -5707 1026 -5669
rect 980 -5741 986 -5707
rect 1020 -5741 1026 -5707
rect 980 -5779 1026 -5741
rect 980 -5813 986 -5779
rect 1020 -5813 1026 -5779
rect 980 -5851 1026 -5813
rect 980 -5885 986 -5851
rect 1020 -5885 1026 -5851
rect 980 -5923 1026 -5885
rect 980 -5957 986 -5923
rect 1020 -5957 1026 -5923
rect 980 -5995 1026 -5957
rect 980 -6029 986 -5995
rect 1020 -6029 1026 -5995
rect 980 -6067 1026 -6029
rect 980 -6101 986 -6067
rect 1020 -6101 1026 -6067
rect 980 -6139 1026 -6101
rect 980 -6173 986 -6139
rect 1020 -6173 1026 -6139
rect 980 -6211 1026 -6173
rect 980 -6245 986 -6211
rect 1020 -6245 1026 -6211
rect 980 -6283 1026 -6245
rect 980 -6317 986 -6283
rect 1020 -6317 1026 -6283
rect 980 -6355 1026 -6317
rect 980 -6389 986 -6355
rect 1020 -6389 1026 -6355
rect 980 -6427 1026 -6389
rect 980 -6461 986 -6427
rect 1020 -6461 1026 -6427
rect 980 -6499 1026 -6461
rect 980 -6533 986 -6499
rect 1020 -6533 1026 -6499
rect 980 -6571 1026 -6533
rect 980 -6605 986 -6571
rect 1020 -6605 1026 -6571
rect 980 -6643 1026 -6605
rect 980 -6677 986 -6643
rect 1020 -6677 1026 -6643
rect 980 -6715 1026 -6677
rect 980 -6749 986 -6715
rect 1020 -6749 1026 -6715
rect 980 -6787 1026 -6749
rect 980 -6821 986 -6787
rect 1020 -6821 1026 -6787
rect 980 -6859 1026 -6821
rect 980 -6893 986 -6859
rect 1020 -6893 1026 -6859
rect 980 -6931 1026 -6893
rect 980 -6965 986 -6931
rect 1020 -6965 1026 -6931
rect 980 -7003 1026 -6965
rect 980 -7037 986 -7003
rect 1020 -7037 1026 -7003
rect 980 -7075 1026 -7037
rect 980 -7109 986 -7075
rect 1020 -7109 1026 -7075
rect 980 -7147 1026 -7109
rect 980 -7181 986 -7147
rect 1020 -7181 1026 -7147
rect 980 -7219 1026 -7181
rect 980 -7253 986 -7219
rect 1020 -7253 1026 -7219
rect 980 -7291 1026 -7253
rect 980 -7325 986 -7291
rect 1020 -7325 1026 -7291
rect 980 -7363 1026 -7325
rect 980 -7397 986 -7363
rect 1020 -7397 1026 -7363
rect 980 -7435 1026 -7397
rect 980 -7469 986 -7435
rect 1020 -7469 1026 -7435
rect 980 -7507 1026 -7469
rect 980 -7541 986 -7507
rect 1020 -7541 1026 -7507
rect 980 -7579 1026 -7541
rect 980 -7613 986 -7579
rect 1020 -7613 1026 -7579
rect 980 -7651 1026 -7613
rect 980 -7685 986 -7651
rect 1020 -7685 1026 -7651
rect 980 -7723 1026 -7685
rect 980 -7757 986 -7723
rect 1020 -7757 1026 -7723
rect 980 -7795 1026 -7757
rect 980 -7829 986 -7795
rect 1020 -7829 1026 -7795
rect 980 -7867 1026 -7829
rect 980 -7901 986 -7867
rect 1020 -7901 1026 -7867
rect 980 -7939 1026 -7901
rect 980 -7973 986 -7939
rect 1020 -7973 1026 -7939
rect 980 -8011 1026 -7973
rect 980 -8045 986 -8011
rect 1020 -8045 1026 -8011
rect 980 -8083 1026 -8045
rect 980 -8117 986 -8083
rect 1020 -8117 1026 -8083
rect 980 -8155 1026 -8117
rect 980 -8189 986 -8155
rect 1020 -8189 1026 -8155
rect 980 -8227 1026 -8189
rect 980 -8261 986 -8227
rect 1020 -8261 1026 -8227
rect 980 -8299 1026 -8261
rect 980 -8333 986 -8299
rect 1020 -8333 1026 -8299
rect 980 -8371 1026 -8333
rect 980 -8405 986 -8371
rect 1020 -8405 1026 -8371
rect 980 -8443 1026 -8405
rect 980 -8477 986 -8443
rect 1020 -8477 1026 -8443
rect 980 -8515 1026 -8477
rect 980 -8549 986 -8515
rect 1020 -8549 1026 -8515
rect 980 -8587 1026 -8549
rect 980 -8621 986 -8587
rect 1020 -8621 1026 -8587
rect 980 -8659 1026 -8621
rect 980 -8693 986 -8659
rect 1020 -8693 1026 -8659
rect 980 -8731 1026 -8693
rect 980 -8765 986 -8731
rect 1020 -8765 1026 -8731
rect 980 -8803 1026 -8765
rect 980 -8837 986 -8803
rect 1020 -8837 1026 -8803
rect 980 -8875 1026 -8837
rect 980 -8909 986 -8875
rect 1020 -8909 1026 -8875
rect 980 -8947 1026 -8909
rect 980 -8981 986 -8947
rect 1020 -8981 1026 -8947
rect 980 -9019 1026 -8981
rect 980 -9053 986 -9019
rect 1020 -9053 1026 -9019
rect 980 -9091 1026 -9053
rect 980 -9125 986 -9091
rect 1020 -9125 1026 -9091
rect 980 -9163 1026 -9125
rect 980 -9197 986 -9163
rect 1020 -9197 1026 -9163
rect 980 -9235 1026 -9197
rect 980 -9269 986 -9235
rect 1020 -9269 1026 -9235
rect 980 -9307 1026 -9269
rect 980 -9341 986 -9307
rect 1020 -9341 1026 -9307
rect 980 -9379 1026 -9341
rect 980 -9413 986 -9379
rect 1020 -9413 1026 -9379
rect 980 -9451 1026 -9413
rect 980 -9485 986 -9451
rect 1020 -9485 1026 -9451
rect 980 -9523 1026 -9485
rect 980 -9557 986 -9523
rect 1020 -9557 1026 -9523
rect 980 -9600 1026 -9557
rect 1098 9557 1144 9600
rect 1098 9523 1104 9557
rect 1138 9523 1144 9557
rect 1098 9485 1144 9523
rect 1098 9451 1104 9485
rect 1138 9451 1144 9485
rect 1098 9413 1144 9451
rect 1098 9379 1104 9413
rect 1138 9379 1144 9413
rect 1098 9341 1144 9379
rect 1098 9307 1104 9341
rect 1138 9307 1144 9341
rect 1098 9269 1144 9307
rect 1098 9235 1104 9269
rect 1138 9235 1144 9269
rect 1098 9197 1144 9235
rect 1098 9163 1104 9197
rect 1138 9163 1144 9197
rect 1098 9125 1144 9163
rect 1098 9091 1104 9125
rect 1138 9091 1144 9125
rect 1098 9053 1144 9091
rect 1098 9019 1104 9053
rect 1138 9019 1144 9053
rect 1098 8981 1144 9019
rect 1098 8947 1104 8981
rect 1138 8947 1144 8981
rect 1098 8909 1144 8947
rect 1098 8875 1104 8909
rect 1138 8875 1144 8909
rect 1098 8837 1144 8875
rect 1098 8803 1104 8837
rect 1138 8803 1144 8837
rect 1098 8765 1144 8803
rect 1098 8731 1104 8765
rect 1138 8731 1144 8765
rect 1098 8693 1144 8731
rect 1098 8659 1104 8693
rect 1138 8659 1144 8693
rect 1098 8621 1144 8659
rect 1098 8587 1104 8621
rect 1138 8587 1144 8621
rect 1098 8549 1144 8587
rect 1098 8515 1104 8549
rect 1138 8515 1144 8549
rect 1098 8477 1144 8515
rect 1098 8443 1104 8477
rect 1138 8443 1144 8477
rect 1098 8405 1144 8443
rect 1098 8371 1104 8405
rect 1138 8371 1144 8405
rect 1098 8333 1144 8371
rect 1098 8299 1104 8333
rect 1138 8299 1144 8333
rect 1098 8261 1144 8299
rect 1098 8227 1104 8261
rect 1138 8227 1144 8261
rect 1098 8189 1144 8227
rect 1098 8155 1104 8189
rect 1138 8155 1144 8189
rect 1098 8117 1144 8155
rect 1098 8083 1104 8117
rect 1138 8083 1144 8117
rect 1098 8045 1144 8083
rect 1098 8011 1104 8045
rect 1138 8011 1144 8045
rect 1098 7973 1144 8011
rect 1098 7939 1104 7973
rect 1138 7939 1144 7973
rect 1098 7901 1144 7939
rect 1098 7867 1104 7901
rect 1138 7867 1144 7901
rect 1098 7829 1144 7867
rect 1098 7795 1104 7829
rect 1138 7795 1144 7829
rect 1098 7757 1144 7795
rect 1098 7723 1104 7757
rect 1138 7723 1144 7757
rect 1098 7685 1144 7723
rect 1098 7651 1104 7685
rect 1138 7651 1144 7685
rect 1098 7613 1144 7651
rect 1098 7579 1104 7613
rect 1138 7579 1144 7613
rect 1098 7541 1144 7579
rect 1098 7507 1104 7541
rect 1138 7507 1144 7541
rect 1098 7469 1144 7507
rect 1098 7435 1104 7469
rect 1138 7435 1144 7469
rect 1098 7397 1144 7435
rect 1098 7363 1104 7397
rect 1138 7363 1144 7397
rect 1098 7325 1144 7363
rect 1098 7291 1104 7325
rect 1138 7291 1144 7325
rect 1098 7253 1144 7291
rect 1098 7219 1104 7253
rect 1138 7219 1144 7253
rect 1098 7181 1144 7219
rect 1098 7147 1104 7181
rect 1138 7147 1144 7181
rect 1098 7109 1144 7147
rect 1098 7075 1104 7109
rect 1138 7075 1144 7109
rect 1098 7037 1144 7075
rect 1098 7003 1104 7037
rect 1138 7003 1144 7037
rect 1098 6965 1144 7003
rect 1098 6931 1104 6965
rect 1138 6931 1144 6965
rect 1098 6893 1144 6931
rect 1098 6859 1104 6893
rect 1138 6859 1144 6893
rect 1098 6821 1144 6859
rect 1098 6787 1104 6821
rect 1138 6787 1144 6821
rect 1098 6749 1144 6787
rect 1098 6715 1104 6749
rect 1138 6715 1144 6749
rect 1098 6677 1144 6715
rect 1098 6643 1104 6677
rect 1138 6643 1144 6677
rect 1098 6605 1144 6643
rect 1098 6571 1104 6605
rect 1138 6571 1144 6605
rect 1098 6533 1144 6571
rect 1098 6499 1104 6533
rect 1138 6499 1144 6533
rect 1098 6461 1144 6499
rect 1098 6427 1104 6461
rect 1138 6427 1144 6461
rect 1098 6389 1144 6427
rect 1098 6355 1104 6389
rect 1138 6355 1144 6389
rect 1098 6317 1144 6355
rect 1098 6283 1104 6317
rect 1138 6283 1144 6317
rect 1098 6245 1144 6283
rect 1098 6211 1104 6245
rect 1138 6211 1144 6245
rect 1098 6173 1144 6211
rect 1098 6139 1104 6173
rect 1138 6139 1144 6173
rect 1098 6101 1144 6139
rect 1098 6067 1104 6101
rect 1138 6067 1144 6101
rect 1098 6029 1144 6067
rect 1098 5995 1104 6029
rect 1138 5995 1144 6029
rect 1098 5957 1144 5995
rect 1098 5923 1104 5957
rect 1138 5923 1144 5957
rect 1098 5885 1144 5923
rect 1098 5851 1104 5885
rect 1138 5851 1144 5885
rect 1098 5813 1144 5851
rect 1098 5779 1104 5813
rect 1138 5779 1144 5813
rect 1098 5741 1144 5779
rect 1098 5707 1104 5741
rect 1138 5707 1144 5741
rect 1098 5669 1144 5707
rect 1098 5635 1104 5669
rect 1138 5635 1144 5669
rect 1098 5597 1144 5635
rect 1098 5563 1104 5597
rect 1138 5563 1144 5597
rect 1098 5525 1144 5563
rect 1098 5491 1104 5525
rect 1138 5491 1144 5525
rect 1098 5453 1144 5491
rect 1098 5419 1104 5453
rect 1138 5419 1144 5453
rect 1098 5381 1144 5419
rect 1098 5347 1104 5381
rect 1138 5347 1144 5381
rect 1098 5309 1144 5347
rect 1098 5275 1104 5309
rect 1138 5275 1144 5309
rect 1098 5237 1144 5275
rect 1098 5203 1104 5237
rect 1138 5203 1144 5237
rect 1098 5165 1144 5203
rect 1098 5131 1104 5165
rect 1138 5131 1144 5165
rect 1098 5093 1144 5131
rect 1098 5059 1104 5093
rect 1138 5059 1144 5093
rect 1098 5021 1144 5059
rect 1098 4987 1104 5021
rect 1138 4987 1144 5021
rect 1098 4949 1144 4987
rect 1098 4915 1104 4949
rect 1138 4915 1144 4949
rect 1098 4877 1144 4915
rect 1098 4843 1104 4877
rect 1138 4843 1144 4877
rect 1098 4805 1144 4843
rect 1098 4771 1104 4805
rect 1138 4771 1144 4805
rect 1098 4733 1144 4771
rect 1098 4699 1104 4733
rect 1138 4699 1144 4733
rect 1098 4661 1144 4699
rect 1098 4627 1104 4661
rect 1138 4627 1144 4661
rect 1098 4589 1144 4627
rect 1098 4555 1104 4589
rect 1138 4555 1144 4589
rect 1098 4517 1144 4555
rect 1098 4483 1104 4517
rect 1138 4483 1144 4517
rect 1098 4445 1144 4483
rect 1098 4411 1104 4445
rect 1138 4411 1144 4445
rect 1098 4373 1144 4411
rect 1098 4339 1104 4373
rect 1138 4339 1144 4373
rect 1098 4301 1144 4339
rect 1098 4267 1104 4301
rect 1138 4267 1144 4301
rect 1098 4229 1144 4267
rect 1098 4195 1104 4229
rect 1138 4195 1144 4229
rect 1098 4157 1144 4195
rect 1098 4123 1104 4157
rect 1138 4123 1144 4157
rect 1098 4085 1144 4123
rect 1098 4051 1104 4085
rect 1138 4051 1144 4085
rect 1098 4013 1144 4051
rect 1098 3979 1104 4013
rect 1138 3979 1144 4013
rect 1098 3941 1144 3979
rect 1098 3907 1104 3941
rect 1138 3907 1144 3941
rect 1098 3869 1144 3907
rect 1098 3835 1104 3869
rect 1138 3835 1144 3869
rect 1098 3797 1144 3835
rect 1098 3763 1104 3797
rect 1138 3763 1144 3797
rect 1098 3725 1144 3763
rect 1098 3691 1104 3725
rect 1138 3691 1144 3725
rect 1098 3653 1144 3691
rect 1098 3619 1104 3653
rect 1138 3619 1144 3653
rect 1098 3581 1144 3619
rect 1098 3547 1104 3581
rect 1138 3547 1144 3581
rect 1098 3509 1144 3547
rect 1098 3475 1104 3509
rect 1138 3475 1144 3509
rect 1098 3437 1144 3475
rect 1098 3403 1104 3437
rect 1138 3403 1144 3437
rect 1098 3365 1144 3403
rect 1098 3331 1104 3365
rect 1138 3331 1144 3365
rect 1098 3293 1144 3331
rect 1098 3259 1104 3293
rect 1138 3259 1144 3293
rect 1098 3221 1144 3259
rect 1098 3187 1104 3221
rect 1138 3187 1144 3221
rect 1098 3149 1144 3187
rect 1098 3115 1104 3149
rect 1138 3115 1144 3149
rect 1098 3077 1144 3115
rect 1098 3043 1104 3077
rect 1138 3043 1144 3077
rect 1098 3005 1144 3043
rect 1098 2971 1104 3005
rect 1138 2971 1144 3005
rect 1098 2933 1144 2971
rect 1098 2899 1104 2933
rect 1138 2899 1144 2933
rect 1098 2861 1144 2899
rect 1098 2827 1104 2861
rect 1138 2827 1144 2861
rect 1098 2789 1144 2827
rect 1098 2755 1104 2789
rect 1138 2755 1144 2789
rect 1098 2717 1144 2755
rect 1098 2683 1104 2717
rect 1138 2683 1144 2717
rect 1098 2645 1144 2683
rect 1098 2611 1104 2645
rect 1138 2611 1144 2645
rect 1098 2573 1144 2611
rect 1098 2539 1104 2573
rect 1138 2539 1144 2573
rect 1098 2501 1144 2539
rect 1098 2467 1104 2501
rect 1138 2467 1144 2501
rect 1098 2429 1144 2467
rect 1098 2395 1104 2429
rect 1138 2395 1144 2429
rect 1098 2357 1144 2395
rect 1098 2323 1104 2357
rect 1138 2323 1144 2357
rect 1098 2285 1144 2323
rect 1098 2251 1104 2285
rect 1138 2251 1144 2285
rect 1098 2213 1144 2251
rect 1098 2179 1104 2213
rect 1138 2179 1144 2213
rect 1098 2141 1144 2179
rect 1098 2107 1104 2141
rect 1138 2107 1144 2141
rect 1098 2069 1144 2107
rect 1098 2035 1104 2069
rect 1138 2035 1144 2069
rect 1098 1997 1144 2035
rect 1098 1963 1104 1997
rect 1138 1963 1144 1997
rect 1098 1925 1144 1963
rect 1098 1891 1104 1925
rect 1138 1891 1144 1925
rect 1098 1853 1144 1891
rect 1098 1819 1104 1853
rect 1138 1819 1144 1853
rect 1098 1781 1144 1819
rect 1098 1747 1104 1781
rect 1138 1747 1144 1781
rect 1098 1709 1144 1747
rect 1098 1675 1104 1709
rect 1138 1675 1144 1709
rect 1098 1637 1144 1675
rect 1098 1603 1104 1637
rect 1138 1603 1144 1637
rect 1098 1565 1144 1603
rect 1098 1531 1104 1565
rect 1138 1531 1144 1565
rect 1098 1493 1144 1531
rect 1098 1459 1104 1493
rect 1138 1459 1144 1493
rect 1098 1421 1144 1459
rect 1098 1387 1104 1421
rect 1138 1387 1144 1421
rect 1098 1349 1144 1387
rect 1098 1315 1104 1349
rect 1138 1315 1144 1349
rect 1098 1277 1144 1315
rect 1098 1243 1104 1277
rect 1138 1243 1144 1277
rect 1098 1205 1144 1243
rect 1098 1171 1104 1205
rect 1138 1171 1144 1205
rect 1098 1133 1144 1171
rect 1098 1099 1104 1133
rect 1138 1099 1144 1133
rect 1098 1061 1144 1099
rect 1098 1027 1104 1061
rect 1138 1027 1144 1061
rect 1098 989 1144 1027
rect 1098 955 1104 989
rect 1138 955 1144 989
rect 1098 917 1144 955
rect 1098 883 1104 917
rect 1138 883 1144 917
rect 1098 845 1144 883
rect 1098 811 1104 845
rect 1138 811 1144 845
rect 1098 773 1144 811
rect 1098 739 1104 773
rect 1138 739 1144 773
rect 1098 701 1144 739
rect 1098 667 1104 701
rect 1138 667 1144 701
rect 1098 629 1144 667
rect 1098 595 1104 629
rect 1138 595 1144 629
rect 1098 557 1144 595
rect 1098 523 1104 557
rect 1138 523 1144 557
rect 1098 485 1144 523
rect 1098 451 1104 485
rect 1138 451 1144 485
rect 1098 413 1144 451
rect 1098 379 1104 413
rect 1138 379 1144 413
rect 1098 341 1144 379
rect 1098 307 1104 341
rect 1138 307 1144 341
rect 1098 269 1144 307
rect 1098 235 1104 269
rect 1138 235 1144 269
rect 1098 197 1144 235
rect 1098 163 1104 197
rect 1138 163 1144 197
rect 1098 125 1144 163
rect 1098 91 1104 125
rect 1138 91 1144 125
rect 1098 53 1144 91
rect 1098 19 1104 53
rect 1138 19 1144 53
rect 1098 -19 1144 19
rect 1098 -53 1104 -19
rect 1138 -53 1144 -19
rect 1098 -91 1144 -53
rect 1098 -125 1104 -91
rect 1138 -125 1144 -91
rect 1098 -163 1144 -125
rect 1098 -197 1104 -163
rect 1138 -197 1144 -163
rect 1098 -235 1144 -197
rect 1098 -269 1104 -235
rect 1138 -269 1144 -235
rect 1098 -307 1144 -269
rect 1098 -341 1104 -307
rect 1138 -341 1144 -307
rect 1098 -379 1144 -341
rect 1098 -413 1104 -379
rect 1138 -413 1144 -379
rect 1098 -451 1144 -413
rect 1098 -485 1104 -451
rect 1138 -485 1144 -451
rect 1098 -523 1144 -485
rect 1098 -557 1104 -523
rect 1138 -557 1144 -523
rect 1098 -595 1144 -557
rect 1098 -629 1104 -595
rect 1138 -629 1144 -595
rect 1098 -667 1144 -629
rect 1098 -701 1104 -667
rect 1138 -701 1144 -667
rect 1098 -739 1144 -701
rect 1098 -773 1104 -739
rect 1138 -773 1144 -739
rect 1098 -811 1144 -773
rect 1098 -845 1104 -811
rect 1138 -845 1144 -811
rect 1098 -883 1144 -845
rect 1098 -917 1104 -883
rect 1138 -917 1144 -883
rect 1098 -955 1144 -917
rect 1098 -989 1104 -955
rect 1138 -989 1144 -955
rect 1098 -1027 1144 -989
rect 1098 -1061 1104 -1027
rect 1138 -1061 1144 -1027
rect 1098 -1099 1144 -1061
rect 1098 -1133 1104 -1099
rect 1138 -1133 1144 -1099
rect 1098 -1171 1144 -1133
rect 1098 -1205 1104 -1171
rect 1138 -1205 1144 -1171
rect 1098 -1243 1144 -1205
rect 1098 -1277 1104 -1243
rect 1138 -1277 1144 -1243
rect 1098 -1315 1144 -1277
rect 1098 -1349 1104 -1315
rect 1138 -1349 1144 -1315
rect 1098 -1387 1144 -1349
rect 1098 -1421 1104 -1387
rect 1138 -1421 1144 -1387
rect 1098 -1459 1144 -1421
rect 1098 -1493 1104 -1459
rect 1138 -1493 1144 -1459
rect 1098 -1531 1144 -1493
rect 1098 -1565 1104 -1531
rect 1138 -1565 1144 -1531
rect 1098 -1603 1144 -1565
rect 1098 -1637 1104 -1603
rect 1138 -1637 1144 -1603
rect 1098 -1675 1144 -1637
rect 1098 -1709 1104 -1675
rect 1138 -1709 1144 -1675
rect 1098 -1747 1144 -1709
rect 1098 -1781 1104 -1747
rect 1138 -1781 1144 -1747
rect 1098 -1819 1144 -1781
rect 1098 -1853 1104 -1819
rect 1138 -1853 1144 -1819
rect 1098 -1891 1144 -1853
rect 1098 -1925 1104 -1891
rect 1138 -1925 1144 -1891
rect 1098 -1963 1144 -1925
rect 1098 -1997 1104 -1963
rect 1138 -1997 1144 -1963
rect 1098 -2035 1144 -1997
rect 1098 -2069 1104 -2035
rect 1138 -2069 1144 -2035
rect 1098 -2107 1144 -2069
rect 1098 -2141 1104 -2107
rect 1138 -2141 1144 -2107
rect 1098 -2179 1144 -2141
rect 1098 -2213 1104 -2179
rect 1138 -2213 1144 -2179
rect 1098 -2251 1144 -2213
rect 1098 -2285 1104 -2251
rect 1138 -2285 1144 -2251
rect 1098 -2323 1144 -2285
rect 1098 -2357 1104 -2323
rect 1138 -2357 1144 -2323
rect 1098 -2395 1144 -2357
rect 1098 -2429 1104 -2395
rect 1138 -2429 1144 -2395
rect 1098 -2467 1144 -2429
rect 1098 -2501 1104 -2467
rect 1138 -2501 1144 -2467
rect 1098 -2539 1144 -2501
rect 1098 -2573 1104 -2539
rect 1138 -2573 1144 -2539
rect 1098 -2611 1144 -2573
rect 1098 -2645 1104 -2611
rect 1138 -2645 1144 -2611
rect 1098 -2683 1144 -2645
rect 1098 -2717 1104 -2683
rect 1138 -2717 1144 -2683
rect 1098 -2755 1144 -2717
rect 1098 -2789 1104 -2755
rect 1138 -2789 1144 -2755
rect 1098 -2827 1144 -2789
rect 1098 -2861 1104 -2827
rect 1138 -2861 1144 -2827
rect 1098 -2899 1144 -2861
rect 1098 -2933 1104 -2899
rect 1138 -2933 1144 -2899
rect 1098 -2971 1144 -2933
rect 1098 -3005 1104 -2971
rect 1138 -3005 1144 -2971
rect 1098 -3043 1144 -3005
rect 1098 -3077 1104 -3043
rect 1138 -3077 1144 -3043
rect 1098 -3115 1144 -3077
rect 1098 -3149 1104 -3115
rect 1138 -3149 1144 -3115
rect 1098 -3187 1144 -3149
rect 1098 -3221 1104 -3187
rect 1138 -3221 1144 -3187
rect 1098 -3259 1144 -3221
rect 1098 -3293 1104 -3259
rect 1138 -3293 1144 -3259
rect 1098 -3331 1144 -3293
rect 1098 -3365 1104 -3331
rect 1138 -3365 1144 -3331
rect 1098 -3403 1144 -3365
rect 1098 -3437 1104 -3403
rect 1138 -3437 1144 -3403
rect 1098 -3475 1144 -3437
rect 1098 -3509 1104 -3475
rect 1138 -3509 1144 -3475
rect 1098 -3547 1144 -3509
rect 1098 -3581 1104 -3547
rect 1138 -3581 1144 -3547
rect 1098 -3619 1144 -3581
rect 1098 -3653 1104 -3619
rect 1138 -3653 1144 -3619
rect 1098 -3691 1144 -3653
rect 1098 -3725 1104 -3691
rect 1138 -3725 1144 -3691
rect 1098 -3763 1144 -3725
rect 1098 -3797 1104 -3763
rect 1138 -3797 1144 -3763
rect 1098 -3835 1144 -3797
rect 1098 -3869 1104 -3835
rect 1138 -3869 1144 -3835
rect 1098 -3907 1144 -3869
rect 1098 -3941 1104 -3907
rect 1138 -3941 1144 -3907
rect 1098 -3979 1144 -3941
rect 1098 -4013 1104 -3979
rect 1138 -4013 1144 -3979
rect 1098 -4051 1144 -4013
rect 1098 -4085 1104 -4051
rect 1138 -4085 1144 -4051
rect 1098 -4123 1144 -4085
rect 1098 -4157 1104 -4123
rect 1138 -4157 1144 -4123
rect 1098 -4195 1144 -4157
rect 1098 -4229 1104 -4195
rect 1138 -4229 1144 -4195
rect 1098 -4267 1144 -4229
rect 1098 -4301 1104 -4267
rect 1138 -4301 1144 -4267
rect 1098 -4339 1144 -4301
rect 1098 -4373 1104 -4339
rect 1138 -4373 1144 -4339
rect 1098 -4411 1144 -4373
rect 1098 -4445 1104 -4411
rect 1138 -4445 1144 -4411
rect 1098 -4483 1144 -4445
rect 1098 -4517 1104 -4483
rect 1138 -4517 1144 -4483
rect 1098 -4555 1144 -4517
rect 1098 -4589 1104 -4555
rect 1138 -4589 1144 -4555
rect 1098 -4627 1144 -4589
rect 1098 -4661 1104 -4627
rect 1138 -4661 1144 -4627
rect 1098 -4699 1144 -4661
rect 1098 -4733 1104 -4699
rect 1138 -4733 1144 -4699
rect 1098 -4771 1144 -4733
rect 1098 -4805 1104 -4771
rect 1138 -4805 1144 -4771
rect 1098 -4843 1144 -4805
rect 1098 -4877 1104 -4843
rect 1138 -4877 1144 -4843
rect 1098 -4915 1144 -4877
rect 1098 -4949 1104 -4915
rect 1138 -4949 1144 -4915
rect 1098 -4987 1144 -4949
rect 1098 -5021 1104 -4987
rect 1138 -5021 1144 -4987
rect 1098 -5059 1144 -5021
rect 1098 -5093 1104 -5059
rect 1138 -5093 1144 -5059
rect 1098 -5131 1144 -5093
rect 1098 -5165 1104 -5131
rect 1138 -5165 1144 -5131
rect 1098 -5203 1144 -5165
rect 1098 -5237 1104 -5203
rect 1138 -5237 1144 -5203
rect 1098 -5275 1144 -5237
rect 1098 -5309 1104 -5275
rect 1138 -5309 1144 -5275
rect 1098 -5347 1144 -5309
rect 1098 -5381 1104 -5347
rect 1138 -5381 1144 -5347
rect 1098 -5419 1144 -5381
rect 1098 -5453 1104 -5419
rect 1138 -5453 1144 -5419
rect 1098 -5491 1144 -5453
rect 1098 -5525 1104 -5491
rect 1138 -5525 1144 -5491
rect 1098 -5563 1144 -5525
rect 1098 -5597 1104 -5563
rect 1138 -5597 1144 -5563
rect 1098 -5635 1144 -5597
rect 1098 -5669 1104 -5635
rect 1138 -5669 1144 -5635
rect 1098 -5707 1144 -5669
rect 1098 -5741 1104 -5707
rect 1138 -5741 1144 -5707
rect 1098 -5779 1144 -5741
rect 1098 -5813 1104 -5779
rect 1138 -5813 1144 -5779
rect 1098 -5851 1144 -5813
rect 1098 -5885 1104 -5851
rect 1138 -5885 1144 -5851
rect 1098 -5923 1144 -5885
rect 1098 -5957 1104 -5923
rect 1138 -5957 1144 -5923
rect 1098 -5995 1144 -5957
rect 1098 -6029 1104 -5995
rect 1138 -6029 1144 -5995
rect 1098 -6067 1144 -6029
rect 1098 -6101 1104 -6067
rect 1138 -6101 1144 -6067
rect 1098 -6139 1144 -6101
rect 1098 -6173 1104 -6139
rect 1138 -6173 1144 -6139
rect 1098 -6211 1144 -6173
rect 1098 -6245 1104 -6211
rect 1138 -6245 1144 -6211
rect 1098 -6283 1144 -6245
rect 1098 -6317 1104 -6283
rect 1138 -6317 1144 -6283
rect 1098 -6355 1144 -6317
rect 1098 -6389 1104 -6355
rect 1138 -6389 1144 -6355
rect 1098 -6427 1144 -6389
rect 1098 -6461 1104 -6427
rect 1138 -6461 1144 -6427
rect 1098 -6499 1144 -6461
rect 1098 -6533 1104 -6499
rect 1138 -6533 1144 -6499
rect 1098 -6571 1144 -6533
rect 1098 -6605 1104 -6571
rect 1138 -6605 1144 -6571
rect 1098 -6643 1144 -6605
rect 1098 -6677 1104 -6643
rect 1138 -6677 1144 -6643
rect 1098 -6715 1144 -6677
rect 1098 -6749 1104 -6715
rect 1138 -6749 1144 -6715
rect 1098 -6787 1144 -6749
rect 1098 -6821 1104 -6787
rect 1138 -6821 1144 -6787
rect 1098 -6859 1144 -6821
rect 1098 -6893 1104 -6859
rect 1138 -6893 1144 -6859
rect 1098 -6931 1144 -6893
rect 1098 -6965 1104 -6931
rect 1138 -6965 1144 -6931
rect 1098 -7003 1144 -6965
rect 1098 -7037 1104 -7003
rect 1138 -7037 1144 -7003
rect 1098 -7075 1144 -7037
rect 1098 -7109 1104 -7075
rect 1138 -7109 1144 -7075
rect 1098 -7147 1144 -7109
rect 1098 -7181 1104 -7147
rect 1138 -7181 1144 -7147
rect 1098 -7219 1144 -7181
rect 1098 -7253 1104 -7219
rect 1138 -7253 1144 -7219
rect 1098 -7291 1144 -7253
rect 1098 -7325 1104 -7291
rect 1138 -7325 1144 -7291
rect 1098 -7363 1144 -7325
rect 1098 -7397 1104 -7363
rect 1138 -7397 1144 -7363
rect 1098 -7435 1144 -7397
rect 1098 -7469 1104 -7435
rect 1138 -7469 1144 -7435
rect 1098 -7507 1144 -7469
rect 1098 -7541 1104 -7507
rect 1138 -7541 1144 -7507
rect 1098 -7579 1144 -7541
rect 1098 -7613 1104 -7579
rect 1138 -7613 1144 -7579
rect 1098 -7651 1144 -7613
rect 1098 -7685 1104 -7651
rect 1138 -7685 1144 -7651
rect 1098 -7723 1144 -7685
rect 1098 -7757 1104 -7723
rect 1138 -7757 1144 -7723
rect 1098 -7795 1144 -7757
rect 1098 -7829 1104 -7795
rect 1138 -7829 1144 -7795
rect 1098 -7867 1144 -7829
rect 1098 -7901 1104 -7867
rect 1138 -7901 1144 -7867
rect 1098 -7939 1144 -7901
rect 1098 -7973 1104 -7939
rect 1138 -7973 1144 -7939
rect 1098 -8011 1144 -7973
rect 1098 -8045 1104 -8011
rect 1138 -8045 1144 -8011
rect 1098 -8083 1144 -8045
rect 1098 -8117 1104 -8083
rect 1138 -8117 1144 -8083
rect 1098 -8155 1144 -8117
rect 1098 -8189 1104 -8155
rect 1138 -8189 1144 -8155
rect 1098 -8227 1144 -8189
rect 1098 -8261 1104 -8227
rect 1138 -8261 1144 -8227
rect 1098 -8299 1144 -8261
rect 1098 -8333 1104 -8299
rect 1138 -8333 1144 -8299
rect 1098 -8371 1144 -8333
rect 1098 -8405 1104 -8371
rect 1138 -8405 1144 -8371
rect 1098 -8443 1144 -8405
rect 1098 -8477 1104 -8443
rect 1138 -8477 1144 -8443
rect 1098 -8515 1144 -8477
rect 1098 -8549 1104 -8515
rect 1138 -8549 1144 -8515
rect 1098 -8587 1144 -8549
rect 1098 -8621 1104 -8587
rect 1138 -8621 1144 -8587
rect 1098 -8659 1144 -8621
rect 1098 -8693 1104 -8659
rect 1138 -8693 1144 -8659
rect 1098 -8731 1144 -8693
rect 1098 -8765 1104 -8731
rect 1138 -8765 1144 -8731
rect 1098 -8803 1144 -8765
rect 1098 -8837 1104 -8803
rect 1138 -8837 1144 -8803
rect 1098 -8875 1144 -8837
rect 1098 -8909 1104 -8875
rect 1138 -8909 1144 -8875
rect 1098 -8947 1144 -8909
rect 1098 -8981 1104 -8947
rect 1138 -8981 1144 -8947
rect 1098 -9019 1144 -8981
rect 1098 -9053 1104 -9019
rect 1138 -9053 1144 -9019
rect 1098 -9091 1144 -9053
rect 1098 -9125 1104 -9091
rect 1138 -9125 1144 -9091
rect 1098 -9163 1144 -9125
rect 1098 -9197 1104 -9163
rect 1138 -9197 1144 -9163
rect 1098 -9235 1144 -9197
rect 1098 -9269 1104 -9235
rect 1138 -9269 1144 -9235
rect 1098 -9307 1144 -9269
rect 1098 -9341 1104 -9307
rect 1138 -9341 1144 -9307
rect 1098 -9379 1144 -9341
rect 1098 -9413 1104 -9379
rect 1138 -9413 1144 -9379
rect 1098 -9451 1144 -9413
rect 1098 -9485 1104 -9451
rect 1138 -9485 1144 -9451
rect 1098 -9523 1144 -9485
rect 1098 -9557 1104 -9523
rect 1138 -9557 1144 -9523
rect 1098 -9600 1144 -9557
rect 1216 9557 1262 9600
rect 1216 9523 1222 9557
rect 1256 9523 1262 9557
rect 1216 9485 1262 9523
rect 1216 9451 1222 9485
rect 1256 9451 1262 9485
rect 1216 9413 1262 9451
rect 1216 9379 1222 9413
rect 1256 9379 1262 9413
rect 1216 9341 1262 9379
rect 1216 9307 1222 9341
rect 1256 9307 1262 9341
rect 1216 9269 1262 9307
rect 1216 9235 1222 9269
rect 1256 9235 1262 9269
rect 1216 9197 1262 9235
rect 1216 9163 1222 9197
rect 1256 9163 1262 9197
rect 1216 9125 1262 9163
rect 1216 9091 1222 9125
rect 1256 9091 1262 9125
rect 1216 9053 1262 9091
rect 1216 9019 1222 9053
rect 1256 9019 1262 9053
rect 1216 8981 1262 9019
rect 1216 8947 1222 8981
rect 1256 8947 1262 8981
rect 1216 8909 1262 8947
rect 1216 8875 1222 8909
rect 1256 8875 1262 8909
rect 1216 8837 1262 8875
rect 1216 8803 1222 8837
rect 1256 8803 1262 8837
rect 1216 8765 1262 8803
rect 1216 8731 1222 8765
rect 1256 8731 1262 8765
rect 1216 8693 1262 8731
rect 1216 8659 1222 8693
rect 1256 8659 1262 8693
rect 1216 8621 1262 8659
rect 1216 8587 1222 8621
rect 1256 8587 1262 8621
rect 1216 8549 1262 8587
rect 1216 8515 1222 8549
rect 1256 8515 1262 8549
rect 1216 8477 1262 8515
rect 1216 8443 1222 8477
rect 1256 8443 1262 8477
rect 1216 8405 1262 8443
rect 1216 8371 1222 8405
rect 1256 8371 1262 8405
rect 1216 8333 1262 8371
rect 1216 8299 1222 8333
rect 1256 8299 1262 8333
rect 1216 8261 1262 8299
rect 1216 8227 1222 8261
rect 1256 8227 1262 8261
rect 1216 8189 1262 8227
rect 1216 8155 1222 8189
rect 1256 8155 1262 8189
rect 1216 8117 1262 8155
rect 1216 8083 1222 8117
rect 1256 8083 1262 8117
rect 1216 8045 1262 8083
rect 1216 8011 1222 8045
rect 1256 8011 1262 8045
rect 1216 7973 1262 8011
rect 1216 7939 1222 7973
rect 1256 7939 1262 7973
rect 1216 7901 1262 7939
rect 1216 7867 1222 7901
rect 1256 7867 1262 7901
rect 1216 7829 1262 7867
rect 1216 7795 1222 7829
rect 1256 7795 1262 7829
rect 1216 7757 1262 7795
rect 1216 7723 1222 7757
rect 1256 7723 1262 7757
rect 1216 7685 1262 7723
rect 1216 7651 1222 7685
rect 1256 7651 1262 7685
rect 1216 7613 1262 7651
rect 1216 7579 1222 7613
rect 1256 7579 1262 7613
rect 1216 7541 1262 7579
rect 1216 7507 1222 7541
rect 1256 7507 1262 7541
rect 1216 7469 1262 7507
rect 1216 7435 1222 7469
rect 1256 7435 1262 7469
rect 1216 7397 1262 7435
rect 1216 7363 1222 7397
rect 1256 7363 1262 7397
rect 1216 7325 1262 7363
rect 1216 7291 1222 7325
rect 1256 7291 1262 7325
rect 1216 7253 1262 7291
rect 1216 7219 1222 7253
rect 1256 7219 1262 7253
rect 1216 7181 1262 7219
rect 1216 7147 1222 7181
rect 1256 7147 1262 7181
rect 1216 7109 1262 7147
rect 1216 7075 1222 7109
rect 1256 7075 1262 7109
rect 1216 7037 1262 7075
rect 1216 7003 1222 7037
rect 1256 7003 1262 7037
rect 1216 6965 1262 7003
rect 1216 6931 1222 6965
rect 1256 6931 1262 6965
rect 1216 6893 1262 6931
rect 1216 6859 1222 6893
rect 1256 6859 1262 6893
rect 1216 6821 1262 6859
rect 1216 6787 1222 6821
rect 1256 6787 1262 6821
rect 1216 6749 1262 6787
rect 1216 6715 1222 6749
rect 1256 6715 1262 6749
rect 1216 6677 1262 6715
rect 1216 6643 1222 6677
rect 1256 6643 1262 6677
rect 1216 6605 1262 6643
rect 1216 6571 1222 6605
rect 1256 6571 1262 6605
rect 1216 6533 1262 6571
rect 1216 6499 1222 6533
rect 1256 6499 1262 6533
rect 1216 6461 1262 6499
rect 1216 6427 1222 6461
rect 1256 6427 1262 6461
rect 1216 6389 1262 6427
rect 1216 6355 1222 6389
rect 1256 6355 1262 6389
rect 1216 6317 1262 6355
rect 1216 6283 1222 6317
rect 1256 6283 1262 6317
rect 1216 6245 1262 6283
rect 1216 6211 1222 6245
rect 1256 6211 1262 6245
rect 1216 6173 1262 6211
rect 1216 6139 1222 6173
rect 1256 6139 1262 6173
rect 1216 6101 1262 6139
rect 1216 6067 1222 6101
rect 1256 6067 1262 6101
rect 1216 6029 1262 6067
rect 1216 5995 1222 6029
rect 1256 5995 1262 6029
rect 1216 5957 1262 5995
rect 1216 5923 1222 5957
rect 1256 5923 1262 5957
rect 1216 5885 1262 5923
rect 1216 5851 1222 5885
rect 1256 5851 1262 5885
rect 1216 5813 1262 5851
rect 1216 5779 1222 5813
rect 1256 5779 1262 5813
rect 1216 5741 1262 5779
rect 1216 5707 1222 5741
rect 1256 5707 1262 5741
rect 1216 5669 1262 5707
rect 1216 5635 1222 5669
rect 1256 5635 1262 5669
rect 1216 5597 1262 5635
rect 1216 5563 1222 5597
rect 1256 5563 1262 5597
rect 1216 5525 1262 5563
rect 1216 5491 1222 5525
rect 1256 5491 1262 5525
rect 1216 5453 1262 5491
rect 1216 5419 1222 5453
rect 1256 5419 1262 5453
rect 1216 5381 1262 5419
rect 1216 5347 1222 5381
rect 1256 5347 1262 5381
rect 1216 5309 1262 5347
rect 1216 5275 1222 5309
rect 1256 5275 1262 5309
rect 1216 5237 1262 5275
rect 1216 5203 1222 5237
rect 1256 5203 1262 5237
rect 1216 5165 1262 5203
rect 1216 5131 1222 5165
rect 1256 5131 1262 5165
rect 1216 5093 1262 5131
rect 1216 5059 1222 5093
rect 1256 5059 1262 5093
rect 1216 5021 1262 5059
rect 1216 4987 1222 5021
rect 1256 4987 1262 5021
rect 1216 4949 1262 4987
rect 1216 4915 1222 4949
rect 1256 4915 1262 4949
rect 1216 4877 1262 4915
rect 1216 4843 1222 4877
rect 1256 4843 1262 4877
rect 1216 4805 1262 4843
rect 1216 4771 1222 4805
rect 1256 4771 1262 4805
rect 1216 4733 1262 4771
rect 1216 4699 1222 4733
rect 1256 4699 1262 4733
rect 1216 4661 1262 4699
rect 1216 4627 1222 4661
rect 1256 4627 1262 4661
rect 1216 4589 1262 4627
rect 1216 4555 1222 4589
rect 1256 4555 1262 4589
rect 1216 4517 1262 4555
rect 1216 4483 1222 4517
rect 1256 4483 1262 4517
rect 1216 4445 1262 4483
rect 1216 4411 1222 4445
rect 1256 4411 1262 4445
rect 1216 4373 1262 4411
rect 1216 4339 1222 4373
rect 1256 4339 1262 4373
rect 1216 4301 1262 4339
rect 1216 4267 1222 4301
rect 1256 4267 1262 4301
rect 1216 4229 1262 4267
rect 1216 4195 1222 4229
rect 1256 4195 1262 4229
rect 1216 4157 1262 4195
rect 1216 4123 1222 4157
rect 1256 4123 1262 4157
rect 1216 4085 1262 4123
rect 1216 4051 1222 4085
rect 1256 4051 1262 4085
rect 1216 4013 1262 4051
rect 1216 3979 1222 4013
rect 1256 3979 1262 4013
rect 1216 3941 1262 3979
rect 1216 3907 1222 3941
rect 1256 3907 1262 3941
rect 1216 3869 1262 3907
rect 1216 3835 1222 3869
rect 1256 3835 1262 3869
rect 1216 3797 1262 3835
rect 1216 3763 1222 3797
rect 1256 3763 1262 3797
rect 1216 3725 1262 3763
rect 1216 3691 1222 3725
rect 1256 3691 1262 3725
rect 1216 3653 1262 3691
rect 1216 3619 1222 3653
rect 1256 3619 1262 3653
rect 1216 3581 1262 3619
rect 1216 3547 1222 3581
rect 1256 3547 1262 3581
rect 1216 3509 1262 3547
rect 1216 3475 1222 3509
rect 1256 3475 1262 3509
rect 1216 3437 1262 3475
rect 1216 3403 1222 3437
rect 1256 3403 1262 3437
rect 1216 3365 1262 3403
rect 1216 3331 1222 3365
rect 1256 3331 1262 3365
rect 1216 3293 1262 3331
rect 1216 3259 1222 3293
rect 1256 3259 1262 3293
rect 1216 3221 1262 3259
rect 1216 3187 1222 3221
rect 1256 3187 1262 3221
rect 1216 3149 1262 3187
rect 1216 3115 1222 3149
rect 1256 3115 1262 3149
rect 1216 3077 1262 3115
rect 1216 3043 1222 3077
rect 1256 3043 1262 3077
rect 1216 3005 1262 3043
rect 1216 2971 1222 3005
rect 1256 2971 1262 3005
rect 1216 2933 1262 2971
rect 1216 2899 1222 2933
rect 1256 2899 1262 2933
rect 1216 2861 1262 2899
rect 1216 2827 1222 2861
rect 1256 2827 1262 2861
rect 1216 2789 1262 2827
rect 1216 2755 1222 2789
rect 1256 2755 1262 2789
rect 1216 2717 1262 2755
rect 1216 2683 1222 2717
rect 1256 2683 1262 2717
rect 1216 2645 1262 2683
rect 1216 2611 1222 2645
rect 1256 2611 1262 2645
rect 1216 2573 1262 2611
rect 1216 2539 1222 2573
rect 1256 2539 1262 2573
rect 1216 2501 1262 2539
rect 1216 2467 1222 2501
rect 1256 2467 1262 2501
rect 1216 2429 1262 2467
rect 1216 2395 1222 2429
rect 1256 2395 1262 2429
rect 1216 2357 1262 2395
rect 1216 2323 1222 2357
rect 1256 2323 1262 2357
rect 1216 2285 1262 2323
rect 1216 2251 1222 2285
rect 1256 2251 1262 2285
rect 1216 2213 1262 2251
rect 1216 2179 1222 2213
rect 1256 2179 1262 2213
rect 1216 2141 1262 2179
rect 1216 2107 1222 2141
rect 1256 2107 1262 2141
rect 1216 2069 1262 2107
rect 1216 2035 1222 2069
rect 1256 2035 1262 2069
rect 1216 1997 1262 2035
rect 1216 1963 1222 1997
rect 1256 1963 1262 1997
rect 1216 1925 1262 1963
rect 1216 1891 1222 1925
rect 1256 1891 1262 1925
rect 1216 1853 1262 1891
rect 1216 1819 1222 1853
rect 1256 1819 1262 1853
rect 1216 1781 1262 1819
rect 1216 1747 1222 1781
rect 1256 1747 1262 1781
rect 1216 1709 1262 1747
rect 1216 1675 1222 1709
rect 1256 1675 1262 1709
rect 1216 1637 1262 1675
rect 1216 1603 1222 1637
rect 1256 1603 1262 1637
rect 1216 1565 1262 1603
rect 1216 1531 1222 1565
rect 1256 1531 1262 1565
rect 1216 1493 1262 1531
rect 1216 1459 1222 1493
rect 1256 1459 1262 1493
rect 1216 1421 1262 1459
rect 1216 1387 1222 1421
rect 1256 1387 1262 1421
rect 1216 1349 1262 1387
rect 1216 1315 1222 1349
rect 1256 1315 1262 1349
rect 1216 1277 1262 1315
rect 1216 1243 1222 1277
rect 1256 1243 1262 1277
rect 1216 1205 1262 1243
rect 1216 1171 1222 1205
rect 1256 1171 1262 1205
rect 1216 1133 1262 1171
rect 1216 1099 1222 1133
rect 1256 1099 1262 1133
rect 1216 1061 1262 1099
rect 1216 1027 1222 1061
rect 1256 1027 1262 1061
rect 1216 989 1262 1027
rect 1216 955 1222 989
rect 1256 955 1262 989
rect 1216 917 1262 955
rect 1216 883 1222 917
rect 1256 883 1262 917
rect 1216 845 1262 883
rect 1216 811 1222 845
rect 1256 811 1262 845
rect 1216 773 1262 811
rect 1216 739 1222 773
rect 1256 739 1262 773
rect 1216 701 1262 739
rect 1216 667 1222 701
rect 1256 667 1262 701
rect 1216 629 1262 667
rect 1216 595 1222 629
rect 1256 595 1262 629
rect 1216 557 1262 595
rect 1216 523 1222 557
rect 1256 523 1262 557
rect 1216 485 1262 523
rect 1216 451 1222 485
rect 1256 451 1262 485
rect 1216 413 1262 451
rect 1216 379 1222 413
rect 1256 379 1262 413
rect 1216 341 1262 379
rect 1216 307 1222 341
rect 1256 307 1262 341
rect 1216 269 1262 307
rect 1216 235 1222 269
rect 1256 235 1262 269
rect 1216 197 1262 235
rect 1216 163 1222 197
rect 1256 163 1262 197
rect 1216 125 1262 163
rect 1216 91 1222 125
rect 1256 91 1262 125
rect 1216 53 1262 91
rect 1216 19 1222 53
rect 1256 19 1262 53
rect 1216 -19 1262 19
rect 1216 -53 1222 -19
rect 1256 -53 1262 -19
rect 1216 -91 1262 -53
rect 1216 -125 1222 -91
rect 1256 -125 1262 -91
rect 1216 -163 1262 -125
rect 1216 -197 1222 -163
rect 1256 -197 1262 -163
rect 1216 -235 1262 -197
rect 1216 -269 1222 -235
rect 1256 -269 1262 -235
rect 1216 -307 1262 -269
rect 1216 -341 1222 -307
rect 1256 -341 1262 -307
rect 1216 -379 1262 -341
rect 1216 -413 1222 -379
rect 1256 -413 1262 -379
rect 1216 -451 1262 -413
rect 1216 -485 1222 -451
rect 1256 -485 1262 -451
rect 1216 -523 1262 -485
rect 1216 -557 1222 -523
rect 1256 -557 1262 -523
rect 1216 -595 1262 -557
rect 1216 -629 1222 -595
rect 1256 -629 1262 -595
rect 1216 -667 1262 -629
rect 1216 -701 1222 -667
rect 1256 -701 1262 -667
rect 1216 -739 1262 -701
rect 1216 -773 1222 -739
rect 1256 -773 1262 -739
rect 1216 -811 1262 -773
rect 1216 -845 1222 -811
rect 1256 -845 1262 -811
rect 1216 -883 1262 -845
rect 1216 -917 1222 -883
rect 1256 -917 1262 -883
rect 1216 -955 1262 -917
rect 1216 -989 1222 -955
rect 1256 -989 1262 -955
rect 1216 -1027 1262 -989
rect 1216 -1061 1222 -1027
rect 1256 -1061 1262 -1027
rect 1216 -1099 1262 -1061
rect 1216 -1133 1222 -1099
rect 1256 -1133 1262 -1099
rect 1216 -1171 1262 -1133
rect 1216 -1205 1222 -1171
rect 1256 -1205 1262 -1171
rect 1216 -1243 1262 -1205
rect 1216 -1277 1222 -1243
rect 1256 -1277 1262 -1243
rect 1216 -1315 1262 -1277
rect 1216 -1349 1222 -1315
rect 1256 -1349 1262 -1315
rect 1216 -1387 1262 -1349
rect 1216 -1421 1222 -1387
rect 1256 -1421 1262 -1387
rect 1216 -1459 1262 -1421
rect 1216 -1493 1222 -1459
rect 1256 -1493 1262 -1459
rect 1216 -1531 1262 -1493
rect 1216 -1565 1222 -1531
rect 1256 -1565 1262 -1531
rect 1216 -1603 1262 -1565
rect 1216 -1637 1222 -1603
rect 1256 -1637 1262 -1603
rect 1216 -1675 1262 -1637
rect 1216 -1709 1222 -1675
rect 1256 -1709 1262 -1675
rect 1216 -1747 1262 -1709
rect 1216 -1781 1222 -1747
rect 1256 -1781 1262 -1747
rect 1216 -1819 1262 -1781
rect 1216 -1853 1222 -1819
rect 1256 -1853 1262 -1819
rect 1216 -1891 1262 -1853
rect 1216 -1925 1222 -1891
rect 1256 -1925 1262 -1891
rect 1216 -1963 1262 -1925
rect 1216 -1997 1222 -1963
rect 1256 -1997 1262 -1963
rect 1216 -2035 1262 -1997
rect 1216 -2069 1222 -2035
rect 1256 -2069 1262 -2035
rect 1216 -2107 1262 -2069
rect 1216 -2141 1222 -2107
rect 1256 -2141 1262 -2107
rect 1216 -2179 1262 -2141
rect 1216 -2213 1222 -2179
rect 1256 -2213 1262 -2179
rect 1216 -2251 1262 -2213
rect 1216 -2285 1222 -2251
rect 1256 -2285 1262 -2251
rect 1216 -2323 1262 -2285
rect 1216 -2357 1222 -2323
rect 1256 -2357 1262 -2323
rect 1216 -2395 1262 -2357
rect 1216 -2429 1222 -2395
rect 1256 -2429 1262 -2395
rect 1216 -2467 1262 -2429
rect 1216 -2501 1222 -2467
rect 1256 -2501 1262 -2467
rect 1216 -2539 1262 -2501
rect 1216 -2573 1222 -2539
rect 1256 -2573 1262 -2539
rect 1216 -2611 1262 -2573
rect 1216 -2645 1222 -2611
rect 1256 -2645 1262 -2611
rect 1216 -2683 1262 -2645
rect 1216 -2717 1222 -2683
rect 1256 -2717 1262 -2683
rect 1216 -2755 1262 -2717
rect 1216 -2789 1222 -2755
rect 1256 -2789 1262 -2755
rect 1216 -2827 1262 -2789
rect 1216 -2861 1222 -2827
rect 1256 -2861 1262 -2827
rect 1216 -2899 1262 -2861
rect 1216 -2933 1222 -2899
rect 1256 -2933 1262 -2899
rect 1216 -2971 1262 -2933
rect 1216 -3005 1222 -2971
rect 1256 -3005 1262 -2971
rect 1216 -3043 1262 -3005
rect 1216 -3077 1222 -3043
rect 1256 -3077 1262 -3043
rect 1216 -3115 1262 -3077
rect 1216 -3149 1222 -3115
rect 1256 -3149 1262 -3115
rect 1216 -3187 1262 -3149
rect 1216 -3221 1222 -3187
rect 1256 -3221 1262 -3187
rect 1216 -3259 1262 -3221
rect 1216 -3293 1222 -3259
rect 1256 -3293 1262 -3259
rect 1216 -3331 1262 -3293
rect 1216 -3365 1222 -3331
rect 1256 -3365 1262 -3331
rect 1216 -3403 1262 -3365
rect 1216 -3437 1222 -3403
rect 1256 -3437 1262 -3403
rect 1216 -3475 1262 -3437
rect 1216 -3509 1222 -3475
rect 1256 -3509 1262 -3475
rect 1216 -3547 1262 -3509
rect 1216 -3581 1222 -3547
rect 1256 -3581 1262 -3547
rect 1216 -3619 1262 -3581
rect 1216 -3653 1222 -3619
rect 1256 -3653 1262 -3619
rect 1216 -3691 1262 -3653
rect 1216 -3725 1222 -3691
rect 1256 -3725 1262 -3691
rect 1216 -3763 1262 -3725
rect 1216 -3797 1222 -3763
rect 1256 -3797 1262 -3763
rect 1216 -3835 1262 -3797
rect 1216 -3869 1222 -3835
rect 1256 -3869 1262 -3835
rect 1216 -3907 1262 -3869
rect 1216 -3941 1222 -3907
rect 1256 -3941 1262 -3907
rect 1216 -3979 1262 -3941
rect 1216 -4013 1222 -3979
rect 1256 -4013 1262 -3979
rect 1216 -4051 1262 -4013
rect 1216 -4085 1222 -4051
rect 1256 -4085 1262 -4051
rect 1216 -4123 1262 -4085
rect 1216 -4157 1222 -4123
rect 1256 -4157 1262 -4123
rect 1216 -4195 1262 -4157
rect 1216 -4229 1222 -4195
rect 1256 -4229 1262 -4195
rect 1216 -4267 1262 -4229
rect 1216 -4301 1222 -4267
rect 1256 -4301 1262 -4267
rect 1216 -4339 1262 -4301
rect 1216 -4373 1222 -4339
rect 1256 -4373 1262 -4339
rect 1216 -4411 1262 -4373
rect 1216 -4445 1222 -4411
rect 1256 -4445 1262 -4411
rect 1216 -4483 1262 -4445
rect 1216 -4517 1222 -4483
rect 1256 -4517 1262 -4483
rect 1216 -4555 1262 -4517
rect 1216 -4589 1222 -4555
rect 1256 -4589 1262 -4555
rect 1216 -4627 1262 -4589
rect 1216 -4661 1222 -4627
rect 1256 -4661 1262 -4627
rect 1216 -4699 1262 -4661
rect 1216 -4733 1222 -4699
rect 1256 -4733 1262 -4699
rect 1216 -4771 1262 -4733
rect 1216 -4805 1222 -4771
rect 1256 -4805 1262 -4771
rect 1216 -4843 1262 -4805
rect 1216 -4877 1222 -4843
rect 1256 -4877 1262 -4843
rect 1216 -4915 1262 -4877
rect 1216 -4949 1222 -4915
rect 1256 -4949 1262 -4915
rect 1216 -4987 1262 -4949
rect 1216 -5021 1222 -4987
rect 1256 -5021 1262 -4987
rect 1216 -5059 1262 -5021
rect 1216 -5093 1222 -5059
rect 1256 -5093 1262 -5059
rect 1216 -5131 1262 -5093
rect 1216 -5165 1222 -5131
rect 1256 -5165 1262 -5131
rect 1216 -5203 1262 -5165
rect 1216 -5237 1222 -5203
rect 1256 -5237 1262 -5203
rect 1216 -5275 1262 -5237
rect 1216 -5309 1222 -5275
rect 1256 -5309 1262 -5275
rect 1216 -5347 1262 -5309
rect 1216 -5381 1222 -5347
rect 1256 -5381 1262 -5347
rect 1216 -5419 1262 -5381
rect 1216 -5453 1222 -5419
rect 1256 -5453 1262 -5419
rect 1216 -5491 1262 -5453
rect 1216 -5525 1222 -5491
rect 1256 -5525 1262 -5491
rect 1216 -5563 1262 -5525
rect 1216 -5597 1222 -5563
rect 1256 -5597 1262 -5563
rect 1216 -5635 1262 -5597
rect 1216 -5669 1222 -5635
rect 1256 -5669 1262 -5635
rect 1216 -5707 1262 -5669
rect 1216 -5741 1222 -5707
rect 1256 -5741 1262 -5707
rect 1216 -5779 1262 -5741
rect 1216 -5813 1222 -5779
rect 1256 -5813 1262 -5779
rect 1216 -5851 1262 -5813
rect 1216 -5885 1222 -5851
rect 1256 -5885 1262 -5851
rect 1216 -5923 1262 -5885
rect 1216 -5957 1222 -5923
rect 1256 -5957 1262 -5923
rect 1216 -5995 1262 -5957
rect 1216 -6029 1222 -5995
rect 1256 -6029 1262 -5995
rect 1216 -6067 1262 -6029
rect 1216 -6101 1222 -6067
rect 1256 -6101 1262 -6067
rect 1216 -6139 1262 -6101
rect 1216 -6173 1222 -6139
rect 1256 -6173 1262 -6139
rect 1216 -6211 1262 -6173
rect 1216 -6245 1222 -6211
rect 1256 -6245 1262 -6211
rect 1216 -6283 1262 -6245
rect 1216 -6317 1222 -6283
rect 1256 -6317 1262 -6283
rect 1216 -6355 1262 -6317
rect 1216 -6389 1222 -6355
rect 1256 -6389 1262 -6355
rect 1216 -6427 1262 -6389
rect 1216 -6461 1222 -6427
rect 1256 -6461 1262 -6427
rect 1216 -6499 1262 -6461
rect 1216 -6533 1222 -6499
rect 1256 -6533 1262 -6499
rect 1216 -6571 1262 -6533
rect 1216 -6605 1222 -6571
rect 1256 -6605 1262 -6571
rect 1216 -6643 1262 -6605
rect 1216 -6677 1222 -6643
rect 1256 -6677 1262 -6643
rect 1216 -6715 1262 -6677
rect 1216 -6749 1222 -6715
rect 1256 -6749 1262 -6715
rect 1216 -6787 1262 -6749
rect 1216 -6821 1222 -6787
rect 1256 -6821 1262 -6787
rect 1216 -6859 1262 -6821
rect 1216 -6893 1222 -6859
rect 1256 -6893 1262 -6859
rect 1216 -6931 1262 -6893
rect 1216 -6965 1222 -6931
rect 1256 -6965 1262 -6931
rect 1216 -7003 1262 -6965
rect 1216 -7037 1222 -7003
rect 1256 -7037 1262 -7003
rect 1216 -7075 1262 -7037
rect 1216 -7109 1222 -7075
rect 1256 -7109 1262 -7075
rect 1216 -7147 1262 -7109
rect 1216 -7181 1222 -7147
rect 1256 -7181 1262 -7147
rect 1216 -7219 1262 -7181
rect 1216 -7253 1222 -7219
rect 1256 -7253 1262 -7219
rect 1216 -7291 1262 -7253
rect 1216 -7325 1222 -7291
rect 1256 -7325 1262 -7291
rect 1216 -7363 1262 -7325
rect 1216 -7397 1222 -7363
rect 1256 -7397 1262 -7363
rect 1216 -7435 1262 -7397
rect 1216 -7469 1222 -7435
rect 1256 -7469 1262 -7435
rect 1216 -7507 1262 -7469
rect 1216 -7541 1222 -7507
rect 1256 -7541 1262 -7507
rect 1216 -7579 1262 -7541
rect 1216 -7613 1222 -7579
rect 1256 -7613 1262 -7579
rect 1216 -7651 1262 -7613
rect 1216 -7685 1222 -7651
rect 1256 -7685 1262 -7651
rect 1216 -7723 1262 -7685
rect 1216 -7757 1222 -7723
rect 1256 -7757 1262 -7723
rect 1216 -7795 1262 -7757
rect 1216 -7829 1222 -7795
rect 1256 -7829 1262 -7795
rect 1216 -7867 1262 -7829
rect 1216 -7901 1222 -7867
rect 1256 -7901 1262 -7867
rect 1216 -7939 1262 -7901
rect 1216 -7973 1222 -7939
rect 1256 -7973 1262 -7939
rect 1216 -8011 1262 -7973
rect 1216 -8045 1222 -8011
rect 1256 -8045 1262 -8011
rect 1216 -8083 1262 -8045
rect 1216 -8117 1222 -8083
rect 1256 -8117 1262 -8083
rect 1216 -8155 1262 -8117
rect 1216 -8189 1222 -8155
rect 1256 -8189 1262 -8155
rect 1216 -8227 1262 -8189
rect 1216 -8261 1222 -8227
rect 1256 -8261 1262 -8227
rect 1216 -8299 1262 -8261
rect 1216 -8333 1222 -8299
rect 1256 -8333 1262 -8299
rect 1216 -8371 1262 -8333
rect 1216 -8405 1222 -8371
rect 1256 -8405 1262 -8371
rect 1216 -8443 1262 -8405
rect 1216 -8477 1222 -8443
rect 1256 -8477 1262 -8443
rect 1216 -8515 1262 -8477
rect 1216 -8549 1222 -8515
rect 1256 -8549 1262 -8515
rect 1216 -8587 1262 -8549
rect 1216 -8621 1222 -8587
rect 1256 -8621 1262 -8587
rect 1216 -8659 1262 -8621
rect 1216 -8693 1222 -8659
rect 1256 -8693 1262 -8659
rect 1216 -8731 1262 -8693
rect 1216 -8765 1222 -8731
rect 1256 -8765 1262 -8731
rect 1216 -8803 1262 -8765
rect 1216 -8837 1222 -8803
rect 1256 -8837 1262 -8803
rect 1216 -8875 1262 -8837
rect 1216 -8909 1222 -8875
rect 1256 -8909 1262 -8875
rect 1216 -8947 1262 -8909
rect 1216 -8981 1222 -8947
rect 1256 -8981 1262 -8947
rect 1216 -9019 1262 -8981
rect 1216 -9053 1222 -9019
rect 1256 -9053 1262 -9019
rect 1216 -9091 1262 -9053
rect 1216 -9125 1222 -9091
rect 1256 -9125 1262 -9091
rect 1216 -9163 1262 -9125
rect 1216 -9197 1222 -9163
rect 1256 -9197 1262 -9163
rect 1216 -9235 1262 -9197
rect 1216 -9269 1222 -9235
rect 1256 -9269 1262 -9235
rect 1216 -9307 1262 -9269
rect 1216 -9341 1222 -9307
rect 1256 -9341 1262 -9307
rect 1216 -9379 1262 -9341
rect 1216 -9413 1222 -9379
rect 1256 -9413 1262 -9379
rect 1216 -9451 1262 -9413
rect 1216 -9485 1222 -9451
rect 1256 -9485 1262 -9451
rect 1216 -9523 1262 -9485
rect 1216 -9557 1222 -9523
rect 1256 -9557 1262 -9523
rect 1216 -9600 1262 -9557
rect 1334 9557 1380 9600
rect 1334 9523 1340 9557
rect 1374 9523 1380 9557
rect 1334 9485 1380 9523
rect 1334 9451 1340 9485
rect 1374 9451 1380 9485
rect 1334 9413 1380 9451
rect 1334 9379 1340 9413
rect 1374 9379 1380 9413
rect 1334 9341 1380 9379
rect 1334 9307 1340 9341
rect 1374 9307 1380 9341
rect 1334 9269 1380 9307
rect 1334 9235 1340 9269
rect 1374 9235 1380 9269
rect 1334 9197 1380 9235
rect 1334 9163 1340 9197
rect 1374 9163 1380 9197
rect 1334 9125 1380 9163
rect 1334 9091 1340 9125
rect 1374 9091 1380 9125
rect 1334 9053 1380 9091
rect 1334 9019 1340 9053
rect 1374 9019 1380 9053
rect 1334 8981 1380 9019
rect 1334 8947 1340 8981
rect 1374 8947 1380 8981
rect 1334 8909 1380 8947
rect 1334 8875 1340 8909
rect 1374 8875 1380 8909
rect 1334 8837 1380 8875
rect 1334 8803 1340 8837
rect 1374 8803 1380 8837
rect 1334 8765 1380 8803
rect 1334 8731 1340 8765
rect 1374 8731 1380 8765
rect 1334 8693 1380 8731
rect 1334 8659 1340 8693
rect 1374 8659 1380 8693
rect 1334 8621 1380 8659
rect 1334 8587 1340 8621
rect 1374 8587 1380 8621
rect 1334 8549 1380 8587
rect 1334 8515 1340 8549
rect 1374 8515 1380 8549
rect 1334 8477 1380 8515
rect 1334 8443 1340 8477
rect 1374 8443 1380 8477
rect 1334 8405 1380 8443
rect 1334 8371 1340 8405
rect 1374 8371 1380 8405
rect 1334 8333 1380 8371
rect 1334 8299 1340 8333
rect 1374 8299 1380 8333
rect 1334 8261 1380 8299
rect 1334 8227 1340 8261
rect 1374 8227 1380 8261
rect 1334 8189 1380 8227
rect 1334 8155 1340 8189
rect 1374 8155 1380 8189
rect 1334 8117 1380 8155
rect 1334 8083 1340 8117
rect 1374 8083 1380 8117
rect 1334 8045 1380 8083
rect 1334 8011 1340 8045
rect 1374 8011 1380 8045
rect 1334 7973 1380 8011
rect 1334 7939 1340 7973
rect 1374 7939 1380 7973
rect 1334 7901 1380 7939
rect 1334 7867 1340 7901
rect 1374 7867 1380 7901
rect 1334 7829 1380 7867
rect 1334 7795 1340 7829
rect 1374 7795 1380 7829
rect 1334 7757 1380 7795
rect 1334 7723 1340 7757
rect 1374 7723 1380 7757
rect 1334 7685 1380 7723
rect 1334 7651 1340 7685
rect 1374 7651 1380 7685
rect 1334 7613 1380 7651
rect 1334 7579 1340 7613
rect 1374 7579 1380 7613
rect 1334 7541 1380 7579
rect 1334 7507 1340 7541
rect 1374 7507 1380 7541
rect 1334 7469 1380 7507
rect 1334 7435 1340 7469
rect 1374 7435 1380 7469
rect 1334 7397 1380 7435
rect 1334 7363 1340 7397
rect 1374 7363 1380 7397
rect 1334 7325 1380 7363
rect 1334 7291 1340 7325
rect 1374 7291 1380 7325
rect 1334 7253 1380 7291
rect 1334 7219 1340 7253
rect 1374 7219 1380 7253
rect 1334 7181 1380 7219
rect 1334 7147 1340 7181
rect 1374 7147 1380 7181
rect 1334 7109 1380 7147
rect 1334 7075 1340 7109
rect 1374 7075 1380 7109
rect 1334 7037 1380 7075
rect 1334 7003 1340 7037
rect 1374 7003 1380 7037
rect 1334 6965 1380 7003
rect 1334 6931 1340 6965
rect 1374 6931 1380 6965
rect 1334 6893 1380 6931
rect 1334 6859 1340 6893
rect 1374 6859 1380 6893
rect 1334 6821 1380 6859
rect 1334 6787 1340 6821
rect 1374 6787 1380 6821
rect 1334 6749 1380 6787
rect 1334 6715 1340 6749
rect 1374 6715 1380 6749
rect 1334 6677 1380 6715
rect 1334 6643 1340 6677
rect 1374 6643 1380 6677
rect 1334 6605 1380 6643
rect 1334 6571 1340 6605
rect 1374 6571 1380 6605
rect 1334 6533 1380 6571
rect 1334 6499 1340 6533
rect 1374 6499 1380 6533
rect 1334 6461 1380 6499
rect 1334 6427 1340 6461
rect 1374 6427 1380 6461
rect 1334 6389 1380 6427
rect 1334 6355 1340 6389
rect 1374 6355 1380 6389
rect 1334 6317 1380 6355
rect 1334 6283 1340 6317
rect 1374 6283 1380 6317
rect 1334 6245 1380 6283
rect 1334 6211 1340 6245
rect 1374 6211 1380 6245
rect 1334 6173 1380 6211
rect 1334 6139 1340 6173
rect 1374 6139 1380 6173
rect 1334 6101 1380 6139
rect 1334 6067 1340 6101
rect 1374 6067 1380 6101
rect 1334 6029 1380 6067
rect 1334 5995 1340 6029
rect 1374 5995 1380 6029
rect 1334 5957 1380 5995
rect 1334 5923 1340 5957
rect 1374 5923 1380 5957
rect 1334 5885 1380 5923
rect 1334 5851 1340 5885
rect 1374 5851 1380 5885
rect 1334 5813 1380 5851
rect 1334 5779 1340 5813
rect 1374 5779 1380 5813
rect 1334 5741 1380 5779
rect 1334 5707 1340 5741
rect 1374 5707 1380 5741
rect 1334 5669 1380 5707
rect 1334 5635 1340 5669
rect 1374 5635 1380 5669
rect 1334 5597 1380 5635
rect 1334 5563 1340 5597
rect 1374 5563 1380 5597
rect 1334 5525 1380 5563
rect 1334 5491 1340 5525
rect 1374 5491 1380 5525
rect 1334 5453 1380 5491
rect 1334 5419 1340 5453
rect 1374 5419 1380 5453
rect 1334 5381 1380 5419
rect 1334 5347 1340 5381
rect 1374 5347 1380 5381
rect 1334 5309 1380 5347
rect 1334 5275 1340 5309
rect 1374 5275 1380 5309
rect 1334 5237 1380 5275
rect 1334 5203 1340 5237
rect 1374 5203 1380 5237
rect 1334 5165 1380 5203
rect 1334 5131 1340 5165
rect 1374 5131 1380 5165
rect 1334 5093 1380 5131
rect 1334 5059 1340 5093
rect 1374 5059 1380 5093
rect 1334 5021 1380 5059
rect 1334 4987 1340 5021
rect 1374 4987 1380 5021
rect 1334 4949 1380 4987
rect 1334 4915 1340 4949
rect 1374 4915 1380 4949
rect 1334 4877 1380 4915
rect 1334 4843 1340 4877
rect 1374 4843 1380 4877
rect 1334 4805 1380 4843
rect 1334 4771 1340 4805
rect 1374 4771 1380 4805
rect 1334 4733 1380 4771
rect 1334 4699 1340 4733
rect 1374 4699 1380 4733
rect 1334 4661 1380 4699
rect 1334 4627 1340 4661
rect 1374 4627 1380 4661
rect 1334 4589 1380 4627
rect 1334 4555 1340 4589
rect 1374 4555 1380 4589
rect 1334 4517 1380 4555
rect 1334 4483 1340 4517
rect 1374 4483 1380 4517
rect 1334 4445 1380 4483
rect 1334 4411 1340 4445
rect 1374 4411 1380 4445
rect 1334 4373 1380 4411
rect 1334 4339 1340 4373
rect 1374 4339 1380 4373
rect 1334 4301 1380 4339
rect 1334 4267 1340 4301
rect 1374 4267 1380 4301
rect 1334 4229 1380 4267
rect 1334 4195 1340 4229
rect 1374 4195 1380 4229
rect 1334 4157 1380 4195
rect 1334 4123 1340 4157
rect 1374 4123 1380 4157
rect 1334 4085 1380 4123
rect 1334 4051 1340 4085
rect 1374 4051 1380 4085
rect 1334 4013 1380 4051
rect 1334 3979 1340 4013
rect 1374 3979 1380 4013
rect 1334 3941 1380 3979
rect 1334 3907 1340 3941
rect 1374 3907 1380 3941
rect 1334 3869 1380 3907
rect 1334 3835 1340 3869
rect 1374 3835 1380 3869
rect 1334 3797 1380 3835
rect 1334 3763 1340 3797
rect 1374 3763 1380 3797
rect 1334 3725 1380 3763
rect 1334 3691 1340 3725
rect 1374 3691 1380 3725
rect 1334 3653 1380 3691
rect 1334 3619 1340 3653
rect 1374 3619 1380 3653
rect 1334 3581 1380 3619
rect 1334 3547 1340 3581
rect 1374 3547 1380 3581
rect 1334 3509 1380 3547
rect 1334 3475 1340 3509
rect 1374 3475 1380 3509
rect 1334 3437 1380 3475
rect 1334 3403 1340 3437
rect 1374 3403 1380 3437
rect 1334 3365 1380 3403
rect 1334 3331 1340 3365
rect 1374 3331 1380 3365
rect 1334 3293 1380 3331
rect 1334 3259 1340 3293
rect 1374 3259 1380 3293
rect 1334 3221 1380 3259
rect 1334 3187 1340 3221
rect 1374 3187 1380 3221
rect 1334 3149 1380 3187
rect 1334 3115 1340 3149
rect 1374 3115 1380 3149
rect 1334 3077 1380 3115
rect 1334 3043 1340 3077
rect 1374 3043 1380 3077
rect 1334 3005 1380 3043
rect 1334 2971 1340 3005
rect 1374 2971 1380 3005
rect 1334 2933 1380 2971
rect 1334 2899 1340 2933
rect 1374 2899 1380 2933
rect 1334 2861 1380 2899
rect 1334 2827 1340 2861
rect 1374 2827 1380 2861
rect 1334 2789 1380 2827
rect 1334 2755 1340 2789
rect 1374 2755 1380 2789
rect 1334 2717 1380 2755
rect 1334 2683 1340 2717
rect 1374 2683 1380 2717
rect 1334 2645 1380 2683
rect 1334 2611 1340 2645
rect 1374 2611 1380 2645
rect 1334 2573 1380 2611
rect 1334 2539 1340 2573
rect 1374 2539 1380 2573
rect 1334 2501 1380 2539
rect 1334 2467 1340 2501
rect 1374 2467 1380 2501
rect 1334 2429 1380 2467
rect 1334 2395 1340 2429
rect 1374 2395 1380 2429
rect 1334 2357 1380 2395
rect 1334 2323 1340 2357
rect 1374 2323 1380 2357
rect 1334 2285 1380 2323
rect 1334 2251 1340 2285
rect 1374 2251 1380 2285
rect 1334 2213 1380 2251
rect 1334 2179 1340 2213
rect 1374 2179 1380 2213
rect 1334 2141 1380 2179
rect 1334 2107 1340 2141
rect 1374 2107 1380 2141
rect 1334 2069 1380 2107
rect 1334 2035 1340 2069
rect 1374 2035 1380 2069
rect 1334 1997 1380 2035
rect 1334 1963 1340 1997
rect 1374 1963 1380 1997
rect 1334 1925 1380 1963
rect 1334 1891 1340 1925
rect 1374 1891 1380 1925
rect 1334 1853 1380 1891
rect 1334 1819 1340 1853
rect 1374 1819 1380 1853
rect 1334 1781 1380 1819
rect 1334 1747 1340 1781
rect 1374 1747 1380 1781
rect 1334 1709 1380 1747
rect 1334 1675 1340 1709
rect 1374 1675 1380 1709
rect 1334 1637 1380 1675
rect 1334 1603 1340 1637
rect 1374 1603 1380 1637
rect 1334 1565 1380 1603
rect 1334 1531 1340 1565
rect 1374 1531 1380 1565
rect 1334 1493 1380 1531
rect 1334 1459 1340 1493
rect 1374 1459 1380 1493
rect 1334 1421 1380 1459
rect 1334 1387 1340 1421
rect 1374 1387 1380 1421
rect 1334 1349 1380 1387
rect 1334 1315 1340 1349
rect 1374 1315 1380 1349
rect 1334 1277 1380 1315
rect 1334 1243 1340 1277
rect 1374 1243 1380 1277
rect 1334 1205 1380 1243
rect 1334 1171 1340 1205
rect 1374 1171 1380 1205
rect 1334 1133 1380 1171
rect 1334 1099 1340 1133
rect 1374 1099 1380 1133
rect 1334 1061 1380 1099
rect 1334 1027 1340 1061
rect 1374 1027 1380 1061
rect 1334 989 1380 1027
rect 1334 955 1340 989
rect 1374 955 1380 989
rect 1334 917 1380 955
rect 1334 883 1340 917
rect 1374 883 1380 917
rect 1334 845 1380 883
rect 1334 811 1340 845
rect 1374 811 1380 845
rect 1334 773 1380 811
rect 1334 739 1340 773
rect 1374 739 1380 773
rect 1334 701 1380 739
rect 1334 667 1340 701
rect 1374 667 1380 701
rect 1334 629 1380 667
rect 1334 595 1340 629
rect 1374 595 1380 629
rect 1334 557 1380 595
rect 1334 523 1340 557
rect 1374 523 1380 557
rect 1334 485 1380 523
rect 1334 451 1340 485
rect 1374 451 1380 485
rect 1334 413 1380 451
rect 1334 379 1340 413
rect 1374 379 1380 413
rect 1334 341 1380 379
rect 1334 307 1340 341
rect 1374 307 1380 341
rect 1334 269 1380 307
rect 1334 235 1340 269
rect 1374 235 1380 269
rect 1334 197 1380 235
rect 1334 163 1340 197
rect 1374 163 1380 197
rect 1334 125 1380 163
rect 1334 91 1340 125
rect 1374 91 1380 125
rect 1334 53 1380 91
rect 1334 19 1340 53
rect 1374 19 1380 53
rect 1334 -19 1380 19
rect 1334 -53 1340 -19
rect 1374 -53 1380 -19
rect 1334 -91 1380 -53
rect 1334 -125 1340 -91
rect 1374 -125 1380 -91
rect 1334 -163 1380 -125
rect 1334 -197 1340 -163
rect 1374 -197 1380 -163
rect 1334 -235 1380 -197
rect 1334 -269 1340 -235
rect 1374 -269 1380 -235
rect 1334 -307 1380 -269
rect 1334 -341 1340 -307
rect 1374 -341 1380 -307
rect 1334 -379 1380 -341
rect 1334 -413 1340 -379
rect 1374 -413 1380 -379
rect 1334 -451 1380 -413
rect 1334 -485 1340 -451
rect 1374 -485 1380 -451
rect 1334 -523 1380 -485
rect 1334 -557 1340 -523
rect 1374 -557 1380 -523
rect 1334 -595 1380 -557
rect 1334 -629 1340 -595
rect 1374 -629 1380 -595
rect 1334 -667 1380 -629
rect 1334 -701 1340 -667
rect 1374 -701 1380 -667
rect 1334 -739 1380 -701
rect 1334 -773 1340 -739
rect 1374 -773 1380 -739
rect 1334 -811 1380 -773
rect 1334 -845 1340 -811
rect 1374 -845 1380 -811
rect 1334 -883 1380 -845
rect 1334 -917 1340 -883
rect 1374 -917 1380 -883
rect 1334 -955 1380 -917
rect 1334 -989 1340 -955
rect 1374 -989 1380 -955
rect 1334 -1027 1380 -989
rect 1334 -1061 1340 -1027
rect 1374 -1061 1380 -1027
rect 1334 -1099 1380 -1061
rect 1334 -1133 1340 -1099
rect 1374 -1133 1380 -1099
rect 1334 -1171 1380 -1133
rect 1334 -1205 1340 -1171
rect 1374 -1205 1380 -1171
rect 1334 -1243 1380 -1205
rect 1334 -1277 1340 -1243
rect 1374 -1277 1380 -1243
rect 1334 -1315 1380 -1277
rect 1334 -1349 1340 -1315
rect 1374 -1349 1380 -1315
rect 1334 -1387 1380 -1349
rect 1334 -1421 1340 -1387
rect 1374 -1421 1380 -1387
rect 1334 -1459 1380 -1421
rect 1334 -1493 1340 -1459
rect 1374 -1493 1380 -1459
rect 1334 -1531 1380 -1493
rect 1334 -1565 1340 -1531
rect 1374 -1565 1380 -1531
rect 1334 -1603 1380 -1565
rect 1334 -1637 1340 -1603
rect 1374 -1637 1380 -1603
rect 1334 -1675 1380 -1637
rect 1334 -1709 1340 -1675
rect 1374 -1709 1380 -1675
rect 1334 -1747 1380 -1709
rect 1334 -1781 1340 -1747
rect 1374 -1781 1380 -1747
rect 1334 -1819 1380 -1781
rect 1334 -1853 1340 -1819
rect 1374 -1853 1380 -1819
rect 1334 -1891 1380 -1853
rect 1334 -1925 1340 -1891
rect 1374 -1925 1380 -1891
rect 1334 -1963 1380 -1925
rect 1334 -1997 1340 -1963
rect 1374 -1997 1380 -1963
rect 1334 -2035 1380 -1997
rect 1334 -2069 1340 -2035
rect 1374 -2069 1380 -2035
rect 1334 -2107 1380 -2069
rect 1334 -2141 1340 -2107
rect 1374 -2141 1380 -2107
rect 1334 -2179 1380 -2141
rect 1334 -2213 1340 -2179
rect 1374 -2213 1380 -2179
rect 1334 -2251 1380 -2213
rect 1334 -2285 1340 -2251
rect 1374 -2285 1380 -2251
rect 1334 -2323 1380 -2285
rect 1334 -2357 1340 -2323
rect 1374 -2357 1380 -2323
rect 1334 -2395 1380 -2357
rect 1334 -2429 1340 -2395
rect 1374 -2429 1380 -2395
rect 1334 -2467 1380 -2429
rect 1334 -2501 1340 -2467
rect 1374 -2501 1380 -2467
rect 1334 -2539 1380 -2501
rect 1334 -2573 1340 -2539
rect 1374 -2573 1380 -2539
rect 1334 -2611 1380 -2573
rect 1334 -2645 1340 -2611
rect 1374 -2645 1380 -2611
rect 1334 -2683 1380 -2645
rect 1334 -2717 1340 -2683
rect 1374 -2717 1380 -2683
rect 1334 -2755 1380 -2717
rect 1334 -2789 1340 -2755
rect 1374 -2789 1380 -2755
rect 1334 -2827 1380 -2789
rect 1334 -2861 1340 -2827
rect 1374 -2861 1380 -2827
rect 1334 -2899 1380 -2861
rect 1334 -2933 1340 -2899
rect 1374 -2933 1380 -2899
rect 1334 -2971 1380 -2933
rect 1334 -3005 1340 -2971
rect 1374 -3005 1380 -2971
rect 1334 -3043 1380 -3005
rect 1334 -3077 1340 -3043
rect 1374 -3077 1380 -3043
rect 1334 -3115 1380 -3077
rect 1334 -3149 1340 -3115
rect 1374 -3149 1380 -3115
rect 1334 -3187 1380 -3149
rect 1334 -3221 1340 -3187
rect 1374 -3221 1380 -3187
rect 1334 -3259 1380 -3221
rect 1334 -3293 1340 -3259
rect 1374 -3293 1380 -3259
rect 1334 -3331 1380 -3293
rect 1334 -3365 1340 -3331
rect 1374 -3365 1380 -3331
rect 1334 -3403 1380 -3365
rect 1334 -3437 1340 -3403
rect 1374 -3437 1380 -3403
rect 1334 -3475 1380 -3437
rect 1334 -3509 1340 -3475
rect 1374 -3509 1380 -3475
rect 1334 -3547 1380 -3509
rect 1334 -3581 1340 -3547
rect 1374 -3581 1380 -3547
rect 1334 -3619 1380 -3581
rect 1334 -3653 1340 -3619
rect 1374 -3653 1380 -3619
rect 1334 -3691 1380 -3653
rect 1334 -3725 1340 -3691
rect 1374 -3725 1380 -3691
rect 1334 -3763 1380 -3725
rect 1334 -3797 1340 -3763
rect 1374 -3797 1380 -3763
rect 1334 -3835 1380 -3797
rect 1334 -3869 1340 -3835
rect 1374 -3869 1380 -3835
rect 1334 -3907 1380 -3869
rect 1334 -3941 1340 -3907
rect 1374 -3941 1380 -3907
rect 1334 -3979 1380 -3941
rect 1334 -4013 1340 -3979
rect 1374 -4013 1380 -3979
rect 1334 -4051 1380 -4013
rect 1334 -4085 1340 -4051
rect 1374 -4085 1380 -4051
rect 1334 -4123 1380 -4085
rect 1334 -4157 1340 -4123
rect 1374 -4157 1380 -4123
rect 1334 -4195 1380 -4157
rect 1334 -4229 1340 -4195
rect 1374 -4229 1380 -4195
rect 1334 -4267 1380 -4229
rect 1334 -4301 1340 -4267
rect 1374 -4301 1380 -4267
rect 1334 -4339 1380 -4301
rect 1334 -4373 1340 -4339
rect 1374 -4373 1380 -4339
rect 1334 -4411 1380 -4373
rect 1334 -4445 1340 -4411
rect 1374 -4445 1380 -4411
rect 1334 -4483 1380 -4445
rect 1334 -4517 1340 -4483
rect 1374 -4517 1380 -4483
rect 1334 -4555 1380 -4517
rect 1334 -4589 1340 -4555
rect 1374 -4589 1380 -4555
rect 1334 -4627 1380 -4589
rect 1334 -4661 1340 -4627
rect 1374 -4661 1380 -4627
rect 1334 -4699 1380 -4661
rect 1334 -4733 1340 -4699
rect 1374 -4733 1380 -4699
rect 1334 -4771 1380 -4733
rect 1334 -4805 1340 -4771
rect 1374 -4805 1380 -4771
rect 1334 -4843 1380 -4805
rect 1334 -4877 1340 -4843
rect 1374 -4877 1380 -4843
rect 1334 -4915 1380 -4877
rect 1334 -4949 1340 -4915
rect 1374 -4949 1380 -4915
rect 1334 -4987 1380 -4949
rect 1334 -5021 1340 -4987
rect 1374 -5021 1380 -4987
rect 1334 -5059 1380 -5021
rect 1334 -5093 1340 -5059
rect 1374 -5093 1380 -5059
rect 1334 -5131 1380 -5093
rect 1334 -5165 1340 -5131
rect 1374 -5165 1380 -5131
rect 1334 -5203 1380 -5165
rect 1334 -5237 1340 -5203
rect 1374 -5237 1380 -5203
rect 1334 -5275 1380 -5237
rect 1334 -5309 1340 -5275
rect 1374 -5309 1380 -5275
rect 1334 -5347 1380 -5309
rect 1334 -5381 1340 -5347
rect 1374 -5381 1380 -5347
rect 1334 -5419 1380 -5381
rect 1334 -5453 1340 -5419
rect 1374 -5453 1380 -5419
rect 1334 -5491 1380 -5453
rect 1334 -5525 1340 -5491
rect 1374 -5525 1380 -5491
rect 1334 -5563 1380 -5525
rect 1334 -5597 1340 -5563
rect 1374 -5597 1380 -5563
rect 1334 -5635 1380 -5597
rect 1334 -5669 1340 -5635
rect 1374 -5669 1380 -5635
rect 1334 -5707 1380 -5669
rect 1334 -5741 1340 -5707
rect 1374 -5741 1380 -5707
rect 1334 -5779 1380 -5741
rect 1334 -5813 1340 -5779
rect 1374 -5813 1380 -5779
rect 1334 -5851 1380 -5813
rect 1334 -5885 1340 -5851
rect 1374 -5885 1380 -5851
rect 1334 -5923 1380 -5885
rect 1334 -5957 1340 -5923
rect 1374 -5957 1380 -5923
rect 1334 -5995 1380 -5957
rect 1334 -6029 1340 -5995
rect 1374 -6029 1380 -5995
rect 1334 -6067 1380 -6029
rect 1334 -6101 1340 -6067
rect 1374 -6101 1380 -6067
rect 1334 -6139 1380 -6101
rect 1334 -6173 1340 -6139
rect 1374 -6173 1380 -6139
rect 1334 -6211 1380 -6173
rect 1334 -6245 1340 -6211
rect 1374 -6245 1380 -6211
rect 1334 -6283 1380 -6245
rect 1334 -6317 1340 -6283
rect 1374 -6317 1380 -6283
rect 1334 -6355 1380 -6317
rect 1334 -6389 1340 -6355
rect 1374 -6389 1380 -6355
rect 1334 -6427 1380 -6389
rect 1334 -6461 1340 -6427
rect 1374 -6461 1380 -6427
rect 1334 -6499 1380 -6461
rect 1334 -6533 1340 -6499
rect 1374 -6533 1380 -6499
rect 1334 -6571 1380 -6533
rect 1334 -6605 1340 -6571
rect 1374 -6605 1380 -6571
rect 1334 -6643 1380 -6605
rect 1334 -6677 1340 -6643
rect 1374 -6677 1380 -6643
rect 1334 -6715 1380 -6677
rect 1334 -6749 1340 -6715
rect 1374 -6749 1380 -6715
rect 1334 -6787 1380 -6749
rect 1334 -6821 1340 -6787
rect 1374 -6821 1380 -6787
rect 1334 -6859 1380 -6821
rect 1334 -6893 1340 -6859
rect 1374 -6893 1380 -6859
rect 1334 -6931 1380 -6893
rect 1334 -6965 1340 -6931
rect 1374 -6965 1380 -6931
rect 1334 -7003 1380 -6965
rect 1334 -7037 1340 -7003
rect 1374 -7037 1380 -7003
rect 1334 -7075 1380 -7037
rect 1334 -7109 1340 -7075
rect 1374 -7109 1380 -7075
rect 1334 -7147 1380 -7109
rect 1334 -7181 1340 -7147
rect 1374 -7181 1380 -7147
rect 1334 -7219 1380 -7181
rect 1334 -7253 1340 -7219
rect 1374 -7253 1380 -7219
rect 1334 -7291 1380 -7253
rect 1334 -7325 1340 -7291
rect 1374 -7325 1380 -7291
rect 1334 -7363 1380 -7325
rect 1334 -7397 1340 -7363
rect 1374 -7397 1380 -7363
rect 1334 -7435 1380 -7397
rect 1334 -7469 1340 -7435
rect 1374 -7469 1380 -7435
rect 1334 -7507 1380 -7469
rect 1334 -7541 1340 -7507
rect 1374 -7541 1380 -7507
rect 1334 -7579 1380 -7541
rect 1334 -7613 1340 -7579
rect 1374 -7613 1380 -7579
rect 1334 -7651 1380 -7613
rect 1334 -7685 1340 -7651
rect 1374 -7685 1380 -7651
rect 1334 -7723 1380 -7685
rect 1334 -7757 1340 -7723
rect 1374 -7757 1380 -7723
rect 1334 -7795 1380 -7757
rect 1334 -7829 1340 -7795
rect 1374 -7829 1380 -7795
rect 1334 -7867 1380 -7829
rect 1334 -7901 1340 -7867
rect 1374 -7901 1380 -7867
rect 1334 -7939 1380 -7901
rect 1334 -7973 1340 -7939
rect 1374 -7973 1380 -7939
rect 1334 -8011 1380 -7973
rect 1334 -8045 1340 -8011
rect 1374 -8045 1380 -8011
rect 1334 -8083 1380 -8045
rect 1334 -8117 1340 -8083
rect 1374 -8117 1380 -8083
rect 1334 -8155 1380 -8117
rect 1334 -8189 1340 -8155
rect 1374 -8189 1380 -8155
rect 1334 -8227 1380 -8189
rect 1334 -8261 1340 -8227
rect 1374 -8261 1380 -8227
rect 1334 -8299 1380 -8261
rect 1334 -8333 1340 -8299
rect 1374 -8333 1380 -8299
rect 1334 -8371 1380 -8333
rect 1334 -8405 1340 -8371
rect 1374 -8405 1380 -8371
rect 1334 -8443 1380 -8405
rect 1334 -8477 1340 -8443
rect 1374 -8477 1380 -8443
rect 1334 -8515 1380 -8477
rect 1334 -8549 1340 -8515
rect 1374 -8549 1380 -8515
rect 1334 -8587 1380 -8549
rect 1334 -8621 1340 -8587
rect 1374 -8621 1380 -8587
rect 1334 -8659 1380 -8621
rect 1334 -8693 1340 -8659
rect 1374 -8693 1380 -8659
rect 1334 -8731 1380 -8693
rect 1334 -8765 1340 -8731
rect 1374 -8765 1380 -8731
rect 1334 -8803 1380 -8765
rect 1334 -8837 1340 -8803
rect 1374 -8837 1380 -8803
rect 1334 -8875 1380 -8837
rect 1334 -8909 1340 -8875
rect 1374 -8909 1380 -8875
rect 1334 -8947 1380 -8909
rect 1334 -8981 1340 -8947
rect 1374 -8981 1380 -8947
rect 1334 -9019 1380 -8981
rect 1334 -9053 1340 -9019
rect 1374 -9053 1380 -9019
rect 1334 -9091 1380 -9053
rect 1334 -9125 1340 -9091
rect 1374 -9125 1380 -9091
rect 1334 -9163 1380 -9125
rect 1334 -9197 1340 -9163
rect 1374 -9197 1380 -9163
rect 1334 -9235 1380 -9197
rect 1334 -9269 1340 -9235
rect 1374 -9269 1380 -9235
rect 1334 -9307 1380 -9269
rect 1334 -9341 1340 -9307
rect 1374 -9341 1380 -9307
rect 1334 -9379 1380 -9341
rect 1334 -9413 1340 -9379
rect 1374 -9413 1380 -9379
rect 1334 -9451 1380 -9413
rect 1334 -9485 1340 -9451
rect 1374 -9485 1380 -9451
rect 1334 -9523 1380 -9485
rect 1334 -9557 1340 -9523
rect 1374 -9557 1380 -9523
rect 1334 -9600 1380 -9557
rect 1452 9557 1498 9600
rect 1452 9523 1458 9557
rect 1492 9523 1498 9557
rect 1452 9485 1498 9523
rect 1452 9451 1458 9485
rect 1492 9451 1498 9485
rect 1452 9413 1498 9451
rect 1452 9379 1458 9413
rect 1492 9379 1498 9413
rect 1452 9341 1498 9379
rect 1452 9307 1458 9341
rect 1492 9307 1498 9341
rect 1452 9269 1498 9307
rect 1452 9235 1458 9269
rect 1492 9235 1498 9269
rect 1452 9197 1498 9235
rect 1452 9163 1458 9197
rect 1492 9163 1498 9197
rect 1452 9125 1498 9163
rect 1452 9091 1458 9125
rect 1492 9091 1498 9125
rect 1452 9053 1498 9091
rect 1452 9019 1458 9053
rect 1492 9019 1498 9053
rect 1452 8981 1498 9019
rect 1452 8947 1458 8981
rect 1492 8947 1498 8981
rect 1452 8909 1498 8947
rect 1452 8875 1458 8909
rect 1492 8875 1498 8909
rect 1452 8837 1498 8875
rect 1452 8803 1458 8837
rect 1492 8803 1498 8837
rect 1452 8765 1498 8803
rect 1452 8731 1458 8765
rect 1492 8731 1498 8765
rect 1452 8693 1498 8731
rect 1452 8659 1458 8693
rect 1492 8659 1498 8693
rect 1452 8621 1498 8659
rect 1452 8587 1458 8621
rect 1492 8587 1498 8621
rect 1452 8549 1498 8587
rect 1452 8515 1458 8549
rect 1492 8515 1498 8549
rect 1452 8477 1498 8515
rect 1452 8443 1458 8477
rect 1492 8443 1498 8477
rect 1452 8405 1498 8443
rect 1452 8371 1458 8405
rect 1492 8371 1498 8405
rect 1452 8333 1498 8371
rect 1452 8299 1458 8333
rect 1492 8299 1498 8333
rect 1452 8261 1498 8299
rect 1452 8227 1458 8261
rect 1492 8227 1498 8261
rect 1452 8189 1498 8227
rect 1452 8155 1458 8189
rect 1492 8155 1498 8189
rect 1452 8117 1498 8155
rect 1452 8083 1458 8117
rect 1492 8083 1498 8117
rect 1452 8045 1498 8083
rect 1452 8011 1458 8045
rect 1492 8011 1498 8045
rect 1452 7973 1498 8011
rect 1452 7939 1458 7973
rect 1492 7939 1498 7973
rect 1452 7901 1498 7939
rect 1452 7867 1458 7901
rect 1492 7867 1498 7901
rect 1452 7829 1498 7867
rect 1452 7795 1458 7829
rect 1492 7795 1498 7829
rect 1452 7757 1498 7795
rect 1452 7723 1458 7757
rect 1492 7723 1498 7757
rect 1452 7685 1498 7723
rect 1452 7651 1458 7685
rect 1492 7651 1498 7685
rect 1452 7613 1498 7651
rect 1452 7579 1458 7613
rect 1492 7579 1498 7613
rect 1452 7541 1498 7579
rect 1452 7507 1458 7541
rect 1492 7507 1498 7541
rect 1452 7469 1498 7507
rect 1452 7435 1458 7469
rect 1492 7435 1498 7469
rect 1452 7397 1498 7435
rect 1452 7363 1458 7397
rect 1492 7363 1498 7397
rect 1452 7325 1498 7363
rect 1452 7291 1458 7325
rect 1492 7291 1498 7325
rect 1452 7253 1498 7291
rect 1452 7219 1458 7253
rect 1492 7219 1498 7253
rect 1452 7181 1498 7219
rect 1452 7147 1458 7181
rect 1492 7147 1498 7181
rect 1452 7109 1498 7147
rect 1452 7075 1458 7109
rect 1492 7075 1498 7109
rect 1452 7037 1498 7075
rect 1452 7003 1458 7037
rect 1492 7003 1498 7037
rect 1452 6965 1498 7003
rect 1452 6931 1458 6965
rect 1492 6931 1498 6965
rect 1452 6893 1498 6931
rect 1452 6859 1458 6893
rect 1492 6859 1498 6893
rect 1452 6821 1498 6859
rect 1452 6787 1458 6821
rect 1492 6787 1498 6821
rect 1452 6749 1498 6787
rect 1452 6715 1458 6749
rect 1492 6715 1498 6749
rect 1452 6677 1498 6715
rect 1452 6643 1458 6677
rect 1492 6643 1498 6677
rect 1452 6605 1498 6643
rect 1452 6571 1458 6605
rect 1492 6571 1498 6605
rect 1452 6533 1498 6571
rect 1452 6499 1458 6533
rect 1492 6499 1498 6533
rect 1452 6461 1498 6499
rect 1452 6427 1458 6461
rect 1492 6427 1498 6461
rect 1452 6389 1498 6427
rect 1452 6355 1458 6389
rect 1492 6355 1498 6389
rect 1452 6317 1498 6355
rect 1452 6283 1458 6317
rect 1492 6283 1498 6317
rect 1452 6245 1498 6283
rect 1452 6211 1458 6245
rect 1492 6211 1498 6245
rect 1452 6173 1498 6211
rect 1452 6139 1458 6173
rect 1492 6139 1498 6173
rect 1452 6101 1498 6139
rect 1452 6067 1458 6101
rect 1492 6067 1498 6101
rect 1452 6029 1498 6067
rect 1452 5995 1458 6029
rect 1492 5995 1498 6029
rect 1452 5957 1498 5995
rect 1452 5923 1458 5957
rect 1492 5923 1498 5957
rect 1452 5885 1498 5923
rect 1452 5851 1458 5885
rect 1492 5851 1498 5885
rect 1452 5813 1498 5851
rect 1452 5779 1458 5813
rect 1492 5779 1498 5813
rect 1452 5741 1498 5779
rect 1452 5707 1458 5741
rect 1492 5707 1498 5741
rect 1452 5669 1498 5707
rect 1452 5635 1458 5669
rect 1492 5635 1498 5669
rect 1452 5597 1498 5635
rect 1452 5563 1458 5597
rect 1492 5563 1498 5597
rect 1452 5525 1498 5563
rect 1452 5491 1458 5525
rect 1492 5491 1498 5525
rect 1452 5453 1498 5491
rect 1452 5419 1458 5453
rect 1492 5419 1498 5453
rect 1452 5381 1498 5419
rect 1452 5347 1458 5381
rect 1492 5347 1498 5381
rect 1452 5309 1498 5347
rect 1452 5275 1458 5309
rect 1492 5275 1498 5309
rect 1452 5237 1498 5275
rect 1452 5203 1458 5237
rect 1492 5203 1498 5237
rect 1452 5165 1498 5203
rect 1452 5131 1458 5165
rect 1492 5131 1498 5165
rect 1452 5093 1498 5131
rect 1452 5059 1458 5093
rect 1492 5059 1498 5093
rect 1452 5021 1498 5059
rect 1452 4987 1458 5021
rect 1492 4987 1498 5021
rect 1452 4949 1498 4987
rect 1452 4915 1458 4949
rect 1492 4915 1498 4949
rect 1452 4877 1498 4915
rect 1452 4843 1458 4877
rect 1492 4843 1498 4877
rect 1452 4805 1498 4843
rect 1452 4771 1458 4805
rect 1492 4771 1498 4805
rect 1452 4733 1498 4771
rect 1452 4699 1458 4733
rect 1492 4699 1498 4733
rect 1452 4661 1498 4699
rect 1452 4627 1458 4661
rect 1492 4627 1498 4661
rect 1452 4589 1498 4627
rect 1452 4555 1458 4589
rect 1492 4555 1498 4589
rect 1452 4517 1498 4555
rect 1452 4483 1458 4517
rect 1492 4483 1498 4517
rect 1452 4445 1498 4483
rect 1452 4411 1458 4445
rect 1492 4411 1498 4445
rect 1452 4373 1498 4411
rect 1452 4339 1458 4373
rect 1492 4339 1498 4373
rect 1452 4301 1498 4339
rect 1452 4267 1458 4301
rect 1492 4267 1498 4301
rect 1452 4229 1498 4267
rect 1452 4195 1458 4229
rect 1492 4195 1498 4229
rect 1452 4157 1498 4195
rect 1452 4123 1458 4157
rect 1492 4123 1498 4157
rect 1452 4085 1498 4123
rect 1452 4051 1458 4085
rect 1492 4051 1498 4085
rect 1452 4013 1498 4051
rect 1452 3979 1458 4013
rect 1492 3979 1498 4013
rect 1452 3941 1498 3979
rect 1452 3907 1458 3941
rect 1492 3907 1498 3941
rect 1452 3869 1498 3907
rect 1452 3835 1458 3869
rect 1492 3835 1498 3869
rect 1452 3797 1498 3835
rect 1452 3763 1458 3797
rect 1492 3763 1498 3797
rect 1452 3725 1498 3763
rect 1452 3691 1458 3725
rect 1492 3691 1498 3725
rect 1452 3653 1498 3691
rect 1452 3619 1458 3653
rect 1492 3619 1498 3653
rect 1452 3581 1498 3619
rect 1452 3547 1458 3581
rect 1492 3547 1498 3581
rect 1452 3509 1498 3547
rect 1452 3475 1458 3509
rect 1492 3475 1498 3509
rect 1452 3437 1498 3475
rect 1452 3403 1458 3437
rect 1492 3403 1498 3437
rect 1452 3365 1498 3403
rect 1452 3331 1458 3365
rect 1492 3331 1498 3365
rect 1452 3293 1498 3331
rect 1452 3259 1458 3293
rect 1492 3259 1498 3293
rect 1452 3221 1498 3259
rect 1452 3187 1458 3221
rect 1492 3187 1498 3221
rect 1452 3149 1498 3187
rect 1452 3115 1458 3149
rect 1492 3115 1498 3149
rect 1452 3077 1498 3115
rect 1452 3043 1458 3077
rect 1492 3043 1498 3077
rect 1452 3005 1498 3043
rect 1452 2971 1458 3005
rect 1492 2971 1498 3005
rect 1452 2933 1498 2971
rect 1452 2899 1458 2933
rect 1492 2899 1498 2933
rect 1452 2861 1498 2899
rect 1452 2827 1458 2861
rect 1492 2827 1498 2861
rect 1452 2789 1498 2827
rect 1452 2755 1458 2789
rect 1492 2755 1498 2789
rect 1452 2717 1498 2755
rect 1452 2683 1458 2717
rect 1492 2683 1498 2717
rect 1452 2645 1498 2683
rect 1452 2611 1458 2645
rect 1492 2611 1498 2645
rect 1452 2573 1498 2611
rect 1452 2539 1458 2573
rect 1492 2539 1498 2573
rect 1452 2501 1498 2539
rect 1452 2467 1458 2501
rect 1492 2467 1498 2501
rect 1452 2429 1498 2467
rect 1452 2395 1458 2429
rect 1492 2395 1498 2429
rect 1452 2357 1498 2395
rect 1452 2323 1458 2357
rect 1492 2323 1498 2357
rect 1452 2285 1498 2323
rect 1452 2251 1458 2285
rect 1492 2251 1498 2285
rect 1452 2213 1498 2251
rect 1452 2179 1458 2213
rect 1492 2179 1498 2213
rect 1452 2141 1498 2179
rect 1452 2107 1458 2141
rect 1492 2107 1498 2141
rect 1452 2069 1498 2107
rect 1452 2035 1458 2069
rect 1492 2035 1498 2069
rect 1452 1997 1498 2035
rect 1452 1963 1458 1997
rect 1492 1963 1498 1997
rect 1452 1925 1498 1963
rect 1452 1891 1458 1925
rect 1492 1891 1498 1925
rect 1452 1853 1498 1891
rect 1452 1819 1458 1853
rect 1492 1819 1498 1853
rect 1452 1781 1498 1819
rect 1452 1747 1458 1781
rect 1492 1747 1498 1781
rect 1452 1709 1498 1747
rect 1452 1675 1458 1709
rect 1492 1675 1498 1709
rect 1452 1637 1498 1675
rect 1452 1603 1458 1637
rect 1492 1603 1498 1637
rect 1452 1565 1498 1603
rect 1452 1531 1458 1565
rect 1492 1531 1498 1565
rect 1452 1493 1498 1531
rect 1452 1459 1458 1493
rect 1492 1459 1498 1493
rect 1452 1421 1498 1459
rect 1452 1387 1458 1421
rect 1492 1387 1498 1421
rect 1452 1349 1498 1387
rect 1452 1315 1458 1349
rect 1492 1315 1498 1349
rect 1452 1277 1498 1315
rect 1452 1243 1458 1277
rect 1492 1243 1498 1277
rect 1452 1205 1498 1243
rect 1452 1171 1458 1205
rect 1492 1171 1498 1205
rect 1452 1133 1498 1171
rect 1452 1099 1458 1133
rect 1492 1099 1498 1133
rect 1452 1061 1498 1099
rect 1452 1027 1458 1061
rect 1492 1027 1498 1061
rect 1452 989 1498 1027
rect 1452 955 1458 989
rect 1492 955 1498 989
rect 1452 917 1498 955
rect 1452 883 1458 917
rect 1492 883 1498 917
rect 1452 845 1498 883
rect 1452 811 1458 845
rect 1492 811 1498 845
rect 1452 773 1498 811
rect 1452 739 1458 773
rect 1492 739 1498 773
rect 1452 701 1498 739
rect 1452 667 1458 701
rect 1492 667 1498 701
rect 1452 629 1498 667
rect 1452 595 1458 629
rect 1492 595 1498 629
rect 1452 557 1498 595
rect 1452 523 1458 557
rect 1492 523 1498 557
rect 1452 485 1498 523
rect 1452 451 1458 485
rect 1492 451 1498 485
rect 1452 413 1498 451
rect 1452 379 1458 413
rect 1492 379 1498 413
rect 1452 341 1498 379
rect 1452 307 1458 341
rect 1492 307 1498 341
rect 1452 269 1498 307
rect 1452 235 1458 269
rect 1492 235 1498 269
rect 1452 197 1498 235
rect 1452 163 1458 197
rect 1492 163 1498 197
rect 1452 125 1498 163
rect 1452 91 1458 125
rect 1492 91 1498 125
rect 1452 53 1498 91
rect 1452 19 1458 53
rect 1492 19 1498 53
rect 1452 -19 1498 19
rect 1452 -53 1458 -19
rect 1492 -53 1498 -19
rect 1452 -91 1498 -53
rect 1452 -125 1458 -91
rect 1492 -125 1498 -91
rect 1452 -163 1498 -125
rect 1452 -197 1458 -163
rect 1492 -197 1498 -163
rect 1452 -235 1498 -197
rect 1452 -269 1458 -235
rect 1492 -269 1498 -235
rect 1452 -307 1498 -269
rect 1452 -341 1458 -307
rect 1492 -341 1498 -307
rect 1452 -379 1498 -341
rect 1452 -413 1458 -379
rect 1492 -413 1498 -379
rect 1452 -451 1498 -413
rect 1452 -485 1458 -451
rect 1492 -485 1498 -451
rect 1452 -523 1498 -485
rect 1452 -557 1458 -523
rect 1492 -557 1498 -523
rect 1452 -595 1498 -557
rect 1452 -629 1458 -595
rect 1492 -629 1498 -595
rect 1452 -667 1498 -629
rect 1452 -701 1458 -667
rect 1492 -701 1498 -667
rect 1452 -739 1498 -701
rect 1452 -773 1458 -739
rect 1492 -773 1498 -739
rect 1452 -811 1498 -773
rect 1452 -845 1458 -811
rect 1492 -845 1498 -811
rect 1452 -883 1498 -845
rect 1452 -917 1458 -883
rect 1492 -917 1498 -883
rect 1452 -955 1498 -917
rect 1452 -989 1458 -955
rect 1492 -989 1498 -955
rect 1452 -1027 1498 -989
rect 1452 -1061 1458 -1027
rect 1492 -1061 1498 -1027
rect 1452 -1099 1498 -1061
rect 1452 -1133 1458 -1099
rect 1492 -1133 1498 -1099
rect 1452 -1171 1498 -1133
rect 1452 -1205 1458 -1171
rect 1492 -1205 1498 -1171
rect 1452 -1243 1498 -1205
rect 1452 -1277 1458 -1243
rect 1492 -1277 1498 -1243
rect 1452 -1315 1498 -1277
rect 1452 -1349 1458 -1315
rect 1492 -1349 1498 -1315
rect 1452 -1387 1498 -1349
rect 1452 -1421 1458 -1387
rect 1492 -1421 1498 -1387
rect 1452 -1459 1498 -1421
rect 1452 -1493 1458 -1459
rect 1492 -1493 1498 -1459
rect 1452 -1531 1498 -1493
rect 1452 -1565 1458 -1531
rect 1492 -1565 1498 -1531
rect 1452 -1603 1498 -1565
rect 1452 -1637 1458 -1603
rect 1492 -1637 1498 -1603
rect 1452 -1675 1498 -1637
rect 1452 -1709 1458 -1675
rect 1492 -1709 1498 -1675
rect 1452 -1747 1498 -1709
rect 1452 -1781 1458 -1747
rect 1492 -1781 1498 -1747
rect 1452 -1819 1498 -1781
rect 1452 -1853 1458 -1819
rect 1492 -1853 1498 -1819
rect 1452 -1891 1498 -1853
rect 1452 -1925 1458 -1891
rect 1492 -1925 1498 -1891
rect 1452 -1963 1498 -1925
rect 1452 -1997 1458 -1963
rect 1492 -1997 1498 -1963
rect 1452 -2035 1498 -1997
rect 1452 -2069 1458 -2035
rect 1492 -2069 1498 -2035
rect 1452 -2107 1498 -2069
rect 1452 -2141 1458 -2107
rect 1492 -2141 1498 -2107
rect 1452 -2179 1498 -2141
rect 1452 -2213 1458 -2179
rect 1492 -2213 1498 -2179
rect 1452 -2251 1498 -2213
rect 1452 -2285 1458 -2251
rect 1492 -2285 1498 -2251
rect 1452 -2323 1498 -2285
rect 1452 -2357 1458 -2323
rect 1492 -2357 1498 -2323
rect 1452 -2395 1498 -2357
rect 1452 -2429 1458 -2395
rect 1492 -2429 1498 -2395
rect 1452 -2467 1498 -2429
rect 1452 -2501 1458 -2467
rect 1492 -2501 1498 -2467
rect 1452 -2539 1498 -2501
rect 1452 -2573 1458 -2539
rect 1492 -2573 1498 -2539
rect 1452 -2611 1498 -2573
rect 1452 -2645 1458 -2611
rect 1492 -2645 1498 -2611
rect 1452 -2683 1498 -2645
rect 1452 -2717 1458 -2683
rect 1492 -2717 1498 -2683
rect 1452 -2755 1498 -2717
rect 1452 -2789 1458 -2755
rect 1492 -2789 1498 -2755
rect 1452 -2827 1498 -2789
rect 1452 -2861 1458 -2827
rect 1492 -2861 1498 -2827
rect 1452 -2899 1498 -2861
rect 1452 -2933 1458 -2899
rect 1492 -2933 1498 -2899
rect 1452 -2971 1498 -2933
rect 1452 -3005 1458 -2971
rect 1492 -3005 1498 -2971
rect 1452 -3043 1498 -3005
rect 1452 -3077 1458 -3043
rect 1492 -3077 1498 -3043
rect 1452 -3115 1498 -3077
rect 1452 -3149 1458 -3115
rect 1492 -3149 1498 -3115
rect 1452 -3187 1498 -3149
rect 1452 -3221 1458 -3187
rect 1492 -3221 1498 -3187
rect 1452 -3259 1498 -3221
rect 1452 -3293 1458 -3259
rect 1492 -3293 1498 -3259
rect 1452 -3331 1498 -3293
rect 1452 -3365 1458 -3331
rect 1492 -3365 1498 -3331
rect 1452 -3403 1498 -3365
rect 1452 -3437 1458 -3403
rect 1492 -3437 1498 -3403
rect 1452 -3475 1498 -3437
rect 1452 -3509 1458 -3475
rect 1492 -3509 1498 -3475
rect 1452 -3547 1498 -3509
rect 1452 -3581 1458 -3547
rect 1492 -3581 1498 -3547
rect 1452 -3619 1498 -3581
rect 1452 -3653 1458 -3619
rect 1492 -3653 1498 -3619
rect 1452 -3691 1498 -3653
rect 1452 -3725 1458 -3691
rect 1492 -3725 1498 -3691
rect 1452 -3763 1498 -3725
rect 1452 -3797 1458 -3763
rect 1492 -3797 1498 -3763
rect 1452 -3835 1498 -3797
rect 1452 -3869 1458 -3835
rect 1492 -3869 1498 -3835
rect 1452 -3907 1498 -3869
rect 1452 -3941 1458 -3907
rect 1492 -3941 1498 -3907
rect 1452 -3979 1498 -3941
rect 1452 -4013 1458 -3979
rect 1492 -4013 1498 -3979
rect 1452 -4051 1498 -4013
rect 1452 -4085 1458 -4051
rect 1492 -4085 1498 -4051
rect 1452 -4123 1498 -4085
rect 1452 -4157 1458 -4123
rect 1492 -4157 1498 -4123
rect 1452 -4195 1498 -4157
rect 1452 -4229 1458 -4195
rect 1492 -4229 1498 -4195
rect 1452 -4267 1498 -4229
rect 1452 -4301 1458 -4267
rect 1492 -4301 1498 -4267
rect 1452 -4339 1498 -4301
rect 1452 -4373 1458 -4339
rect 1492 -4373 1498 -4339
rect 1452 -4411 1498 -4373
rect 1452 -4445 1458 -4411
rect 1492 -4445 1498 -4411
rect 1452 -4483 1498 -4445
rect 1452 -4517 1458 -4483
rect 1492 -4517 1498 -4483
rect 1452 -4555 1498 -4517
rect 1452 -4589 1458 -4555
rect 1492 -4589 1498 -4555
rect 1452 -4627 1498 -4589
rect 1452 -4661 1458 -4627
rect 1492 -4661 1498 -4627
rect 1452 -4699 1498 -4661
rect 1452 -4733 1458 -4699
rect 1492 -4733 1498 -4699
rect 1452 -4771 1498 -4733
rect 1452 -4805 1458 -4771
rect 1492 -4805 1498 -4771
rect 1452 -4843 1498 -4805
rect 1452 -4877 1458 -4843
rect 1492 -4877 1498 -4843
rect 1452 -4915 1498 -4877
rect 1452 -4949 1458 -4915
rect 1492 -4949 1498 -4915
rect 1452 -4987 1498 -4949
rect 1452 -5021 1458 -4987
rect 1492 -5021 1498 -4987
rect 1452 -5059 1498 -5021
rect 1452 -5093 1458 -5059
rect 1492 -5093 1498 -5059
rect 1452 -5131 1498 -5093
rect 1452 -5165 1458 -5131
rect 1492 -5165 1498 -5131
rect 1452 -5203 1498 -5165
rect 1452 -5237 1458 -5203
rect 1492 -5237 1498 -5203
rect 1452 -5275 1498 -5237
rect 1452 -5309 1458 -5275
rect 1492 -5309 1498 -5275
rect 1452 -5347 1498 -5309
rect 1452 -5381 1458 -5347
rect 1492 -5381 1498 -5347
rect 1452 -5419 1498 -5381
rect 1452 -5453 1458 -5419
rect 1492 -5453 1498 -5419
rect 1452 -5491 1498 -5453
rect 1452 -5525 1458 -5491
rect 1492 -5525 1498 -5491
rect 1452 -5563 1498 -5525
rect 1452 -5597 1458 -5563
rect 1492 -5597 1498 -5563
rect 1452 -5635 1498 -5597
rect 1452 -5669 1458 -5635
rect 1492 -5669 1498 -5635
rect 1452 -5707 1498 -5669
rect 1452 -5741 1458 -5707
rect 1492 -5741 1498 -5707
rect 1452 -5779 1498 -5741
rect 1452 -5813 1458 -5779
rect 1492 -5813 1498 -5779
rect 1452 -5851 1498 -5813
rect 1452 -5885 1458 -5851
rect 1492 -5885 1498 -5851
rect 1452 -5923 1498 -5885
rect 1452 -5957 1458 -5923
rect 1492 -5957 1498 -5923
rect 1452 -5995 1498 -5957
rect 1452 -6029 1458 -5995
rect 1492 -6029 1498 -5995
rect 1452 -6067 1498 -6029
rect 1452 -6101 1458 -6067
rect 1492 -6101 1498 -6067
rect 1452 -6139 1498 -6101
rect 1452 -6173 1458 -6139
rect 1492 -6173 1498 -6139
rect 1452 -6211 1498 -6173
rect 1452 -6245 1458 -6211
rect 1492 -6245 1498 -6211
rect 1452 -6283 1498 -6245
rect 1452 -6317 1458 -6283
rect 1492 -6317 1498 -6283
rect 1452 -6355 1498 -6317
rect 1452 -6389 1458 -6355
rect 1492 -6389 1498 -6355
rect 1452 -6427 1498 -6389
rect 1452 -6461 1458 -6427
rect 1492 -6461 1498 -6427
rect 1452 -6499 1498 -6461
rect 1452 -6533 1458 -6499
rect 1492 -6533 1498 -6499
rect 1452 -6571 1498 -6533
rect 1452 -6605 1458 -6571
rect 1492 -6605 1498 -6571
rect 1452 -6643 1498 -6605
rect 1452 -6677 1458 -6643
rect 1492 -6677 1498 -6643
rect 1452 -6715 1498 -6677
rect 1452 -6749 1458 -6715
rect 1492 -6749 1498 -6715
rect 1452 -6787 1498 -6749
rect 1452 -6821 1458 -6787
rect 1492 -6821 1498 -6787
rect 1452 -6859 1498 -6821
rect 1452 -6893 1458 -6859
rect 1492 -6893 1498 -6859
rect 1452 -6931 1498 -6893
rect 1452 -6965 1458 -6931
rect 1492 -6965 1498 -6931
rect 1452 -7003 1498 -6965
rect 1452 -7037 1458 -7003
rect 1492 -7037 1498 -7003
rect 1452 -7075 1498 -7037
rect 1452 -7109 1458 -7075
rect 1492 -7109 1498 -7075
rect 1452 -7147 1498 -7109
rect 1452 -7181 1458 -7147
rect 1492 -7181 1498 -7147
rect 1452 -7219 1498 -7181
rect 1452 -7253 1458 -7219
rect 1492 -7253 1498 -7219
rect 1452 -7291 1498 -7253
rect 1452 -7325 1458 -7291
rect 1492 -7325 1498 -7291
rect 1452 -7363 1498 -7325
rect 1452 -7397 1458 -7363
rect 1492 -7397 1498 -7363
rect 1452 -7435 1498 -7397
rect 1452 -7469 1458 -7435
rect 1492 -7469 1498 -7435
rect 1452 -7507 1498 -7469
rect 1452 -7541 1458 -7507
rect 1492 -7541 1498 -7507
rect 1452 -7579 1498 -7541
rect 1452 -7613 1458 -7579
rect 1492 -7613 1498 -7579
rect 1452 -7651 1498 -7613
rect 1452 -7685 1458 -7651
rect 1492 -7685 1498 -7651
rect 1452 -7723 1498 -7685
rect 1452 -7757 1458 -7723
rect 1492 -7757 1498 -7723
rect 1452 -7795 1498 -7757
rect 1452 -7829 1458 -7795
rect 1492 -7829 1498 -7795
rect 1452 -7867 1498 -7829
rect 1452 -7901 1458 -7867
rect 1492 -7901 1498 -7867
rect 1452 -7939 1498 -7901
rect 1452 -7973 1458 -7939
rect 1492 -7973 1498 -7939
rect 1452 -8011 1498 -7973
rect 1452 -8045 1458 -8011
rect 1492 -8045 1498 -8011
rect 1452 -8083 1498 -8045
rect 1452 -8117 1458 -8083
rect 1492 -8117 1498 -8083
rect 1452 -8155 1498 -8117
rect 1452 -8189 1458 -8155
rect 1492 -8189 1498 -8155
rect 1452 -8227 1498 -8189
rect 1452 -8261 1458 -8227
rect 1492 -8261 1498 -8227
rect 1452 -8299 1498 -8261
rect 1452 -8333 1458 -8299
rect 1492 -8333 1498 -8299
rect 1452 -8371 1498 -8333
rect 1452 -8405 1458 -8371
rect 1492 -8405 1498 -8371
rect 1452 -8443 1498 -8405
rect 1452 -8477 1458 -8443
rect 1492 -8477 1498 -8443
rect 1452 -8515 1498 -8477
rect 1452 -8549 1458 -8515
rect 1492 -8549 1498 -8515
rect 1452 -8587 1498 -8549
rect 1452 -8621 1458 -8587
rect 1492 -8621 1498 -8587
rect 1452 -8659 1498 -8621
rect 1452 -8693 1458 -8659
rect 1492 -8693 1498 -8659
rect 1452 -8731 1498 -8693
rect 1452 -8765 1458 -8731
rect 1492 -8765 1498 -8731
rect 1452 -8803 1498 -8765
rect 1452 -8837 1458 -8803
rect 1492 -8837 1498 -8803
rect 1452 -8875 1498 -8837
rect 1452 -8909 1458 -8875
rect 1492 -8909 1498 -8875
rect 1452 -8947 1498 -8909
rect 1452 -8981 1458 -8947
rect 1492 -8981 1498 -8947
rect 1452 -9019 1498 -8981
rect 1452 -9053 1458 -9019
rect 1492 -9053 1498 -9019
rect 1452 -9091 1498 -9053
rect 1452 -9125 1458 -9091
rect 1492 -9125 1498 -9091
rect 1452 -9163 1498 -9125
rect 1452 -9197 1458 -9163
rect 1492 -9197 1498 -9163
rect 1452 -9235 1498 -9197
rect 1452 -9269 1458 -9235
rect 1492 -9269 1498 -9235
rect 1452 -9307 1498 -9269
rect 1452 -9341 1458 -9307
rect 1492 -9341 1498 -9307
rect 1452 -9379 1498 -9341
rect 1452 -9413 1458 -9379
rect 1492 -9413 1498 -9379
rect 1452 -9451 1498 -9413
rect 1452 -9485 1458 -9451
rect 1492 -9485 1498 -9451
rect 1452 -9523 1498 -9485
rect 1452 -9557 1458 -9523
rect 1492 -9557 1498 -9523
rect 1452 -9600 1498 -9557
<< end >>
