magic
tech sky130A
timestamp 1666811438
<< error_p >>
rect -16 939 16 942
rect -16 922 -10 939
rect -16 919 16 922
rect -16 -922 16 -919
rect -16 -939 -10 -922
rect -16 -942 16 -939
<< nmos >>
rect -18 -903 18 903
<< ndiff >>
rect -47 897 -18 903
rect -47 -897 -41 897
rect -24 -897 -18 897
rect -47 -903 -18 -897
rect 18 897 47 903
rect 18 -897 24 897
rect 41 -897 47 897
rect 18 -903 47 -897
<< ndiffc >>
rect -41 -897 -24 897
rect 24 -897 41 897
<< poly >>
rect -18 939 18 947
rect -18 922 -10 939
rect 10 922 18 939
rect -18 903 18 922
rect -18 -922 18 -903
rect -18 -939 -10 -922
rect 10 -939 18 -922
rect -18 -947 18 -939
<< polycont >>
rect -10 922 10 939
rect -10 -939 10 -922
<< locali >>
rect -18 922 -10 939
rect 10 922 18 939
rect -41 897 -24 905
rect -41 -905 -24 -897
rect 24 897 41 905
rect 24 -905 41 -897
rect -18 -939 -10 -922
rect 10 -939 18 -922
<< viali >>
rect -10 922 10 939
rect -41 -897 -24 897
rect 24 -897 41 897
rect -10 -939 10 -922
<< metal1 >>
rect -16 939 16 942
rect -16 922 -10 939
rect 10 922 16 939
rect -16 919 16 922
rect -44 897 -21 903
rect -44 -897 -41 897
rect -24 -897 -21 897
rect -44 -903 -21 -897
rect 21 897 44 903
rect 21 -897 24 897
rect 41 -897 44 897
rect 21 -903 44 -897
rect -16 -922 16 -919
rect -16 -939 -10 -922
rect 10 -939 16 -922
rect -16 -942 16 -939
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 18.055 l 0.361 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
