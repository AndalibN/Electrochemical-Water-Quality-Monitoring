magic
tech sky130A
magscale 1 2
timestamp 1668032717
<< xpolycontact >>
rect -35 2457 35 2889
rect -35 -2889 35 -2457
<< xpolyres >>
rect -35 -2457 35 2457
<< viali >>
rect -19 2474 19 2871
rect -19 -2871 19 -2474
<< metal1 >>
rect -25 2871 25 2883
rect -25 2474 -19 2871
rect 19 2474 25 2871
rect -25 2462 25 2474
rect -25 -2474 25 -2462
rect -25 -2871 -19 -2474
rect 19 -2871 25 -2474
rect -25 -2883 25 -2871
<< res0p35 >>
rect -37 -2459 37 2459
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 24.57 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 141.475k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
