magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 2457 35 2889
rect -35 -2889 35 -2457
<< xpolyres >>
rect -35 -2457 35 2457
<< viali >>
rect -17 2835 17 2869
rect -17 2763 17 2797
rect -17 2691 17 2725
rect -17 2619 17 2653
rect -17 2547 17 2581
rect -17 2475 17 2509
rect -17 -2510 17 -2476
rect -17 -2582 17 -2548
rect -17 -2654 17 -2620
rect -17 -2726 17 -2692
rect -17 -2798 17 -2764
rect -17 -2870 17 -2836
<< metal1 >>
rect -25 2869 25 2883
rect -25 2835 -17 2869
rect 17 2835 25 2869
rect -25 2797 25 2835
rect -25 2763 -17 2797
rect 17 2763 25 2797
rect -25 2725 25 2763
rect -25 2691 -17 2725
rect 17 2691 25 2725
rect -25 2653 25 2691
rect -25 2619 -17 2653
rect 17 2619 25 2653
rect -25 2581 25 2619
rect -25 2547 -17 2581
rect 17 2547 25 2581
rect -25 2509 25 2547
rect -25 2475 -17 2509
rect 17 2475 25 2509
rect -25 2462 25 2475
rect -25 -2476 25 -2462
rect -25 -2510 -17 -2476
rect 17 -2510 25 -2476
rect -25 -2548 25 -2510
rect -25 -2582 -17 -2548
rect 17 -2582 25 -2548
rect -25 -2620 25 -2582
rect -25 -2654 -17 -2620
rect 17 -2654 25 -2620
rect -25 -2692 25 -2654
rect -25 -2726 -17 -2692
rect 17 -2726 25 -2692
rect -25 -2764 25 -2726
rect -25 -2798 -17 -2764
rect 17 -2798 25 -2764
rect -25 -2836 25 -2798
rect -25 -2870 -17 -2836
rect 17 -2870 25 -2836
rect -25 -2883 25 -2870
<< end >>
