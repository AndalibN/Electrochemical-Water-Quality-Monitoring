magic
tech sky130A
magscale 1 2
timestamp 1668369016
<< error_p >>
rect -1073 6072 -1015 6078
rect -841 6072 -783 6078
rect -609 6072 -551 6078
rect -377 6072 -319 6078
rect -145 6072 -87 6078
rect 87 6072 145 6078
rect 319 6072 377 6078
rect 551 6072 609 6078
rect 783 6072 841 6078
rect 1015 6072 1073 6078
rect -1073 6038 -1061 6072
rect -841 6038 -829 6072
rect -609 6038 -597 6072
rect -377 6038 -365 6072
rect -145 6038 -133 6072
rect 87 6038 99 6072
rect 319 6038 331 6072
rect 551 6038 563 6072
rect 783 6038 795 6072
rect 1015 6038 1027 6072
rect -1073 6032 -1015 6038
rect -841 6032 -783 6038
rect -609 6032 -551 6038
rect -377 6032 -319 6038
rect -145 6032 -87 6038
rect 87 6032 145 6038
rect 319 6032 377 6038
rect 551 6032 609 6038
rect 783 6032 841 6038
rect 1015 6032 1073 6038
rect -1073 -6038 -1015 -6032
rect -841 -6038 -783 -6032
rect -609 -6038 -551 -6032
rect -377 -6038 -319 -6032
rect -145 -6038 -87 -6032
rect 87 -6038 145 -6032
rect 319 -6038 377 -6032
rect 551 -6038 609 -6032
rect 783 -6038 841 -6032
rect 1015 -6038 1073 -6032
rect -1073 -6072 -1061 -6038
rect -841 -6072 -829 -6038
rect -609 -6072 -597 -6038
rect -377 -6072 -365 -6038
rect -145 -6072 -133 -6038
rect 87 -6072 99 -6038
rect 319 -6072 331 -6038
rect 551 -6072 563 -6038
rect 783 -6072 795 -6038
rect 1015 -6072 1027 -6038
rect -1073 -6078 -1015 -6072
rect -841 -6078 -783 -6072
rect -609 -6078 -551 -6072
rect -377 -6078 -319 -6072
rect -145 -6078 -87 -6072
rect 87 -6078 145 -6072
rect 319 -6078 377 -6072
rect 551 -6078 609 -6072
rect 783 -6078 841 -6072
rect 1015 -6078 1073 -6072
<< nmos >>
rect -1074 -6000 -1014 6000
rect -842 -6000 -782 6000
rect -610 -6000 -550 6000
rect -378 -6000 -318 6000
rect -146 -6000 -86 6000
rect 86 -6000 146 6000
rect 318 -6000 378 6000
rect 550 -6000 610 6000
rect 782 -6000 842 6000
rect 1014 -6000 1074 6000
<< ndiff >>
rect -1132 5988 -1074 6000
rect -1132 -5988 -1120 5988
rect -1086 -5988 -1074 5988
rect -1132 -6000 -1074 -5988
rect -1014 5988 -956 6000
rect -1014 -5988 -1002 5988
rect -968 -5988 -956 5988
rect -1014 -6000 -956 -5988
rect -900 5988 -842 6000
rect -900 -5988 -888 5988
rect -854 -5988 -842 5988
rect -900 -6000 -842 -5988
rect -782 5988 -724 6000
rect -782 -5988 -770 5988
rect -736 -5988 -724 5988
rect -782 -6000 -724 -5988
rect -668 5988 -610 6000
rect -668 -5988 -656 5988
rect -622 -5988 -610 5988
rect -668 -6000 -610 -5988
rect -550 5988 -492 6000
rect -550 -5988 -538 5988
rect -504 -5988 -492 5988
rect -550 -6000 -492 -5988
rect -436 5988 -378 6000
rect -436 -5988 -424 5988
rect -390 -5988 -378 5988
rect -436 -6000 -378 -5988
rect -318 5988 -260 6000
rect -318 -5988 -306 5988
rect -272 -5988 -260 5988
rect -318 -6000 -260 -5988
rect -204 5988 -146 6000
rect -204 -5988 -192 5988
rect -158 -5988 -146 5988
rect -204 -6000 -146 -5988
rect -86 5988 -28 6000
rect -86 -5988 -74 5988
rect -40 -5988 -28 5988
rect -86 -6000 -28 -5988
rect 28 5988 86 6000
rect 28 -5988 40 5988
rect 74 -5988 86 5988
rect 28 -6000 86 -5988
rect 146 5988 204 6000
rect 146 -5988 158 5988
rect 192 -5988 204 5988
rect 146 -6000 204 -5988
rect 260 5988 318 6000
rect 260 -5988 272 5988
rect 306 -5988 318 5988
rect 260 -6000 318 -5988
rect 378 5988 436 6000
rect 378 -5988 390 5988
rect 424 -5988 436 5988
rect 378 -6000 436 -5988
rect 492 5988 550 6000
rect 492 -5988 504 5988
rect 538 -5988 550 5988
rect 492 -6000 550 -5988
rect 610 5988 668 6000
rect 610 -5988 622 5988
rect 656 -5988 668 5988
rect 610 -6000 668 -5988
rect 724 5988 782 6000
rect 724 -5988 736 5988
rect 770 -5988 782 5988
rect 724 -6000 782 -5988
rect 842 5988 900 6000
rect 842 -5988 854 5988
rect 888 -5988 900 5988
rect 842 -6000 900 -5988
rect 956 5988 1014 6000
rect 956 -5988 968 5988
rect 1002 -5988 1014 5988
rect 956 -6000 1014 -5988
rect 1074 5988 1132 6000
rect 1074 -5988 1086 5988
rect 1120 -5988 1132 5988
rect 1074 -6000 1132 -5988
<< ndiffc >>
rect -1120 -5988 -1086 5988
rect -1002 -5988 -968 5988
rect -888 -5988 -854 5988
rect -770 -5988 -736 5988
rect -656 -5988 -622 5988
rect -538 -5988 -504 5988
rect -424 -5988 -390 5988
rect -306 -5988 -272 5988
rect -192 -5988 -158 5988
rect -74 -5988 -40 5988
rect 40 -5988 74 5988
rect 158 -5988 192 5988
rect 272 -5988 306 5988
rect 390 -5988 424 5988
rect 504 -5988 538 5988
rect 622 -5988 656 5988
rect 736 -5988 770 5988
rect 854 -5988 888 5988
rect 968 -5988 1002 5988
rect 1086 -5988 1120 5988
<< poly >>
rect -1077 6072 -1011 6088
rect -1077 6038 -1061 6072
rect -1027 6038 -1011 6072
rect -1077 6022 -1011 6038
rect -845 6072 -779 6088
rect -845 6038 -829 6072
rect -795 6038 -779 6072
rect -845 6022 -779 6038
rect -613 6072 -547 6088
rect -613 6038 -597 6072
rect -563 6038 -547 6072
rect -613 6022 -547 6038
rect -381 6072 -315 6088
rect -381 6038 -365 6072
rect -331 6038 -315 6072
rect -381 6022 -315 6038
rect -149 6072 -83 6088
rect -149 6038 -133 6072
rect -99 6038 -83 6072
rect -149 6022 -83 6038
rect 83 6072 149 6088
rect 83 6038 99 6072
rect 133 6038 149 6072
rect 83 6022 149 6038
rect 315 6072 381 6088
rect 315 6038 331 6072
rect 365 6038 381 6072
rect 315 6022 381 6038
rect 547 6072 613 6088
rect 547 6038 563 6072
rect 597 6038 613 6072
rect 547 6022 613 6038
rect 779 6072 845 6088
rect 779 6038 795 6072
rect 829 6038 845 6072
rect 779 6022 845 6038
rect 1011 6072 1077 6088
rect 1011 6038 1027 6072
rect 1061 6038 1077 6072
rect 1011 6022 1077 6038
rect -1074 6000 -1014 6022
rect -842 6000 -782 6022
rect -610 6000 -550 6022
rect -378 6000 -318 6022
rect -146 6000 -86 6022
rect 86 6000 146 6022
rect 318 6000 378 6022
rect 550 6000 610 6022
rect 782 6000 842 6022
rect 1014 6000 1074 6022
rect -1074 -6022 -1014 -6000
rect -842 -6022 -782 -6000
rect -610 -6022 -550 -6000
rect -378 -6022 -318 -6000
rect -146 -6022 -86 -6000
rect 86 -6022 146 -6000
rect 318 -6022 378 -6000
rect 550 -6022 610 -6000
rect 782 -6022 842 -6000
rect 1014 -6022 1074 -6000
rect -1077 -6038 -1011 -6022
rect -1077 -6072 -1061 -6038
rect -1027 -6072 -1011 -6038
rect -1077 -6088 -1011 -6072
rect -845 -6038 -779 -6022
rect -845 -6072 -829 -6038
rect -795 -6072 -779 -6038
rect -845 -6088 -779 -6072
rect -613 -6038 -547 -6022
rect -613 -6072 -597 -6038
rect -563 -6072 -547 -6038
rect -613 -6088 -547 -6072
rect -381 -6038 -315 -6022
rect -381 -6072 -365 -6038
rect -331 -6072 -315 -6038
rect -381 -6088 -315 -6072
rect -149 -6038 -83 -6022
rect -149 -6072 -133 -6038
rect -99 -6072 -83 -6038
rect -149 -6088 -83 -6072
rect 83 -6038 149 -6022
rect 83 -6072 99 -6038
rect 133 -6072 149 -6038
rect 83 -6088 149 -6072
rect 315 -6038 381 -6022
rect 315 -6072 331 -6038
rect 365 -6072 381 -6038
rect 315 -6088 381 -6072
rect 547 -6038 613 -6022
rect 547 -6072 563 -6038
rect 597 -6072 613 -6038
rect 547 -6088 613 -6072
rect 779 -6038 845 -6022
rect 779 -6072 795 -6038
rect 829 -6072 845 -6038
rect 779 -6088 845 -6072
rect 1011 -6038 1077 -6022
rect 1011 -6072 1027 -6038
rect 1061 -6072 1077 -6038
rect 1011 -6088 1077 -6072
<< polycont >>
rect -1061 6038 -1027 6072
rect -829 6038 -795 6072
rect -597 6038 -563 6072
rect -365 6038 -331 6072
rect -133 6038 -99 6072
rect 99 6038 133 6072
rect 331 6038 365 6072
rect 563 6038 597 6072
rect 795 6038 829 6072
rect 1027 6038 1061 6072
rect -1061 -6072 -1027 -6038
rect -829 -6072 -795 -6038
rect -597 -6072 -563 -6038
rect -365 -6072 -331 -6038
rect -133 -6072 -99 -6038
rect 99 -6072 133 -6038
rect 331 -6072 365 -6038
rect 563 -6072 597 -6038
rect 795 -6072 829 -6038
rect 1027 -6072 1061 -6038
<< locali >>
rect -1077 6038 -1061 6072
rect -1027 6038 -1011 6072
rect -845 6038 -829 6072
rect -795 6038 -779 6072
rect -613 6038 -597 6072
rect -563 6038 -547 6072
rect -381 6038 -365 6072
rect -331 6038 -315 6072
rect -149 6038 -133 6072
rect -99 6038 -83 6072
rect 83 6038 99 6072
rect 133 6038 149 6072
rect 315 6038 331 6072
rect 365 6038 381 6072
rect 547 6038 563 6072
rect 597 6038 613 6072
rect 779 6038 795 6072
rect 829 6038 845 6072
rect 1011 6038 1027 6072
rect 1061 6038 1077 6072
rect -1120 5988 -1086 6004
rect -1120 -6004 -1086 -5988
rect -1002 5988 -968 6004
rect -1002 -6004 -968 -5988
rect -888 5988 -854 6004
rect -888 -6004 -854 -5988
rect -770 5988 -736 6004
rect -770 -6004 -736 -5988
rect -656 5988 -622 6004
rect -656 -6004 -622 -5988
rect -538 5988 -504 6004
rect -538 -6004 -504 -5988
rect -424 5988 -390 6004
rect -424 -6004 -390 -5988
rect -306 5988 -272 6004
rect -306 -6004 -272 -5988
rect -192 5988 -158 6004
rect -192 -6004 -158 -5988
rect -74 5988 -40 6004
rect -74 -6004 -40 -5988
rect 40 5988 74 6004
rect 40 -6004 74 -5988
rect 158 5988 192 6004
rect 158 -6004 192 -5988
rect 272 5988 306 6004
rect 272 -6004 306 -5988
rect 390 5988 424 6004
rect 390 -6004 424 -5988
rect 504 5988 538 6004
rect 504 -6004 538 -5988
rect 622 5988 656 6004
rect 622 -6004 656 -5988
rect 736 5988 770 6004
rect 736 -6004 770 -5988
rect 854 5988 888 6004
rect 854 -6004 888 -5988
rect 968 5988 1002 6004
rect 968 -6004 1002 -5988
rect 1086 5988 1120 6004
rect 1086 -6004 1120 -5988
rect -1077 -6072 -1061 -6038
rect -1027 -6072 -1011 -6038
rect -845 -6072 -829 -6038
rect -795 -6072 -779 -6038
rect -613 -6072 -597 -6038
rect -563 -6072 -547 -6038
rect -381 -6072 -365 -6038
rect -331 -6072 -315 -6038
rect -149 -6072 -133 -6038
rect -99 -6072 -83 -6038
rect 83 -6072 99 -6038
rect 133 -6072 149 -6038
rect 315 -6072 331 -6038
rect 365 -6072 381 -6038
rect 547 -6072 563 -6038
rect 597 -6072 613 -6038
rect 779 -6072 795 -6038
rect 829 -6072 845 -6038
rect 1011 -6072 1027 -6038
rect 1061 -6072 1077 -6038
<< viali >>
rect -1061 6038 -1027 6072
rect -829 6038 -795 6072
rect -597 6038 -563 6072
rect -365 6038 -331 6072
rect -133 6038 -99 6072
rect 99 6038 133 6072
rect 331 6038 365 6072
rect 563 6038 597 6072
rect 795 6038 829 6072
rect 1027 6038 1061 6072
rect -1120 -5988 -1086 5988
rect -1002 -5988 -968 5988
rect -888 -5988 -854 5988
rect -770 -5988 -736 5988
rect -656 -5988 -622 5988
rect -538 -5988 -504 5988
rect -424 -5988 -390 5988
rect -306 -5988 -272 5988
rect -192 -5988 -158 5988
rect -74 -5988 -40 5988
rect 40 -5988 74 5988
rect 158 -5988 192 5988
rect 272 -5988 306 5988
rect 390 -5988 424 5988
rect 504 -5988 538 5988
rect 622 -5988 656 5988
rect 736 -5988 770 5988
rect 854 -5988 888 5988
rect 968 -5988 1002 5988
rect 1086 -5988 1120 5988
rect -1061 -6072 -1027 -6038
rect -829 -6072 -795 -6038
rect -597 -6072 -563 -6038
rect -365 -6072 -331 -6038
rect -133 -6072 -99 -6038
rect 99 -6072 133 -6038
rect 331 -6072 365 -6038
rect 563 -6072 597 -6038
rect 795 -6072 829 -6038
rect 1027 -6072 1061 -6038
<< metal1 >>
rect -1073 6072 -1015 6078
rect -1073 6038 -1061 6072
rect -1027 6038 -1015 6072
rect -1073 6032 -1015 6038
rect -841 6072 -783 6078
rect -841 6038 -829 6072
rect -795 6038 -783 6072
rect -841 6032 -783 6038
rect -609 6072 -551 6078
rect -609 6038 -597 6072
rect -563 6038 -551 6072
rect -609 6032 -551 6038
rect -377 6072 -319 6078
rect -377 6038 -365 6072
rect -331 6038 -319 6072
rect -377 6032 -319 6038
rect -145 6072 -87 6078
rect -145 6038 -133 6072
rect -99 6038 -87 6072
rect -145 6032 -87 6038
rect 87 6072 145 6078
rect 87 6038 99 6072
rect 133 6038 145 6072
rect 87 6032 145 6038
rect 319 6072 377 6078
rect 319 6038 331 6072
rect 365 6038 377 6072
rect 319 6032 377 6038
rect 551 6072 609 6078
rect 551 6038 563 6072
rect 597 6038 609 6072
rect 551 6032 609 6038
rect 783 6072 841 6078
rect 783 6038 795 6072
rect 829 6038 841 6072
rect 783 6032 841 6038
rect 1015 6072 1073 6078
rect 1015 6038 1027 6072
rect 1061 6038 1073 6072
rect 1015 6032 1073 6038
rect -1126 5988 -1080 6000
rect -1126 -5988 -1120 5988
rect -1086 -5988 -1080 5988
rect -1126 -6000 -1080 -5988
rect -1008 5988 -962 6000
rect -1008 -5988 -1002 5988
rect -968 -5988 -962 5988
rect -1008 -6000 -962 -5988
rect -894 5988 -848 6000
rect -894 -5988 -888 5988
rect -854 -5988 -848 5988
rect -894 -6000 -848 -5988
rect -776 5988 -730 6000
rect -776 -5988 -770 5988
rect -736 -5988 -730 5988
rect -776 -6000 -730 -5988
rect -662 5988 -616 6000
rect -662 -5988 -656 5988
rect -622 -5988 -616 5988
rect -662 -6000 -616 -5988
rect -544 5988 -498 6000
rect -544 -5988 -538 5988
rect -504 -5988 -498 5988
rect -544 -6000 -498 -5988
rect -430 5988 -384 6000
rect -430 -5988 -424 5988
rect -390 -5988 -384 5988
rect -430 -6000 -384 -5988
rect -312 5988 -266 6000
rect -312 -5988 -306 5988
rect -272 -5988 -266 5988
rect -312 -6000 -266 -5988
rect -198 5988 -152 6000
rect -198 -5988 -192 5988
rect -158 -5988 -152 5988
rect -198 -6000 -152 -5988
rect -80 5988 -34 6000
rect -80 -5988 -74 5988
rect -40 -5988 -34 5988
rect -80 -6000 -34 -5988
rect 34 5988 80 6000
rect 34 -5988 40 5988
rect 74 -5988 80 5988
rect 34 -6000 80 -5988
rect 152 5988 198 6000
rect 152 -5988 158 5988
rect 192 -5988 198 5988
rect 152 -6000 198 -5988
rect 266 5988 312 6000
rect 266 -5988 272 5988
rect 306 -5988 312 5988
rect 266 -6000 312 -5988
rect 384 5988 430 6000
rect 384 -5988 390 5988
rect 424 -5988 430 5988
rect 384 -6000 430 -5988
rect 498 5988 544 6000
rect 498 -5988 504 5988
rect 538 -5988 544 5988
rect 498 -6000 544 -5988
rect 616 5988 662 6000
rect 616 -5988 622 5988
rect 656 -5988 662 5988
rect 616 -6000 662 -5988
rect 730 5988 776 6000
rect 730 -5988 736 5988
rect 770 -5988 776 5988
rect 730 -6000 776 -5988
rect 848 5988 894 6000
rect 848 -5988 854 5988
rect 888 -5988 894 5988
rect 848 -6000 894 -5988
rect 962 5988 1008 6000
rect 962 -5988 968 5988
rect 1002 -5988 1008 5988
rect 962 -6000 1008 -5988
rect 1080 5988 1126 6000
rect 1080 -5988 1086 5988
rect 1120 -5988 1126 5988
rect 1080 -6000 1126 -5988
rect -1073 -6038 -1015 -6032
rect -1073 -6072 -1061 -6038
rect -1027 -6072 -1015 -6038
rect -1073 -6078 -1015 -6072
rect -841 -6038 -783 -6032
rect -841 -6072 -829 -6038
rect -795 -6072 -783 -6038
rect -841 -6078 -783 -6072
rect -609 -6038 -551 -6032
rect -609 -6072 -597 -6038
rect -563 -6072 -551 -6038
rect -609 -6078 -551 -6072
rect -377 -6038 -319 -6032
rect -377 -6072 -365 -6038
rect -331 -6072 -319 -6038
rect -377 -6078 -319 -6072
rect -145 -6038 -87 -6032
rect -145 -6072 -133 -6038
rect -99 -6072 -87 -6038
rect -145 -6078 -87 -6072
rect 87 -6038 145 -6032
rect 87 -6072 99 -6038
rect 133 -6072 145 -6038
rect 87 -6078 145 -6072
rect 319 -6038 377 -6032
rect 319 -6072 331 -6038
rect 365 -6072 377 -6038
rect 319 -6078 377 -6072
rect 551 -6038 609 -6032
rect 551 -6072 563 -6038
rect 597 -6072 609 -6038
rect 551 -6078 609 -6072
rect 783 -6038 841 -6032
rect 783 -6072 795 -6038
rect 829 -6072 841 -6038
rect 783 -6078 841 -6072
rect 1015 -6038 1073 -6032
rect 1015 -6072 1027 -6038
rect 1061 -6072 1073 -6038
rect 1015 -6078 1073 -6072
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 60 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
