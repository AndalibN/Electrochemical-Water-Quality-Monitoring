magic
tech sky130A
magscale 1 2
timestamp 1666625676
<< xpolycontact >>
rect -3851 190 -3781 622
rect -3851 -622 -3781 -190
rect -3533 190 -3463 622
rect -3533 -622 -3463 -190
rect -3215 190 -3145 622
rect -3215 -622 -3145 -190
rect -2897 190 -2827 622
rect -2897 -622 -2827 -190
rect -2579 190 -2509 622
rect -2579 -622 -2509 -190
rect -2261 190 -2191 622
rect -2261 -622 -2191 -190
rect -1943 190 -1873 622
rect -1943 -622 -1873 -190
rect -1625 190 -1555 622
rect -1625 -622 -1555 -190
rect -1307 190 -1237 622
rect -1307 -622 -1237 -190
rect -989 190 -919 622
rect -989 -622 -919 -190
rect -671 190 -601 622
rect -671 -622 -601 -190
rect -353 190 -283 622
rect -353 -622 -283 -190
rect -35 190 35 622
rect -35 -622 35 -190
rect 283 190 353 622
rect 283 -622 353 -190
rect 601 190 671 622
rect 601 -622 671 -190
rect 919 190 989 622
rect 919 -622 989 -190
rect 1237 190 1307 622
rect 1237 -622 1307 -190
rect 1555 190 1625 622
rect 1555 -622 1625 -190
rect 1873 190 1943 622
rect 1873 -622 1943 -190
rect 2191 190 2261 622
rect 2191 -622 2261 -190
rect 2509 190 2579 622
rect 2509 -622 2579 -190
rect 2827 190 2897 622
rect 2827 -622 2897 -190
rect 3145 190 3215 622
rect 3145 -622 3215 -190
rect 3463 190 3533 622
rect 3463 -622 3533 -190
rect 3781 190 3851 622
rect 3781 -622 3851 -190
<< xpolyres >>
rect -3851 -190 -3781 190
rect -3533 -190 -3463 190
rect -3215 -190 -3145 190
rect -2897 -190 -2827 190
rect -2579 -190 -2509 190
rect -2261 -190 -2191 190
rect -1943 -190 -1873 190
rect -1625 -190 -1555 190
rect -1307 -190 -1237 190
rect -989 -190 -919 190
rect -671 -190 -601 190
rect -353 -190 -283 190
rect -35 -190 35 190
rect 283 -190 353 190
rect 601 -190 671 190
rect 919 -190 989 190
rect 1237 -190 1307 190
rect 1555 -190 1625 190
rect 1873 -190 1943 190
rect 2191 -190 2261 190
rect 2509 -190 2579 190
rect 2827 -190 2897 190
rect 3145 -190 3215 190
rect 3463 -190 3533 190
rect 3781 -190 3851 190
<< viali >>
rect -3835 207 -3797 604
rect -3517 207 -3479 604
rect -3199 207 -3161 604
rect -2881 207 -2843 604
rect -2563 207 -2525 604
rect -2245 207 -2207 604
rect -1927 207 -1889 604
rect -1609 207 -1571 604
rect -1291 207 -1253 604
rect -973 207 -935 604
rect -655 207 -617 604
rect -337 207 -299 604
rect -19 207 19 604
rect 299 207 337 604
rect 617 207 655 604
rect 935 207 973 604
rect 1253 207 1291 604
rect 1571 207 1609 604
rect 1889 207 1927 604
rect 2207 207 2245 604
rect 2525 207 2563 604
rect 2843 207 2881 604
rect 3161 207 3199 604
rect 3479 207 3517 604
rect 3797 207 3835 604
rect -3835 -604 -3797 -207
rect -3517 -604 -3479 -207
rect -3199 -604 -3161 -207
rect -2881 -604 -2843 -207
rect -2563 -604 -2525 -207
rect -2245 -604 -2207 -207
rect -1927 -604 -1889 -207
rect -1609 -604 -1571 -207
rect -1291 -604 -1253 -207
rect -973 -604 -935 -207
rect -655 -604 -617 -207
rect -337 -604 -299 -207
rect -19 -604 19 -207
rect 299 -604 337 -207
rect 617 -604 655 -207
rect 935 -604 973 -207
rect 1253 -604 1291 -207
rect 1571 -604 1609 -207
rect 1889 -604 1927 -207
rect 2207 -604 2245 -207
rect 2525 -604 2563 -207
rect 2843 -604 2881 -207
rect 3161 -604 3199 -207
rect 3479 -604 3517 -207
rect 3797 -604 3835 -207
<< metal1 >>
rect -3841 604 -3791 616
rect -3841 207 -3835 604
rect -3797 207 -3791 604
rect -3841 195 -3791 207
rect -3523 604 -3473 616
rect -3523 207 -3517 604
rect -3479 207 -3473 604
rect -3523 195 -3473 207
rect -3205 604 -3155 616
rect -3205 207 -3199 604
rect -3161 207 -3155 604
rect -3205 195 -3155 207
rect -2887 604 -2837 616
rect -2887 207 -2881 604
rect -2843 207 -2837 604
rect -2887 195 -2837 207
rect -2569 604 -2519 616
rect -2569 207 -2563 604
rect -2525 207 -2519 604
rect -2569 195 -2519 207
rect -2251 604 -2201 616
rect -2251 207 -2245 604
rect -2207 207 -2201 604
rect -2251 195 -2201 207
rect -1933 604 -1883 616
rect -1933 207 -1927 604
rect -1889 207 -1883 604
rect -1933 195 -1883 207
rect -1615 604 -1565 616
rect -1615 207 -1609 604
rect -1571 207 -1565 604
rect -1615 195 -1565 207
rect -1297 604 -1247 616
rect -1297 207 -1291 604
rect -1253 207 -1247 604
rect -1297 195 -1247 207
rect -979 604 -929 616
rect -979 207 -973 604
rect -935 207 -929 604
rect -979 195 -929 207
rect -661 604 -611 616
rect -661 207 -655 604
rect -617 207 -611 604
rect -661 195 -611 207
rect -343 604 -293 616
rect -343 207 -337 604
rect -299 207 -293 604
rect -343 195 -293 207
rect -25 604 25 616
rect -25 207 -19 604
rect 19 207 25 604
rect -25 195 25 207
rect 293 604 343 616
rect 293 207 299 604
rect 337 207 343 604
rect 293 195 343 207
rect 611 604 661 616
rect 611 207 617 604
rect 655 207 661 604
rect 611 195 661 207
rect 929 604 979 616
rect 929 207 935 604
rect 973 207 979 604
rect 929 195 979 207
rect 1247 604 1297 616
rect 1247 207 1253 604
rect 1291 207 1297 604
rect 1247 195 1297 207
rect 1565 604 1615 616
rect 1565 207 1571 604
rect 1609 207 1615 604
rect 1565 195 1615 207
rect 1883 604 1933 616
rect 1883 207 1889 604
rect 1927 207 1933 604
rect 1883 195 1933 207
rect 2201 604 2251 616
rect 2201 207 2207 604
rect 2245 207 2251 604
rect 2201 195 2251 207
rect 2519 604 2569 616
rect 2519 207 2525 604
rect 2563 207 2569 604
rect 2519 195 2569 207
rect 2837 604 2887 616
rect 2837 207 2843 604
rect 2881 207 2887 604
rect 2837 195 2887 207
rect 3155 604 3205 616
rect 3155 207 3161 604
rect 3199 207 3205 604
rect 3155 195 3205 207
rect 3473 604 3523 616
rect 3473 207 3479 604
rect 3517 207 3523 604
rect 3473 195 3523 207
rect 3791 604 3841 616
rect 3791 207 3797 604
rect 3835 207 3841 604
rect 3791 195 3841 207
rect -3841 -207 -3791 -195
rect -3841 -604 -3835 -207
rect -3797 -604 -3791 -207
rect -3841 -616 -3791 -604
rect -3523 -207 -3473 -195
rect -3523 -604 -3517 -207
rect -3479 -604 -3473 -207
rect -3523 -616 -3473 -604
rect -3205 -207 -3155 -195
rect -3205 -604 -3199 -207
rect -3161 -604 -3155 -207
rect -3205 -616 -3155 -604
rect -2887 -207 -2837 -195
rect -2887 -604 -2881 -207
rect -2843 -604 -2837 -207
rect -2887 -616 -2837 -604
rect -2569 -207 -2519 -195
rect -2569 -604 -2563 -207
rect -2525 -604 -2519 -207
rect -2569 -616 -2519 -604
rect -2251 -207 -2201 -195
rect -2251 -604 -2245 -207
rect -2207 -604 -2201 -207
rect -2251 -616 -2201 -604
rect -1933 -207 -1883 -195
rect -1933 -604 -1927 -207
rect -1889 -604 -1883 -207
rect -1933 -616 -1883 -604
rect -1615 -207 -1565 -195
rect -1615 -604 -1609 -207
rect -1571 -604 -1565 -207
rect -1615 -616 -1565 -604
rect -1297 -207 -1247 -195
rect -1297 -604 -1291 -207
rect -1253 -604 -1247 -207
rect -1297 -616 -1247 -604
rect -979 -207 -929 -195
rect -979 -604 -973 -207
rect -935 -604 -929 -207
rect -979 -616 -929 -604
rect -661 -207 -611 -195
rect -661 -604 -655 -207
rect -617 -604 -611 -207
rect -661 -616 -611 -604
rect -343 -207 -293 -195
rect -343 -604 -337 -207
rect -299 -604 -293 -207
rect -343 -616 -293 -604
rect -25 -207 25 -195
rect -25 -604 -19 -207
rect 19 -604 25 -207
rect -25 -616 25 -604
rect 293 -207 343 -195
rect 293 -604 299 -207
rect 337 -604 343 -207
rect 293 -616 343 -604
rect 611 -207 661 -195
rect 611 -604 617 -207
rect 655 -604 661 -207
rect 611 -616 661 -604
rect 929 -207 979 -195
rect 929 -604 935 -207
rect 973 -604 979 -207
rect 929 -616 979 -604
rect 1247 -207 1297 -195
rect 1247 -604 1253 -207
rect 1291 -604 1297 -207
rect 1247 -616 1297 -604
rect 1565 -207 1615 -195
rect 1565 -604 1571 -207
rect 1609 -604 1615 -207
rect 1565 -616 1615 -604
rect 1883 -207 1933 -195
rect 1883 -604 1889 -207
rect 1927 -604 1933 -207
rect 1883 -616 1933 -604
rect 2201 -207 2251 -195
rect 2201 -604 2207 -207
rect 2245 -604 2251 -207
rect 2201 -616 2251 -604
rect 2519 -207 2569 -195
rect 2519 -604 2525 -207
rect 2563 -604 2569 -207
rect 2519 -616 2569 -604
rect 2837 -207 2887 -195
rect 2837 -604 2843 -207
rect 2881 -604 2887 -207
rect 2837 -616 2887 -604
rect 3155 -207 3205 -195
rect 3155 -604 3161 -207
rect 3199 -604 3205 -207
rect 3155 -616 3205 -604
rect 3473 -207 3523 -195
rect 3473 -604 3479 -207
rect 3517 -604 3523 -207
rect 3473 -616 3523 -604
rect 3791 -207 3841 -195
rect 3791 -604 3797 -207
rect 3835 -604 3841 -207
rect 3791 -616 3841 -604
<< res0p35 >>
rect -3853 -192 -3779 192
rect -3535 -192 -3461 192
rect -3217 -192 -3143 192
rect -2899 -192 -2825 192
rect -2581 -192 -2507 192
rect -2263 -192 -2189 192
rect -1945 -192 -1871 192
rect -1627 -192 -1553 192
rect -1309 -192 -1235 192
rect -991 -192 -917 192
rect -673 -192 -599 192
rect -355 -192 -281 192
rect -37 -192 37 192
rect 281 -192 355 192
rect 599 -192 673 192
rect 917 -192 991 192
rect 1235 -192 1309 192
rect 1553 -192 1627 192
rect 1871 -192 1945 192
rect 2189 -192 2263 192
rect 2507 -192 2581 192
rect 2825 -192 2899 192
rect 3143 -192 3217 192
rect 3461 -192 3535 192
rect 3779 -192 3853 192
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 1.9 m 1 nx 25 wmin 0.350 lmin 0.50 rho 2000 val 11.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
