magic
tech sky130A
magscale 1 2
timestamp 1669742938
<< error_p >>
rect -819000 -60480 -806400 -60094
rect -819000 -80640 -786240 -60480
rect -729800 -64600 -729000 -64200
rect -730600 -65200 -729800 -64600
rect -729000 -65200 -707600 -64600
rect -734387 -67762 -730600 -65200
rect -771400 -80640 -734387 -67762
rect -819000 -92800 -779630 -80640
rect -771400 -92800 -745920 -80640
rect -707600 -92800 -707400 -65200
rect -819000 -98400 -771400 -92800
rect -709400 -93072 -707400 -92800
rect -709460 -93132 -707400 -93072
rect -710387 -93800 -707400 -93132
rect -822562 -100800 -806400 -98400
rect -788600 -99400 -771400 -98400
rect -788600 -100800 -766080 -99400
rect -822562 -104267 -745920 -100800
rect -725853 -104267 -710387 -93800
rect -822562 -104932 -786240 -104267
rect -851600 -120960 -786240 -104932
rect -778567 -104932 -745920 -104267
rect -726836 -104932 -725853 -104267
rect -778567 -120960 -726836 -104932
rect -851600 -135091 -782287 -120960
rect -778567 -135091 -736813 -120960
rect -851600 -137577 -736813 -135091
rect -851600 -141120 -806400 -137577
rect -788595 -140201 -736813 -137577
rect -851600 -147200 -826560 -141120
rect -788595 -142200 -771400 -140201
rect -736813 -141200 -735791 -140201
rect -788595 -146728 -745920 -142200
rect -788664 -146734 -788628 -146728
rect -788604 -146734 -788544 -146728
rect -789301 -147200 -788636 -146734
rect -853094 -148362 -851600 -147200
rect -790825 -148239 -789301 -147200
rect -790886 -148267 -789301 -148239
rect -854703 -149613 -853094 -148362
rect -792876 -149613 -790886 -148267
rect -826313 -161280 -792876 -149613
rect -777547 -161280 -745920 -146728
rect -826313 -172238 -806400 -161280
rect -831044 -175439 -826313 -172238
rect -831044 -175460 -831030 -175439
rect -831483 -175800 -831030 -175460
rect -832000 -176059 -831483 -175800
rect -777547 -179400 -739153 -161280
rect -739153 -179548 -739000 -179400
<< metal4 >>
tri -729800 -64600 -729200 -64200 se
tri -729200 -64600 -729000 -64200 sw
tri -730600 -65200 -729800 -64600 se
rect -729800 -65200 -729000 -64600
tri -729000 -65200 -707600 -64600 sw
tri -734387 -67762 -730600 -65200 se
rect -730600 -67762 -707600 -65200
tri -771400 -92800 -734387 -67762 se
rect -734387 -92438 -733038 -67762
rect -708162 -92438 -707600 -67762
rect -734387 -92800 -707600 -92438
tri -707600 -92800 -707400 -65200 sw
tri -788600 -104267 -771400 -92800 se
rect -771400 -93132 -709400 -92800
rect -771400 -93800 -710387 -93132
tri -710387 -93800 -709400 -93132 nw
tri -709400 -93800 -707400 -92800 nw
rect -771400 -104267 -725853 -93800
tri -725853 -104267 -710387 -93800 nw
tri -788883 -104456 -788600 -104267 se
rect -788600 -104456 -726836 -104267
tri -788902 -104468 -788883 -104456 se
rect -788883 -104468 -726836 -104456
tri -789301 -104932 -788618 -104468 se
rect -788618 -104932 -726836 -104468
tri -726836 -104932 -725853 -104267 nw
tri -851600 -147200 -789301 -104932 se
rect -789301 -135091 -771400 -104932
tri -771400 -135091 -726836 -104932 nw
rect -789301 -146728 -788595 -135091
tri -788595 -146728 -771400 -135091 nw
rect -789301 -146734 -788636 -146728
tri -788636 -146734 -788628 -146728 nw
tri -788604 -146734 -788595 -146728 nw
tri -789301 -147200 -788636 -146734 nw
tri -853094 -148362 -851600 -147200 se
rect -851600 -148239 -790825 -147200
rect -851600 -148267 -790886 -148239
tri -790886 -148267 -790844 -148239 nw
tri -790844 -148267 -790825 -148239 ne
tri -790825 -148267 -789301 -147200 nw
rect -851600 -148362 -792876 -148267
tri -854703 -149613 -853094 -148362 se
rect -853094 -149613 -853038 -148362
rect -854703 -172238 -853038 -149613
rect -828362 -149613 -792876 -148362
tri -792876 -149613 -790886 -148267 nw
rect -828362 -172238 -826313 -149613
tri -826313 -172238 -792876 -149613 nw
rect -854703 -175460 -831044 -172238
tri -831044 -175439 -826313 -172238 nw
tri -831044 -175460 -831030 -175439 sw
rect -854703 -175800 -831483 -175460
tri -831483 -175800 -831030 -175460 nw
tri -832000 -176059 -831828 -175800 ne
tri -831828 -176059 -831483 -175800 nw
<< via4 >>
rect -733038 -92438 -708162 -67762
rect -853038 -172238 -828362 -148362
<< metal5 >>
rect -1058800 -60000 -1022000 -59934
rect -1058800 -98400 -819000 -60000
tri -819000 -98400 -779630 -60094 sw
rect -540800 -61000 -498737 -60951
rect -743200 -67762 -498737 -61000
rect -743200 -92438 -733038 -67762
rect -708162 -92438 -498737 -67762
tri -779610 -98400 -779591 -98381 sw
rect -1058800 -581200 -1020400 -98400
tri -822562 -137577 -782287 -98400 ne
rect -782287 -99400 -779591 -98400
tri -779591 -99400 -778567 -98400 sw
rect -743200 -99400 -498737 -92438
tri -782317 -137607 -782287 -137577 ne
rect -782287 -137607 -778567 -99400
tri -782287 -137637 -782256 -137607 ne
rect -782256 -137637 -778567 -137607
tri -782256 -137666 -782226 -137637 ne
rect -782226 -137666 -778567 -137637
tri -782226 -137695 -782196 -137666 ne
rect -782196 -137695 -778567 -137666
tri -782196 -137725 -782166 -137695 ne
rect -782166 -137725 -778567 -137695
tri -782166 -137741 -782149 -137725 ne
rect -782149 -137741 -778567 -137725
tri -782149 -137770 -782119 -137741 ne
rect -782119 -137770 -778567 -137741
tri -782119 -137799 -782089 -137770 ne
rect -782089 -137799 -778567 -137770
tri -782089 -137828 -782059 -137799 ne
rect -782059 -137828 -778567 -137799
tri -782059 -137856 -782030 -137828 ne
rect -782030 -137856 -778567 -137828
tri -782030 -140201 -779610 -137856 ne
rect -779610 -140201 -778567 -137856
tri -778567 -140201 -736813 -99400 sw
tri -779610 -141200 -778579 -140201 ne
rect -778579 -141200 -736813 -140201
tri -736813 -141200 -735791 -140201 sw
tri -778579 -142200 -777547 -141200 ne
rect -777547 -142200 -580939 -141200
rect -940000 -142250 -819800 -142200
rect -978400 -148362 -819800 -142250
rect -978400 -172238 -853038 -148362
rect -828362 -172238 -819800 -148362
rect -978400 -179400 -819800 -172238
tri -777547 -179400 -739153 -142200 ne
rect -739153 -179400 -580939 -142200
rect -978400 -500800 -940000 -179400
tri -739153 -179548 -739000 -179400 ne
rect -739000 -179600 -580939 -179400
rect -619000 -500800 -580939 -179600
rect -978800 -539600 -581036 -500800
rect -540800 -580200 -498737 -99400
rect -739000 -581200 -498737 -580200
rect -1058800 -623000 -819000 -581200
rect -739000 -621800 -498549 -581200
rect -1058800 -623200 -818800 -623000
rect -850600 -649800 -818800 -623200
rect -738800 -650400 -710000 -621800
<< end >>
