magic
tech sky130A
magscale 1 2
timestamp 1668228285
<< error_p >>
rect -70 50 -10 950
rect 10 50 70 950
rect 818 810 841 811
rect 878 810 921 891
rect 925 850 956 866
rect 940 151 956 850
rect 925 150 956 151
rect 995 78 1005 922
rect -70 -950 -10 -50
rect 10 -950 70 -50
rect 925 -150 956 -134
rect 818 -811 841 -810
rect 878 -891 921 -810
rect 940 -849 956 -150
rect 925 -850 956 -849
rect 995 -922 1005 -78
<< metal3 >>
rect -1009 922 -10 950
rect -1009 78 -94 922
rect -30 78 -10 922
rect -1009 50 -10 78
rect 10 922 1138 950
rect 10 78 925 922
rect 989 78 995 922
rect 1118 78 1138 922
rect 10 50 1138 78
rect -1009 -78 -10 -50
rect -1009 -922 -94 -78
rect -30 -922 -10 -78
rect -1009 -950 -10 -922
rect 10 -78 1138 -50
rect 10 -922 925 -78
rect 989 -922 995 -78
rect 1118 -922 1138 -78
rect 10 -950 1138 -922
<< via3 >>
rect -94 78 -30 922
rect 925 78 989 922
rect 995 78 1118 922
rect -94 -922 -30 -78
rect 925 -922 989 -78
rect 995 -922 1118 -78
<< mimcap >>
rect -909 810 -208 850
rect -909 190 -869 810
rect -248 190 -208 810
rect -909 150 -208 190
rect 110 810 940 850
rect 110 190 150 810
rect 900 190 940 810
rect 110 150 940 190
rect -909 -190 -208 -150
rect -909 -810 -869 -190
rect -248 -810 -208 -190
rect -909 -850 -208 -810
rect 110 -190 940 -150
rect 110 -810 150 -190
rect 900 -810 940 -190
rect 110 -850 940 -810
<< mimcapcontact >>
rect -869 190 -248 810
rect 150 190 900 810
rect -869 -810 -248 -190
rect 150 -810 900 -190
<< metal4 >>
rect -611 811 -506 1000
rect -141 938 -36 1000
rect -141 922 -14 938
rect -870 810 -248 811
rect -870 190 -869 810
rect -870 188 -248 190
rect -611 -188 -506 188
rect -141 78 -94 922
rect -30 78 -14 922
rect 408 811 642 1000
rect 878 938 1112 1000
rect 878 922 1134 938
rect 149 810 841 811
rect 878 810 925 922
rect 149 190 150 810
rect 900 190 925 810
rect 149 189 925 190
rect 278 188 925 189
rect -141 62 -14 78
rect -141 -62 -36 62
rect -141 -78 -14 -62
rect -870 -190 -248 -188
rect -870 -810 -869 -190
rect -870 -811 -248 -810
rect -611 -1000 -506 -811
rect -141 -922 -94 -78
rect -30 -922 -14 -78
rect 408 -188 642 188
rect 878 78 925 188
rect 989 78 995 922
rect 1118 78 1134 922
rect 878 62 1134 78
rect 878 -62 1112 62
rect 878 -78 1134 -62
rect 878 -188 925 -78
rect 278 -189 925 -188
rect 149 -190 925 -189
rect 149 -810 150 -190
rect 900 -810 925 -190
rect 149 -811 841 -810
rect -141 -938 -14 -922
rect -141 -1000 -36 -938
rect 408 -1000 642 -811
rect 878 -922 925 -810
rect 989 -922 995 -78
rect 1118 -922 1134 -78
rect 878 -938 1134 -922
rect 878 -1000 1112 -938
<< properties >>
string FIXED_BBOX 10 50 910 950
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.5 l 3.5 val 27.16 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
