magic
tech sky130A
magscale 1 2
timestamp 1668022138
<< nwell >>
rect -184 -580 184 580
<< pmos >>
rect -90 -480 90 480
<< pdiff >>
rect -148 468 -90 480
rect -148 -468 -136 468
rect -102 -468 -90 468
rect -148 -480 -90 -468
rect 90 468 148 480
rect 90 -468 102 468
rect 136 -468 148 468
rect 90 -480 148 -468
<< pdiffc >>
rect -136 -468 -102 468
rect 102 -468 136 468
<< poly >>
rect -90 561 90 577
rect -90 527 -74 561
rect 74 527 90 561
rect -90 480 90 527
rect -90 -527 90 -480
rect -90 -561 -74 -527
rect 74 -561 90 -527
rect -90 -577 90 -561
<< polycont >>
rect -74 527 74 561
rect -74 -561 74 -527
<< locali >>
rect -90 527 -74 561
rect 74 527 90 561
rect -136 468 -102 484
rect -136 -484 -102 -468
rect 102 468 136 484
rect 102 -484 136 -468
rect -90 -561 -74 -527
rect 74 -561 90 -527
<< viali >>
rect -74 527 74 561
rect -136 -468 -102 468
rect 102 -468 136 468
rect -74 -561 74 -527
<< metal1 >>
rect -86 561 86 567
rect -86 527 -74 561
rect 74 527 86 561
rect -86 521 86 527
rect -142 468 -96 480
rect -142 -468 -136 468
rect -102 -468 -96 468
rect -142 -480 -96 -468
rect 96 468 142 480
rect 96 -468 102 468
rect 136 -468 142 468
rect 96 -480 142 -468
rect -86 -527 86 -521
rect -86 -561 -74 -527
rect 74 -561 86 -527
rect -86 -567 86 -561
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.9 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
