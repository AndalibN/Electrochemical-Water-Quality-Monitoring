magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_s >>
rect 5231 4326 5683 4438
rect 5308 4163 5486 4184
rect 5562 4126 5740 4163
<< pwell >>
rect 6385 4190 6955 4319
<< psubdiff >>
rect 6411 4271 6929 4293
rect 6411 4237 6449 4271
rect 6483 4237 6517 4271
rect 6551 4237 6585 4271
rect 6619 4237 6653 4271
rect 6687 4237 6721 4271
rect 6755 4237 6789 4271
rect 6823 4237 6857 4271
rect 6891 4237 6929 4271
rect 6411 4216 6929 4237
<< psubdiffcont >>
rect 6449 4237 6483 4271
rect 6517 4237 6551 4271
rect 6585 4237 6619 4271
rect 6653 4237 6687 4271
rect 6721 4237 6755 4271
rect 6789 4237 6823 4271
rect 6857 4237 6891 4271
<< poly >>
rect 6672 4542 6713 4608
rect 6445 4094 6504 4095
<< locali >>
rect 6662 4552 6712 4598
rect 5435 4454 5481 4503
rect 6418 4271 6923 4288
rect 6418 4237 6449 4271
rect 6483 4237 6517 4271
rect 6551 4237 6585 4271
rect 6619 4237 6653 4271
rect 6687 4237 6721 4271
rect 6755 4237 6789 4271
rect 6823 4237 6857 4271
rect 6891 4237 6923 4271
rect 6418 4221 6923 4237
<< metal1 >>
rect 5103 4462 5381 4497
rect 5289 4402 5386 4410
rect 5428 4404 5486 4552
rect 5532 4462 5609 4741
rect 6611 4549 6763 4601
rect 6534 4476 6622 4491
rect 6534 4424 6554 4476
rect 6606 4424 6622 4476
rect 5519 4412 5624 4417
rect 5289 4350 5312 4402
rect 5364 4350 5386 4402
rect 5519 4360 5546 4412
rect 5598 4360 5624 4412
rect 6534 4408 6622 4424
rect 5519 4352 5624 4360
rect 5289 4342 5386 4350
rect 5297 4177 5376 4184
rect 5297 4125 5318 4177
rect 5370 4125 5376 4177
rect 5297 4117 5376 4125
rect 5316 3614 5350 4052
rect 5404 3692 5438 4272
rect 6670 4236 6704 4489
rect 6753 4476 6826 4498
rect 6753 4424 6762 4476
rect 6814 4424 6826 4476
rect 6753 4407 6826 4424
rect 5640 4155 5708 4163
rect 5640 4103 5648 4155
rect 5700 4103 5708 4155
rect 5640 4097 5708 4103
rect 6438 4147 6510 4159
rect 6438 4095 6448 4147
rect 6500 4095 6510 4147
rect 6438 4091 6510 4095
rect 5492 3802 5644 4052
rect 6503 4051 6538 4052
rect 6627 4039 6693 4051
rect 5492 3750 5502 3802
rect 5554 3750 5644 3802
rect 5492 3692 5644 3750
rect 5422 3620 5509 3635
rect 5422 3614 5438 3620
rect 5316 3578 5438 3614
rect 5422 3568 5438 3578
rect 5490 3568 5509 3620
rect 5422 3558 5509 3568
rect 5610 3356 5644 3692
rect 5697 4004 5774 4034
rect 5697 3952 5708 4004
rect 5760 3952 5774 4004
rect 5697 3940 5774 3952
rect 5697 3888 5708 3940
rect 5760 3888 5774 3940
rect 5697 3876 5774 3888
rect 5697 3824 5708 3876
rect 5760 3824 5774 3876
rect 5697 3812 5774 3824
rect 5697 3760 5708 3812
rect 5760 3760 5774 3812
rect 5697 3748 5774 3760
rect 5697 3696 5708 3748
rect 5760 3696 5774 3748
rect 5697 3684 5774 3696
rect 5697 3632 5708 3684
rect 5760 3632 5774 3684
rect 5697 3620 5774 3632
rect 5697 3568 5708 3620
rect 5760 3568 5774 3620
rect 5697 3556 5774 3568
rect 5697 3504 5708 3556
rect 5760 3504 5774 3556
rect 5697 3492 5774 3504
rect 5697 3440 5708 3492
rect 5760 3440 5774 3492
rect 5697 3428 5774 3440
rect 5697 3376 5708 3428
rect 5760 3376 5774 3428
rect 5697 3350 5774 3376
rect 6374 4004 6451 4034
rect 6374 3952 6387 4004
rect 6439 3952 6451 4004
rect 6627 3987 6633 4039
rect 6685 3987 6693 4039
rect 6627 3975 6693 3987
rect 6741 3975 6775 4273
rect 6805 4148 6877 4153
rect 6805 4096 6815 4148
rect 6867 4096 6877 4148
rect 6805 4091 6877 4096
rect 6374 3940 6451 3952
rect 6374 3888 6387 3940
rect 6439 3888 6451 3940
rect 6374 3876 6451 3888
rect 6374 3824 6387 3876
rect 6439 3824 6451 3876
rect 6503 3830 6538 3975
rect 6671 3916 6759 3929
rect 6826 3916 6867 4051
rect 6671 3913 6867 3916
rect 6671 3861 6687 3913
rect 6739 3861 6867 3913
rect 6671 3847 6759 3861
rect 6826 3860 6867 3861
rect 6374 3812 6451 3824
rect 6374 3760 6387 3812
rect 6439 3760 6451 3812
rect 6374 3748 6451 3760
rect 6374 3696 6387 3748
rect 6439 3696 6451 3748
rect 6502 3803 6603 3830
rect 6502 3751 6529 3803
rect 6581 3751 6603 3803
rect 6502 3726 6603 3751
rect 6374 3684 6451 3696
rect 6374 3632 6387 3684
rect 6439 3632 6451 3684
rect 6374 3620 6451 3632
rect 6374 3568 6387 3620
rect 6439 3568 6451 3620
rect 6374 3556 6451 3568
rect 6374 3504 6387 3556
rect 6439 3504 6451 3556
rect 6374 3492 6451 3504
rect 6374 3440 6387 3492
rect 6439 3440 6451 3492
rect 6374 3428 6451 3440
rect 6374 3376 6387 3428
rect 6439 3376 6451 3428
rect 6374 3351 6451 3376
rect 6503 3355 6538 3726
rect 6401 3350 6451 3351
<< via1 >>
rect 6554 4424 6606 4476
rect 5312 4350 5364 4402
rect 5546 4360 5598 4412
rect 5318 4125 5370 4177
rect 6762 4424 6814 4476
rect 5648 4103 5700 4155
rect 6448 4095 6500 4147
rect 5502 3750 5554 3802
rect 5438 3568 5490 3620
rect 5708 3952 5760 4004
rect 5708 3888 5760 3940
rect 5708 3824 5760 3876
rect 5708 3760 5760 3812
rect 5708 3696 5760 3748
rect 5708 3632 5760 3684
rect 5708 3568 5760 3620
rect 5708 3504 5760 3556
rect 5708 3440 5760 3492
rect 5708 3376 5760 3428
rect 6387 3952 6439 4004
rect 6633 3987 6685 4039
rect 6815 4096 6867 4148
rect 6387 3888 6439 3940
rect 6387 3824 6439 3876
rect 6687 3861 6739 3913
rect 6387 3760 6439 3812
rect 6387 3696 6439 3748
rect 6529 3751 6581 3803
rect 6387 3632 6439 3684
rect 6387 3568 6439 3620
rect 6387 3504 6439 3556
rect 6387 3440 6439 3492
rect 6387 3376 6439 3428
<< metal2 >>
rect 6438 4476 6622 4491
rect 6438 4424 6554 4476
rect 6606 4424 6622 4476
rect 5515 4412 5719 4418
rect 5285 4402 5391 4412
rect 5285 4350 5312 4402
rect 5364 4350 5391 4402
rect 5285 4177 5391 4350
rect 5515 4360 5546 4412
rect 5598 4360 5719 4412
rect 5515 4348 5719 4360
rect 6438 4408 6622 4424
rect 6751 4476 6881 4498
rect 6751 4424 6762 4476
rect 6814 4424 6881 4476
rect 5285 4125 5318 4177
rect 5370 4125 5391 4177
rect 5285 4116 5391 4125
rect 5641 4155 5718 4348
rect 5641 4103 5648 4155
rect 5700 4103 5718 4155
rect 5641 4096 5718 4103
rect 6438 4147 6509 4408
rect 6751 4406 6881 4424
rect 6438 4095 6448 4147
rect 6500 4095 6509 4147
rect 6438 4089 6509 4095
rect 6803 4148 6881 4406
rect 6803 4096 6815 4148
rect 6867 4096 6881 4148
rect 6803 4089 6881 4096
rect 6368 4039 6693 4051
rect 6368 4033 6633 4039
rect 5697 4004 6633 4033
rect 5697 3952 5708 4004
rect 5760 3952 6387 4004
rect 6439 3987 6633 4004
rect 6685 3987 6693 4039
rect 6439 3975 6693 3987
rect 6439 3952 6451 3975
rect 5697 3940 6451 3952
rect 5697 3888 5708 3940
rect 5760 3888 6387 3940
rect 6439 3888 6451 3940
rect 5697 3876 6451 3888
rect 5491 3804 5565 3828
rect 5491 3748 5500 3804
rect 5556 3748 5565 3804
rect 5491 3726 5565 3748
rect 5697 3824 5708 3876
rect 5760 3824 6387 3876
rect 6439 3824 6451 3876
rect 6667 3915 6759 3930
rect 6667 3859 6685 3915
rect 6741 3859 6759 3915
rect 6667 3844 6759 3859
rect 5697 3812 6451 3824
rect 5697 3760 5708 3812
rect 5760 3760 6387 3812
rect 6439 3760 6451 3812
rect 5697 3748 6451 3760
rect 5697 3696 5708 3748
rect 5760 3696 6387 3748
rect 6439 3696 6451 3748
rect 6507 3805 6604 3831
rect 6507 3749 6527 3805
rect 6583 3749 6604 3805
rect 6507 3726 6604 3749
rect 5697 3684 6451 3696
rect 5416 3622 5511 3640
rect 5416 3566 5435 3622
rect 5491 3566 5511 3622
rect 5416 3550 5511 3566
rect 5697 3632 5708 3684
rect 5760 3632 6387 3684
rect 6439 3632 6451 3684
rect 5697 3620 6451 3632
rect 5697 3568 5708 3620
rect 5760 3568 6387 3620
rect 6439 3568 6451 3620
rect 5697 3556 6451 3568
rect 5697 3504 5708 3556
rect 5760 3504 6387 3556
rect 6439 3504 6451 3556
rect 5697 3492 6451 3504
rect 5697 3440 5708 3492
rect 5760 3440 6387 3492
rect 6439 3440 6451 3492
rect 5697 3428 6451 3440
rect 5697 3376 5708 3428
rect 5760 3376 6387 3428
rect 6439 3376 6451 3428
rect 5697 3350 6451 3376
<< via2 >>
rect 5500 3802 5556 3804
rect 5500 3750 5502 3802
rect 5502 3750 5554 3802
rect 5554 3750 5556 3802
rect 5500 3748 5556 3750
rect 6685 3913 6741 3915
rect 6685 3861 6687 3913
rect 6687 3861 6739 3913
rect 6739 3861 6741 3913
rect 6685 3859 6741 3861
rect 6527 3803 6583 3805
rect 6527 3751 6529 3803
rect 6529 3751 6581 3803
rect 6581 3751 6583 3803
rect 6527 3749 6583 3751
rect 5435 3620 5491 3622
rect 5435 3568 5438 3620
rect 5438 3568 5490 3620
rect 5490 3568 5491 3620
rect 5435 3566 5491 3568
<< metal3 >>
rect 6671 3915 6759 3929
rect 6671 3859 6685 3915
rect 6741 3859 6759 3915
rect 6671 3847 6759 3859
rect 5491 3805 6604 3829
rect 5491 3804 6527 3805
rect 5491 3748 5500 3804
rect 5556 3749 6527 3804
rect 6583 3749 6604 3805
rect 5556 3748 6604 3749
rect 5491 3726 6604 3748
rect 5417 3635 5512 3637
rect 6674 3635 6754 3847
rect 5417 3622 6754 3635
rect 5417 3566 5435 3622
rect 5491 3566 6754 3622
rect 5417 3559 6754 3566
rect 5417 3557 6753 3559
rect 5417 3553 5512 3557
use sky130_fd_pr__nfet_01v8_JBX99N  XM2
timestamp 1669522153
transform 1 0 6802 0 1 4044
box -99 -107 99 107
use sky130_fd_pr__pfet_01v8_L42X7S  XM3
timestamp 1669522153
transform 1 0 5465 0 1 3836
box -109 -274 109 290
use sky130_fd_pr__nfet_01v8_JB6ZCM  XM4
timestamp 1669522153
transform 1 0 6714 0 1 3982
box -99 -127 99 107
use sky130_fd_pr__pfet_01v8_SCSK2Z  XM5
timestamp 1669522153
transform 1 0 5674 0 1 3739
box -112 -458 112 424
use sky130_fd_pr__nfet_01v8_C9ME4G  XM6
timestamp 1669522153
transform 1 0 6474 0 1 3734
box -102 -417 102 417
use sky130_fd_pr__pfet_01v8_LJPFBL  XM8
timestamp 1669522153
transform 0 -1 5379 1 0 4523
box -109 -114 109 148
use sky130_fd_pr__pfet_01v8_MJPFBN  XM9
timestamp 1669522153
transform 0 1 5379 1 0 4435
box -109 -148 109 114
use sky130_fd_pr__nfet_01v8_JB6ZCM  XM10
timestamp 1669522153
transform -1 0 6731 0 -1 4481
box -99 -127 99 107
use sky130_fd_pr__nfet_01v8_JB6ZCM  sky130_fd_pr__nfet_01v8_JB6ZCM_0
timestamp 1669522153
transform -1 0 6643 0 -1 4481
box -99 -127 99 107
use sky130_fd_pr__pfet_01v8_M42X7L  sky130_fd_pr__pfet_01v8_M42X7L_0
timestamp 1669522153
transform 1 0 5377 0 1 3908
box -109 -290 109 276
use sky130_fd_pr__pfet_01v8_MJPFFN  sky130_fd_pr__pfet_01v8_MJPFFN_0
timestamp 1669522153
transform 0 -1 5535 1 0 4435
box -109 -148 109 114
<< end >>
