magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< error_p >>
rect -29 5081 29 5087
rect -29 5047 -17 5081
rect -29 5041 29 5047
rect -29 -5047 29 -5041
rect -29 -5081 -17 -5047
rect -29 -5087 29 -5081
<< nwell >>
rect -114 -5100 114 5100
<< pmos >>
rect -20 -5000 20 5000
<< pdiff >>
rect -78 4988 -20 5000
rect -78 -4988 -66 4988
rect -32 -4988 -20 4988
rect -78 -5000 -20 -4988
rect 20 4988 78 5000
rect 20 -4988 32 4988
rect 66 -4988 78 4988
rect 20 -5000 78 -4988
<< pdiffc >>
rect -66 -4988 -32 4988
rect 32 -4988 66 4988
<< poly >>
rect -33 5081 33 5097
rect -33 5047 -17 5081
rect 17 5047 33 5081
rect -33 5031 33 5047
rect -20 5000 20 5031
rect -20 -5031 20 -5000
rect -33 -5047 33 -5031
rect -33 -5081 -17 -5047
rect 17 -5081 33 -5047
rect -33 -5097 33 -5081
<< polycont >>
rect -17 5047 17 5081
rect -17 -5081 17 -5047
<< locali >>
rect -33 5047 -17 5081
rect 17 5047 33 5081
rect -66 4988 -32 5004
rect -66 -5004 -32 -4988
rect 32 4988 66 5004
rect 32 -5004 66 -4988
rect -33 -5081 -17 -5047
rect 17 -5081 33 -5047
<< viali >>
rect -17 5047 17 5081
rect -66 -4988 -32 4988
rect 32 -4988 66 4988
rect -17 -5081 17 -5047
<< metal1 >>
rect -29 5081 29 5087
rect -29 5047 -17 5081
rect 17 5047 29 5081
rect -29 5041 29 5047
rect -72 4988 -26 5000
rect -72 -4988 -66 4988
rect -32 -4988 -26 4988
rect -72 -5000 -26 -4988
rect 26 4988 72 5000
rect 26 -4988 32 4988
rect 66 -4988 72 4988
rect 26 -5000 72 -4988
rect -29 -5047 29 -5041
rect -29 -5081 -17 -5047
rect 17 -5081 29 -5047
rect -29 -5087 29 -5081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 50.0 l 0.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
