magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nmos >>
rect -287 -2500 -187 2500
rect -129 -2500 -29 2500
rect 29 -2500 129 2500
rect 187 -2500 287 2500
<< ndiff >>
rect -345 2488 -287 2500
rect -345 -2488 -333 2488
rect -299 -2488 -287 2488
rect -345 -2500 -287 -2488
rect -187 2488 -129 2500
rect -187 -2488 -175 2488
rect -141 -2488 -129 2488
rect -187 -2500 -129 -2488
rect -29 2488 29 2500
rect -29 -2488 -17 2488
rect 17 -2488 29 2488
rect -29 -2500 29 -2488
rect 129 2488 187 2500
rect 129 -2488 141 2488
rect 175 -2488 187 2488
rect 129 -2500 187 -2488
rect 287 2488 345 2500
rect 287 -2488 299 2488
rect 333 -2488 345 2488
rect 287 -2500 345 -2488
<< ndiffc >>
rect -333 -2488 -299 2488
rect -175 -2488 -141 2488
rect -17 -2488 17 2488
rect 141 -2488 175 2488
rect 299 -2488 333 2488
<< poly >>
rect -287 2572 -187 2588
rect -287 2538 -271 2572
rect -203 2538 -187 2572
rect -287 2500 -187 2538
rect -129 2572 -29 2588
rect -129 2538 -113 2572
rect -45 2538 -29 2572
rect -129 2500 -29 2538
rect 29 2572 129 2588
rect 29 2538 45 2572
rect 113 2538 129 2572
rect 29 2500 129 2538
rect 187 2572 287 2588
rect 187 2538 203 2572
rect 271 2538 287 2572
rect 187 2500 287 2538
rect -287 -2538 -187 -2500
rect -287 -2572 -271 -2538
rect -203 -2572 -187 -2538
rect -287 -2588 -187 -2572
rect -129 -2538 -29 -2500
rect -129 -2572 -113 -2538
rect -45 -2572 -29 -2538
rect -129 -2588 -29 -2572
rect 29 -2538 129 -2500
rect 29 -2572 45 -2538
rect 113 -2572 129 -2538
rect 29 -2588 129 -2572
rect 187 -2538 287 -2500
rect 187 -2572 203 -2538
rect 271 -2572 287 -2538
rect 187 -2588 287 -2572
<< polycont >>
rect -271 2538 -203 2572
rect -113 2538 -45 2572
rect 45 2538 113 2572
rect 203 2538 271 2572
rect -271 -2572 -203 -2538
rect -113 -2572 -45 -2538
rect 45 -2572 113 -2538
rect 203 -2572 271 -2538
<< locali >>
rect -287 2538 -271 2572
rect -203 2538 -187 2572
rect -129 2538 -113 2572
rect -45 2538 -29 2572
rect 29 2538 45 2572
rect 113 2538 129 2572
rect 187 2538 203 2572
rect 271 2538 287 2572
rect -333 2488 -299 2504
rect -333 -2504 -299 -2488
rect -175 2488 -141 2504
rect -175 -2504 -141 -2488
rect -17 2488 17 2504
rect -17 -2504 17 -2488
rect 141 2488 175 2504
rect 141 -2504 175 -2488
rect 299 2488 333 2504
rect 299 -2504 333 -2488
rect -287 -2572 -271 -2538
rect -203 -2572 -187 -2538
rect -129 -2572 -113 -2538
rect -45 -2572 -29 -2538
rect 29 -2572 45 -2538
rect 113 -2572 129 -2538
rect 187 -2572 203 -2538
rect 271 -2572 287 -2538
<< viali >>
rect -271 2538 -203 2572
rect -113 2538 -45 2572
rect 45 2538 113 2572
rect 203 2538 271 2572
rect -333 -2488 -299 2488
rect -175 -2488 -141 2488
rect -17 -2488 17 2488
rect 141 -2488 175 2488
rect 299 -2488 333 2488
rect -271 -2572 -203 -2538
rect -113 -2572 -45 -2538
rect 45 -2572 113 -2538
rect 203 -2572 271 -2538
<< metal1 >>
rect -283 2572 -191 2578
rect -283 2538 -271 2572
rect -203 2538 -191 2572
rect -283 2532 -191 2538
rect -125 2572 -33 2578
rect -125 2538 -113 2572
rect -45 2538 -33 2572
rect -125 2532 -33 2538
rect 33 2572 125 2578
rect 33 2538 45 2572
rect 113 2538 125 2572
rect 33 2532 125 2538
rect 191 2572 283 2578
rect 191 2538 203 2572
rect 271 2538 283 2572
rect 191 2532 283 2538
rect -339 2488 -293 2500
rect -339 -2488 -333 2488
rect -299 -2488 -293 2488
rect -339 -2500 -293 -2488
rect -181 2488 -135 2500
rect -181 -2488 -175 2488
rect -141 -2488 -135 2488
rect -181 -2500 -135 -2488
rect -23 2488 23 2500
rect -23 -2488 -17 2488
rect 17 -2488 23 2488
rect -23 -2500 23 -2488
rect 135 2488 181 2500
rect 135 -2488 141 2488
rect 175 -2488 181 2488
rect 135 -2500 181 -2488
rect 293 2488 339 2500
rect 293 -2488 299 2488
rect 333 -2488 339 2488
rect 293 -2500 339 -2488
rect -283 -2538 -191 -2532
rect -283 -2572 -271 -2538
rect -203 -2572 -191 -2538
rect -283 -2578 -191 -2572
rect -125 -2538 -33 -2532
rect -125 -2572 -113 -2538
rect -45 -2572 -33 -2538
rect -125 -2578 -33 -2572
rect 33 -2538 125 -2532
rect 33 -2572 45 -2538
rect 113 -2572 125 -2538
rect 33 -2578 125 -2572
rect 191 -2538 283 -2532
rect 191 -2572 203 -2538
rect 271 -2572 283 -2538
rect 191 -2578 283 -2572
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 25 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
