magic
tech sky130A
magscale 1 2
timestamp 1669742938
<< error_p >>
rect 239800 589920 252400 590306
rect 239800 569760 272560 589920
rect 329000 585800 329800 586200
rect 328200 585200 329000 585800
rect 329800 585200 351200 585800
rect 324413 582638 328200 585200
rect 287400 569760 324413 582638
rect 239800 557600 279170 569760
rect 287400 557600 312880 569760
rect 351200 557600 351400 585200
rect 239800 552000 287400 557600
rect 349400 557328 351400 557600
rect 349340 557268 351400 557328
rect 348413 556600 351400 557268
rect 236238 549600 252400 552000
rect 270200 551000 287400 552000
rect 270200 549600 292720 551000
rect 236238 546133 312880 549600
rect 332947 546133 348413 556600
rect 236238 545468 272560 546133
rect 207200 529440 272560 545468
rect 280233 545468 312880 546133
rect 331964 545468 332947 546133
rect 280233 529440 331964 545468
rect 207200 515309 276513 529440
rect 280233 515309 321987 529440
rect 207200 512823 321987 515309
rect 207200 509280 252400 512823
rect 270205 510199 321987 512823
rect 207200 503200 232240 509280
rect 270205 508200 287400 510199
rect 321987 509200 323009 510199
rect 270205 503672 312880 508200
rect 270136 503666 270172 503672
rect 270196 503666 270256 503672
rect 269499 503200 270164 503666
rect 205706 502038 207200 503200
rect 267975 502161 269499 503200
rect 267914 502133 269499 502161
rect 204097 500787 205706 502038
rect 265924 500787 267914 502133
rect 232487 489120 265924 500787
rect 281253 489120 312880 503672
rect 232487 478162 252400 489120
rect 227756 474961 232487 478162
rect 227756 474940 227770 474961
rect 227317 474600 227770 474940
rect 226800 474341 227317 474600
rect 281253 471000 319647 489120
rect 319647 470852 319800 471000
use diffind_sam_bk  diffind_sam_bk_0
timestamp 1669742938
transform 1 0 1058800 0 1 650400
box -1058800 -650400 -498549 -59934
<< end >>
