magic
tech sky130A
magscale 1 2
timestamp 1668094176
<< error_p >>
rect -29 1041 29 1047
rect -29 1007 -17 1041
rect -29 1001 29 1007
rect -29 -1007 29 -1001
rect -29 -1041 -17 -1007
rect -29 -1047 29 -1041
<< nwell >>
rect -124 -1060 124 1060
<< pmos >>
rect -30 -960 30 960
<< pdiff >>
rect -88 948 -30 960
rect -88 -948 -76 948
rect -42 -948 -30 948
rect -88 -960 -30 -948
rect 30 948 88 960
rect 30 -948 42 948
rect 76 -948 88 948
rect 30 -960 88 -948
<< pdiffc >>
rect -76 -948 -42 948
rect 42 -948 76 948
<< poly >>
rect -33 1041 33 1057
rect -33 1007 -17 1041
rect 17 1007 33 1041
rect -33 991 33 1007
rect -30 960 30 991
rect -30 -991 30 -960
rect -33 -1007 33 -991
rect -33 -1041 -17 -1007
rect 17 -1041 33 -1007
rect -33 -1057 33 -1041
<< polycont >>
rect -17 1007 17 1041
rect -17 -1041 17 -1007
<< locali >>
rect -33 1007 -17 1041
rect 17 1007 33 1041
rect -76 948 -42 964
rect -76 -964 -42 -948
rect 42 948 76 964
rect 42 -964 76 -948
rect -33 -1041 -17 -1007
rect 17 -1041 33 -1007
<< viali >>
rect -17 1007 17 1041
rect -76 -948 -42 948
rect 42 -948 76 948
rect -17 -1041 17 -1007
<< metal1 >>
rect -29 1041 29 1047
rect -29 1007 -17 1041
rect 17 1007 29 1041
rect -29 1001 29 1007
rect -82 948 -36 960
rect -82 -948 -76 948
rect -42 -948 -36 948
rect -82 -960 -36 -948
rect 36 948 82 960
rect 36 -948 42 948
rect 76 -948 82 948
rect 36 -960 82 -948
rect -29 -1007 29 -1001
rect -29 -1041 -17 -1007
rect 17 -1041 29 -1007
rect -29 -1047 29 -1041
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9.6 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
