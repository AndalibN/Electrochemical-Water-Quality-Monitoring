magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -4276 20533 -3605 20836
rect 12158 20631 12815 20809
rect 12158 20533 12744 20631
rect -4316 20314 12744 20533
rect -4196 -496 -3660 20314
rect 12208 -448 12744 20314
rect -4286 -606 -3517 -496
rect 12121 -606 12887 -448
rect -4286 -825 12887 -606
rect -4286 -988 -3517 -825
rect 12121 -889 12887 -825
<< psubdiff >>
rect -4250 20787 -3631 20810
rect -4250 20507 -4198 20787
rect -4290 20447 -4198 20507
rect -3688 20507 -3631 20787
rect 12184 20719 12789 20783
rect 12184 20657 12258 20719
rect 12234 20507 12258 20657
rect -3688 20447 12258 20507
rect 12700 20657 12789 20719
rect -4290 20345 -4266 20447
rect -4290 20340 -4130 20345
rect -4170 -522 -4130 20340
rect -4260 -565 -4130 -522
rect -3688 20340 12258 20345
rect -3688 -522 -3686 20340
rect 12234 -474 12258 20340
rect 12147 -497 12258 -474
rect 12700 -474 12718 20657
rect 12700 -497 12861 -474
rect -3688 -565 -3543 -522
rect -4260 -939 -4198 -565
rect -3620 -632 -3543 -565
rect 12147 -632 12190 -497
rect -3620 -633 12190 -632
rect -3620 -799 12190 -735
rect -3620 -939 -3543 -799
rect 12147 -803 12190 -799
rect 12836 -803 12861 -497
rect 12147 -863 12861 -803
rect -4260 -962 -3543 -939
<< psubdiffcont >>
rect -4198 20447 -3688 20787
rect 12258 20447 12700 20719
rect -4266 20345 12700 20447
rect -4130 -565 -3688 20345
rect 12258 -497 12700 20345
rect -4198 -633 -3620 -565
rect 12190 -633 12836 -497
rect -4198 -735 12836 -633
rect -4198 -939 -3620 -735
rect 12190 -803 12836 -735
<< poly >>
rect 2953 20233 5250 20235
rect 2892 20190 5250 20233
rect 2892 20179 2965 20190
rect 3120 20180 5250 20190
rect 2892 20143 2958 20179
rect 5219 20104 5250 20180
rect 5219 20057 5388 20104
rect 8189 20102 8255 20113
rect 8189 20068 8205 20102
rect 8239 20068 8255 20102
rect 8189 20052 8255 20068
<< polycont >>
rect 8205 20068 8239 20102
<< locali >>
rect -4242 20787 -3639 20810
rect -4242 20507 -4198 20787
rect -4282 20447 -4198 20507
rect -3688 20507 -3639 20787
rect 12192 20719 12781 20783
rect 12192 20657 12258 20719
rect 12234 20507 12258 20657
rect -3688 20447 12258 20507
rect 12700 20657 12781 20719
rect -4282 20345 -4266 20447
rect -4282 20340 -4130 20345
rect -4170 -522 -4130 20340
rect -4252 -565 -4130 -522
rect -3688 20340 12258 20345
rect -3688 -522 -3686 20340
rect 8189 20130 8480 20147
rect 8189 20102 8432 20130
rect 8189 20068 8205 20102
rect 8239 20096 8432 20102
rect 8466 20096 8480 20130
rect 8239 20079 8480 20096
rect 8239 20068 8255 20079
rect 8189 20065 8255 20068
rect -2534 760 -2500 920
rect -2298 760 -2264 919
rect -2062 760 -2028 919
rect -1826 760 -1792 919
rect -1590 760 -1556 919
rect -1354 760 -1320 921
rect -2535 756 -1320 760
rect -2535 729 -1316 756
rect 253 729 287 869
rect -2535 722 287 729
rect -1350 710 287 722
rect 489 710 523 869
rect 725 710 759 870
rect 961 710 995 870
rect 1197 710 1231 869
rect 1433 710 1467 871
rect 1669 710 1703 870
rect 1905 710 1939 872
rect 2141 710 2175 870
rect 2377 710 2411 871
rect 2613 710 2647 870
rect 2849 710 2883 870
rect 3085 710 3119 871
rect -1350 687 3119 710
rect 253 681 3119 687
rect 253 676 3118 681
rect 5432 680 5466 839
rect 5668 680 5702 839
rect 5904 680 5938 840
rect 6140 680 6174 840
rect 6376 680 6410 839
rect 6612 680 6646 841
rect 6848 680 6882 840
rect 7084 680 7118 842
rect 7320 680 7354 840
rect 7556 680 7590 841
rect 7792 680 7826 840
rect 8028 680 8062 840
rect 8264 740 8298 841
rect 10072 754 10106 914
rect 10308 754 10342 913
rect 10544 754 10578 913
rect 10780 754 10814 913
rect 11016 754 11050 913
rect 11252 754 11286 915
rect 10071 740 11286 754
rect 8264 733 11286 740
rect 8264 716 11284 733
rect 8264 680 10108 716
rect 5432 646 10108 680
rect 8264 645 10108 646
rect 4416 -141 4485 -129
rect 4416 -175 4432 -141
rect 4466 -175 4485 -141
rect 4416 -181 4485 -175
rect -3688 -565 -3551 -522
rect -4252 -939 -4198 -565
rect -3620 -632 -3551 -565
rect 4424 -632 4473 -181
rect 12234 -474 12258 20340
rect 12155 -497 12258 -474
rect 12700 -474 12718 20657
rect 12700 -497 12853 -474
rect 12155 -632 12190 -497
rect -3620 -633 12190 -632
rect -3620 -799 12190 -735
rect -3620 -939 -3551 -799
rect -4252 -962 -3551 -939
rect 4404 -958 4479 -799
rect 12155 -803 12190 -799
rect 12836 -803 12853 -497
rect 12155 -863 12853 -803
rect 4162 -1382 4716 -958
<< viali >>
rect 8205 20068 8239 20102
rect 8432 20096 8466 20130
rect -2475 12944 -2441 12978
rect 4432 -175 4466 -141
<< metal1 >>
rect 1013 21003 1290 21034
rect 1013 20887 1033 21003
rect 1277 20887 1290 21003
rect 1013 20635 1290 20887
rect 7388 20987 7665 21018
rect 7388 20871 7408 20987
rect 7652 20871 7665 20987
rect 7388 20775 7665 20871
rect 1082 20265 1217 20635
rect 134 20185 1217 20265
rect -5344 12983 -5276 13020
rect -5344 12981 -4228 12983
rect -2526 12981 -2425 12984
rect -5344 12978 -2425 12981
rect -5344 12944 -2475 12978
rect -2441 12944 -2425 12978
rect -5344 12941 -2425 12944
rect -5344 12940 -4228 12941
rect -5344 12910 -5276 12940
rect -2526 12938 -2425 12941
rect -2416 671 -2382 12894
rect -2180 671 -2146 12894
rect -1944 671 -1910 12894
rect -1708 671 -1674 12894
rect -1472 671 -1438 12894
rect -2416 642 -1438 671
rect -2416 641 -1439 642
rect -2180 639 -2146 641
rect -1676 434 -1639 641
rect 135 519 169 20185
rect 371 519 405 20046
rect 607 519 641 20046
rect 843 519 877 20046
rect 1079 519 1113 20046
rect 1315 519 1349 20046
rect 1551 519 1585 20046
rect 1787 519 1821 20046
rect 2023 519 2057 20046
rect 2259 519 2293 20046
rect 2495 519 2529 20046
rect 2731 519 2765 20046
rect 2967 519 3001 20046
rect 5314 554 5348 20255
rect 7459 20198 7599 20775
rect 15446 20160 15862 20368
rect 12132 20155 15862 20160
rect 8412 20130 15862 20155
rect 8189 20102 8255 20117
rect 8189 20068 8205 20102
rect 8239 20068 8255 20102
rect 8189 20062 8255 20068
rect 8412 20096 8432 20130
rect 8466 20096 15862 20130
rect 8412 20072 15862 20096
rect 8412 20067 12157 20072
rect 5550 554 5584 20015
rect 5786 554 5820 20015
rect 6022 554 6056 20015
rect 6258 554 6292 20015
rect 6494 554 6528 20015
rect 6730 554 6764 20015
rect 6966 554 7000 20015
rect 7202 554 7236 20015
rect 7438 554 7472 20015
rect 7674 554 7708 20015
rect 7910 554 7944 20015
rect 8146 554 8180 20015
rect 15446 19928 15862 20072
rect 10125 13103 11384 13131
rect 10115 13058 11384 13103
rect 10115 12932 10178 13058
rect 11322 12974 11383 13058
rect 13040 12974 13108 13008
rect 11322 12956 13108 12974
rect 11330 12933 13108 12956
rect 13040 12898 13108 12933
rect 10190 657 10224 12888
rect 10426 657 10460 12888
rect 10662 657 10696 12888
rect 10898 657 10932 12888
rect 11134 657 11168 12888
rect 10189 623 11169 657
rect 135 485 3001 519
rect 5311 494 8182 554
rect 135 478 169 485
rect 371 479 405 485
rect 607 484 641 485
rect 1079 483 1113 485
rect 1315 484 1349 485
rect 1551 480 1585 485
rect 1787 481 1821 485
rect 2023 480 2057 485
rect 2259 482 2293 485
rect 2731 482 2765 485
rect 2967 481 3001 485
rect 10371 437 10416 623
rect 10371 436 10415 437
rect 9410 435 10415 436
rect 3876 434 10415 435
rect -1676 413 10415 434
rect -1668 400 10415 413
rect -1668 399 3884 400
rect 4420 -129 4476 400
rect 4416 -141 4485 -129
rect 4416 -175 4432 -141
rect 4466 -175 4485 -141
rect 4416 -181 4485 -175
<< via1 >>
rect 1033 20887 1277 21003
rect 7408 20871 7652 20987
<< metal2 >>
rect 992 21422 1310 21504
rect 992 21286 1043 21422
rect 1259 21286 1310 21422
rect 992 21003 1310 21286
rect 992 20887 1033 21003
rect 1277 20887 1310 21003
rect 992 20842 1310 20887
rect 7367 21406 7685 21488
rect 7367 21270 7418 21406
rect 7634 21270 7685 21406
rect 7367 20987 7685 21270
rect 7367 20871 7408 20987
rect 7652 20871 7685 20987
rect 7367 20826 7685 20871
<< via2 >>
rect 1043 21286 1259 21422
rect 7418 21270 7634 21406
<< metal3 >>
rect 957 22046 1336 22151
rect 957 21902 1030 22046
rect 1254 21902 1336 22046
rect 957 21422 1336 21902
rect 957 21286 1043 21422
rect 1259 21286 1336 21422
rect 957 21177 1336 21286
rect 7332 22030 7711 22135
rect 7332 21886 7405 22030
rect 7629 21886 7711 22030
rect 7332 21406 7711 21886
rect 7332 21270 7418 21406
rect 7634 21270 7711 21406
rect 7332 21161 7711 21270
<< via3 >>
rect 1030 21902 1254 22046
rect 7405 21886 7629 22030
<< metal4 >>
rect 914 22700 1362 22746
rect 914 22464 1024 22700
rect 1260 22464 1362 22700
rect 914 22046 1362 22464
rect 914 21902 1030 22046
rect 1254 21902 1362 22046
rect 914 21177 1362 21902
rect 7289 22684 7737 22730
rect 7289 22448 7399 22684
rect 7635 22448 7737 22684
rect 7289 22030 7737 22448
rect 7289 21886 7405 22030
rect 7629 21886 7737 22030
rect 7289 21178 7737 21886
rect 15656 21038 16374 21738
<< via4 >>
rect 1024 22464 1260 22700
rect 7399 22448 7635 22684
<< metal5 >>
rect 6820 23914 8416 24392
rect 6816 23910 8416 23914
rect 462 23894 1256 23908
rect 462 23536 2012 23894
rect 6364 23552 8416 23910
rect 6816 23550 8416 23552
rect 462 22908 1388 23536
rect 6820 23098 8416 23550
rect 888 22700 1388 22908
rect 7262 22762 7763 23098
rect 888 22464 1024 22700
rect 1260 22464 1388 22700
rect 888 22375 1388 22464
rect 7263 22684 7763 22762
rect 7263 22448 7399 22684
rect 7635 22448 7763 22684
rect 7263 22359 7763 22448
use sky130_fd_pr__nfet_01v8_MWCSZB  XM2
timestamp 1669522153
transform 1 0 10679 0 1 6900
box -645 -6088 645 6088
use sky130_fd_pr__nfet_01v8_TXCS3D  XM4
timestamp 1669522153
transform 1 0 6806 0 1 10426
box -1530 -9688 1530 9688
use ind_PA  ind_PA_0
timestamp 1669522153
transform -1 0 1668 0 -1 20710
box 1200 -12000 11600 -2200
use ind_PA  ind_PA_1
timestamp 1669522153
transform 1 0 7180 0 -1 21188
box 1200 -12000 11600 -2200
use sky130_fd_pr__nfet_01v8_MWCSZB  sky130_fd_pr__nfet_01v8_MWCSZB_0
timestamp 1669522153
transform 1 0 -1927 0 1 6906
box -645 -6088 645 6088
use sky130_fd_pr__nfet_01v8_TXCS3D  sky130_fd_pr__nfet_01v8_TXCS3D_0
timestamp 1669522153
transform 1 0 1627 0 1 10457
box -1530 -9688 1530 9688
<< labels >>
rlabel locali s 4162 -1382 4716 -958 4 GND
port 1 nsew
rlabel metal1 s -5344 12910 -5276 13020 4 Vin
port 2 nsew
rlabel metal1 s 13040 12898 13108 13008 4 Vina
port 3 nsew
rlabel metal1 s 15446 19928 15862 20368 4 Vb
port 4 nsew
rlabel metal4 s 15656 21038 16374 21738 4 VDD
port 5 nsew
<< end >>
