magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -213 -780 213 847
<< pmos >>
rect -119 47 -29 647
rect 29 47 119 647
rect -119 -718 -29 -118
rect 29 -718 119 -118
<< pdiff >>
rect -177 602 -119 647
rect -177 568 -165 602
rect -131 568 -119 602
rect -177 534 -119 568
rect -177 500 -165 534
rect -131 500 -119 534
rect -177 466 -119 500
rect -177 432 -165 466
rect -131 432 -119 466
rect -177 398 -119 432
rect -177 364 -165 398
rect -131 364 -119 398
rect -177 330 -119 364
rect -177 296 -165 330
rect -131 296 -119 330
rect -177 262 -119 296
rect -177 228 -165 262
rect -131 228 -119 262
rect -177 194 -119 228
rect -177 160 -165 194
rect -131 160 -119 194
rect -177 126 -119 160
rect -177 92 -165 126
rect -131 92 -119 126
rect -177 47 -119 92
rect -29 602 29 647
rect -29 568 -17 602
rect 17 568 29 602
rect -29 534 29 568
rect -29 500 -17 534
rect 17 500 29 534
rect -29 466 29 500
rect -29 432 -17 466
rect 17 432 29 466
rect -29 398 29 432
rect -29 364 -17 398
rect 17 364 29 398
rect -29 330 29 364
rect -29 296 -17 330
rect 17 296 29 330
rect -29 262 29 296
rect -29 228 -17 262
rect 17 228 29 262
rect -29 194 29 228
rect -29 160 -17 194
rect 17 160 29 194
rect -29 126 29 160
rect -29 92 -17 126
rect 17 92 29 126
rect -29 47 29 92
rect 119 602 177 647
rect 119 568 131 602
rect 165 568 177 602
rect 119 534 177 568
rect 119 500 131 534
rect 165 500 177 534
rect 119 466 177 500
rect 119 432 131 466
rect 165 432 177 466
rect 119 398 177 432
rect 119 364 131 398
rect 165 364 177 398
rect 119 330 177 364
rect 119 296 131 330
rect 165 296 177 330
rect 119 262 177 296
rect 119 228 131 262
rect 165 228 177 262
rect 119 194 177 228
rect 119 160 131 194
rect 165 160 177 194
rect 119 126 177 160
rect 119 92 131 126
rect 165 92 177 126
rect 119 47 177 92
rect -177 -163 -119 -118
rect -177 -197 -165 -163
rect -131 -197 -119 -163
rect -177 -231 -119 -197
rect -177 -265 -165 -231
rect -131 -265 -119 -231
rect -177 -299 -119 -265
rect -177 -333 -165 -299
rect -131 -333 -119 -299
rect -177 -367 -119 -333
rect -177 -401 -165 -367
rect -131 -401 -119 -367
rect -177 -435 -119 -401
rect -177 -469 -165 -435
rect -131 -469 -119 -435
rect -177 -503 -119 -469
rect -177 -537 -165 -503
rect -131 -537 -119 -503
rect -177 -571 -119 -537
rect -177 -605 -165 -571
rect -131 -605 -119 -571
rect -177 -639 -119 -605
rect -177 -673 -165 -639
rect -131 -673 -119 -639
rect -177 -718 -119 -673
rect -29 -163 29 -118
rect -29 -197 -17 -163
rect 17 -197 29 -163
rect -29 -231 29 -197
rect -29 -265 -17 -231
rect 17 -265 29 -231
rect -29 -299 29 -265
rect -29 -333 -17 -299
rect 17 -333 29 -299
rect -29 -367 29 -333
rect -29 -401 -17 -367
rect 17 -401 29 -367
rect -29 -435 29 -401
rect -29 -469 -17 -435
rect 17 -469 29 -435
rect -29 -503 29 -469
rect -29 -537 -17 -503
rect 17 -537 29 -503
rect -29 -571 29 -537
rect -29 -605 -17 -571
rect 17 -605 29 -571
rect -29 -639 29 -605
rect -29 -673 -17 -639
rect 17 -673 29 -639
rect -29 -718 29 -673
rect 119 -163 177 -118
rect 119 -197 131 -163
rect 165 -197 177 -163
rect 119 -231 177 -197
rect 119 -265 131 -231
rect 165 -265 177 -231
rect 119 -299 177 -265
rect 119 -333 131 -299
rect 165 -333 177 -299
rect 119 -367 177 -333
rect 119 -401 131 -367
rect 165 -401 177 -367
rect 119 -435 177 -401
rect 119 -469 131 -435
rect 165 -469 177 -435
rect 119 -503 177 -469
rect 119 -537 131 -503
rect 165 -537 177 -503
rect 119 -571 177 -537
rect 119 -605 131 -571
rect 165 -605 177 -571
rect 119 -639 177 -605
rect 119 -673 131 -639
rect 165 -673 177 -639
rect 119 -718 177 -673
<< pdiffc >>
rect -165 568 -131 602
rect -165 500 -131 534
rect -165 432 -131 466
rect -165 364 -131 398
rect -165 296 -131 330
rect -165 228 -131 262
rect -165 160 -131 194
rect -165 92 -131 126
rect -17 568 17 602
rect -17 500 17 534
rect -17 432 17 466
rect -17 364 17 398
rect -17 296 17 330
rect -17 228 17 262
rect -17 160 17 194
rect -17 92 17 126
rect 131 568 165 602
rect 131 500 165 534
rect 131 432 165 466
rect 131 364 165 398
rect 131 296 165 330
rect 131 228 165 262
rect 131 160 165 194
rect 131 92 165 126
rect -165 -197 -131 -163
rect -165 -265 -131 -231
rect -165 -333 -131 -299
rect -165 -401 -131 -367
rect -165 -469 -131 -435
rect -165 -537 -131 -503
rect -165 -605 -131 -571
rect -165 -673 -131 -639
rect -17 -197 17 -163
rect -17 -265 17 -231
rect -17 -333 17 -299
rect -17 -401 17 -367
rect -17 -469 17 -435
rect -17 -537 17 -503
rect -17 -605 17 -571
rect -17 -673 17 -639
rect 131 -197 165 -163
rect 131 -265 165 -231
rect 131 -333 165 -299
rect 131 -401 165 -367
rect 131 -469 165 -435
rect 131 -537 165 -503
rect 131 -605 165 -571
rect 131 -673 165 -639
<< poly >>
rect -119 798 -29 814
rect -119 764 -91 798
rect -57 764 -29 798
rect -119 647 -29 764
rect 29 798 119 814
rect 29 764 57 798
rect 91 764 119 798
rect 29 647 119 764
rect -119 -118 -29 47
rect 29 -118 119 47
rect -119 -741 -29 -718
rect 29 -741 119 -718
rect -119 -780 119 -741
<< polycont >>
rect -91 764 -57 798
rect 57 764 91 798
<< locali >>
rect -119 764 -91 798
rect -57 764 -29 798
rect 29 764 57 798
rect 91 764 119 798
rect -165 616 -131 651
rect -165 544 -131 568
rect -165 472 -131 500
rect -165 400 -131 432
rect -165 330 -131 364
rect -165 262 -131 294
rect -165 194 -131 222
rect -165 126 -131 150
rect -165 43 -131 78
rect -17 616 17 651
rect -17 544 17 568
rect -17 472 17 500
rect -17 400 17 432
rect -17 330 17 364
rect -17 262 17 294
rect -17 194 17 222
rect -17 126 17 150
rect -17 43 17 78
rect 131 616 165 651
rect 131 544 165 568
rect 131 472 165 500
rect 131 400 165 432
rect 131 330 165 364
rect 131 262 165 294
rect 131 194 165 222
rect 131 126 165 150
rect 131 43 165 78
rect -165 -149 -131 -114
rect -165 -221 -131 -197
rect -165 -293 -131 -265
rect -165 -365 -131 -333
rect -165 -435 -131 -401
rect -165 -503 -131 -471
rect -165 -571 -131 -543
rect -165 -639 -131 -615
rect -165 -722 -131 -687
rect -17 -149 17 -114
rect -17 -221 17 -197
rect -17 -293 17 -265
rect -17 -365 17 -333
rect -17 -435 17 -401
rect -17 -503 17 -471
rect -17 -571 17 -543
rect -17 -639 17 -615
rect -17 -722 17 -687
rect 131 -149 165 -114
rect 131 -221 165 -197
rect 131 -293 165 -265
rect 131 -365 165 -333
rect 131 -435 165 -401
rect 131 -503 165 -471
rect 131 -571 165 -543
rect 131 -639 165 -615
rect 131 -722 165 -687
<< viali >>
rect -91 764 -57 798
rect 57 764 91 798
rect -165 602 -131 616
rect -165 582 -131 602
rect -165 534 -131 544
rect -165 510 -131 534
rect -165 466 -131 472
rect -165 438 -131 466
rect -165 398 -131 400
rect -165 366 -131 398
rect -165 296 -131 328
rect -165 294 -131 296
rect -165 228 -131 256
rect -165 222 -131 228
rect -165 160 -131 184
rect -165 150 -131 160
rect -165 92 -131 112
rect -165 78 -131 92
rect -17 602 17 616
rect -17 582 17 602
rect -17 534 17 544
rect -17 510 17 534
rect -17 466 17 472
rect -17 438 17 466
rect -17 398 17 400
rect -17 366 17 398
rect -17 296 17 328
rect -17 294 17 296
rect -17 228 17 256
rect -17 222 17 228
rect -17 160 17 184
rect -17 150 17 160
rect -17 92 17 112
rect -17 78 17 92
rect 131 602 165 616
rect 131 582 165 602
rect 131 534 165 544
rect 131 510 165 534
rect 131 466 165 472
rect 131 438 165 466
rect 131 398 165 400
rect 131 366 165 398
rect 131 296 165 328
rect 131 294 165 296
rect 131 228 165 256
rect 131 222 165 228
rect 131 160 165 184
rect 131 150 165 160
rect 131 92 165 112
rect 131 78 165 92
rect -165 -163 -131 -149
rect -165 -183 -131 -163
rect -165 -231 -131 -221
rect -165 -255 -131 -231
rect -165 -299 -131 -293
rect -165 -327 -131 -299
rect -165 -367 -131 -365
rect -165 -399 -131 -367
rect -165 -469 -131 -437
rect -165 -471 -131 -469
rect -165 -537 -131 -509
rect -165 -543 -131 -537
rect -165 -605 -131 -581
rect -165 -615 -131 -605
rect -165 -673 -131 -653
rect -165 -687 -131 -673
rect -17 -163 17 -149
rect -17 -183 17 -163
rect -17 -231 17 -221
rect -17 -255 17 -231
rect -17 -299 17 -293
rect -17 -327 17 -299
rect -17 -367 17 -365
rect -17 -399 17 -367
rect -17 -469 17 -437
rect -17 -471 17 -469
rect -17 -537 17 -509
rect -17 -543 17 -537
rect -17 -605 17 -581
rect -17 -615 17 -605
rect -17 -673 17 -653
rect -17 -687 17 -673
rect 131 -163 165 -149
rect 131 -183 165 -163
rect 131 -231 165 -221
rect 131 -255 165 -231
rect 131 -299 165 -293
rect 131 -327 165 -299
rect 131 -367 165 -365
rect 131 -399 165 -367
rect 131 -469 165 -437
rect 131 -471 165 -469
rect 131 -537 165 -509
rect 131 -543 165 -537
rect 131 -605 165 -581
rect 131 -615 165 -605
rect 131 -673 165 -653
rect 131 -687 165 -673
<< metal1 >>
rect -115 798 -33 804
rect -115 764 -91 798
rect -57 764 -33 798
rect -115 758 -33 764
rect 33 798 115 804
rect 33 764 57 798
rect 91 764 115 798
rect 33 758 115 764
rect -171 616 -125 647
rect -171 582 -165 616
rect -131 582 -125 616
rect -171 544 -125 582
rect -171 510 -165 544
rect -131 510 -125 544
rect -171 472 -125 510
rect -171 438 -165 472
rect -131 438 -125 472
rect -171 400 -125 438
rect -171 366 -165 400
rect -131 366 -125 400
rect -171 328 -125 366
rect -171 294 -165 328
rect -131 294 -125 328
rect -171 256 -125 294
rect -171 222 -165 256
rect -131 222 -125 256
rect -171 184 -125 222
rect -171 150 -165 184
rect -131 150 -125 184
rect -171 112 -125 150
rect -171 78 -165 112
rect -131 78 -125 112
rect -171 47 -125 78
rect -23 616 23 647
rect -23 582 -17 616
rect 17 582 23 616
rect -23 544 23 582
rect -23 510 -17 544
rect 17 510 23 544
rect -23 472 23 510
rect -23 438 -17 472
rect 17 438 23 472
rect -23 400 23 438
rect -23 366 -17 400
rect 17 366 23 400
rect -23 328 23 366
rect -23 294 -17 328
rect 17 294 23 328
rect -23 256 23 294
rect -23 222 -17 256
rect 17 222 23 256
rect -23 184 23 222
rect -23 150 -17 184
rect 17 150 23 184
rect -23 112 23 150
rect -23 78 -17 112
rect 17 78 23 112
rect -23 47 23 78
rect 125 616 171 647
rect 125 582 131 616
rect 165 582 171 616
rect 125 544 171 582
rect 125 510 131 544
rect 165 510 171 544
rect 125 472 171 510
rect 125 438 131 472
rect 165 438 171 472
rect 125 400 171 438
rect 125 366 131 400
rect 165 366 171 400
rect 125 328 171 366
rect 125 294 131 328
rect 165 294 171 328
rect 125 256 171 294
rect 125 222 131 256
rect 165 222 171 256
rect 125 184 171 222
rect 125 150 131 184
rect 165 150 171 184
rect 125 112 171 150
rect 125 78 131 112
rect 165 78 171 112
rect 125 47 171 78
rect -171 -149 -125 -118
rect -171 -183 -165 -149
rect -131 -183 -125 -149
rect -171 -221 -125 -183
rect -171 -255 -165 -221
rect -131 -255 -125 -221
rect -171 -293 -125 -255
rect -171 -327 -165 -293
rect -131 -327 -125 -293
rect -171 -365 -125 -327
rect -171 -399 -165 -365
rect -131 -399 -125 -365
rect -171 -437 -125 -399
rect -171 -471 -165 -437
rect -131 -471 -125 -437
rect -171 -509 -125 -471
rect -171 -543 -165 -509
rect -131 -543 -125 -509
rect -171 -581 -125 -543
rect -171 -615 -165 -581
rect -131 -615 -125 -581
rect -171 -653 -125 -615
rect -171 -687 -165 -653
rect -131 -687 -125 -653
rect -171 -718 -125 -687
rect -23 -149 23 -118
rect -23 -183 -17 -149
rect 17 -183 23 -149
rect -23 -221 23 -183
rect -23 -255 -17 -221
rect 17 -255 23 -221
rect -23 -293 23 -255
rect -23 -327 -17 -293
rect 17 -327 23 -293
rect -23 -365 23 -327
rect -23 -399 -17 -365
rect 17 -399 23 -365
rect -23 -437 23 -399
rect -23 -471 -17 -437
rect 17 -471 23 -437
rect -23 -509 23 -471
rect -23 -543 -17 -509
rect 17 -543 23 -509
rect -23 -581 23 -543
rect -23 -615 -17 -581
rect 17 -615 23 -581
rect -23 -653 23 -615
rect -23 -687 -17 -653
rect 17 -687 23 -653
rect -23 -718 23 -687
rect 125 -149 171 -118
rect 125 -183 131 -149
rect 165 -183 171 -149
rect 125 -221 171 -183
rect 125 -255 131 -221
rect 165 -255 171 -221
rect 125 -293 171 -255
rect 125 -327 131 -293
rect 165 -327 171 -293
rect 125 -365 171 -327
rect 125 -399 131 -365
rect 165 -399 171 -365
rect 125 -437 171 -399
rect 125 -471 131 -437
rect 165 -471 171 -437
rect 125 -509 171 -471
rect 125 -543 131 -509
rect 165 -543 171 -509
rect 125 -581 171 -543
rect 125 -615 131 -581
rect 165 -615 171 -581
rect 125 -653 171 -615
rect 125 -687 131 -653
rect 165 -687 171 -653
rect 125 -718 171 -687
<< end >>
