magic
tech sky130A
magscale 1 2
timestamp 1667443641
<< nwell >>
rect -194 -2900 194 2900
<< pmos >>
rect -100 -2800 100 2800
<< pdiff >>
rect -158 2788 -100 2800
rect -158 -2788 -146 2788
rect -112 -2788 -100 2788
rect -158 -2800 -100 -2788
rect 100 2788 158 2800
rect 100 -2788 112 2788
rect 146 -2788 158 2788
rect 100 -2800 158 -2788
<< pdiffc >>
rect -146 -2788 -112 2788
rect 112 -2788 146 2788
<< poly >>
rect -100 2881 100 2897
rect -100 2847 -84 2881
rect 84 2847 100 2881
rect -100 2800 100 2847
rect -100 -2847 100 -2800
rect -100 -2881 -84 -2847
rect 84 -2881 100 -2847
rect -100 -2897 100 -2881
<< polycont >>
rect -84 2847 84 2881
rect -84 -2881 84 -2847
<< locali >>
rect -100 2847 -84 2881
rect 84 2847 100 2881
rect -146 2788 -112 2804
rect -146 -2804 -112 -2788
rect 112 2788 146 2804
rect 112 -2804 146 -2788
rect -100 -2881 -84 -2847
rect 84 -2881 100 -2847
<< viali >>
rect -84 2847 84 2881
rect -146 -2788 -112 2788
rect 112 -2788 146 2788
rect -84 -2881 84 -2847
<< metal1 >>
rect -96 2881 96 2887
rect -96 2847 -84 2881
rect 84 2847 96 2881
rect -96 2841 96 2847
rect -152 2788 -106 2800
rect -152 -2788 -146 2788
rect -112 -2788 -106 2788
rect -152 -2800 -106 -2788
rect 106 2788 152 2800
rect 106 -2788 112 2788
rect 146 -2788 152 2788
rect 106 -2800 152 -2788
rect -96 -2847 96 -2841
rect -96 -2881 -84 -2847
rect 84 -2881 96 -2847
rect -96 -2887 96 -2881
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 28 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
