magic
tech sky130A
magscale 1 2
timestamp 1667488624
<< error_p >>
rect -29 273 29 279
rect -29 239 -17 273
rect -29 233 29 239
rect -29 -239 29 -233
rect -29 -273 -17 -239
rect -29 -279 29 -273
<< nwell >>
rect -211 -411 211 411
<< pmos >>
rect -15 -192 15 192
<< pdiff >>
rect -73 180 -15 192
rect -73 -180 -61 180
rect -27 -180 -15 180
rect -73 -192 -15 -180
rect 15 180 73 192
rect 15 -180 27 180
rect 61 -180 73 180
rect 15 -192 73 -180
<< pdiffc >>
rect -61 -180 -27 180
rect 27 -180 61 180
<< nsubdiff >>
rect -175 341 -79 375
rect 79 341 175 375
rect -175 279 -141 341
rect 141 279 175 341
rect -175 -341 -141 -279
rect 141 -341 175 -279
rect -175 -375 -79 -341
rect 79 -375 175 -341
<< nsubdiffcont >>
rect -79 341 79 375
rect -175 -279 -141 279
rect 141 -279 175 279
rect -79 -375 79 -341
<< poly >>
rect -33 273 33 289
rect -33 239 -17 273
rect 17 239 33 273
rect -33 223 33 239
rect -15 192 15 223
rect -15 -223 15 -192
rect -33 -239 33 -223
rect -33 -273 -17 -239
rect 17 -273 33 -239
rect -33 -289 33 -273
<< polycont >>
rect -17 239 17 273
rect -17 -273 17 -239
<< locali >>
rect -175 341 -79 375
rect 79 341 175 375
rect -175 279 -141 341
rect 141 279 175 341
rect -33 239 -17 273
rect 17 239 33 273
rect -61 180 -27 196
rect -61 -196 -27 -180
rect 27 180 61 196
rect 27 -196 61 -180
rect -33 -273 -17 -239
rect 17 -273 33 -239
rect -175 -341 -141 -279
rect 141 -341 175 -279
rect -175 -375 -79 -341
rect 79 -375 175 -341
<< viali >>
rect -17 239 17 273
rect -61 -180 -27 180
rect 27 -180 61 180
rect -17 -273 17 -239
<< metal1 >>
rect -29 273 29 279
rect -29 239 -17 273
rect 17 239 29 273
rect -29 233 29 239
rect -67 180 -21 192
rect -67 -180 -61 180
rect -27 -180 -21 180
rect -67 -192 -21 -180
rect 21 180 67 192
rect 21 -180 27 180
rect 61 -180 67 180
rect 21 -192 67 -180
rect -29 -239 29 -233
rect -29 -273 -17 -239
rect 17 -273 29 -239
rect -29 -279 29 -273
<< properties >>
string FIXED_BBOX -158 -358 158 358
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.92 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
