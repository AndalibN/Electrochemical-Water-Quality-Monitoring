magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -129 -170 129 108
<< nmos >>
rect -45 -144 45 82
<< ndiff >>
rect -103 54 -45 82
rect -103 20 -91 54
rect -57 20 -45 54
rect -103 -14 -45 20
rect -103 -48 -91 -14
rect -57 -48 -45 -14
rect -103 -82 -45 -48
rect -103 -116 -91 -82
rect -57 -116 -45 -82
rect -103 -144 -45 -116
rect 45 54 103 82
rect 45 20 57 54
rect 91 20 103 54
rect 45 -14 103 20
rect 45 -48 57 -14
rect 91 -48 103 -14
rect 45 -82 103 -48
rect 45 -116 57 -82
rect 91 -116 103 -82
rect 45 -144 103 -116
<< ndiffc >>
rect -91 20 -57 54
rect -91 -48 -57 -14
rect -91 -116 -57 -82
rect 57 20 91 54
rect 57 -48 91 -14
rect 57 -116 91 -82
<< poly >>
rect -45 224 45 240
rect -45 190 -17 224
rect 17 190 45 224
rect -45 82 45 190
rect -45 -170 45 -144
<< polycont >>
rect -17 190 17 224
<< locali >>
rect -45 190 -17 224
rect 17 190 45 224
rect -91 58 -57 86
rect -91 -14 -57 20
rect -91 -82 -57 -48
rect -91 -148 -57 -120
rect 57 58 91 86
rect 57 -14 91 20
rect 57 -82 91 -48
rect 57 -148 91 -120
<< viali >>
rect -17 190 17 224
rect -91 54 -57 58
rect -91 24 -57 54
rect -91 -48 -57 -14
rect -91 -116 -57 -86
rect -91 -120 -57 -116
rect 57 54 91 58
rect 57 24 91 54
rect 57 -48 91 -14
rect 57 -116 91 -86
rect 57 -120 91 -116
<< metal1 >>
rect -41 224 41 230
rect -41 190 -17 224
rect 17 190 41 224
rect -41 184 41 190
rect -97 58 -51 82
rect -97 24 -91 58
rect -57 24 -51 58
rect -97 -14 -51 24
rect -97 -48 -91 -14
rect -57 -48 -51 -14
rect -97 -86 -51 -48
rect -97 -120 -91 -86
rect -57 -120 -51 -86
rect -97 -144 -51 -120
rect 51 58 97 82
rect 51 24 57 58
rect 91 24 97 58
rect 51 -14 97 24
rect 51 -48 57 -14
rect 91 -48 97 -14
rect 51 -86 97 -48
rect 51 -120 57 -86
rect 91 -120 97 -86
rect 51 -144 97 -120
<< end >>
