magic
tech sky130A
magscale 1 2
timestamp 1666877676
<< error_s >>
rect 2285 6356 2320 6390
rect 2286 6337 2320 6356
rect 468 3697 503 3731
rect 469 3678 503 3697
rect 488 583 503 3678
rect 522 3644 557 3678
rect 522 583 556 3644
rect 1008 2825 1042 2879
rect 1600 2861 1634 2879
rect 522 549 537 583
rect 1027 530 1042 2825
rect 1061 2791 1096 2825
rect 1061 530 1095 2791
rect 1061 496 1076 530
rect 1564 477 1634 2861
rect 1564 441 1617 477
rect 2305 424 2320 6337
rect 2339 6303 2374 6337
rect 2339 424 2373 6303
rect 3025 3484 3059 3538
rect 2339 390 2354 424
rect 3044 371 3059 3484
rect 3078 3450 3113 3484
rect 3563 3450 3598 3484
rect 3078 371 3112 3450
rect 3564 3431 3598 3450
rect 3078 337 3093 371
rect 3583 318 3598 3431
rect 3617 3397 3652 3431
rect 3617 318 3651 3397
rect 4103 1996 4137 2014
rect 4103 1960 4173 1996
rect 4120 1926 4191 1960
rect 4641 1926 4676 1960
rect 3617 284 3632 318
rect 4120 265 4190 1926
rect 4642 1907 4676 1926
rect 4120 229 4173 265
rect 4661 212 4676 1907
rect 4695 1873 4730 1907
rect 5180 1873 5215 1907
rect 4695 212 4729 1873
rect 5181 1854 5215 1873
rect 4695 178 4710 212
rect 5200 159 5215 1854
rect 5234 1820 5269 1854
rect 5719 1820 5754 1854
rect 5234 159 5268 1820
rect 5720 1801 5754 1820
rect 5234 125 5249 159
rect 5739 106 5754 1801
rect 5773 1767 5808 1801
rect 5773 106 5807 1767
rect 5773 72 5788 106
rect 6278 53 6293 1801
rect 6312 53 6346 1855
rect 6312 19 6327 53
rect 6817 0 6832 2348
rect 6851 0 6885 2402
rect 6851 -34 6866 0
use sky130_fd_pr__cap_mim_m3_1_WYFAV5  XC1
timestamp 1666877501
transform 1 0 7757 0 1 211
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_WYFAV5  XC2
timestamp 1666877501
transform 1 0 8995 0 1 158
box -350 -300 349 300
use sky130_fd_pr__nfet_01v8_RXXQKA  XM1
timestamp 1666877501
transform 1 0 243 0 1 2157
box -296 -1610 296 1610
use sky130_fd_pr__nfet_01v8_RXXQKA  XM2
timestamp 1666877501
transform 1 0 782 0 1 2104
box -296 -1610 296 1610
use sky130_fd_pr__nfet_01v8_6WXQK8  XM3
timestamp 1666877501
transform 1 0 1321 0 1 1651
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_5QDSA6  XM4
timestamp 1666877501
transform 1 0 1960 0 1 3407
box -396 -3019 396 3019
use sky130_fd_pr__pfet_01v8_5QDSA6  XM5
timestamp 1666877501
transform 1 0 2699 0 1 3354
box -396 -3019 396 3019
use sky130_fd_pr__pfet_01v8_GGN3CJ  XM6
timestamp 1666877501
transform 1 0 3338 0 1 1901
box -296 -1619 296 1619
use sky130_fd_pr__pfet_01v8_GGN3CJ  XM7
timestamp 1666877501
transform 1 0 3877 0 1 1848
box -296 -1619 296 1619
use sky130_fd_pr__nfet_01v8_XVAA4Y  XM8
timestamp 1666877501
transform 1 0 4416 0 1 1086
box -296 -910 296 910
use sky130_fd_pr__nfet_01v8_XVAA4Y  XM9
timestamp 1666877501
transform 1 0 4955 0 1 1033
box -296 -910 296 910
use sky130_fd_pr__nfet_01v8_XVAA4Y  XM10
timestamp 1666877501
transform 1 0 5494 0 1 980
box -296 -910 296 910
use sky130_fd_pr__nfet_01v8_XVAA4Y  XM11
timestamp 1666877501
transform 1 0 6033 0 1 927
box -296 -910 296 910
use sky130_fd_pr__nfet_01v8_U7E5KL  XM12
timestamp 1666877501
transform 1 0 7111 0 1 2921
box -296 -3010 296 3010
use sky130_fd_pr__pfet_01v8_3HPSVM  XM13
timestamp 1666877501
transform 1 0 8349 0 1 777
box -296 -919 296 919
use sky130_fd_pr__pfet_01v8_9QH3CS  XM14
timestamp 1666877501
transform 1 0 9687 0 1 1424
box -396 -1619 396 1619
use sky130_fd_pr__nfet_01v8_6WXQK8  XMB1
timestamp 1666877501
transform 1 0 6572 0 1 1174
box -296 -1210 296 1210
<< end >>
