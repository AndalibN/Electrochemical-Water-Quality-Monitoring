magic
tech sky130A
magscale 1 2
timestamp 1667588522
<< nwell >>
rect 6876 7686 7234 7690
rect 5410 7684 7636 7686
rect 478 7242 10376 7684
rect 472 5248 10376 7242
rect 474 5194 10376 5248
rect 474 5156 1062 5194
rect 474 5116 1060 5156
rect 520 5034 560 5102
rect 1320 2370 1708 5194
rect 1966 5168 10376 5194
rect 1966 5166 3012 5168
rect 3314 5166 10376 5168
rect 4360 5148 10376 5166
rect 8270 5112 8544 5148
rect 8540 4738 8544 5112
rect 1452 2368 1708 2370
rect 1454 2364 1708 2368
rect 1458 2248 1708 2364
rect 1630 2174 1708 2248
<< psubdiff >>
rect 6910 -3598 9628 -3596
rect 10018 -3598 10102 -3596
rect 13264 -3598 13664 -3596
rect -1908 -3600 -1878 -3598
rect -920 -3600 -702 -3598
rect 6910 -3600 10504 -3598
rect 11476 -3600 14238 -3598
rect -1908 -3628 14238 -3600
rect -1908 -3850 -1878 -3628
rect -1610 -3632 14238 -3628
rect -1610 -3662 -982 -3632
rect -1610 -3836 -1426 -3662
rect -1038 -3836 -982 -3662
rect -1610 -3848 -982 -3836
rect -628 -3634 14238 -3632
rect -628 -3640 11314 -3634
rect -628 -3646 9652 -3640
rect -628 -3832 2012 -3646
rect 2332 -3648 7540 -3646
rect 2332 -3832 2388 -3648
rect -628 -3840 2388 -3832
rect 2736 -3654 6930 -3648
rect 7080 -3654 7540 -3648
rect 2736 -3834 6022 -3654
rect 6284 -3834 6426 -3654
rect 2736 -3838 6426 -3834
rect 6698 -3834 6742 -3654
rect 7146 -3834 7540 -3654
rect 6698 -3838 7540 -3834
rect 2736 -3840 7540 -3838
rect -628 -3842 7540 -3840
rect 8038 -3838 8092 -3646
rect 8398 -3650 9652 -3646
rect 8398 -3826 8568 -3650
rect 9484 -3826 9652 -3650
rect 10346 -3652 11314 -3640
rect 8398 -3834 9652 -3826
rect 10398 -3834 11314 -3652
rect 11736 -3642 14238 -3634
rect 11736 -3644 13838 -3642
rect 11736 -3832 12412 -3644
rect 12910 -3646 13838 -3644
rect 12910 -3832 13030 -3646
rect 11736 -3834 13030 -3832
rect 13442 -3834 13838 -3646
rect 14164 -3834 14238 -3642
rect 8398 -3838 14238 -3834
rect 8038 -3842 14238 -3838
rect -628 -3848 14238 -3842
rect -1610 -3850 14238 -3848
rect -1908 -3860 14238 -3850
rect -1886 -3862 -876 -3860
<< nsubdiff >>
rect 6876 7596 7234 7602
rect 2940 7594 10336 7596
rect 514 7554 10336 7594
rect 514 7550 5854 7554
rect 514 7534 5310 7550
rect 514 7324 524 7534
rect 974 7520 5310 7534
rect 974 7336 2266 7520
rect 2710 7518 5310 7520
rect 2710 7336 3602 7518
rect 974 7332 3602 7336
rect 4054 7332 5310 7518
rect 974 7324 5310 7332
rect 514 7316 5310 7324
rect 5740 7316 5854 7550
rect 514 7300 5854 7316
rect 6142 7550 10336 7554
rect 6142 7310 6884 7550
rect 7212 7546 10336 7550
rect 7212 7310 7864 7546
rect 6142 7308 7864 7310
rect 8178 7308 8780 7546
rect 9094 7544 10336 7546
rect 9094 7308 9644 7544
rect 6142 7306 9644 7308
rect 9958 7306 10336 7544
rect 6142 7300 10336 7306
rect 514 7264 10336 7300
rect 2940 7262 4304 7264
rect 7584 7262 10336 7264
rect 3858 7260 3890 7262
<< psubdiffcont >>
rect -1878 -3850 -1610 -3628
rect -1426 -3836 -1038 -3662
rect -982 -3848 -628 -3632
rect 2012 -3832 2332 -3646
rect 2388 -3840 2736 -3648
rect 6930 -3654 7080 -3648
rect 6022 -3834 6284 -3654
rect 6426 -3838 6698 -3654
rect 6742 -3834 7146 -3654
rect 7540 -3842 8038 -3646
rect 8092 -3838 8398 -3646
rect 8568 -3826 9484 -3650
rect 9652 -3652 10346 -3640
rect 9652 -3834 10398 -3652
rect 11314 -3834 11736 -3634
rect 12412 -3832 12910 -3644
rect 13030 -3834 13442 -3646
rect 13838 -3834 14164 -3642
<< nsubdiffcont >>
rect 524 7324 974 7534
rect 2266 7336 2710 7520
rect 3602 7332 4054 7518
rect 5310 7316 5740 7550
rect 5854 7300 6142 7554
rect 6884 7310 7212 7550
rect 7864 7308 8178 7546
rect 8780 7308 9094 7546
rect 9644 7306 9958 7544
<< locali >>
rect 6876 7564 7234 7570
rect 524 7554 10320 7564
rect 524 7550 5854 7554
rect 524 7534 5310 7550
rect 974 7520 5310 7534
rect 974 7336 2266 7520
rect 2710 7518 5310 7520
rect 2710 7336 3602 7518
rect 974 7332 3602 7336
rect 4054 7332 5310 7518
rect 974 7324 5310 7332
rect 524 7316 5310 7324
rect 5740 7316 5854 7550
rect 524 7300 5854 7316
rect 6142 7550 10320 7554
rect 6142 7310 6884 7550
rect 7212 7546 10320 7550
rect 7212 7310 7864 7546
rect 6142 7308 7864 7310
rect 8178 7308 8780 7546
rect 9094 7544 10320 7546
rect 9094 7308 9644 7544
rect 6142 7306 9644 7308
rect 9958 7306 10320 7544
rect 6142 7300 10320 7306
rect 524 7294 10320 7300
rect 524 7264 564 7294
rect 522 5444 564 7264
rect 2474 7248 2512 7294
rect 3824 7248 3858 7294
rect 2470 5444 2510 7248
rect 522 5202 560 5444
rect 2470 5220 2508 5444
rect 522 5098 558 5202
rect 2472 5086 2506 5220
rect 3820 5214 3858 7248
rect 5456 7248 5494 7294
rect 5680 7292 7568 7294
rect 5456 7048 5490 7248
rect 5914 7064 5948 7292
rect 6944 7266 6984 7292
rect 6944 7254 6982 7266
rect 6946 7078 6980 7254
rect 5946 7056 5948 7064
rect 8002 7054 8036 7294
rect 8866 7064 8900 7294
rect 9714 7066 9748 7294
rect 8002 7048 8034 7054
rect 8866 7042 8898 7064
rect 9714 7040 9746 7066
rect 3818 5090 3858 5214
rect 5456 5082 5490 5132
rect -1166 4712 -1086 4796
rect 10290 4320 10340 4322
rect 10290 4278 11146 4320
rect 1242 4150 1450 4158
rect 1242 4122 1460 4150
rect -2190 -1660 -2152 1302
rect 1092 1152 1170 1174
rect 1242 1152 1276 4122
rect 4280 3252 5096 3328
rect 4280 3250 4362 3252
rect 4468 3100 4790 3144
rect 3390 1190 3392 1200
rect 1014 1118 1276 1152
rect 1660 1146 2014 1182
rect 1092 1112 1170 1118
rect 968 1012 1372 1048
rect 1092 810 1168 874
rect 1104 630 1152 810
rect 1920 730 1960 1146
rect 2922 1106 2982 1178
rect 3220 1116 3362 1190
rect 3364 1120 3392 1190
rect 2710 1056 3460 1058
rect 2710 1024 3408 1056
rect 2240 950 2310 1024
rect 3562 1008 3676 1082
rect 3980 950 4040 1036
rect 4150 1004 4240 1070
rect 2240 880 4040 950
rect 4468 844 4544 3100
rect 4736 3044 4790 3100
rect 5026 2750 5096 3252
rect 10196 3116 10220 3156
rect 9340 3044 9798 3046
rect 8636 3040 8960 3044
rect 5876 3034 7472 3036
rect 8420 3034 8960 3040
rect 5876 2998 8120 3034
rect 5876 2996 7472 2998
rect 7994 2996 8120 2998
rect 8330 2996 8960 3034
rect 9272 3032 9798 3044
rect 9030 3000 9798 3032
rect 9030 2998 9498 3000
rect 8400 2994 8960 2996
rect 8420 2988 8960 2994
rect 5026 2692 8190 2750
rect 5026 2690 5286 2692
rect 5026 2594 5096 2690
rect 4926 2534 5228 2594
rect 8140 2586 8190 2692
rect 8698 2588 9676 2590
rect 8698 2586 9736 2588
rect 10290 2586 10340 4278
rect 11088 4026 11146 4278
rect 8140 2518 10340 2586
rect 8140 2516 9736 2518
rect 8140 2514 9676 2516
rect 6520 1872 6560 2372
rect 6520 1432 6562 1872
rect 6956 1706 7034 1726
rect 6956 1662 6972 1706
rect 7018 1662 7034 1706
rect 6956 1648 7034 1662
rect 8140 1712 8218 1720
rect 8140 1664 8156 1712
rect 8200 1664 8218 1712
rect 8140 1652 8218 1664
rect 3220 766 4544 844
rect 4700 972 4744 1006
rect 1660 650 1684 720
rect 1920 690 3510 730
rect 3460 636 3510 690
rect 4700 660 4742 972
rect 3930 630 4742 660
rect 1104 594 1268 630
rect 1104 526 1152 594
rect -864 348 -828 466
rect 1232 350 1268 594
rect 3930 608 4740 630
rect 3320 490 3354 580
rect 3930 400 3980 608
rect 3784 352 4094 400
rect 3784 350 4066 352
rect 3784 348 3818 350
rect -910 346 -828 348
rect -910 338 -822 346
rect -910 262 -820 338
rect -2190 -1698 -1980 -1660
rect -2190 -1700 -2152 -1698
rect -2040 -1700 -1980 -1698
rect -2020 -3372 -1980 -1700
rect -1800 -2184 -1742 -1674
rect -1800 -2242 -1118 -2184
rect -2020 -3420 -1732 -3372
rect -1800 -3622 -1732 -3420
rect -1374 -3622 -1314 -2884
rect -1158 -3622 -1090 -3286
rect -910 -3622 -860 262
rect 930 30 974 214
rect 928 -4 1478 30
rect 2512 4 2590 6
rect 1418 -6 1478 -4
rect 2510 -8 2590 4
rect 2510 -60 2524 -8
rect 2574 -60 2590 -8
rect 2510 -68 2590 -60
rect 2512 -70 2590 -68
rect 2104 -142 2164 -140
rect 2096 -220 2168 -142
rect 2104 -1876 2164 -220
rect 6120 -1404 6154 274
rect 2104 -1880 2168 -1876
rect 6120 -1880 6156 -1404
rect 6520 -1880 6560 1432
rect 6796 -1880 6864 1556
rect 7652 1298 7732 1580
rect 6950 1196 7026 1214
rect 6950 1154 6968 1196
rect 7008 1154 7026 1196
rect 6950 1138 7026 1154
rect 8140 1202 8214 1222
rect 8140 1162 8158 1202
rect 8194 1162 8214 1202
rect 8140 1148 8214 1162
rect 7078 928 7246 1088
rect 6948 860 7026 880
rect 6948 814 6970 860
rect 7008 814 7026 860
rect 6948 800 7026 814
rect 8140 864 8216 872
rect 8140 822 8154 864
rect 8196 822 8216 864
rect 8140 806 8216 822
rect 7644 448 7724 730
rect 6948 344 7026 360
rect 6948 304 6966 344
rect 7010 304 7026 344
rect 6948 290 7026 304
rect 8142 348 8218 364
rect 8142 306 8156 348
rect 8194 306 8218 348
rect 8142 292 8218 306
rect 6940 20 7040 42
rect 6940 -46 6954 20
rect 7016 -46 7040 20
rect 6940 -56 7040 -46
rect 8134 8 8214 18
rect 8134 -36 8150 8
rect 8198 -36 8214 8
rect 8134 -50 8214 -36
rect 7642 -400 7722 -118
rect 11462 -416 11532 316
rect 6954 -492 7038 -474
rect 6954 -532 6978 -492
rect 7014 -532 7038 -492
rect 6954 -548 7038 -532
rect 8140 -488 8214 -472
rect 8140 -530 8156 -488
rect 8194 -530 8214 -488
rect 8140 -540 8214 -530
rect 6956 -828 7030 -812
rect 6956 -874 6974 -828
rect 7014 -874 7030 -828
rect 6956 -888 7030 -874
rect 8138 -828 8216 -814
rect 8138 -876 8154 -828
rect 8194 -876 8216 -828
rect 8138 -890 8216 -876
rect 2106 -2494 2168 -1880
rect -1894 -3624 -698 -3622
rect 2106 -3624 2170 -2494
rect 6122 -2500 6156 -1880
rect 6522 -2500 6558 -1880
rect 6798 -2500 6864 -1880
rect 7638 -2496 7724 -980
rect 7640 -2500 7724 -2496
rect 6122 -2558 6158 -2500
rect 6120 -3624 6160 -2558
rect 6522 -3624 6562 -2500
rect 6798 -3624 6866 -2500
rect 7640 -3624 7726 -2500
rect 9380 -2674 9420 -1448
rect 8918 -3624 8974 -3014
rect 9380 -3150 9418 -2674
rect 10440 -2930 10516 -2732
rect 10440 -2968 11026 -2930
rect 10440 -2970 10516 -2968
rect 9380 -3188 9846 -3150
rect 10984 -3162 11026 -2968
rect 9782 -3544 9846 -3188
rect 10200 -3380 10274 -3168
rect 10984 -3202 11024 -3162
rect 10200 -3442 10700 -3380
rect 9782 -3622 9844 -3544
rect 10200 -3546 10258 -3442
rect 10200 -3588 10256 -3546
rect 10200 -3622 10258 -3588
rect 11462 -3622 11520 -416
rect 11610 -1960 12210 -1956
rect 11610 -2010 12218 -1960
rect 12428 -2010 12486 -136
rect 13390 -1932 13448 -574
rect 14172 -1580 14238 -706
rect 14048 -1660 14238 -1580
rect 14048 -1668 14110 -1660
rect 13184 -1984 13448 -1932
rect 13390 -1986 13448 -1984
rect 11610 -2012 12210 -2010
rect 11610 -3622 11676 -2012
rect 12430 -3622 12482 -2010
rect 13132 -2472 13188 -2108
rect 13132 -3622 13186 -2472
rect 13922 -3622 13970 -1968
rect 14050 -3622 14110 -1668
rect 9598 -3624 10504 -3622
rect 11462 -3624 11958 -3622
rect 12400 -3624 14238 -3622
rect -1894 -3628 14238 -3624
rect -1894 -3850 -1878 -3628
rect -1610 -3632 14238 -3628
rect -1610 -3662 -982 -3632
rect -1610 -3836 -1426 -3662
rect -1038 -3836 -982 -3662
rect -1610 -3848 -982 -3836
rect -628 -3634 14238 -3632
rect -628 -3640 11314 -3634
rect -628 -3646 9652 -3640
rect -628 -3832 2012 -3646
rect 2332 -3648 7540 -3646
rect 2332 -3832 2388 -3648
rect 2736 -3654 6930 -3648
rect 7080 -3654 7540 -3648
rect -628 -3840 2388 -3832
rect 2736 -3834 6022 -3654
rect 6284 -3834 6426 -3654
rect 2736 -3838 6426 -3834
rect 6698 -3834 6742 -3654
rect 7146 -3834 7540 -3654
rect 6698 -3838 7540 -3834
rect 2736 -3840 7540 -3838
rect -628 -3842 7540 -3840
rect 8038 -3838 8092 -3646
rect 8398 -3650 9652 -3646
rect 8398 -3826 8568 -3650
rect 9484 -3826 9652 -3650
rect 10346 -3652 11314 -3640
rect 8398 -3834 9652 -3826
rect 10398 -3834 11314 -3652
rect 11736 -3642 14238 -3634
rect 11736 -3644 13838 -3642
rect 11736 -3832 12412 -3644
rect 12910 -3646 13838 -3644
rect 12910 -3832 13030 -3646
rect 11736 -3834 13030 -3832
rect 13442 -3834 13838 -3646
rect 14164 -3834 14238 -3642
rect 8398 -3838 14238 -3834
rect 8038 -3842 14238 -3838
rect -628 -3848 14238 -3842
rect -1610 -3850 14238 -3848
rect -1894 -3852 -872 -3850
<< viali >>
rect 6972 1662 7018 1706
rect 8156 1664 8200 1712
rect 2524 -60 2574 -8
rect 6968 1154 7008 1196
rect 8158 1162 8194 1202
rect 6970 814 7008 860
rect 8154 822 8196 864
rect 6966 304 7010 344
rect 8156 306 8194 348
rect 6954 -46 7016 20
rect 8150 -36 8198 8
rect 6978 -532 7014 -492
rect 8156 -530 8194 -488
rect 6974 -874 7014 -828
rect 8154 -876 8194 -828
rect 2526 -3778 2572 -3728
rect 6970 -3734 7010 -3688
rect 8148 -3768 8200 -3712
<< metal1 >>
rect 524 7264 564 7534
rect 2476 7320 2510 7520
rect 522 5444 564 7264
rect 2474 7248 2512 7320
rect 3824 7248 3858 7518
rect 5460 7328 5494 7550
rect 2470 5444 2510 7248
rect 522 5202 560 5444
rect 2470 5220 2508 5444
rect 522 5070 558 5202
rect 2472 5086 2506 5220
rect 3820 5214 3858 7248
rect 5456 7248 5494 7328
rect 5456 7048 5490 7248
rect 5914 7064 5948 7476
rect 6946 7330 6984 7548
rect 6944 7266 6984 7330
rect 8002 7294 8034 7428
rect 8866 7294 8898 7442
rect 9714 7294 9746 7440
rect 6944 7254 6982 7266
rect 6946 7078 6980 7254
rect 5946 7056 5948 7064
rect 8002 7054 8036 7294
rect 8866 7064 8900 7294
rect 9714 7066 9748 7294
rect 8002 7048 8034 7054
rect 8866 7042 8898 7064
rect 9714 7040 9746 7066
rect 3818 5090 3858 5214
rect 5456 5080 5490 5132
rect -1166 4788 -1086 4796
rect -1166 4786 -1152 4788
rect -1166 4722 -1154 4786
rect -1100 4724 -1086 4788
rect -1102 4722 -1086 4724
rect -1166 4712 -1086 4722
rect 10290 4320 10340 4322
rect 10290 4278 11146 4320
rect 1242 4150 1450 4158
rect 1242 4122 1460 4150
rect -2190 -1660 -2152 1302
rect 1092 1168 1170 1174
rect 1092 1152 1106 1168
rect 980 1118 1106 1152
rect 1092 1116 1106 1118
rect 1158 1152 1170 1168
rect 1242 1152 1276 4122
rect 4280 3252 5096 3328
rect 4280 3250 4362 3252
rect 4468 3100 4790 3144
rect 3390 1190 3392 1200
rect 1158 1118 1276 1152
rect 1626 1146 2048 1184
rect 3220 1180 3362 1190
rect 2922 1172 2982 1178
rect 1158 1116 1170 1118
rect 1092 1112 1170 1116
rect 584 1014 1406 1048
rect 1368 1010 1402 1014
rect 1362 934 1408 950
rect 1362 928 1420 934
rect 1414 876 1420 928
rect 1092 868 1168 874
rect 1092 816 1098 868
rect 1162 816 1168 868
rect 1362 842 1408 876
rect 1092 810 1168 816
rect 1104 630 1152 810
rect 1920 730 1960 1146
rect 2922 1114 2926 1172
rect 2978 1114 2982 1172
rect 3220 1128 3230 1180
rect 3300 1128 3362 1180
rect 3220 1116 3362 1128
rect 3364 1120 3392 1190
rect 2922 1106 2982 1114
rect 3562 1074 3676 1082
rect 2240 1054 2320 1056
rect 2240 950 2310 1054
rect 2706 1024 3468 1058
rect 3562 1016 3584 1074
rect 3656 1016 3676 1074
rect 4150 1064 4240 1070
rect 3562 1008 3676 1016
rect 3980 950 4040 1036
rect 4150 1012 4160 1064
rect 4230 1012 4240 1064
rect 4150 1004 4240 1012
rect 2240 942 4040 950
rect 2240 890 2250 942
rect 2310 890 4040 942
rect 2240 880 4040 890
rect 4468 844 4544 3100
rect 4736 3044 4790 3100
rect 5026 2750 5096 3252
rect 7402 3172 7462 3178
rect 7400 3158 7462 3172
rect 10164 3168 10230 3170
rect 7400 3100 7406 3158
rect 7460 3100 7462 3158
rect 9308 3154 9368 3162
rect 7400 3094 7462 3100
rect 8446 3142 8506 3148
rect 8446 3090 8454 3142
rect 9308 3102 9316 3154
rect 10164 3116 10172 3168
rect 10224 3116 10230 3168
rect 10164 3106 10230 3116
rect 9308 3092 9368 3102
rect 8446 3080 8506 3090
rect 5610 3052 5680 3060
rect 5610 3000 5620 3052
rect 5672 3000 5680 3052
rect 9340 3044 9798 3046
rect 8636 3040 8960 3044
rect 5610 2990 5680 3000
rect 5876 3034 7472 3036
rect 8420 3034 8960 3040
rect 5876 2998 8120 3034
rect 5876 2996 7472 2998
rect 7994 2996 8120 2998
rect 8330 2996 8960 3034
rect 9272 3032 9798 3044
rect 9030 3000 9798 3032
rect 9030 2998 9498 3000
rect 8400 2994 8960 2996
rect 8420 2988 8960 2994
rect 5026 2692 8190 2750
rect 5026 2690 5286 2692
rect 5026 2594 5096 2690
rect 4926 2534 5228 2594
rect 7550 2592 7620 2600
rect 7550 2536 7558 2592
rect 7610 2536 7620 2592
rect 7550 2530 7620 2536
rect 8140 2586 8190 2692
rect 8698 2588 9676 2590
rect 8698 2586 9736 2588
rect 10290 2586 10340 4278
rect 11088 4026 11146 4278
rect 8140 2518 10340 2586
rect 8140 2516 9736 2518
rect 8140 2514 9676 2516
rect 6520 1872 6560 2372
rect 6520 1432 6562 1872
rect 6956 1716 7034 1726
rect 6956 1656 6966 1716
rect 7026 1656 7034 1716
rect 6956 1648 7034 1656
rect 8140 1714 8218 1720
rect 8140 1660 8150 1714
rect 8206 1660 8218 1714
rect 8140 1652 8218 1660
rect 8900 1632 8992 1660
rect 3220 836 4544 844
rect 3220 774 3234 836
rect 3306 774 3570 836
rect 3220 768 3570 774
rect 3672 768 4544 836
rect 3220 766 4544 768
rect 4700 972 4744 1006
rect 1618 712 1684 720
rect 1618 660 1626 712
rect 1678 660 1684 712
rect 1920 690 3510 730
rect 1618 652 1684 660
rect 1660 650 1684 652
rect 3460 636 3510 690
rect 4700 660 4742 972
rect 3930 630 4742 660
rect 1104 594 1268 630
rect 1104 526 1152 594
rect -864 348 -828 466
rect 1232 350 1268 594
rect 3930 608 4740 630
rect 3320 550 3354 580
rect 3300 542 3368 550
rect 3300 490 3310 542
rect 3362 490 3368 542
rect 3300 482 3368 490
rect 3930 400 3980 608
rect 4150 512 4252 514
rect 4150 460 4168 512
rect 4240 460 4252 512
rect 4150 450 4252 460
rect 3784 352 4094 400
rect 3784 350 4066 352
rect 3784 348 3818 350
rect -910 346 -828 348
rect -910 338 -822 346
rect -910 262 -820 338
rect -2190 -1698 -1980 -1660
rect -2190 -1700 -2152 -1698
rect -2040 -1700 -1980 -1698
rect -2020 -3372 -1980 -1700
rect -1800 -2184 -1742 -1674
rect -1800 -2242 -1118 -2184
rect -2020 -3420 -1732 -3372
rect -1800 -3792 -1732 -3420
rect -1374 -3748 -1314 -2884
rect -1158 -3758 -1090 -3286
rect -910 -3828 -860 262
rect -746 226 -744 228
rect -788 202 -744 226
rect 930 30 974 214
rect 1616 180 1690 192
rect 1616 110 1624 180
rect 1676 110 1690 180
rect 1616 88 1690 110
rect 928 -4 1478 30
rect 2512 4 2590 6
rect 1418 -6 1478 -4
rect 2510 -4 2590 4
rect 2510 -64 2520 -4
rect 2580 -64 2590 -4
rect 2510 -68 2590 -64
rect 2512 -70 2590 -68
rect 2096 -142 2164 -140
rect 2096 -220 2168 -142
rect 2104 -1876 2164 -220
rect 6120 -1404 6154 274
rect 2104 -1880 2168 -1876
rect 6120 -1880 6156 -1404
rect 6520 -1880 6560 1432
rect 6796 -1880 6864 1556
rect 7652 1298 7732 1580
rect 8900 1560 8920 1632
rect 8972 1560 8992 1632
rect 8900 1542 8992 1560
rect 12158 1322 12278 1334
rect 12158 1238 12170 1322
rect 12258 1238 12278 1322
rect 12158 1230 12176 1238
rect 12244 1230 12278 1238
rect 6950 1204 7026 1214
rect 6950 1150 6958 1204
rect 7016 1150 7026 1204
rect 6950 1138 7026 1150
rect 8140 1210 8214 1222
rect 12158 1216 12278 1230
rect 8140 1158 8154 1210
rect 8206 1158 8214 1210
rect 8140 1148 8214 1158
rect 7078 1074 7246 1088
rect 7078 942 7092 1074
rect 7226 942 7246 1074
rect 7078 928 7246 942
rect 13110 894 13216 898
rect 13104 892 13216 894
rect 6948 868 7026 880
rect 6948 808 6958 868
rect 7014 808 7026 868
rect 6948 800 7026 808
rect 8140 870 8216 872
rect 8140 818 8150 870
rect 8202 818 8216 870
rect 13104 820 13118 892
rect 8140 806 8216 818
rect 13110 812 13118 820
rect 13206 812 13216 892
rect 13110 804 13216 812
rect 7644 448 7724 730
rect 13900 724 13988 726
rect 13900 670 13910 724
rect 13980 670 13988 724
rect 13900 664 13988 670
rect 6948 352 7026 360
rect 6948 296 6960 352
rect 7014 296 7026 352
rect 6948 290 7026 296
rect 8142 356 8218 364
rect 8142 300 8144 356
rect 8204 300 8218 356
rect 8142 292 8218 300
rect 6940 26 7040 42
rect 6940 -50 6950 26
rect 7024 -50 7040 26
rect 8134 12 8214 18
rect 8134 -40 8142 12
rect 8202 -40 8214 12
rect 8134 -50 8214 -40
rect 6940 -56 7040 -50
rect 7642 -400 7722 -118
rect 11462 -416 11532 316
rect 6954 -484 7038 -474
rect 6954 -538 6970 -484
rect 7022 -538 7038 -484
rect 6954 -548 7038 -538
rect 8140 -480 8214 -472
rect 8140 -532 8152 -480
rect 8204 -532 8214 -480
rect 8140 -540 8214 -532
rect 6956 -822 7030 -812
rect 6956 -880 6968 -822
rect 7020 -880 7030 -822
rect 6956 -888 7030 -880
rect 8138 -824 8216 -814
rect 8138 -884 8148 -824
rect 8202 -884 8216 -824
rect 8138 -890 8216 -884
rect 2106 -2494 2168 -1880
rect 2106 -3822 2170 -2494
rect 6122 -2500 6156 -1880
rect 6522 -2500 6558 -1880
rect 6798 -2500 6864 -1880
rect 7638 -2496 7724 -980
rect 7640 -2500 7724 -2496
rect 6122 -2558 6158 -2500
rect 2512 -3718 2590 -3704
rect 2512 -3784 2524 -3718
rect 2578 -3784 2590 -3718
rect 6120 -3744 6160 -2558
rect 2512 -3792 2590 -3784
rect 6522 -3834 6562 -2500
rect 6798 -3784 6866 -2500
rect 6958 -3680 7030 -3672
rect 6958 -3740 6964 -3680
rect 7018 -3740 7030 -3680
rect 6958 -3748 7030 -3740
rect 7640 -3826 7726 -2500
rect 9380 -2674 9420 -1448
rect 8136 -3700 8230 -3690
rect 8136 -3772 8146 -3700
rect 8206 -3772 8230 -3700
rect 8136 -3778 8230 -3772
rect 8918 -3778 8974 -3014
rect 9380 -3150 9418 -2674
rect 10440 -2930 10516 -2732
rect 10440 -2968 11026 -2930
rect 10440 -2970 10516 -2968
rect 9380 -3188 9846 -3150
rect 10984 -3162 11026 -2968
rect 9782 -3544 9846 -3188
rect 10200 -3380 10274 -3168
rect 10984 -3202 11024 -3162
rect 10200 -3442 10700 -3380
rect 9782 -3640 9844 -3544
rect 10200 -3546 10258 -3442
rect 10200 -3588 10256 -3546
rect 10200 -3640 10258 -3588
rect 9786 -3826 9842 -3640
rect 10202 -3824 10258 -3640
rect 11462 -3766 11520 -416
rect 11610 -1960 12210 -1956
rect 11610 -2010 12218 -1960
rect 12428 -2010 12486 -136
rect 13390 -1932 13448 -574
rect 14172 -1580 14238 -706
rect 14048 -1660 14238 -1580
rect 14048 -1668 14110 -1660
rect 13184 -1984 13448 -1932
rect 13390 -1986 13448 -1984
rect 11610 -2012 12210 -2010
rect 11610 -3776 11676 -2012
rect 12430 -3770 12482 -2010
rect 13132 -2472 13188 -2108
rect 13132 -3814 13186 -2472
rect 13922 -3814 13970 -1968
rect 14050 -3752 14110 -1668
<< via1 >>
rect -1152 4786 -1100 4788
rect -1154 4724 -1100 4786
rect -1154 4722 -1102 4724
rect 1106 1116 1158 1168
rect 1362 876 1414 928
rect 1098 816 1162 868
rect 2926 1114 2978 1172
rect 3230 1128 3300 1180
rect 3584 1016 3656 1074
rect 4160 1012 4230 1064
rect 2250 890 2310 942
rect 7406 3100 7460 3158
rect 8454 3090 8506 3142
rect 9316 3102 9368 3154
rect 10172 3116 10224 3168
rect 5620 3000 5672 3052
rect 7558 2536 7610 2592
rect 7114 1806 7218 1912
rect 7960 1808 8058 1914
rect 6966 1706 7026 1716
rect 6966 1662 6972 1706
rect 6972 1662 7018 1706
rect 7018 1662 7026 1706
rect 6966 1656 7026 1662
rect 8150 1712 8206 1714
rect 8150 1664 8156 1712
rect 8156 1664 8200 1712
rect 8200 1664 8206 1712
rect 8150 1660 8206 1664
rect 3234 774 3306 836
rect 3570 768 3672 836
rect 1626 660 1678 712
rect 3310 490 3362 542
rect 4168 460 4240 512
rect 1624 110 1676 180
rect 2334 94 2434 190
rect 2520 -8 2580 -4
rect 2520 -60 2524 -8
rect 2524 -60 2574 -8
rect 2574 -60 2580 -8
rect 2520 -64 2580 -60
rect 8920 1560 8972 1632
rect 12170 1238 12258 1322
rect 12176 1230 12244 1238
rect 6958 1196 7016 1204
rect 6958 1154 6968 1196
rect 6968 1154 7008 1196
rect 7008 1154 7016 1196
rect 6958 1150 7016 1154
rect 8154 1202 8206 1210
rect 8154 1162 8158 1202
rect 8158 1162 8194 1202
rect 8194 1162 8206 1202
rect 8154 1158 8206 1162
rect 7092 942 7226 1074
rect 7954 962 8052 1068
rect 6958 860 7014 868
rect 6958 814 6970 860
rect 6970 814 7008 860
rect 7008 814 7014 860
rect 6958 808 7014 814
rect 8150 864 8202 870
rect 8150 822 8154 864
rect 8154 822 8196 864
rect 8196 822 8202 864
rect 8150 818 8202 822
rect 13118 812 13206 892
rect 13910 670 13980 724
rect 6960 344 7014 352
rect 6960 304 6966 344
rect 6966 304 7010 344
rect 7010 304 7014 344
rect 6960 296 7014 304
rect 8144 348 8204 356
rect 8144 306 8156 348
rect 8156 306 8194 348
rect 8194 306 8204 348
rect 8144 300 8204 306
rect 7108 106 7210 208
rect 7954 106 8052 212
rect 6950 20 7024 26
rect 6950 -46 6954 20
rect 6954 -46 7016 20
rect 7016 -46 7024 20
rect 6950 -50 7024 -46
rect 8142 8 8202 12
rect 8142 -36 8150 8
rect 8150 -36 8198 8
rect 8198 -36 8202 8
rect 8142 -40 8202 -36
rect 6970 -492 7022 -484
rect 6970 -532 6978 -492
rect 6978 -532 7014 -492
rect 7014 -532 7022 -492
rect 6970 -538 7022 -532
rect 8152 -488 8204 -480
rect 8152 -530 8156 -488
rect 8156 -530 8194 -488
rect 8194 -530 8204 -488
rect 8152 -532 8204 -530
rect 7112 -734 7214 -632
rect 7954 -732 8056 -630
rect 6968 -828 7020 -822
rect 6968 -874 6974 -828
rect 6974 -874 7014 -828
rect 7014 -874 7020 -828
rect 6968 -880 7020 -874
rect 8148 -828 8202 -824
rect 8148 -876 8154 -828
rect 8154 -876 8194 -828
rect 8194 -876 8202 -828
rect 8148 -884 8202 -876
rect 2524 -3728 2578 -3718
rect 2524 -3778 2526 -3728
rect 2526 -3778 2572 -3728
rect 2572 -3778 2578 -3728
rect 2524 -3784 2578 -3778
rect 6964 -3688 7018 -3680
rect 6964 -3734 6970 -3688
rect 6970 -3734 7010 -3688
rect 7010 -3734 7018 -3688
rect 6964 -3740 7018 -3734
rect 8146 -3712 8206 -3700
rect 8146 -3768 8148 -3712
rect 8148 -3768 8200 -3712
rect 8200 -3768 8206 -3712
rect 8146 -3772 8206 -3768
<< metal2 >>
rect -1168 4788 -522 4798
rect -1168 4786 -1152 4788
rect -1168 4722 -1154 4786
rect -1100 4724 -522 4788
rect -1102 4722 -522 4724
rect -1168 4712 -522 4722
rect -580 2966 -522 4712
rect 10164 3174 10388 3176
rect 10164 3168 10390 3174
rect 7400 3162 7462 3168
rect 7398 3160 7462 3162
rect 7398 3158 7932 3160
rect 7398 3100 7406 3158
rect 7460 3100 7932 3158
rect 9308 3154 9496 3162
rect 7398 3096 7932 3100
rect 7398 3094 7462 3096
rect 5610 3052 5680 3060
rect 5610 3000 5620 3052
rect 5672 3000 5680 3052
rect -580 722 -510 2966
rect 5610 2920 5680 3000
rect 4382 2880 5680 2920
rect 2924 1180 2966 1182
rect 3220 1180 3310 1190
rect 1092 1168 1170 1174
rect 1092 1116 1106 1168
rect 1158 1116 1170 1168
rect 1092 874 1170 1116
rect 2924 1172 3120 1180
rect 2924 1114 2926 1172
rect 2978 1114 3120 1172
rect 2924 1102 3120 1114
rect 2924 1100 2966 1102
rect 3050 950 3120 1102
rect 1348 948 3120 950
rect 3220 1128 3230 1180
rect 3300 1128 3310 1180
rect 1348 942 3122 948
rect 1348 928 2250 942
rect 1348 876 1362 928
rect 1414 890 2250 928
rect 2310 890 3122 942
rect 1414 876 3122 890
rect 1092 868 1168 874
rect 1092 816 1098 868
rect 1162 816 1168 868
rect 1348 846 3122 876
rect 3220 926 3310 1128
rect 3560 1074 3680 1082
rect 3560 1016 3584 1074
rect 3656 1016 3680 1074
rect 1348 842 3120 846
rect 1092 810 1168 816
rect -580 712 1684 722
rect -580 660 1626 712
rect 1678 660 1684 712
rect -580 650 1684 660
rect 3050 550 3120 842
rect 3220 836 3312 926
rect 3220 774 3234 836
rect 3306 774 3312 836
rect 3220 766 3312 774
rect 3560 836 3680 1016
rect 4150 1064 4240 1070
rect 4150 1012 4160 1064
rect 4230 1012 4240 1064
rect 4150 970 4240 1012
rect 4382 970 4420 2880
rect 7550 2592 7630 2600
rect 7550 2536 7558 2592
rect 7610 2536 7630 2592
rect 7550 2400 7630 2536
rect 7102 2350 7630 2400
rect 7892 2422 7932 3096
rect 8446 3142 8636 3150
rect 8446 3090 8454 3142
rect 8506 3090 8636 3142
rect 9308 3102 9316 3154
rect 9368 3102 9496 3154
rect 10164 3116 10172 3168
rect 10224 3116 10390 3168
rect 10164 3106 10390 3116
rect 9308 3092 9496 3102
rect 8446 3080 8636 3090
rect 8596 2770 8636 3080
rect 9456 2902 9496 3092
rect 9456 2900 9642 2902
rect 9456 2860 10160 2900
rect 8596 2730 10020 2770
rect 8290 2424 8330 2426
rect 8290 2422 8650 2424
rect 7892 2382 8650 2422
rect 7102 1920 7222 2350
rect 8574 2156 8650 2382
rect 9980 2288 10020 2730
rect 8574 2054 9012 2156
rect 8570 2052 9012 2054
rect 8570 2038 8690 2052
rect 8570 1956 8582 2038
rect 8670 1956 8690 2038
rect 8570 1934 8690 1956
rect 7102 1912 7226 1920
rect 7102 1806 7114 1912
rect 7218 1806 7226 1912
rect 7102 1798 7226 1806
rect 7100 1796 7226 1798
rect 7942 1914 8072 1926
rect 7942 1808 7960 1914
rect 8058 1808 8072 1914
rect 6956 1716 7034 1726
rect 6956 1658 6966 1716
rect 6950 1656 6966 1658
rect 7026 1656 7034 1716
rect 6950 1648 7034 1656
rect 6950 1204 7026 1648
rect 6950 1150 6958 1204
rect 7016 1150 7026 1204
rect 6950 1138 7026 1150
rect 7100 1094 7224 1796
rect 4150 930 4420 970
rect 7078 1074 7246 1094
rect 7078 942 7092 1074
rect 7226 942 7246 1074
rect 7078 928 7246 942
rect 7942 1068 8072 1808
rect 8140 1714 8218 1720
rect 8140 1660 8150 1714
rect 8206 1660 8218 1714
rect 8140 1652 8218 1660
rect 8142 1222 8210 1652
rect 8890 1632 9012 2052
rect 8890 1560 8920 1632
rect 8972 1560 9012 1632
rect 8890 1542 9012 1560
rect 9980 1262 10018 2288
rect 10120 1452 10160 2860
rect 10346 1570 10390 3106
rect 10346 1530 13610 1570
rect 10346 1528 10390 1530
rect 12328 1452 12872 1454
rect 10120 1408 12872 1452
rect 10120 1406 10160 1408
rect 12158 1322 12278 1334
rect 12158 1262 12170 1322
rect 9980 1238 12170 1262
rect 12258 1238 12278 1322
rect 9980 1230 12176 1238
rect 12244 1230 12278 1238
rect 8140 1210 8214 1222
rect 9980 1220 12278 1230
rect 12158 1216 12278 1220
rect 8140 1158 8154 1210
rect 8206 1158 8214 1210
rect 8140 1148 8214 1158
rect 12778 1210 12872 1408
rect 7942 962 7954 1068
rect 8052 962 8072 1068
rect 3560 768 3570 836
rect 3672 800 3680 836
rect 6948 868 7026 880
rect 6948 808 6958 868
rect 7014 808 7026 868
rect 6948 800 7026 808
rect 3672 768 4260 800
rect 3560 740 4260 768
rect 3926 738 4260 740
rect 3050 542 3368 550
rect 3050 490 3310 542
rect 3362 490 3368 542
rect 3050 480 3368 490
rect 4150 512 4260 738
rect 4150 460 4168 512
rect 4240 460 4260 512
rect 4150 450 4260 460
rect 6948 360 7024 800
rect 6948 352 7026 360
rect 6948 296 6960 352
rect 7014 296 7026 352
rect 6948 290 7026 296
rect 7102 208 7224 928
rect 2318 190 2450 206
rect 1616 180 2334 190
rect 1616 110 1624 180
rect 1676 110 2334 180
rect 1616 94 2334 110
rect 2434 94 2450 190
rect 1616 88 2450 94
rect 2318 74 2450 88
rect 7102 106 7108 208
rect 7210 106 7224 208
rect 6940 26 7040 42
rect 2508 -4 2592 6
rect 2508 -64 2520 -4
rect 2580 -64 2592 -4
rect 6940 -50 6950 26
rect 7024 -50 7040 26
rect 6940 -56 7040 -50
rect 2508 -68 2592 -64
rect 2512 -3718 2592 -68
rect 6950 -474 7030 -56
rect 6950 -476 7038 -474
rect 6954 -484 7038 -476
rect 6954 -538 6970 -484
rect 7022 -538 7038 -484
rect 6954 -548 7038 -538
rect 7102 -616 7224 106
rect 7942 212 8072 962
rect 12778 922 12870 1210
rect 12778 900 13198 922
rect 12778 892 13220 900
rect 8140 870 8216 872
rect 8140 818 8150 870
rect 8202 818 8216 870
rect 12778 832 13118 892
rect 8140 806 8216 818
rect 13102 810 13118 832
rect 13206 810 13220 892
rect 8142 364 8216 806
rect 13106 788 13220 810
rect 13500 752 13610 1530
rect 13890 752 14000 754
rect 13500 744 14002 752
rect 13500 662 13900 744
rect 13988 662 14002 744
rect 13500 644 14002 662
rect 13888 642 14002 644
rect 8142 356 8218 364
rect 8142 300 8144 356
rect 8204 300 8218 356
rect 8142 292 8218 300
rect 7942 106 7954 212
rect 8052 106 8072 212
rect 7942 -616 8072 106
rect 8134 12 8214 18
rect 8134 -40 8142 12
rect 8202 -40 8214 12
rect 8134 -50 8214 -40
rect 8140 -480 8214 -50
rect 8140 -532 8152 -480
rect 8204 -532 8214 -480
rect 8140 -540 8214 -532
rect 7100 -630 8072 -616
rect 7100 -632 7954 -630
rect 7100 -734 7112 -632
rect 7214 -732 7954 -632
rect 8056 -732 8072 -630
rect 7214 -734 8072 -732
rect 7100 -750 8072 -734
rect 6956 -822 7030 -812
rect 6956 -880 6968 -822
rect 7020 -880 7030 -822
rect 6956 -888 7030 -880
rect 2512 -3784 2524 -3718
rect 2578 -3784 2592 -3718
rect 6958 -3680 7030 -888
rect 8138 -824 8216 -814
rect 8138 -884 8148 -824
rect 8202 -884 8216 -824
rect 8138 -890 8216 -884
rect 6958 -3740 6964 -3680
rect 7018 -3740 7030 -3680
rect 8140 -3690 8216 -890
rect 6958 -3748 7030 -3740
rect 8136 -3700 8230 -3690
rect 8136 -3772 8146 -3700
rect 8206 -3772 8230 -3700
rect 8136 -3778 8230 -3772
rect 2512 -3794 2592 -3784
<< via2 >>
rect 8582 1956 8670 2038
rect 12170 1238 12258 1320
rect 13118 812 13206 892
rect 13118 810 13206 812
rect 13900 724 13988 744
rect 13900 670 13910 724
rect 13910 670 13980 724
rect 13980 670 13988 724
rect 13900 662 13988 670
<< metal3 >>
rect 8572 2040 8684 2046
rect 8572 1956 8582 2040
rect 8670 1956 8684 2040
rect 8572 1944 8684 1956
rect 12160 1322 12272 1328
rect 12160 1238 12170 1322
rect 12258 1238 12272 1322
rect 12160 1226 12272 1238
rect 13108 894 13220 900
rect 13108 810 13118 894
rect 13206 810 13220 894
rect 13108 798 13220 810
rect 13890 746 14002 752
rect 13890 662 13900 746
rect 13988 662 14002 746
rect 13890 650 14002 662
<< via3 >>
rect 8582 2038 8670 2040
rect 8582 1956 8670 2038
rect 12170 1320 12258 1322
rect 12170 1238 12258 1320
rect 13118 892 13206 894
rect 13118 810 13206 892
rect 13900 744 13988 746
rect 13900 662 13988 744
<< metal4 >>
rect 8572 2040 8684 2046
rect 8572 1956 8582 2040
rect 8670 1956 8684 2040
rect 8572 1948 8684 1956
rect 8570 1858 8684 1948
rect 13978 1858 14200 2120
rect 8570 1798 14200 1858
rect 14280 1328 14530 1612
rect 12158 1322 14530 1328
rect 12158 1238 12170 1322
rect 12258 1238 14530 1322
rect 12158 1216 14530 1238
rect 14970 920 15220 1244
rect 13106 894 15220 920
rect 13106 810 13118 894
rect 13206 860 15220 894
rect 13206 858 13810 860
rect 13206 810 13220 858
rect 13106 788 13220 810
rect 13888 746 14002 752
rect 13888 662 13900 746
rect 13988 702 14002 746
rect 15462 702 15700 956
rect 13988 662 15700 702
rect 13888 642 15700 662
use 298k  R1 /research/mlab/chipathon/magic_design_files
timestamp 1666627716
transform 1 0 6899 0 1 335
box 0 0 1 1
use 52k  R2 /research/mlab/chipathon/magic_design_files
timestamp 1666627716
transform 1 0 6895 0 1 335
box 0 0 1 1
use 485k  R3 /research/mlab/chipathon/magic_design_files
timestamp 1666627716
transform 1 0 6896 0 1 335
box 0 0 1 1
use 520k  R4 /research/mlab/chipathon/magic_design_files
timestamp 1666627716
transform 1 0 6897 0 1 335
box 0 0 1 1
use 520k  R5
timestamp 1666627716
transform 1 0 6898 0 1 335
box 0 0 1 1
use 295k  R6 /research/mlab/chipathon/magic_design_files
timestamp 1666627716
transform 1 0 8517 0 1 176
box 0 0 1 1
use 298k  R7
timestamp 1666627716
transform 1 0 8518 0 1 176
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_E8XWE6  XM7 /research/mlab/chipathon/magic_design_files
timestamp 1666896002
transform 1 0 4066 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__nfet_01v8_VYYYB6  XM8 /research/mlab/chipathon/magic_design_files
timestamp 1666901352
transform 1 0 3568 0 1 -387
box -258 -1057 258 1057
use sky130_fd_pr__nfet_01v8_2HQT3D  XM10 /research/mlab/chipathon/magic_design_files
timestamp 1667411627
transform 1 0 5106 0 1 361
box -1058 -157 1058 157
use sky130_fd_pr__pfet_01v8_6PERLV  XM11 /research/mlab/chipathon/magic_design_files
timestamp 1667408630
transform 1 0 7194 0 1 5054
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  XM12 /research/mlab/chipathon/magic_design_files
timestamp 1666810850
transform 1 0 2260 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1653785680
transform 1 0 1986 0 1 -258
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ2
timestamp 1653785680
transform 1 0 6768 0 1 1458
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ3
timestamp 1653785680
transform 1 0 6762 0 1 610
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ4
timestamp 1653785680
transform 1 0 6762 0 1 -242
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ5
timestamp 1653785680
transform 1 0 6766 0 1 -1080
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ6
timestamp 1653785680
transform 1 0 7608 0 1 -1078
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ7
timestamp 1653785680
transform 1 0 7608 0 1 -242
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ8
timestamp 1653785680
transform 1 0 7608 0 1 614
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ10
timestamp 1653785680
transform 1 0 7612 0 1 1462
box 0 0 796 796
use res2_529K  res2_529K_0 /research/mlab/chipathon/magic_design_files
timestamp 1667425878
transform 0 -1 11356 1 0 -3218
box -258 0 74 1174
use res2_529K  res2_529K_1
timestamp 1667425878
transform 1 0 -1160 0 1 -3322
box -258 0 74 1174
use res52_504  res52_504_0 /research/mlab/chipathon/magic_design_files
timestamp 1667019087
transform 0 -1 7872 1 0 2530
box -202 0 74 2664
use res54_789k  res54_789k_0 /research/mlab/chipathon/magic_design_files
timestamp 1667400688
transform -1 0 10486 0 -1 3662
box -3806 2918 -3420 5662
use res63_92k  res63_92k_0 /research/mlab/chipathon/magic_design_files
timestamp 1667400564
transform -1 0 9706 0 -1 3838
box -3806 2918 -3420 6106
use res298k  res298k_0 /research/mlab/chipathon/magic_design_files
timestamp 1667400309
transform -1 0 8744 0 -1 4252
box -3806 2918 -3420 6312
use res484_3K  res484_3K_0 /research/mlab/chipathon/magic_design_files
timestamp 1667399187
transform -1 0 8984 0 -1 1656
box -654 0 74 4764
use res517_512K  res517_512K_0 /research/mlab/chipathon/magic_design_files
timestamp 1667019531
transform 1 0 -1806 0 1 -1726
box -608 0 710 6864
use res517_512K  res517_512K_1
timestamp 1667019531
transform -1 0 11156 0 -1 4084
box -608 0 710 6864
use sky130_fd_pr__nfet_01v8_7ZFCMD  sky130_fd_pr__nfet_01v8_7ZFCMD_0 /research/mlab/chipathon/magic_design_files
timestamp 1666810850
transform 1 0 188 0 1 366
box -1058 -188 1058 188
use sky130_fd_pr__nfet_01v8_7ZFCMD  sky130_fd_pr__nfet_01v8_7ZFCMD_1
timestamp 1666810850
transform 0 -1 4786 1 0 2020
box -1058 -188 1058 188
use sky130_fd_pr__pfet_01v8_6HAMAW  sky130_fd_pr__pfet_01v8_6HAMAW_0 /research/mlab/chipathon/magic_design_files
timestamp 1667404707
transform 1 0 1514 0 1 2074
box -194 -2100 194 2100
use sky130_fd_pr__pfet_01v8_A42UEE  sky130_fd_pr__pfet_01v8_A42UEE_0 /research/mlab/chipathon/magic_design_files
timestamp 1666810850
transform 1 0 768 0 1 3058
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_0
timestamp 1666810850
transform 1 0 2718 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_1
timestamp 1666810850
transform 1 0 3608 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_2
timestamp 1666810850
transform 1 0 5702 0 1 5044
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_3
timestamp 1666810850
transform 1 0 8248 0 1 5042
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_4
timestamp 1666810850
transform 1 0 9112 0 1 5050
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_5
timestamp 1666810850
transform 1 0 9960 0 1 5054
box -294 -2064 294 2098
use sky130_fd_pr__res_xhigh_po_0p35_L4QNDW  sky130_fd_pr__res_xhigh_po_0p35_L4QNDW_0
timestamp 1667588522
transform 1 0 15204 0 1 8563
box -196 -4977 196 4977
<< labels >>
rlabel metal1 3792 894 3914 942 1 G11
rlabel locali 4382 7394 4704 7548 1 Vdd
rlabel metal1 4570 3258 4762 3312 1 SM7
rlabel metal2 7130 2248 7198 2372 1 Q2
rlabel metal1 4334 616 4406 648 1 SM9
rlabel metal2 4174 678 4244 750 1 G10
rlabel metal4 14018 1848 14140 2008 1 Vout
rlabel metal4 15036 912 15128 1078 1 Vref2
rlabel metal4 15500 672 15620 828 1 Vref3
rlabel locali 3472 -3784 3790 -3664 1 GND
rlabel metal4 13996 1240 14198 1326 1 Vref1
rlabel metal1 1118 596 1194 624 1 G1
rlabel metal1 2388 702 2476 726 1 G9
rlabel metal1 10634 -2954 10676 -2936 1 R2
rlabel metal1 -1588 -2224 -1486 -2196 1 R7
<< end >>
