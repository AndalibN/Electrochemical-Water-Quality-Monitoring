magic
tech sky130A
magscale 1 2
timestamp 1668369161
<< error_p >>
rect -3277 6072 -3219 6078
rect -3045 6072 -2987 6078
rect -2813 6072 -2755 6078
rect -2581 6072 -2523 6078
rect -2349 6072 -2291 6078
rect -2117 6072 -2059 6078
rect -1885 6072 -1827 6078
rect -1653 6072 -1595 6078
rect -1421 6072 -1363 6078
rect -1189 6072 -1131 6078
rect -957 6072 -899 6078
rect -725 6072 -667 6078
rect -493 6072 -435 6078
rect -261 6072 -203 6078
rect -29 6072 29 6078
rect 203 6072 261 6078
rect 435 6072 493 6078
rect 667 6072 725 6078
rect 899 6072 957 6078
rect 1131 6072 1189 6078
rect 1363 6072 1421 6078
rect 1595 6072 1653 6078
rect 1827 6072 1885 6078
rect 2059 6072 2117 6078
rect 2291 6072 2349 6078
rect 2523 6072 2581 6078
rect 2755 6072 2813 6078
rect 2987 6072 3045 6078
rect 3219 6072 3277 6078
rect -3277 6038 -3265 6072
rect -3045 6038 -3033 6072
rect -2813 6038 -2801 6072
rect -2581 6038 -2569 6072
rect -2349 6038 -2337 6072
rect -2117 6038 -2105 6072
rect -1885 6038 -1873 6072
rect -1653 6038 -1641 6072
rect -1421 6038 -1409 6072
rect -1189 6038 -1177 6072
rect -957 6038 -945 6072
rect -725 6038 -713 6072
rect -493 6038 -481 6072
rect -261 6038 -249 6072
rect -29 6038 -17 6072
rect 203 6038 215 6072
rect 435 6038 447 6072
rect 667 6038 679 6072
rect 899 6038 911 6072
rect 1131 6038 1143 6072
rect 1363 6038 1375 6072
rect 1595 6038 1607 6072
rect 1827 6038 1839 6072
rect 2059 6038 2071 6072
rect 2291 6038 2303 6072
rect 2523 6038 2535 6072
rect 2755 6038 2767 6072
rect 2987 6038 2999 6072
rect 3219 6038 3231 6072
rect -3277 6032 -3219 6038
rect -3045 6032 -2987 6038
rect -2813 6032 -2755 6038
rect -2581 6032 -2523 6038
rect -2349 6032 -2291 6038
rect -2117 6032 -2059 6038
rect -1885 6032 -1827 6038
rect -1653 6032 -1595 6038
rect -1421 6032 -1363 6038
rect -1189 6032 -1131 6038
rect -957 6032 -899 6038
rect -725 6032 -667 6038
rect -493 6032 -435 6038
rect -261 6032 -203 6038
rect -29 6032 29 6038
rect 203 6032 261 6038
rect 435 6032 493 6038
rect 667 6032 725 6038
rect 899 6032 957 6038
rect 1131 6032 1189 6038
rect 1363 6032 1421 6038
rect 1595 6032 1653 6038
rect 1827 6032 1885 6038
rect 2059 6032 2117 6038
rect 2291 6032 2349 6038
rect 2523 6032 2581 6038
rect 2755 6032 2813 6038
rect 2987 6032 3045 6038
rect 3219 6032 3277 6038
rect -3277 -6038 -3219 -6032
rect -3045 -6038 -2987 -6032
rect -2813 -6038 -2755 -6032
rect -2581 -6038 -2523 -6032
rect -2349 -6038 -2291 -6032
rect -2117 -6038 -2059 -6032
rect -1885 -6038 -1827 -6032
rect -1653 -6038 -1595 -6032
rect -1421 -6038 -1363 -6032
rect -1189 -6038 -1131 -6032
rect -957 -6038 -899 -6032
rect -725 -6038 -667 -6032
rect -493 -6038 -435 -6032
rect -261 -6038 -203 -6032
rect -29 -6038 29 -6032
rect 203 -6038 261 -6032
rect 435 -6038 493 -6032
rect 667 -6038 725 -6032
rect 899 -6038 957 -6032
rect 1131 -6038 1189 -6032
rect 1363 -6038 1421 -6032
rect 1595 -6038 1653 -6032
rect 1827 -6038 1885 -6032
rect 2059 -6038 2117 -6032
rect 2291 -6038 2349 -6032
rect 2523 -6038 2581 -6032
rect 2755 -6038 2813 -6032
rect 2987 -6038 3045 -6032
rect 3219 -6038 3277 -6032
rect -3277 -6072 -3265 -6038
rect -3045 -6072 -3033 -6038
rect -2813 -6072 -2801 -6038
rect -2581 -6072 -2569 -6038
rect -2349 -6072 -2337 -6038
rect -2117 -6072 -2105 -6038
rect -1885 -6072 -1873 -6038
rect -1653 -6072 -1641 -6038
rect -1421 -6072 -1409 -6038
rect -1189 -6072 -1177 -6038
rect -957 -6072 -945 -6038
rect -725 -6072 -713 -6038
rect -493 -6072 -481 -6038
rect -261 -6072 -249 -6038
rect -29 -6072 -17 -6038
rect 203 -6072 215 -6038
rect 435 -6072 447 -6038
rect 667 -6072 679 -6038
rect 899 -6072 911 -6038
rect 1131 -6072 1143 -6038
rect 1363 -6072 1375 -6038
rect 1595 -6072 1607 -6038
rect 1827 -6072 1839 -6038
rect 2059 -6072 2071 -6038
rect 2291 -6072 2303 -6038
rect 2523 -6072 2535 -6038
rect 2755 -6072 2767 -6038
rect 2987 -6072 2999 -6038
rect 3219 -6072 3231 -6038
rect -3277 -6078 -3219 -6072
rect -3045 -6078 -2987 -6072
rect -2813 -6078 -2755 -6072
rect -2581 -6078 -2523 -6072
rect -2349 -6078 -2291 -6072
rect -2117 -6078 -2059 -6072
rect -1885 -6078 -1827 -6072
rect -1653 -6078 -1595 -6072
rect -1421 -6078 -1363 -6072
rect -1189 -6078 -1131 -6072
rect -957 -6078 -899 -6072
rect -725 -6078 -667 -6072
rect -493 -6078 -435 -6072
rect -261 -6078 -203 -6072
rect -29 -6078 29 -6072
rect 203 -6078 261 -6072
rect 435 -6078 493 -6072
rect 667 -6078 725 -6072
rect 899 -6078 957 -6072
rect 1131 -6078 1189 -6072
rect 1363 -6078 1421 -6072
rect 1595 -6078 1653 -6072
rect 1827 -6078 1885 -6072
rect 2059 -6078 2117 -6072
rect 2291 -6078 2349 -6072
rect 2523 -6078 2581 -6072
rect 2755 -6078 2813 -6072
rect 2987 -6078 3045 -6072
rect 3219 -6078 3277 -6072
<< nmos >>
rect -3278 -6000 -3218 6000
rect -3046 -6000 -2986 6000
rect -2814 -6000 -2754 6000
rect -2582 -6000 -2522 6000
rect -2350 -6000 -2290 6000
rect -2118 -6000 -2058 6000
rect -1886 -6000 -1826 6000
rect -1654 -6000 -1594 6000
rect -1422 -6000 -1362 6000
rect -1190 -6000 -1130 6000
rect -958 -6000 -898 6000
rect -726 -6000 -666 6000
rect -494 -6000 -434 6000
rect -262 -6000 -202 6000
rect -30 -6000 30 6000
rect 202 -6000 262 6000
rect 434 -6000 494 6000
rect 666 -6000 726 6000
rect 898 -6000 958 6000
rect 1130 -6000 1190 6000
rect 1362 -6000 1422 6000
rect 1594 -6000 1654 6000
rect 1826 -6000 1886 6000
rect 2058 -6000 2118 6000
rect 2290 -6000 2350 6000
rect 2522 -6000 2582 6000
rect 2754 -6000 2814 6000
rect 2986 -6000 3046 6000
rect 3218 -6000 3278 6000
<< ndiff >>
rect -3336 5988 -3278 6000
rect -3336 -5988 -3324 5988
rect -3290 -5988 -3278 5988
rect -3336 -6000 -3278 -5988
rect -3218 5988 -3160 6000
rect -3218 -5988 -3206 5988
rect -3172 -5988 -3160 5988
rect -3218 -6000 -3160 -5988
rect -3104 5988 -3046 6000
rect -3104 -5988 -3092 5988
rect -3058 -5988 -3046 5988
rect -3104 -6000 -3046 -5988
rect -2986 5988 -2928 6000
rect -2986 -5988 -2974 5988
rect -2940 -5988 -2928 5988
rect -2986 -6000 -2928 -5988
rect -2872 5988 -2814 6000
rect -2872 -5988 -2860 5988
rect -2826 -5988 -2814 5988
rect -2872 -6000 -2814 -5988
rect -2754 5988 -2696 6000
rect -2754 -5988 -2742 5988
rect -2708 -5988 -2696 5988
rect -2754 -6000 -2696 -5988
rect -2640 5988 -2582 6000
rect -2640 -5988 -2628 5988
rect -2594 -5988 -2582 5988
rect -2640 -6000 -2582 -5988
rect -2522 5988 -2464 6000
rect -2522 -5988 -2510 5988
rect -2476 -5988 -2464 5988
rect -2522 -6000 -2464 -5988
rect -2408 5988 -2350 6000
rect -2408 -5988 -2396 5988
rect -2362 -5988 -2350 5988
rect -2408 -6000 -2350 -5988
rect -2290 5988 -2232 6000
rect -2290 -5988 -2278 5988
rect -2244 -5988 -2232 5988
rect -2290 -6000 -2232 -5988
rect -2176 5988 -2118 6000
rect -2176 -5988 -2164 5988
rect -2130 -5988 -2118 5988
rect -2176 -6000 -2118 -5988
rect -2058 5988 -2000 6000
rect -2058 -5988 -2046 5988
rect -2012 -5988 -2000 5988
rect -2058 -6000 -2000 -5988
rect -1944 5988 -1886 6000
rect -1944 -5988 -1932 5988
rect -1898 -5988 -1886 5988
rect -1944 -6000 -1886 -5988
rect -1826 5988 -1768 6000
rect -1826 -5988 -1814 5988
rect -1780 -5988 -1768 5988
rect -1826 -6000 -1768 -5988
rect -1712 5988 -1654 6000
rect -1712 -5988 -1700 5988
rect -1666 -5988 -1654 5988
rect -1712 -6000 -1654 -5988
rect -1594 5988 -1536 6000
rect -1594 -5988 -1582 5988
rect -1548 -5988 -1536 5988
rect -1594 -6000 -1536 -5988
rect -1480 5988 -1422 6000
rect -1480 -5988 -1468 5988
rect -1434 -5988 -1422 5988
rect -1480 -6000 -1422 -5988
rect -1362 5988 -1304 6000
rect -1362 -5988 -1350 5988
rect -1316 -5988 -1304 5988
rect -1362 -6000 -1304 -5988
rect -1248 5988 -1190 6000
rect -1248 -5988 -1236 5988
rect -1202 -5988 -1190 5988
rect -1248 -6000 -1190 -5988
rect -1130 5988 -1072 6000
rect -1130 -5988 -1118 5988
rect -1084 -5988 -1072 5988
rect -1130 -6000 -1072 -5988
rect -1016 5988 -958 6000
rect -1016 -5988 -1004 5988
rect -970 -5988 -958 5988
rect -1016 -6000 -958 -5988
rect -898 5988 -840 6000
rect -898 -5988 -886 5988
rect -852 -5988 -840 5988
rect -898 -6000 -840 -5988
rect -784 5988 -726 6000
rect -784 -5988 -772 5988
rect -738 -5988 -726 5988
rect -784 -6000 -726 -5988
rect -666 5988 -608 6000
rect -666 -5988 -654 5988
rect -620 -5988 -608 5988
rect -666 -6000 -608 -5988
rect -552 5988 -494 6000
rect -552 -5988 -540 5988
rect -506 -5988 -494 5988
rect -552 -6000 -494 -5988
rect -434 5988 -376 6000
rect -434 -5988 -422 5988
rect -388 -5988 -376 5988
rect -434 -6000 -376 -5988
rect -320 5988 -262 6000
rect -320 -5988 -308 5988
rect -274 -5988 -262 5988
rect -320 -6000 -262 -5988
rect -202 5988 -144 6000
rect -202 -5988 -190 5988
rect -156 -5988 -144 5988
rect -202 -6000 -144 -5988
rect -88 5988 -30 6000
rect -88 -5988 -76 5988
rect -42 -5988 -30 5988
rect -88 -6000 -30 -5988
rect 30 5988 88 6000
rect 30 -5988 42 5988
rect 76 -5988 88 5988
rect 30 -6000 88 -5988
rect 144 5988 202 6000
rect 144 -5988 156 5988
rect 190 -5988 202 5988
rect 144 -6000 202 -5988
rect 262 5988 320 6000
rect 262 -5988 274 5988
rect 308 -5988 320 5988
rect 262 -6000 320 -5988
rect 376 5988 434 6000
rect 376 -5988 388 5988
rect 422 -5988 434 5988
rect 376 -6000 434 -5988
rect 494 5988 552 6000
rect 494 -5988 506 5988
rect 540 -5988 552 5988
rect 494 -6000 552 -5988
rect 608 5988 666 6000
rect 608 -5988 620 5988
rect 654 -5988 666 5988
rect 608 -6000 666 -5988
rect 726 5988 784 6000
rect 726 -5988 738 5988
rect 772 -5988 784 5988
rect 726 -6000 784 -5988
rect 840 5988 898 6000
rect 840 -5988 852 5988
rect 886 -5988 898 5988
rect 840 -6000 898 -5988
rect 958 5988 1016 6000
rect 958 -5988 970 5988
rect 1004 -5988 1016 5988
rect 958 -6000 1016 -5988
rect 1072 5988 1130 6000
rect 1072 -5988 1084 5988
rect 1118 -5988 1130 5988
rect 1072 -6000 1130 -5988
rect 1190 5988 1248 6000
rect 1190 -5988 1202 5988
rect 1236 -5988 1248 5988
rect 1190 -6000 1248 -5988
rect 1304 5988 1362 6000
rect 1304 -5988 1316 5988
rect 1350 -5988 1362 5988
rect 1304 -6000 1362 -5988
rect 1422 5988 1480 6000
rect 1422 -5988 1434 5988
rect 1468 -5988 1480 5988
rect 1422 -6000 1480 -5988
rect 1536 5988 1594 6000
rect 1536 -5988 1548 5988
rect 1582 -5988 1594 5988
rect 1536 -6000 1594 -5988
rect 1654 5988 1712 6000
rect 1654 -5988 1666 5988
rect 1700 -5988 1712 5988
rect 1654 -6000 1712 -5988
rect 1768 5988 1826 6000
rect 1768 -5988 1780 5988
rect 1814 -5988 1826 5988
rect 1768 -6000 1826 -5988
rect 1886 5988 1944 6000
rect 1886 -5988 1898 5988
rect 1932 -5988 1944 5988
rect 1886 -6000 1944 -5988
rect 2000 5988 2058 6000
rect 2000 -5988 2012 5988
rect 2046 -5988 2058 5988
rect 2000 -6000 2058 -5988
rect 2118 5988 2176 6000
rect 2118 -5988 2130 5988
rect 2164 -5988 2176 5988
rect 2118 -6000 2176 -5988
rect 2232 5988 2290 6000
rect 2232 -5988 2244 5988
rect 2278 -5988 2290 5988
rect 2232 -6000 2290 -5988
rect 2350 5988 2408 6000
rect 2350 -5988 2362 5988
rect 2396 -5988 2408 5988
rect 2350 -6000 2408 -5988
rect 2464 5988 2522 6000
rect 2464 -5988 2476 5988
rect 2510 -5988 2522 5988
rect 2464 -6000 2522 -5988
rect 2582 5988 2640 6000
rect 2582 -5988 2594 5988
rect 2628 -5988 2640 5988
rect 2582 -6000 2640 -5988
rect 2696 5988 2754 6000
rect 2696 -5988 2708 5988
rect 2742 -5988 2754 5988
rect 2696 -6000 2754 -5988
rect 2814 5988 2872 6000
rect 2814 -5988 2826 5988
rect 2860 -5988 2872 5988
rect 2814 -6000 2872 -5988
rect 2928 5988 2986 6000
rect 2928 -5988 2940 5988
rect 2974 -5988 2986 5988
rect 2928 -6000 2986 -5988
rect 3046 5988 3104 6000
rect 3046 -5988 3058 5988
rect 3092 -5988 3104 5988
rect 3046 -6000 3104 -5988
rect 3160 5988 3218 6000
rect 3160 -5988 3172 5988
rect 3206 -5988 3218 5988
rect 3160 -6000 3218 -5988
rect 3278 5988 3336 6000
rect 3278 -5988 3290 5988
rect 3324 -5988 3336 5988
rect 3278 -6000 3336 -5988
<< ndiffc >>
rect -3324 -5988 -3290 5988
rect -3206 -5988 -3172 5988
rect -3092 -5988 -3058 5988
rect -2974 -5988 -2940 5988
rect -2860 -5988 -2826 5988
rect -2742 -5988 -2708 5988
rect -2628 -5988 -2594 5988
rect -2510 -5988 -2476 5988
rect -2396 -5988 -2362 5988
rect -2278 -5988 -2244 5988
rect -2164 -5988 -2130 5988
rect -2046 -5988 -2012 5988
rect -1932 -5988 -1898 5988
rect -1814 -5988 -1780 5988
rect -1700 -5988 -1666 5988
rect -1582 -5988 -1548 5988
rect -1468 -5988 -1434 5988
rect -1350 -5988 -1316 5988
rect -1236 -5988 -1202 5988
rect -1118 -5988 -1084 5988
rect -1004 -5988 -970 5988
rect -886 -5988 -852 5988
rect -772 -5988 -738 5988
rect -654 -5988 -620 5988
rect -540 -5988 -506 5988
rect -422 -5988 -388 5988
rect -308 -5988 -274 5988
rect -190 -5988 -156 5988
rect -76 -5988 -42 5988
rect 42 -5988 76 5988
rect 156 -5988 190 5988
rect 274 -5988 308 5988
rect 388 -5988 422 5988
rect 506 -5988 540 5988
rect 620 -5988 654 5988
rect 738 -5988 772 5988
rect 852 -5988 886 5988
rect 970 -5988 1004 5988
rect 1084 -5988 1118 5988
rect 1202 -5988 1236 5988
rect 1316 -5988 1350 5988
rect 1434 -5988 1468 5988
rect 1548 -5988 1582 5988
rect 1666 -5988 1700 5988
rect 1780 -5988 1814 5988
rect 1898 -5988 1932 5988
rect 2012 -5988 2046 5988
rect 2130 -5988 2164 5988
rect 2244 -5988 2278 5988
rect 2362 -5988 2396 5988
rect 2476 -5988 2510 5988
rect 2594 -5988 2628 5988
rect 2708 -5988 2742 5988
rect 2826 -5988 2860 5988
rect 2940 -5988 2974 5988
rect 3058 -5988 3092 5988
rect 3172 -5988 3206 5988
rect 3290 -5988 3324 5988
<< poly >>
rect -3281 6072 -3215 6088
rect -3281 6038 -3265 6072
rect -3231 6038 -3215 6072
rect -3281 6022 -3215 6038
rect -3049 6072 -2983 6088
rect -3049 6038 -3033 6072
rect -2999 6038 -2983 6072
rect -3049 6022 -2983 6038
rect -2817 6072 -2751 6088
rect -2817 6038 -2801 6072
rect -2767 6038 -2751 6072
rect -2817 6022 -2751 6038
rect -2585 6072 -2519 6088
rect -2585 6038 -2569 6072
rect -2535 6038 -2519 6072
rect -2585 6022 -2519 6038
rect -2353 6072 -2287 6088
rect -2353 6038 -2337 6072
rect -2303 6038 -2287 6072
rect -2353 6022 -2287 6038
rect -2121 6072 -2055 6088
rect -2121 6038 -2105 6072
rect -2071 6038 -2055 6072
rect -2121 6022 -2055 6038
rect -1889 6072 -1823 6088
rect -1889 6038 -1873 6072
rect -1839 6038 -1823 6072
rect -1889 6022 -1823 6038
rect -1657 6072 -1591 6088
rect -1657 6038 -1641 6072
rect -1607 6038 -1591 6072
rect -1657 6022 -1591 6038
rect -1425 6072 -1359 6088
rect -1425 6038 -1409 6072
rect -1375 6038 -1359 6072
rect -1425 6022 -1359 6038
rect -1193 6072 -1127 6088
rect -1193 6038 -1177 6072
rect -1143 6038 -1127 6072
rect -1193 6022 -1127 6038
rect -961 6072 -895 6088
rect -961 6038 -945 6072
rect -911 6038 -895 6072
rect -961 6022 -895 6038
rect -729 6072 -663 6088
rect -729 6038 -713 6072
rect -679 6038 -663 6072
rect -729 6022 -663 6038
rect -497 6072 -431 6088
rect -497 6038 -481 6072
rect -447 6038 -431 6072
rect -497 6022 -431 6038
rect -265 6072 -199 6088
rect -265 6038 -249 6072
rect -215 6038 -199 6072
rect -265 6022 -199 6038
rect -33 6072 33 6088
rect -33 6038 -17 6072
rect 17 6038 33 6072
rect -33 6022 33 6038
rect 199 6072 265 6088
rect 199 6038 215 6072
rect 249 6038 265 6072
rect 199 6022 265 6038
rect 431 6072 497 6088
rect 431 6038 447 6072
rect 481 6038 497 6072
rect 431 6022 497 6038
rect 663 6072 729 6088
rect 663 6038 679 6072
rect 713 6038 729 6072
rect 663 6022 729 6038
rect 895 6072 961 6088
rect 895 6038 911 6072
rect 945 6038 961 6072
rect 895 6022 961 6038
rect 1127 6072 1193 6088
rect 1127 6038 1143 6072
rect 1177 6038 1193 6072
rect 1127 6022 1193 6038
rect 1359 6072 1425 6088
rect 1359 6038 1375 6072
rect 1409 6038 1425 6072
rect 1359 6022 1425 6038
rect 1591 6072 1657 6088
rect 1591 6038 1607 6072
rect 1641 6038 1657 6072
rect 1591 6022 1657 6038
rect 1823 6072 1889 6088
rect 1823 6038 1839 6072
rect 1873 6038 1889 6072
rect 1823 6022 1889 6038
rect 2055 6072 2121 6088
rect 2055 6038 2071 6072
rect 2105 6038 2121 6072
rect 2055 6022 2121 6038
rect 2287 6072 2353 6088
rect 2287 6038 2303 6072
rect 2337 6038 2353 6072
rect 2287 6022 2353 6038
rect 2519 6072 2585 6088
rect 2519 6038 2535 6072
rect 2569 6038 2585 6072
rect 2519 6022 2585 6038
rect 2751 6072 2817 6088
rect 2751 6038 2767 6072
rect 2801 6038 2817 6072
rect 2751 6022 2817 6038
rect 2983 6072 3049 6088
rect 2983 6038 2999 6072
rect 3033 6038 3049 6072
rect 2983 6022 3049 6038
rect 3215 6072 3281 6088
rect 3215 6038 3231 6072
rect 3265 6038 3281 6072
rect 3215 6022 3281 6038
rect -3278 6000 -3218 6022
rect -3046 6000 -2986 6022
rect -2814 6000 -2754 6022
rect -2582 6000 -2522 6022
rect -2350 6000 -2290 6022
rect -2118 6000 -2058 6022
rect -1886 6000 -1826 6022
rect -1654 6000 -1594 6022
rect -1422 6000 -1362 6022
rect -1190 6000 -1130 6022
rect -958 6000 -898 6022
rect -726 6000 -666 6022
rect -494 6000 -434 6022
rect -262 6000 -202 6022
rect -30 6000 30 6022
rect 202 6000 262 6022
rect 434 6000 494 6022
rect 666 6000 726 6022
rect 898 6000 958 6022
rect 1130 6000 1190 6022
rect 1362 6000 1422 6022
rect 1594 6000 1654 6022
rect 1826 6000 1886 6022
rect 2058 6000 2118 6022
rect 2290 6000 2350 6022
rect 2522 6000 2582 6022
rect 2754 6000 2814 6022
rect 2986 6000 3046 6022
rect 3218 6000 3278 6022
rect -3278 -6022 -3218 -6000
rect -3046 -6022 -2986 -6000
rect -2814 -6022 -2754 -6000
rect -2582 -6022 -2522 -6000
rect -2350 -6022 -2290 -6000
rect -2118 -6022 -2058 -6000
rect -1886 -6022 -1826 -6000
rect -1654 -6022 -1594 -6000
rect -1422 -6022 -1362 -6000
rect -1190 -6022 -1130 -6000
rect -958 -6022 -898 -6000
rect -726 -6022 -666 -6000
rect -494 -6022 -434 -6000
rect -262 -6022 -202 -6000
rect -30 -6022 30 -6000
rect 202 -6022 262 -6000
rect 434 -6022 494 -6000
rect 666 -6022 726 -6000
rect 898 -6022 958 -6000
rect 1130 -6022 1190 -6000
rect 1362 -6022 1422 -6000
rect 1594 -6022 1654 -6000
rect 1826 -6022 1886 -6000
rect 2058 -6022 2118 -6000
rect 2290 -6022 2350 -6000
rect 2522 -6022 2582 -6000
rect 2754 -6022 2814 -6000
rect 2986 -6022 3046 -6000
rect 3218 -6022 3278 -6000
rect -3281 -6038 -3215 -6022
rect -3281 -6072 -3265 -6038
rect -3231 -6072 -3215 -6038
rect -3281 -6088 -3215 -6072
rect -3049 -6038 -2983 -6022
rect -3049 -6072 -3033 -6038
rect -2999 -6072 -2983 -6038
rect -3049 -6088 -2983 -6072
rect -2817 -6038 -2751 -6022
rect -2817 -6072 -2801 -6038
rect -2767 -6072 -2751 -6038
rect -2817 -6088 -2751 -6072
rect -2585 -6038 -2519 -6022
rect -2585 -6072 -2569 -6038
rect -2535 -6072 -2519 -6038
rect -2585 -6088 -2519 -6072
rect -2353 -6038 -2287 -6022
rect -2353 -6072 -2337 -6038
rect -2303 -6072 -2287 -6038
rect -2353 -6088 -2287 -6072
rect -2121 -6038 -2055 -6022
rect -2121 -6072 -2105 -6038
rect -2071 -6072 -2055 -6038
rect -2121 -6088 -2055 -6072
rect -1889 -6038 -1823 -6022
rect -1889 -6072 -1873 -6038
rect -1839 -6072 -1823 -6038
rect -1889 -6088 -1823 -6072
rect -1657 -6038 -1591 -6022
rect -1657 -6072 -1641 -6038
rect -1607 -6072 -1591 -6038
rect -1657 -6088 -1591 -6072
rect -1425 -6038 -1359 -6022
rect -1425 -6072 -1409 -6038
rect -1375 -6072 -1359 -6038
rect -1425 -6088 -1359 -6072
rect -1193 -6038 -1127 -6022
rect -1193 -6072 -1177 -6038
rect -1143 -6072 -1127 -6038
rect -1193 -6088 -1127 -6072
rect -961 -6038 -895 -6022
rect -961 -6072 -945 -6038
rect -911 -6072 -895 -6038
rect -961 -6088 -895 -6072
rect -729 -6038 -663 -6022
rect -729 -6072 -713 -6038
rect -679 -6072 -663 -6038
rect -729 -6088 -663 -6072
rect -497 -6038 -431 -6022
rect -497 -6072 -481 -6038
rect -447 -6072 -431 -6038
rect -497 -6088 -431 -6072
rect -265 -6038 -199 -6022
rect -265 -6072 -249 -6038
rect -215 -6072 -199 -6038
rect -265 -6088 -199 -6072
rect -33 -6038 33 -6022
rect -33 -6072 -17 -6038
rect 17 -6072 33 -6038
rect -33 -6088 33 -6072
rect 199 -6038 265 -6022
rect 199 -6072 215 -6038
rect 249 -6072 265 -6038
rect 199 -6088 265 -6072
rect 431 -6038 497 -6022
rect 431 -6072 447 -6038
rect 481 -6072 497 -6038
rect 431 -6088 497 -6072
rect 663 -6038 729 -6022
rect 663 -6072 679 -6038
rect 713 -6072 729 -6038
rect 663 -6088 729 -6072
rect 895 -6038 961 -6022
rect 895 -6072 911 -6038
rect 945 -6072 961 -6038
rect 895 -6088 961 -6072
rect 1127 -6038 1193 -6022
rect 1127 -6072 1143 -6038
rect 1177 -6072 1193 -6038
rect 1127 -6088 1193 -6072
rect 1359 -6038 1425 -6022
rect 1359 -6072 1375 -6038
rect 1409 -6072 1425 -6038
rect 1359 -6088 1425 -6072
rect 1591 -6038 1657 -6022
rect 1591 -6072 1607 -6038
rect 1641 -6072 1657 -6038
rect 1591 -6088 1657 -6072
rect 1823 -6038 1889 -6022
rect 1823 -6072 1839 -6038
rect 1873 -6072 1889 -6038
rect 1823 -6088 1889 -6072
rect 2055 -6038 2121 -6022
rect 2055 -6072 2071 -6038
rect 2105 -6072 2121 -6038
rect 2055 -6088 2121 -6072
rect 2287 -6038 2353 -6022
rect 2287 -6072 2303 -6038
rect 2337 -6072 2353 -6038
rect 2287 -6088 2353 -6072
rect 2519 -6038 2585 -6022
rect 2519 -6072 2535 -6038
rect 2569 -6072 2585 -6038
rect 2519 -6088 2585 -6072
rect 2751 -6038 2817 -6022
rect 2751 -6072 2767 -6038
rect 2801 -6072 2817 -6038
rect 2751 -6088 2817 -6072
rect 2983 -6038 3049 -6022
rect 2983 -6072 2999 -6038
rect 3033 -6072 3049 -6038
rect 2983 -6088 3049 -6072
rect 3215 -6038 3281 -6022
rect 3215 -6072 3231 -6038
rect 3265 -6072 3281 -6038
rect 3215 -6088 3281 -6072
<< polycont >>
rect -3265 6038 -3231 6072
rect -3033 6038 -2999 6072
rect -2801 6038 -2767 6072
rect -2569 6038 -2535 6072
rect -2337 6038 -2303 6072
rect -2105 6038 -2071 6072
rect -1873 6038 -1839 6072
rect -1641 6038 -1607 6072
rect -1409 6038 -1375 6072
rect -1177 6038 -1143 6072
rect -945 6038 -911 6072
rect -713 6038 -679 6072
rect -481 6038 -447 6072
rect -249 6038 -215 6072
rect -17 6038 17 6072
rect 215 6038 249 6072
rect 447 6038 481 6072
rect 679 6038 713 6072
rect 911 6038 945 6072
rect 1143 6038 1177 6072
rect 1375 6038 1409 6072
rect 1607 6038 1641 6072
rect 1839 6038 1873 6072
rect 2071 6038 2105 6072
rect 2303 6038 2337 6072
rect 2535 6038 2569 6072
rect 2767 6038 2801 6072
rect 2999 6038 3033 6072
rect 3231 6038 3265 6072
rect -3265 -6072 -3231 -6038
rect -3033 -6072 -2999 -6038
rect -2801 -6072 -2767 -6038
rect -2569 -6072 -2535 -6038
rect -2337 -6072 -2303 -6038
rect -2105 -6072 -2071 -6038
rect -1873 -6072 -1839 -6038
rect -1641 -6072 -1607 -6038
rect -1409 -6072 -1375 -6038
rect -1177 -6072 -1143 -6038
rect -945 -6072 -911 -6038
rect -713 -6072 -679 -6038
rect -481 -6072 -447 -6038
rect -249 -6072 -215 -6038
rect -17 -6072 17 -6038
rect 215 -6072 249 -6038
rect 447 -6072 481 -6038
rect 679 -6072 713 -6038
rect 911 -6072 945 -6038
rect 1143 -6072 1177 -6038
rect 1375 -6072 1409 -6038
rect 1607 -6072 1641 -6038
rect 1839 -6072 1873 -6038
rect 2071 -6072 2105 -6038
rect 2303 -6072 2337 -6038
rect 2535 -6072 2569 -6038
rect 2767 -6072 2801 -6038
rect 2999 -6072 3033 -6038
rect 3231 -6072 3265 -6038
<< locali >>
rect -3281 6038 -3265 6072
rect -3231 6038 -3215 6072
rect -3049 6038 -3033 6072
rect -2999 6038 -2983 6072
rect -2817 6038 -2801 6072
rect -2767 6038 -2751 6072
rect -2585 6038 -2569 6072
rect -2535 6038 -2519 6072
rect -2353 6038 -2337 6072
rect -2303 6038 -2287 6072
rect -2121 6038 -2105 6072
rect -2071 6038 -2055 6072
rect -1889 6038 -1873 6072
rect -1839 6038 -1823 6072
rect -1657 6038 -1641 6072
rect -1607 6038 -1591 6072
rect -1425 6038 -1409 6072
rect -1375 6038 -1359 6072
rect -1193 6038 -1177 6072
rect -1143 6038 -1127 6072
rect -961 6038 -945 6072
rect -911 6038 -895 6072
rect -729 6038 -713 6072
rect -679 6038 -663 6072
rect -497 6038 -481 6072
rect -447 6038 -431 6072
rect -265 6038 -249 6072
rect -215 6038 -199 6072
rect -33 6038 -17 6072
rect 17 6038 33 6072
rect 199 6038 215 6072
rect 249 6038 265 6072
rect 431 6038 447 6072
rect 481 6038 497 6072
rect 663 6038 679 6072
rect 713 6038 729 6072
rect 895 6038 911 6072
rect 945 6038 961 6072
rect 1127 6038 1143 6072
rect 1177 6038 1193 6072
rect 1359 6038 1375 6072
rect 1409 6038 1425 6072
rect 1591 6038 1607 6072
rect 1641 6038 1657 6072
rect 1823 6038 1839 6072
rect 1873 6038 1889 6072
rect 2055 6038 2071 6072
rect 2105 6038 2121 6072
rect 2287 6038 2303 6072
rect 2337 6038 2353 6072
rect 2519 6038 2535 6072
rect 2569 6038 2585 6072
rect 2751 6038 2767 6072
rect 2801 6038 2817 6072
rect 2983 6038 2999 6072
rect 3033 6038 3049 6072
rect 3215 6038 3231 6072
rect 3265 6038 3281 6072
rect -3324 5988 -3290 6004
rect -3324 -6004 -3290 -5988
rect -3206 5988 -3172 6004
rect -3206 -6004 -3172 -5988
rect -3092 5988 -3058 6004
rect -3092 -6004 -3058 -5988
rect -2974 5988 -2940 6004
rect -2974 -6004 -2940 -5988
rect -2860 5988 -2826 6004
rect -2860 -6004 -2826 -5988
rect -2742 5988 -2708 6004
rect -2742 -6004 -2708 -5988
rect -2628 5988 -2594 6004
rect -2628 -6004 -2594 -5988
rect -2510 5988 -2476 6004
rect -2510 -6004 -2476 -5988
rect -2396 5988 -2362 6004
rect -2396 -6004 -2362 -5988
rect -2278 5988 -2244 6004
rect -2278 -6004 -2244 -5988
rect -2164 5988 -2130 6004
rect -2164 -6004 -2130 -5988
rect -2046 5988 -2012 6004
rect -2046 -6004 -2012 -5988
rect -1932 5988 -1898 6004
rect -1932 -6004 -1898 -5988
rect -1814 5988 -1780 6004
rect -1814 -6004 -1780 -5988
rect -1700 5988 -1666 6004
rect -1700 -6004 -1666 -5988
rect -1582 5988 -1548 6004
rect -1582 -6004 -1548 -5988
rect -1468 5988 -1434 6004
rect -1468 -6004 -1434 -5988
rect -1350 5988 -1316 6004
rect -1350 -6004 -1316 -5988
rect -1236 5988 -1202 6004
rect -1236 -6004 -1202 -5988
rect -1118 5988 -1084 6004
rect -1118 -6004 -1084 -5988
rect -1004 5988 -970 6004
rect -1004 -6004 -970 -5988
rect -886 5988 -852 6004
rect -886 -6004 -852 -5988
rect -772 5988 -738 6004
rect -772 -6004 -738 -5988
rect -654 5988 -620 6004
rect -654 -6004 -620 -5988
rect -540 5988 -506 6004
rect -540 -6004 -506 -5988
rect -422 5988 -388 6004
rect -422 -6004 -388 -5988
rect -308 5988 -274 6004
rect -308 -6004 -274 -5988
rect -190 5988 -156 6004
rect -190 -6004 -156 -5988
rect -76 5988 -42 6004
rect -76 -6004 -42 -5988
rect 42 5988 76 6004
rect 42 -6004 76 -5988
rect 156 5988 190 6004
rect 156 -6004 190 -5988
rect 274 5988 308 6004
rect 274 -6004 308 -5988
rect 388 5988 422 6004
rect 388 -6004 422 -5988
rect 506 5988 540 6004
rect 506 -6004 540 -5988
rect 620 5988 654 6004
rect 620 -6004 654 -5988
rect 738 5988 772 6004
rect 738 -6004 772 -5988
rect 852 5988 886 6004
rect 852 -6004 886 -5988
rect 970 5988 1004 6004
rect 970 -6004 1004 -5988
rect 1084 5988 1118 6004
rect 1084 -6004 1118 -5988
rect 1202 5988 1236 6004
rect 1202 -6004 1236 -5988
rect 1316 5988 1350 6004
rect 1316 -6004 1350 -5988
rect 1434 5988 1468 6004
rect 1434 -6004 1468 -5988
rect 1548 5988 1582 6004
rect 1548 -6004 1582 -5988
rect 1666 5988 1700 6004
rect 1666 -6004 1700 -5988
rect 1780 5988 1814 6004
rect 1780 -6004 1814 -5988
rect 1898 5988 1932 6004
rect 1898 -6004 1932 -5988
rect 2012 5988 2046 6004
rect 2012 -6004 2046 -5988
rect 2130 5988 2164 6004
rect 2130 -6004 2164 -5988
rect 2244 5988 2278 6004
rect 2244 -6004 2278 -5988
rect 2362 5988 2396 6004
rect 2362 -6004 2396 -5988
rect 2476 5988 2510 6004
rect 2476 -6004 2510 -5988
rect 2594 5988 2628 6004
rect 2594 -6004 2628 -5988
rect 2708 5988 2742 6004
rect 2708 -6004 2742 -5988
rect 2826 5988 2860 6004
rect 2826 -6004 2860 -5988
rect 2940 5988 2974 6004
rect 2940 -6004 2974 -5988
rect 3058 5988 3092 6004
rect 3058 -6004 3092 -5988
rect 3172 5988 3206 6004
rect 3172 -6004 3206 -5988
rect 3290 5988 3324 6004
rect 3290 -6004 3324 -5988
rect -3281 -6072 -3265 -6038
rect -3231 -6072 -3215 -6038
rect -3049 -6072 -3033 -6038
rect -2999 -6072 -2983 -6038
rect -2817 -6072 -2801 -6038
rect -2767 -6072 -2751 -6038
rect -2585 -6072 -2569 -6038
rect -2535 -6072 -2519 -6038
rect -2353 -6072 -2337 -6038
rect -2303 -6072 -2287 -6038
rect -2121 -6072 -2105 -6038
rect -2071 -6072 -2055 -6038
rect -1889 -6072 -1873 -6038
rect -1839 -6072 -1823 -6038
rect -1657 -6072 -1641 -6038
rect -1607 -6072 -1591 -6038
rect -1425 -6072 -1409 -6038
rect -1375 -6072 -1359 -6038
rect -1193 -6072 -1177 -6038
rect -1143 -6072 -1127 -6038
rect -961 -6072 -945 -6038
rect -911 -6072 -895 -6038
rect -729 -6072 -713 -6038
rect -679 -6072 -663 -6038
rect -497 -6072 -481 -6038
rect -447 -6072 -431 -6038
rect -265 -6072 -249 -6038
rect -215 -6072 -199 -6038
rect -33 -6072 -17 -6038
rect 17 -6072 33 -6038
rect 199 -6072 215 -6038
rect 249 -6072 265 -6038
rect 431 -6072 447 -6038
rect 481 -6072 497 -6038
rect 663 -6072 679 -6038
rect 713 -6072 729 -6038
rect 895 -6072 911 -6038
rect 945 -6072 961 -6038
rect 1127 -6072 1143 -6038
rect 1177 -6072 1193 -6038
rect 1359 -6072 1375 -6038
rect 1409 -6072 1425 -6038
rect 1591 -6072 1607 -6038
rect 1641 -6072 1657 -6038
rect 1823 -6072 1839 -6038
rect 1873 -6072 1889 -6038
rect 2055 -6072 2071 -6038
rect 2105 -6072 2121 -6038
rect 2287 -6072 2303 -6038
rect 2337 -6072 2353 -6038
rect 2519 -6072 2535 -6038
rect 2569 -6072 2585 -6038
rect 2751 -6072 2767 -6038
rect 2801 -6072 2817 -6038
rect 2983 -6072 2999 -6038
rect 3033 -6072 3049 -6038
rect 3215 -6072 3231 -6038
rect 3265 -6072 3281 -6038
<< viali >>
rect -3265 6038 -3231 6072
rect -3033 6038 -2999 6072
rect -2801 6038 -2767 6072
rect -2569 6038 -2535 6072
rect -2337 6038 -2303 6072
rect -2105 6038 -2071 6072
rect -1873 6038 -1839 6072
rect -1641 6038 -1607 6072
rect -1409 6038 -1375 6072
rect -1177 6038 -1143 6072
rect -945 6038 -911 6072
rect -713 6038 -679 6072
rect -481 6038 -447 6072
rect -249 6038 -215 6072
rect -17 6038 17 6072
rect 215 6038 249 6072
rect 447 6038 481 6072
rect 679 6038 713 6072
rect 911 6038 945 6072
rect 1143 6038 1177 6072
rect 1375 6038 1409 6072
rect 1607 6038 1641 6072
rect 1839 6038 1873 6072
rect 2071 6038 2105 6072
rect 2303 6038 2337 6072
rect 2535 6038 2569 6072
rect 2767 6038 2801 6072
rect 2999 6038 3033 6072
rect 3231 6038 3265 6072
rect -3324 -5988 -3290 5988
rect -3206 -5988 -3172 5988
rect -3092 -5988 -3058 5988
rect -2974 -5988 -2940 5988
rect -2860 -5988 -2826 5988
rect -2742 -5988 -2708 5988
rect -2628 -5988 -2594 5988
rect -2510 -5988 -2476 5988
rect -2396 -5988 -2362 5988
rect -2278 -5988 -2244 5988
rect -2164 -5988 -2130 5988
rect -2046 -5988 -2012 5988
rect -1932 -5988 -1898 5988
rect -1814 -5988 -1780 5988
rect -1700 -5988 -1666 5988
rect -1582 -5988 -1548 5988
rect -1468 -5988 -1434 5988
rect -1350 -5988 -1316 5988
rect -1236 -5988 -1202 5988
rect -1118 -5988 -1084 5988
rect -1004 -5988 -970 5988
rect -886 -5988 -852 5988
rect -772 -5988 -738 5988
rect -654 -5988 -620 5988
rect -540 -5988 -506 5988
rect -422 -5988 -388 5988
rect -308 -5988 -274 5988
rect -190 -5988 -156 5988
rect -76 -5988 -42 5988
rect 42 -5988 76 5988
rect 156 -5988 190 5988
rect 274 -5988 308 5988
rect 388 -5988 422 5988
rect 506 -5988 540 5988
rect 620 -5988 654 5988
rect 738 -5988 772 5988
rect 852 -5988 886 5988
rect 970 -5988 1004 5988
rect 1084 -5988 1118 5988
rect 1202 -5988 1236 5988
rect 1316 -5988 1350 5988
rect 1434 -5988 1468 5988
rect 1548 -5988 1582 5988
rect 1666 -5988 1700 5988
rect 1780 -5988 1814 5988
rect 1898 -5988 1932 5988
rect 2012 -5988 2046 5988
rect 2130 -5988 2164 5988
rect 2244 -5988 2278 5988
rect 2362 -5988 2396 5988
rect 2476 -5988 2510 5988
rect 2594 -5988 2628 5988
rect 2708 -5988 2742 5988
rect 2826 -5988 2860 5988
rect 2940 -5988 2974 5988
rect 3058 -5988 3092 5988
rect 3172 -5988 3206 5988
rect 3290 -5988 3324 5988
rect -3265 -6072 -3231 -6038
rect -3033 -6072 -2999 -6038
rect -2801 -6072 -2767 -6038
rect -2569 -6072 -2535 -6038
rect -2337 -6072 -2303 -6038
rect -2105 -6072 -2071 -6038
rect -1873 -6072 -1839 -6038
rect -1641 -6072 -1607 -6038
rect -1409 -6072 -1375 -6038
rect -1177 -6072 -1143 -6038
rect -945 -6072 -911 -6038
rect -713 -6072 -679 -6038
rect -481 -6072 -447 -6038
rect -249 -6072 -215 -6038
rect -17 -6072 17 -6038
rect 215 -6072 249 -6038
rect 447 -6072 481 -6038
rect 679 -6072 713 -6038
rect 911 -6072 945 -6038
rect 1143 -6072 1177 -6038
rect 1375 -6072 1409 -6038
rect 1607 -6072 1641 -6038
rect 1839 -6072 1873 -6038
rect 2071 -6072 2105 -6038
rect 2303 -6072 2337 -6038
rect 2535 -6072 2569 -6038
rect 2767 -6072 2801 -6038
rect 2999 -6072 3033 -6038
rect 3231 -6072 3265 -6038
<< metal1 >>
rect -3277 6072 -3219 6078
rect -3277 6038 -3265 6072
rect -3231 6038 -3219 6072
rect -3277 6032 -3219 6038
rect -3045 6072 -2987 6078
rect -3045 6038 -3033 6072
rect -2999 6038 -2987 6072
rect -3045 6032 -2987 6038
rect -2813 6072 -2755 6078
rect -2813 6038 -2801 6072
rect -2767 6038 -2755 6072
rect -2813 6032 -2755 6038
rect -2581 6072 -2523 6078
rect -2581 6038 -2569 6072
rect -2535 6038 -2523 6072
rect -2581 6032 -2523 6038
rect -2349 6072 -2291 6078
rect -2349 6038 -2337 6072
rect -2303 6038 -2291 6072
rect -2349 6032 -2291 6038
rect -2117 6072 -2059 6078
rect -2117 6038 -2105 6072
rect -2071 6038 -2059 6072
rect -2117 6032 -2059 6038
rect -1885 6072 -1827 6078
rect -1885 6038 -1873 6072
rect -1839 6038 -1827 6072
rect -1885 6032 -1827 6038
rect -1653 6072 -1595 6078
rect -1653 6038 -1641 6072
rect -1607 6038 -1595 6072
rect -1653 6032 -1595 6038
rect -1421 6072 -1363 6078
rect -1421 6038 -1409 6072
rect -1375 6038 -1363 6072
rect -1421 6032 -1363 6038
rect -1189 6072 -1131 6078
rect -1189 6038 -1177 6072
rect -1143 6038 -1131 6072
rect -1189 6032 -1131 6038
rect -957 6072 -899 6078
rect -957 6038 -945 6072
rect -911 6038 -899 6072
rect -957 6032 -899 6038
rect -725 6072 -667 6078
rect -725 6038 -713 6072
rect -679 6038 -667 6072
rect -725 6032 -667 6038
rect -493 6072 -435 6078
rect -493 6038 -481 6072
rect -447 6038 -435 6072
rect -493 6032 -435 6038
rect -261 6072 -203 6078
rect -261 6038 -249 6072
rect -215 6038 -203 6072
rect -261 6032 -203 6038
rect -29 6072 29 6078
rect -29 6038 -17 6072
rect 17 6038 29 6072
rect -29 6032 29 6038
rect 203 6072 261 6078
rect 203 6038 215 6072
rect 249 6038 261 6072
rect 203 6032 261 6038
rect 435 6072 493 6078
rect 435 6038 447 6072
rect 481 6038 493 6072
rect 435 6032 493 6038
rect 667 6072 725 6078
rect 667 6038 679 6072
rect 713 6038 725 6072
rect 667 6032 725 6038
rect 899 6072 957 6078
rect 899 6038 911 6072
rect 945 6038 957 6072
rect 899 6032 957 6038
rect 1131 6072 1189 6078
rect 1131 6038 1143 6072
rect 1177 6038 1189 6072
rect 1131 6032 1189 6038
rect 1363 6072 1421 6078
rect 1363 6038 1375 6072
rect 1409 6038 1421 6072
rect 1363 6032 1421 6038
rect 1595 6072 1653 6078
rect 1595 6038 1607 6072
rect 1641 6038 1653 6072
rect 1595 6032 1653 6038
rect 1827 6072 1885 6078
rect 1827 6038 1839 6072
rect 1873 6038 1885 6072
rect 1827 6032 1885 6038
rect 2059 6072 2117 6078
rect 2059 6038 2071 6072
rect 2105 6038 2117 6072
rect 2059 6032 2117 6038
rect 2291 6072 2349 6078
rect 2291 6038 2303 6072
rect 2337 6038 2349 6072
rect 2291 6032 2349 6038
rect 2523 6072 2581 6078
rect 2523 6038 2535 6072
rect 2569 6038 2581 6072
rect 2523 6032 2581 6038
rect 2755 6072 2813 6078
rect 2755 6038 2767 6072
rect 2801 6038 2813 6072
rect 2755 6032 2813 6038
rect 2987 6072 3045 6078
rect 2987 6038 2999 6072
rect 3033 6038 3045 6072
rect 2987 6032 3045 6038
rect 3219 6072 3277 6078
rect 3219 6038 3231 6072
rect 3265 6038 3277 6072
rect 3219 6032 3277 6038
rect -3330 5988 -3284 6000
rect -3330 -5988 -3324 5988
rect -3290 -5988 -3284 5988
rect -3330 -6000 -3284 -5988
rect -3212 5988 -3166 6000
rect -3212 -5988 -3206 5988
rect -3172 -5988 -3166 5988
rect -3212 -6000 -3166 -5988
rect -3098 5988 -3052 6000
rect -3098 -5988 -3092 5988
rect -3058 -5988 -3052 5988
rect -3098 -6000 -3052 -5988
rect -2980 5988 -2934 6000
rect -2980 -5988 -2974 5988
rect -2940 -5988 -2934 5988
rect -2980 -6000 -2934 -5988
rect -2866 5988 -2820 6000
rect -2866 -5988 -2860 5988
rect -2826 -5988 -2820 5988
rect -2866 -6000 -2820 -5988
rect -2748 5988 -2702 6000
rect -2748 -5988 -2742 5988
rect -2708 -5988 -2702 5988
rect -2748 -6000 -2702 -5988
rect -2634 5988 -2588 6000
rect -2634 -5988 -2628 5988
rect -2594 -5988 -2588 5988
rect -2634 -6000 -2588 -5988
rect -2516 5988 -2470 6000
rect -2516 -5988 -2510 5988
rect -2476 -5988 -2470 5988
rect -2516 -6000 -2470 -5988
rect -2402 5988 -2356 6000
rect -2402 -5988 -2396 5988
rect -2362 -5988 -2356 5988
rect -2402 -6000 -2356 -5988
rect -2284 5988 -2238 6000
rect -2284 -5988 -2278 5988
rect -2244 -5988 -2238 5988
rect -2284 -6000 -2238 -5988
rect -2170 5988 -2124 6000
rect -2170 -5988 -2164 5988
rect -2130 -5988 -2124 5988
rect -2170 -6000 -2124 -5988
rect -2052 5988 -2006 6000
rect -2052 -5988 -2046 5988
rect -2012 -5988 -2006 5988
rect -2052 -6000 -2006 -5988
rect -1938 5988 -1892 6000
rect -1938 -5988 -1932 5988
rect -1898 -5988 -1892 5988
rect -1938 -6000 -1892 -5988
rect -1820 5988 -1774 6000
rect -1820 -5988 -1814 5988
rect -1780 -5988 -1774 5988
rect -1820 -6000 -1774 -5988
rect -1706 5988 -1660 6000
rect -1706 -5988 -1700 5988
rect -1666 -5988 -1660 5988
rect -1706 -6000 -1660 -5988
rect -1588 5988 -1542 6000
rect -1588 -5988 -1582 5988
rect -1548 -5988 -1542 5988
rect -1588 -6000 -1542 -5988
rect -1474 5988 -1428 6000
rect -1474 -5988 -1468 5988
rect -1434 -5988 -1428 5988
rect -1474 -6000 -1428 -5988
rect -1356 5988 -1310 6000
rect -1356 -5988 -1350 5988
rect -1316 -5988 -1310 5988
rect -1356 -6000 -1310 -5988
rect -1242 5988 -1196 6000
rect -1242 -5988 -1236 5988
rect -1202 -5988 -1196 5988
rect -1242 -6000 -1196 -5988
rect -1124 5988 -1078 6000
rect -1124 -5988 -1118 5988
rect -1084 -5988 -1078 5988
rect -1124 -6000 -1078 -5988
rect -1010 5988 -964 6000
rect -1010 -5988 -1004 5988
rect -970 -5988 -964 5988
rect -1010 -6000 -964 -5988
rect -892 5988 -846 6000
rect -892 -5988 -886 5988
rect -852 -5988 -846 5988
rect -892 -6000 -846 -5988
rect -778 5988 -732 6000
rect -778 -5988 -772 5988
rect -738 -5988 -732 5988
rect -778 -6000 -732 -5988
rect -660 5988 -614 6000
rect -660 -5988 -654 5988
rect -620 -5988 -614 5988
rect -660 -6000 -614 -5988
rect -546 5988 -500 6000
rect -546 -5988 -540 5988
rect -506 -5988 -500 5988
rect -546 -6000 -500 -5988
rect -428 5988 -382 6000
rect -428 -5988 -422 5988
rect -388 -5988 -382 5988
rect -428 -6000 -382 -5988
rect -314 5988 -268 6000
rect -314 -5988 -308 5988
rect -274 -5988 -268 5988
rect -314 -6000 -268 -5988
rect -196 5988 -150 6000
rect -196 -5988 -190 5988
rect -156 -5988 -150 5988
rect -196 -6000 -150 -5988
rect -82 5988 -36 6000
rect -82 -5988 -76 5988
rect -42 -5988 -36 5988
rect -82 -6000 -36 -5988
rect 36 5988 82 6000
rect 36 -5988 42 5988
rect 76 -5988 82 5988
rect 36 -6000 82 -5988
rect 150 5988 196 6000
rect 150 -5988 156 5988
rect 190 -5988 196 5988
rect 150 -6000 196 -5988
rect 268 5988 314 6000
rect 268 -5988 274 5988
rect 308 -5988 314 5988
rect 268 -6000 314 -5988
rect 382 5988 428 6000
rect 382 -5988 388 5988
rect 422 -5988 428 5988
rect 382 -6000 428 -5988
rect 500 5988 546 6000
rect 500 -5988 506 5988
rect 540 -5988 546 5988
rect 500 -6000 546 -5988
rect 614 5988 660 6000
rect 614 -5988 620 5988
rect 654 -5988 660 5988
rect 614 -6000 660 -5988
rect 732 5988 778 6000
rect 732 -5988 738 5988
rect 772 -5988 778 5988
rect 732 -6000 778 -5988
rect 846 5988 892 6000
rect 846 -5988 852 5988
rect 886 -5988 892 5988
rect 846 -6000 892 -5988
rect 964 5988 1010 6000
rect 964 -5988 970 5988
rect 1004 -5988 1010 5988
rect 964 -6000 1010 -5988
rect 1078 5988 1124 6000
rect 1078 -5988 1084 5988
rect 1118 -5988 1124 5988
rect 1078 -6000 1124 -5988
rect 1196 5988 1242 6000
rect 1196 -5988 1202 5988
rect 1236 -5988 1242 5988
rect 1196 -6000 1242 -5988
rect 1310 5988 1356 6000
rect 1310 -5988 1316 5988
rect 1350 -5988 1356 5988
rect 1310 -6000 1356 -5988
rect 1428 5988 1474 6000
rect 1428 -5988 1434 5988
rect 1468 -5988 1474 5988
rect 1428 -6000 1474 -5988
rect 1542 5988 1588 6000
rect 1542 -5988 1548 5988
rect 1582 -5988 1588 5988
rect 1542 -6000 1588 -5988
rect 1660 5988 1706 6000
rect 1660 -5988 1666 5988
rect 1700 -5988 1706 5988
rect 1660 -6000 1706 -5988
rect 1774 5988 1820 6000
rect 1774 -5988 1780 5988
rect 1814 -5988 1820 5988
rect 1774 -6000 1820 -5988
rect 1892 5988 1938 6000
rect 1892 -5988 1898 5988
rect 1932 -5988 1938 5988
rect 1892 -6000 1938 -5988
rect 2006 5988 2052 6000
rect 2006 -5988 2012 5988
rect 2046 -5988 2052 5988
rect 2006 -6000 2052 -5988
rect 2124 5988 2170 6000
rect 2124 -5988 2130 5988
rect 2164 -5988 2170 5988
rect 2124 -6000 2170 -5988
rect 2238 5988 2284 6000
rect 2238 -5988 2244 5988
rect 2278 -5988 2284 5988
rect 2238 -6000 2284 -5988
rect 2356 5988 2402 6000
rect 2356 -5988 2362 5988
rect 2396 -5988 2402 5988
rect 2356 -6000 2402 -5988
rect 2470 5988 2516 6000
rect 2470 -5988 2476 5988
rect 2510 -5988 2516 5988
rect 2470 -6000 2516 -5988
rect 2588 5988 2634 6000
rect 2588 -5988 2594 5988
rect 2628 -5988 2634 5988
rect 2588 -6000 2634 -5988
rect 2702 5988 2748 6000
rect 2702 -5988 2708 5988
rect 2742 -5988 2748 5988
rect 2702 -6000 2748 -5988
rect 2820 5988 2866 6000
rect 2820 -5988 2826 5988
rect 2860 -5988 2866 5988
rect 2820 -6000 2866 -5988
rect 2934 5988 2980 6000
rect 2934 -5988 2940 5988
rect 2974 -5988 2980 5988
rect 2934 -6000 2980 -5988
rect 3052 5988 3098 6000
rect 3052 -5988 3058 5988
rect 3092 -5988 3098 5988
rect 3052 -6000 3098 -5988
rect 3166 5988 3212 6000
rect 3166 -5988 3172 5988
rect 3206 -5988 3212 5988
rect 3166 -6000 3212 -5988
rect 3284 5988 3330 6000
rect 3284 -5988 3290 5988
rect 3324 -5988 3330 5988
rect 3284 -6000 3330 -5988
rect -3277 -6038 -3219 -6032
rect -3277 -6072 -3265 -6038
rect -3231 -6072 -3219 -6038
rect -3277 -6078 -3219 -6072
rect -3045 -6038 -2987 -6032
rect -3045 -6072 -3033 -6038
rect -2999 -6072 -2987 -6038
rect -3045 -6078 -2987 -6072
rect -2813 -6038 -2755 -6032
rect -2813 -6072 -2801 -6038
rect -2767 -6072 -2755 -6038
rect -2813 -6078 -2755 -6072
rect -2581 -6038 -2523 -6032
rect -2581 -6072 -2569 -6038
rect -2535 -6072 -2523 -6038
rect -2581 -6078 -2523 -6072
rect -2349 -6038 -2291 -6032
rect -2349 -6072 -2337 -6038
rect -2303 -6072 -2291 -6038
rect -2349 -6078 -2291 -6072
rect -2117 -6038 -2059 -6032
rect -2117 -6072 -2105 -6038
rect -2071 -6072 -2059 -6038
rect -2117 -6078 -2059 -6072
rect -1885 -6038 -1827 -6032
rect -1885 -6072 -1873 -6038
rect -1839 -6072 -1827 -6038
rect -1885 -6078 -1827 -6072
rect -1653 -6038 -1595 -6032
rect -1653 -6072 -1641 -6038
rect -1607 -6072 -1595 -6038
rect -1653 -6078 -1595 -6072
rect -1421 -6038 -1363 -6032
rect -1421 -6072 -1409 -6038
rect -1375 -6072 -1363 -6038
rect -1421 -6078 -1363 -6072
rect -1189 -6038 -1131 -6032
rect -1189 -6072 -1177 -6038
rect -1143 -6072 -1131 -6038
rect -1189 -6078 -1131 -6072
rect -957 -6038 -899 -6032
rect -957 -6072 -945 -6038
rect -911 -6072 -899 -6038
rect -957 -6078 -899 -6072
rect -725 -6038 -667 -6032
rect -725 -6072 -713 -6038
rect -679 -6072 -667 -6038
rect -725 -6078 -667 -6072
rect -493 -6038 -435 -6032
rect -493 -6072 -481 -6038
rect -447 -6072 -435 -6038
rect -493 -6078 -435 -6072
rect -261 -6038 -203 -6032
rect -261 -6072 -249 -6038
rect -215 -6072 -203 -6038
rect -261 -6078 -203 -6072
rect -29 -6038 29 -6032
rect -29 -6072 -17 -6038
rect 17 -6072 29 -6038
rect -29 -6078 29 -6072
rect 203 -6038 261 -6032
rect 203 -6072 215 -6038
rect 249 -6072 261 -6038
rect 203 -6078 261 -6072
rect 435 -6038 493 -6032
rect 435 -6072 447 -6038
rect 481 -6072 493 -6038
rect 435 -6078 493 -6072
rect 667 -6038 725 -6032
rect 667 -6072 679 -6038
rect 713 -6072 725 -6038
rect 667 -6078 725 -6072
rect 899 -6038 957 -6032
rect 899 -6072 911 -6038
rect 945 -6072 957 -6038
rect 899 -6078 957 -6072
rect 1131 -6038 1189 -6032
rect 1131 -6072 1143 -6038
rect 1177 -6072 1189 -6038
rect 1131 -6078 1189 -6072
rect 1363 -6038 1421 -6032
rect 1363 -6072 1375 -6038
rect 1409 -6072 1421 -6038
rect 1363 -6078 1421 -6072
rect 1595 -6038 1653 -6032
rect 1595 -6072 1607 -6038
rect 1641 -6072 1653 -6038
rect 1595 -6078 1653 -6072
rect 1827 -6038 1885 -6032
rect 1827 -6072 1839 -6038
rect 1873 -6072 1885 -6038
rect 1827 -6078 1885 -6072
rect 2059 -6038 2117 -6032
rect 2059 -6072 2071 -6038
rect 2105 -6072 2117 -6038
rect 2059 -6078 2117 -6072
rect 2291 -6038 2349 -6032
rect 2291 -6072 2303 -6038
rect 2337 -6072 2349 -6038
rect 2291 -6078 2349 -6072
rect 2523 -6038 2581 -6032
rect 2523 -6072 2535 -6038
rect 2569 -6072 2581 -6038
rect 2523 -6078 2581 -6072
rect 2755 -6038 2813 -6032
rect 2755 -6072 2767 -6038
rect 2801 -6072 2813 -6038
rect 2755 -6078 2813 -6072
rect 2987 -6038 3045 -6032
rect 2987 -6072 2999 -6038
rect 3033 -6072 3045 -6038
rect 2987 -6078 3045 -6072
rect 3219 -6038 3277 -6032
rect 3219 -6072 3231 -6038
rect 3265 -6072 3277 -6038
rect 3219 -6078 3277 -6072
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 60 l 0.3 m 1 nf 29 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
