magic
tech sky130A
magscale 1 2
timestamp 1667776540
<< nwell >>
rect -375 -1500 385 1500
<< pmos >>
rect -229 -1400 -29 1400
rect 39 -1400 239 1400
<< pdiff >>
rect -339 1388 -229 1400
rect -339 -1388 -301 1388
rect -267 -1388 -229 1388
rect -339 -1400 -229 -1388
rect -29 1388 39 1400
rect -29 -1388 -12 1388
rect 22 -1388 39 1388
rect -29 -1400 39 -1388
rect 239 1388 349 1400
rect 239 -1388 277 1388
rect 311 -1388 349 1388
rect 239 -1400 349 -1388
<< pdiffc >>
rect -301 -1388 -267 1388
rect -12 -1388 22 1388
rect 277 -1388 311 1388
<< poly >>
rect -229 1481 240 1497
rect -229 1447 55 1481
rect 223 1447 240 1481
rect -229 1435 240 1447
rect -229 1400 -29 1435
rect 39 1400 239 1435
rect -229 -1447 -29 -1400
rect -229 -1481 -213 -1447
rect -45 -1481 -29 -1447
rect -229 -1497 -29 -1481
rect 39 -1447 239 -1400
rect 39 -1481 55 -1447
rect 223 -1481 239 -1447
rect 39 -1497 239 -1481
<< polycont >>
rect 55 1447 223 1481
rect -213 -1481 -45 -1447
rect 55 -1481 223 -1447
<< locali >>
rect 39 1447 55 1481
rect 223 1447 239 1481
rect -301 1388 -267 1404
rect -301 -1404 -267 -1388
rect -12 1388 22 1404
rect -12 -1404 22 -1388
rect 277 1388 311 1404
rect 277 -1404 311 -1388
rect -229 -1481 -213 -1447
rect -45 -1481 -29 -1447
rect 39 -1481 55 -1447
rect 223 -1481 239 -1447
<< viali >>
rect 55 1447 223 1481
rect -301 -1388 -267 1388
rect -12 -1388 22 1388
rect 277 -1388 311 1388
rect -213 -1481 -45 -1447
rect 55 -1481 223 -1447
<< metal1 >>
rect 43 1481 235 1487
rect 43 1447 55 1481
rect 223 1447 235 1481
rect 43 1441 235 1447
rect -307 1388 -261 1400
rect -307 -1388 -301 1388
rect -267 -1388 -261 1388
rect -307 -1400 -261 -1388
rect -18 1388 28 1400
rect -18 -1388 -12 1388
rect 22 -1388 28 1388
rect -18 -1400 28 -1388
rect 271 1388 317 1400
rect 271 -1388 277 1388
rect 311 -1388 317 1388
rect 271 -1400 317 -1388
rect -225 -1447 -33 -1441
rect -225 -1481 -213 -1447
rect -45 -1481 -33 -1447
rect -225 -1487 -33 -1481
rect 43 -1447 235 -1441
rect 43 -1481 55 -1447
rect 223 -1481 235 -1447
rect 43 -1487 235 -1481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 14 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
