magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -560 6072 -502 6078
rect -560 6038 -548 6072
rect -560 6032 -502 6038
<< pwell >>
rect -645 -6026 645 6026
<< nmos >>
rect -561 -6000 -501 6000
rect -443 -6000 -383 6000
rect -325 -6000 -265 6000
rect -207 -6000 -147 6000
rect -89 -6000 -29 6000
rect 29 -6000 89 6000
rect 147 -6000 207 6000
rect 265 -6000 325 6000
rect 383 -6000 443 6000
rect 501 -6000 561 6000
<< ndiff >>
rect -619 5967 -561 6000
rect -619 5933 -607 5967
rect -573 5933 -561 5967
rect -619 5899 -561 5933
rect -619 5865 -607 5899
rect -573 5865 -561 5899
rect -619 5831 -561 5865
rect -619 5797 -607 5831
rect -573 5797 -561 5831
rect -619 5763 -561 5797
rect -619 5729 -607 5763
rect -573 5729 -561 5763
rect -619 5695 -561 5729
rect -619 5661 -607 5695
rect -573 5661 -561 5695
rect -619 5627 -561 5661
rect -619 5593 -607 5627
rect -573 5593 -561 5627
rect -619 5559 -561 5593
rect -619 5525 -607 5559
rect -573 5525 -561 5559
rect -619 5491 -561 5525
rect -619 5457 -607 5491
rect -573 5457 -561 5491
rect -619 5423 -561 5457
rect -619 5389 -607 5423
rect -573 5389 -561 5423
rect -619 5355 -561 5389
rect -619 5321 -607 5355
rect -573 5321 -561 5355
rect -619 5287 -561 5321
rect -619 5253 -607 5287
rect -573 5253 -561 5287
rect -619 5219 -561 5253
rect -619 5185 -607 5219
rect -573 5185 -561 5219
rect -619 5151 -561 5185
rect -619 5117 -607 5151
rect -573 5117 -561 5151
rect -619 5083 -561 5117
rect -619 5049 -607 5083
rect -573 5049 -561 5083
rect -619 5015 -561 5049
rect -619 4981 -607 5015
rect -573 4981 -561 5015
rect -619 4947 -561 4981
rect -619 4913 -607 4947
rect -573 4913 -561 4947
rect -619 4879 -561 4913
rect -619 4845 -607 4879
rect -573 4845 -561 4879
rect -619 4811 -561 4845
rect -619 4777 -607 4811
rect -573 4777 -561 4811
rect -619 4743 -561 4777
rect -619 4709 -607 4743
rect -573 4709 -561 4743
rect -619 4675 -561 4709
rect -619 4641 -607 4675
rect -573 4641 -561 4675
rect -619 4607 -561 4641
rect -619 4573 -607 4607
rect -573 4573 -561 4607
rect -619 4539 -561 4573
rect -619 4505 -607 4539
rect -573 4505 -561 4539
rect -619 4471 -561 4505
rect -619 4437 -607 4471
rect -573 4437 -561 4471
rect -619 4403 -561 4437
rect -619 4369 -607 4403
rect -573 4369 -561 4403
rect -619 4335 -561 4369
rect -619 4301 -607 4335
rect -573 4301 -561 4335
rect -619 4267 -561 4301
rect -619 4233 -607 4267
rect -573 4233 -561 4267
rect -619 4199 -561 4233
rect -619 4165 -607 4199
rect -573 4165 -561 4199
rect -619 4131 -561 4165
rect -619 4097 -607 4131
rect -573 4097 -561 4131
rect -619 4063 -561 4097
rect -619 4029 -607 4063
rect -573 4029 -561 4063
rect -619 3995 -561 4029
rect -619 3961 -607 3995
rect -573 3961 -561 3995
rect -619 3927 -561 3961
rect -619 3893 -607 3927
rect -573 3893 -561 3927
rect -619 3859 -561 3893
rect -619 3825 -607 3859
rect -573 3825 -561 3859
rect -619 3791 -561 3825
rect -619 3757 -607 3791
rect -573 3757 -561 3791
rect -619 3723 -561 3757
rect -619 3689 -607 3723
rect -573 3689 -561 3723
rect -619 3655 -561 3689
rect -619 3621 -607 3655
rect -573 3621 -561 3655
rect -619 3587 -561 3621
rect -619 3553 -607 3587
rect -573 3553 -561 3587
rect -619 3519 -561 3553
rect -619 3485 -607 3519
rect -573 3485 -561 3519
rect -619 3451 -561 3485
rect -619 3417 -607 3451
rect -573 3417 -561 3451
rect -619 3383 -561 3417
rect -619 3349 -607 3383
rect -573 3349 -561 3383
rect -619 3315 -561 3349
rect -619 3281 -607 3315
rect -573 3281 -561 3315
rect -619 3247 -561 3281
rect -619 3213 -607 3247
rect -573 3213 -561 3247
rect -619 3179 -561 3213
rect -619 3145 -607 3179
rect -573 3145 -561 3179
rect -619 3111 -561 3145
rect -619 3077 -607 3111
rect -573 3077 -561 3111
rect -619 3043 -561 3077
rect -619 3009 -607 3043
rect -573 3009 -561 3043
rect -619 2975 -561 3009
rect -619 2941 -607 2975
rect -573 2941 -561 2975
rect -619 2907 -561 2941
rect -619 2873 -607 2907
rect -573 2873 -561 2907
rect -619 2839 -561 2873
rect -619 2805 -607 2839
rect -573 2805 -561 2839
rect -619 2771 -561 2805
rect -619 2737 -607 2771
rect -573 2737 -561 2771
rect -619 2703 -561 2737
rect -619 2669 -607 2703
rect -573 2669 -561 2703
rect -619 2635 -561 2669
rect -619 2601 -607 2635
rect -573 2601 -561 2635
rect -619 2567 -561 2601
rect -619 2533 -607 2567
rect -573 2533 -561 2567
rect -619 2499 -561 2533
rect -619 2465 -607 2499
rect -573 2465 -561 2499
rect -619 2431 -561 2465
rect -619 2397 -607 2431
rect -573 2397 -561 2431
rect -619 2363 -561 2397
rect -619 2329 -607 2363
rect -573 2329 -561 2363
rect -619 2295 -561 2329
rect -619 2261 -607 2295
rect -573 2261 -561 2295
rect -619 2227 -561 2261
rect -619 2193 -607 2227
rect -573 2193 -561 2227
rect -619 2159 -561 2193
rect -619 2125 -607 2159
rect -573 2125 -561 2159
rect -619 2091 -561 2125
rect -619 2057 -607 2091
rect -573 2057 -561 2091
rect -619 2023 -561 2057
rect -619 1989 -607 2023
rect -573 1989 -561 2023
rect -619 1955 -561 1989
rect -619 1921 -607 1955
rect -573 1921 -561 1955
rect -619 1887 -561 1921
rect -619 1853 -607 1887
rect -573 1853 -561 1887
rect -619 1819 -561 1853
rect -619 1785 -607 1819
rect -573 1785 -561 1819
rect -619 1751 -561 1785
rect -619 1717 -607 1751
rect -573 1717 -561 1751
rect -619 1683 -561 1717
rect -619 1649 -607 1683
rect -573 1649 -561 1683
rect -619 1615 -561 1649
rect -619 1581 -607 1615
rect -573 1581 -561 1615
rect -619 1547 -561 1581
rect -619 1513 -607 1547
rect -573 1513 -561 1547
rect -619 1479 -561 1513
rect -619 1445 -607 1479
rect -573 1445 -561 1479
rect -619 1411 -561 1445
rect -619 1377 -607 1411
rect -573 1377 -561 1411
rect -619 1343 -561 1377
rect -619 1309 -607 1343
rect -573 1309 -561 1343
rect -619 1275 -561 1309
rect -619 1241 -607 1275
rect -573 1241 -561 1275
rect -619 1207 -561 1241
rect -619 1173 -607 1207
rect -573 1173 -561 1207
rect -619 1139 -561 1173
rect -619 1105 -607 1139
rect -573 1105 -561 1139
rect -619 1071 -561 1105
rect -619 1037 -607 1071
rect -573 1037 -561 1071
rect -619 1003 -561 1037
rect -619 969 -607 1003
rect -573 969 -561 1003
rect -619 935 -561 969
rect -619 901 -607 935
rect -573 901 -561 935
rect -619 867 -561 901
rect -619 833 -607 867
rect -573 833 -561 867
rect -619 799 -561 833
rect -619 765 -607 799
rect -573 765 -561 799
rect -619 731 -561 765
rect -619 697 -607 731
rect -573 697 -561 731
rect -619 663 -561 697
rect -619 629 -607 663
rect -573 629 -561 663
rect -619 595 -561 629
rect -619 561 -607 595
rect -573 561 -561 595
rect -619 527 -561 561
rect -619 493 -607 527
rect -573 493 -561 527
rect -619 459 -561 493
rect -619 425 -607 459
rect -573 425 -561 459
rect -619 391 -561 425
rect -619 357 -607 391
rect -573 357 -561 391
rect -619 323 -561 357
rect -619 289 -607 323
rect -573 289 -561 323
rect -619 255 -561 289
rect -619 221 -607 255
rect -573 221 -561 255
rect -619 187 -561 221
rect -619 153 -607 187
rect -573 153 -561 187
rect -619 119 -561 153
rect -619 85 -607 119
rect -573 85 -561 119
rect -619 51 -561 85
rect -619 17 -607 51
rect -573 17 -561 51
rect -619 -17 -561 17
rect -619 -51 -607 -17
rect -573 -51 -561 -17
rect -619 -85 -561 -51
rect -619 -119 -607 -85
rect -573 -119 -561 -85
rect -619 -153 -561 -119
rect -619 -187 -607 -153
rect -573 -187 -561 -153
rect -619 -221 -561 -187
rect -619 -255 -607 -221
rect -573 -255 -561 -221
rect -619 -289 -561 -255
rect -619 -323 -607 -289
rect -573 -323 -561 -289
rect -619 -357 -561 -323
rect -619 -391 -607 -357
rect -573 -391 -561 -357
rect -619 -425 -561 -391
rect -619 -459 -607 -425
rect -573 -459 -561 -425
rect -619 -493 -561 -459
rect -619 -527 -607 -493
rect -573 -527 -561 -493
rect -619 -561 -561 -527
rect -619 -595 -607 -561
rect -573 -595 -561 -561
rect -619 -629 -561 -595
rect -619 -663 -607 -629
rect -573 -663 -561 -629
rect -619 -697 -561 -663
rect -619 -731 -607 -697
rect -573 -731 -561 -697
rect -619 -765 -561 -731
rect -619 -799 -607 -765
rect -573 -799 -561 -765
rect -619 -833 -561 -799
rect -619 -867 -607 -833
rect -573 -867 -561 -833
rect -619 -901 -561 -867
rect -619 -935 -607 -901
rect -573 -935 -561 -901
rect -619 -969 -561 -935
rect -619 -1003 -607 -969
rect -573 -1003 -561 -969
rect -619 -1037 -561 -1003
rect -619 -1071 -607 -1037
rect -573 -1071 -561 -1037
rect -619 -1105 -561 -1071
rect -619 -1139 -607 -1105
rect -573 -1139 -561 -1105
rect -619 -1173 -561 -1139
rect -619 -1207 -607 -1173
rect -573 -1207 -561 -1173
rect -619 -1241 -561 -1207
rect -619 -1275 -607 -1241
rect -573 -1275 -561 -1241
rect -619 -1309 -561 -1275
rect -619 -1343 -607 -1309
rect -573 -1343 -561 -1309
rect -619 -1377 -561 -1343
rect -619 -1411 -607 -1377
rect -573 -1411 -561 -1377
rect -619 -1445 -561 -1411
rect -619 -1479 -607 -1445
rect -573 -1479 -561 -1445
rect -619 -1513 -561 -1479
rect -619 -1547 -607 -1513
rect -573 -1547 -561 -1513
rect -619 -1581 -561 -1547
rect -619 -1615 -607 -1581
rect -573 -1615 -561 -1581
rect -619 -1649 -561 -1615
rect -619 -1683 -607 -1649
rect -573 -1683 -561 -1649
rect -619 -1717 -561 -1683
rect -619 -1751 -607 -1717
rect -573 -1751 -561 -1717
rect -619 -1785 -561 -1751
rect -619 -1819 -607 -1785
rect -573 -1819 -561 -1785
rect -619 -1853 -561 -1819
rect -619 -1887 -607 -1853
rect -573 -1887 -561 -1853
rect -619 -1921 -561 -1887
rect -619 -1955 -607 -1921
rect -573 -1955 -561 -1921
rect -619 -1989 -561 -1955
rect -619 -2023 -607 -1989
rect -573 -2023 -561 -1989
rect -619 -2057 -561 -2023
rect -619 -2091 -607 -2057
rect -573 -2091 -561 -2057
rect -619 -2125 -561 -2091
rect -619 -2159 -607 -2125
rect -573 -2159 -561 -2125
rect -619 -2193 -561 -2159
rect -619 -2227 -607 -2193
rect -573 -2227 -561 -2193
rect -619 -2261 -561 -2227
rect -619 -2295 -607 -2261
rect -573 -2295 -561 -2261
rect -619 -2329 -561 -2295
rect -619 -2363 -607 -2329
rect -573 -2363 -561 -2329
rect -619 -2397 -561 -2363
rect -619 -2431 -607 -2397
rect -573 -2431 -561 -2397
rect -619 -2465 -561 -2431
rect -619 -2499 -607 -2465
rect -573 -2499 -561 -2465
rect -619 -2533 -561 -2499
rect -619 -2567 -607 -2533
rect -573 -2567 -561 -2533
rect -619 -2601 -561 -2567
rect -619 -2635 -607 -2601
rect -573 -2635 -561 -2601
rect -619 -2669 -561 -2635
rect -619 -2703 -607 -2669
rect -573 -2703 -561 -2669
rect -619 -2737 -561 -2703
rect -619 -2771 -607 -2737
rect -573 -2771 -561 -2737
rect -619 -2805 -561 -2771
rect -619 -2839 -607 -2805
rect -573 -2839 -561 -2805
rect -619 -2873 -561 -2839
rect -619 -2907 -607 -2873
rect -573 -2907 -561 -2873
rect -619 -2941 -561 -2907
rect -619 -2975 -607 -2941
rect -573 -2975 -561 -2941
rect -619 -3009 -561 -2975
rect -619 -3043 -607 -3009
rect -573 -3043 -561 -3009
rect -619 -3077 -561 -3043
rect -619 -3111 -607 -3077
rect -573 -3111 -561 -3077
rect -619 -3145 -561 -3111
rect -619 -3179 -607 -3145
rect -573 -3179 -561 -3145
rect -619 -3213 -561 -3179
rect -619 -3247 -607 -3213
rect -573 -3247 -561 -3213
rect -619 -3281 -561 -3247
rect -619 -3315 -607 -3281
rect -573 -3315 -561 -3281
rect -619 -3349 -561 -3315
rect -619 -3383 -607 -3349
rect -573 -3383 -561 -3349
rect -619 -3417 -561 -3383
rect -619 -3451 -607 -3417
rect -573 -3451 -561 -3417
rect -619 -3485 -561 -3451
rect -619 -3519 -607 -3485
rect -573 -3519 -561 -3485
rect -619 -3553 -561 -3519
rect -619 -3587 -607 -3553
rect -573 -3587 -561 -3553
rect -619 -3621 -561 -3587
rect -619 -3655 -607 -3621
rect -573 -3655 -561 -3621
rect -619 -3689 -561 -3655
rect -619 -3723 -607 -3689
rect -573 -3723 -561 -3689
rect -619 -3757 -561 -3723
rect -619 -3791 -607 -3757
rect -573 -3791 -561 -3757
rect -619 -3825 -561 -3791
rect -619 -3859 -607 -3825
rect -573 -3859 -561 -3825
rect -619 -3893 -561 -3859
rect -619 -3927 -607 -3893
rect -573 -3927 -561 -3893
rect -619 -3961 -561 -3927
rect -619 -3995 -607 -3961
rect -573 -3995 -561 -3961
rect -619 -4029 -561 -3995
rect -619 -4063 -607 -4029
rect -573 -4063 -561 -4029
rect -619 -4097 -561 -4063
rect -619 -4131 -607 -4097
rect -573 -4131 -561 -4097
rect -619 -4165 -561 -4131
rect -619 -4199 -607 -4165
rect -573 -4199 -561 -4165
rect -619 -4233 -561 -4199
rect -619 -4267 -607 -4233
rect -573 -4267 -561 -4233
rect -619 -4301 -561 -4267
rect -619 -4335 -607 -4301
rect -573 -4335 -561 -4301
rect -619 -4369 -561 -4335
rect -619 -4403 -607 -4369
rect -573 -4403 -561 -4369
rect -619 -4437 -561 -4403
rect -619 -4471 -607 -4437
rect -573 -4471 -561 -4437
rect -619 -4505 -561 -4471
rect -619 -4539 -607 -4505
rect -573 -4539 -561 -4505
rect -619 -4573 -561 -4539
rect -619 -4607 -607 -4573
rect -573 -4607 -561 -4573
rect -619 -4641 -561 -4607
rect -619 -4675 -607 -4641
rect -573 -4675 -561 -4641
rect -619 -4709 -561 -4675
rect -619 -4743 -607 -4709
rect -573 -4743 -561 -4709
rect -619 -4777 -561 -4743
rect -619 -4811 -607 -4777
rect -573 -4811 -561 -4777
rect -619 -4845 -561 -4811
rect -619 -4879 -607 -4845
rect -573 -4879 -561 -4845
rect -619 -4913 -561 -4879
rect -619 -4947 -607 -4913
rect -573 -4947 -561 -4913
rect -619 -4981 -561 -4947
rect -619 -5015 -607 -4981
rect -573 -5015 -561 -4981
rect -619 -5049 -561 -5015
rect -619 -5083 -607 -5049
rect -573 -5083 -561 -5049
rect -619 -5117 -561 -5083
rect -619 -5151 -607 -5117
rect -573 -5151 -561 -5117
rect -619 -5185 -561 -5151
rect -619 -5219 -607 -5185
rect -573 -5219 -561 -5185
rect -619 -5253 -561 -5219
rect -619 -5287 -607 -5253
rect -573 -5287 -561 -5253
rect -619 -5321 -561 -5287
rect -619 -5355 -607 -5321
rect -573 -5355 -561 -5321
rect -619 -5389 -561 -5355
rect -619 -5423 -607 -5389
rect -573 -5423 -561 -5389
rect -619 -5457 -561 -5423
rect -619 -5491 -607 -5457
rect -573 -5491 -561 -5457
rect -619 -5525 -561 -5491
rect -619 -5559 -607 -5525
rect -573 -5559 -561 -5525
rect -619 -5593 -561 -5559
rect -619 -5627 -607 -5593
rect -573 -5627 -561 -5593
rect -619 -5661 -561 -5627
rect -619 -5695 -607 -5661
rect -573 -5695 -561 -5661
rect -619 -5729 -561 -5695
rect -619 -5763 -607 -5729
rect -573 -5763 -561 -5729
rect -619 -5797 -561 -5763
rect -619 -5831 -607 -5797
rect -573 -5831 -561 -5797
rect -619 -5865 -561 -5831
rect -619 -5899 -607 -5865
rect -573 -5899 -561 -5865
rect -619 -5933 -561 -5899
rect -619 -5967 -607 -5933
rect -573 -5967 -561 -5933
rect -619 -6000 -561 -5967
rect -501 5967 -443 6000
rect -501 5933 -489 5967
rect -455 5933 -443 5967
rect -501 5899 -443 5933
rect -501 5865 -489 5899
rect -455 5865 -443 5899
rect -501 5831 -443 5865
rect -501 5797 -489 5831
rect -455 5797 -443 5831
rect -501 5763 -443 5797
rect -501 5729 -489 5763
rect -455 5729 -443 5763
rect -501 5695 -443 5729
rect -501 5661 -489 5695
rect -455 5661 -443 5695
rect -501 5627 -443 5661
rect -501 5593 -489 5627
rect -455 5593 -443 5627
rect -501 5559 -443 5593
rect -501 5525 -489 5559
rect -455 5525 -443 5559
rect -501 5491 -443 5525
rect -501 5457 -489 5491
rect -455 5457 -443 5491
rect -501 5423 -443 5457
rect -501 5389 -489 5423
rect -455 5389 -443 5423
rect -501 5355 -443 5389
rect -501 5321 -489 5355
rect -455 5321 -443 5355
rect -501 5287 -443 5321
rect -501 5253 -489 5287
rect -455 5253 -443 5287
rect -501 5219 -443 5253
rect -501 5185 -489 5219
rect -455 5185 -443 5219
rect -501 5151 -443 5185
rect -501 5117 -489 5151
rect -455 5117 -443 5151
rect -501 5083 -443 5117
rect -501 5049 -489 5083
rect -455 5049 -443 5083
rect -501 5015 -443 5049
rect -501 4981 -489 5015
rect -455 4981 -443 5015
rect -501 4947 -443 4981
rect -501 4913 -489 4947
rect -455 4913 -443 4947
rect -501 4879 -443 4913
rect -501 4845 -489 4879
rect -455 4845 -443 4879
rect -501 4811 -443 4845
rect -501 4777 -489 4811
rect -455 4777 -443 4811
rect -501 4743 -443 4777
rect -501 4709 -489 4743
rect -455 4709 -443 4743
rect -501 4675 -443 4709
rect -501 4641 -489 4675
rect -455 4641 -443 4675
rect -501 4607 -443 4641
rect -501 4573 -489 4607
rect -455 4573 -443 4607
rect -501 4539 -443 4573
rect -501 4505 -489 4539
rect -455 4505 -443 4539
rect -501 4471 -443 4505
rect -501 4437 -489 4471
rect -455 4437 -443 4471
rect -501 4403 -443 4437
rect -501 4369 -489 4403
rect -455 4369 -443 4403
rect -501 4335 -443 4369
rect -501 4301 -489 4335
rect -455 4301 -443 4335
rect -501 4267 -443 4301
rect -501 4233 -489 4267
rect -455 4233 -443 4267
rect -501 4199 -443 4233
rect -501 4165 -489 4199
rect -455 4165 -443 4199
rect -501 4131 -443 4165
rect -501 4097 -489 4131
rect -455 4097 -443 4131
rect -501 4063 -443 4097
rect -501 4029 -489 4063
rect -455 4029 -443 4063
rect -501 3995 -443 4029
rect -501 3961 -489 3995
rect -455 3961 -443 3995
rect -501 3927 -443 3961
rect -501 3893 -489 3927
rect -455 3893 -443 3927
rect -501 3859 -443 3893
rect -501 3825 -489 3859
rect -455 3825 -443 3859
rect -501 3791 -443 3825
rect -501 3757 -489 3791
rect -455 3757 -443 3791
rect -501 3723 -443 3757
rect -501 3689 -489 3723
rect -455 3689 -443 3723
rect -501 3655 -443 3689
rect -501 3621 -489 3655
rect -455 3621 -443 3655
rect -501 3587 -443 3621
rect -501 3553 -489 3587
rect -455 3553 -443 3587
rect -501 3519 -443 3553
rect -501 3485 -489 3519
rect -455 3485 -443 3519
rect -501 3451 -443 3485
rect -501 3417 -489 3451
rect -455 3417 -443 3451
rect -501 3383 -443 3417
rect -501 3349 -489 3383
rect -455 3349 -443 3383
rect -501 3315 -443 3349
rect -501 3281 -489 3315
rect -455 3281 -443 3315
rect -501 3247 -443 3281
rect -501 3213 -489 3247
rect -455 3213 -443 3247
rect -501 3179 -443 3213
rect -501 3145 -489 3179
rect -455 3145 -443 3179
rect -501 3111 -443 3145
rect -501 3077 -489 3111
rect -455 3077 -443 3111
rect -501 3043 -443 3077
rect -501 3009 -489 3043
rect -455 3009 -443 3043
rect -501 2975 -443 3009
rect -501 2941 -489 2975
rect -455 2941 -443 2975
rect -501 2907 -443 2941
rect -501 2873 -489 2907
rect -455 2873 -443 2907
rect -501 2839 -443 2873
rect -501 2805 -489 2839
rect -455 2805 -443 2839
rect -501 2771 -443 2805
rect -501 2737 -489 2771
rect -455 2737 -443 2771
rect -501 2703 -443 2737
rect -501 2669 -489 2703
rect -455 2669 -443 2703
rect -501 2635 -443 2669
rect -501 2601 -489 2635
rect -455 2601 -443 2635
rect -501 2567 -443 2601
rect -501 2533 -489 2567
rect -455 2533 -443 2567
rect -501 2499 -443 2533
rect -501 2465 -489 2499
rect -455 2465 -443 2499
rect -501 2431 -443 2465
rect -501 2397 -489 2431
rect -455 2397 -443 2431
rect -501 2363 -443 2397
rect -501 2329 -489 2363
rect -455 2329 -443 2363
rect -501 2295 -443 2329
rect -501 2261 -489 2295
rect -455 2261 -443 2295
rect -501 2227 -443 2261
rect -501 2193 -489 2227
rect -455 2193 -443 2227
rect -501 2159 -443 2193
rect -501 2125 -489 2159
rect -455 2125 -443 2159
rect -501 2091 -443 2125
rect -501 2057 -489 2091
rect -455 2057 -443 2091
rect -501 2023 -443 2057
rect -501 1989 -489 2023
rect -455 1989 -443 2023
rect -501 1955 -443 1989
rect -501 1921 -489 1955
rect -455 1921 -443 1955
rect -501 1887 -443 1921
rect -501 1853 -489 1887
rect -455 1853 -443 1887
rect -501 1819 -443 1853
rect -501 1785 -489 1819
rect -455 1785 -443 1819
rect -501 1751 -443 1785
rect -501 1717 -489 1751
rect -455 1717 -443 1751
rect -501 1683 -443 1717
rect -501 1649 -489 1683
rect -455 1649 -443 1683
rect -501 1615 -443 1649
rect -501 1581 -489 1615
rect -455 1581 -443 1615
rect -501 1547 -443 1581
rect -501 1513 -489 1547
rect -455 1513 -443 1547
rect -501 1479 -443 1513
rect -501 1445 -489 1479
rect -455 1445 -443 1479
rect -501 1411 -443 1445
rect -501 1377 -489 1411
rect -455 1377 -443 1411
rect -501 1343 -443 1377
rect -501 1309 -489 1343
rect -455 1309 -443 1343
rect -501 1275 -443 1309
rect -501 1241 -489 1275
rect -455 1241 -443 1275
rect -501 1207 -443 1241
rect -501 1173 -489 1207
rect -455 1173 -443 1207
rect -501 1139 -443 1173
rect -501 1105 -489 1139
rect -455 1105 -443 1139
rect -501 1071 -443 1105
rect -501 1037 -489 1071
rect -455 1037 -443 1071
rect -501 1003 -443 1037
rect -501 969 -489 1003
rect -455 969 -443 1003
rect -501 935 -443 969
rect -501 901 -489 935
rect -455 901 -443 935
rect -501 867 -443 901
rect -501 833 -489 867
rect -455 833 -443 867
rect -501 799 -443 833
rect -501 765 -489 799
rect -455 765 -443 799
rect -501 731 -443 765
rect -501 697 -489 731
rect -455 697 -443 731
rect -501 663 -443 697
rect -501 629 -489 663
rect -455 629 -443 663
rect -501 595 -443 629
rect -501 561 -489 595
rect -455 561 -443 595
rect -501 527 -443 561
rect -501 493 -489 527
rect -455 493 -443 527
rect -501 459 -443 493
rect -501 425 -489 459
rect -455 425 -443 459
rect -501 391 -443 425
rect -501 357 -489 391
rect -455 357 -443 391
rect -501 323 -443 357
rect -501 289 -489 323
rect -455 289 -443 323
rect -501 255 -443 289
rect -501 221 -489 255
rect -455 221 -443 255
rect -501 187 -443 221
rect -501 153 -489 187
rect -455 153 -443 187
rect -501 119 -443 153
rect -501 85 -489 119
rect -455 85 -443 119
rect -501 51 -443 85
rect -501 17 -489 51
rect -455 17 -443 51
rect -501 -17 -443 17
rect -501 -51 -489 -17
rect -455 -51 -443 -17
rect -501 -85 -443 -51
rect -501 -119 -489 -85
rect -455 -119 -443 -85
rect -501 -153 -443 -119
rect -501 -187 -489 -153
rect -455 -187 -443 -153
rect -501 -221 -443 -187
rect -501 -255 -489 -221
rect -455 -255 -443 -221
rect -501 -289 -443 -255
rect -501 -323 -489 -289
rect -455 -323 -443 -289
rect -501 -357 -443 -323
rect -501 -391 -489 -357
rect -455 -391 -443 -357
rect -501 -425 -443 -391
rect -501 -459 -489 -425
rect -455 -459 -443 -425
rect -501 -493 -443 -459
rect -501 -527 -489 -493
rect -455 -527 -443 -493
rect -501 -561 -443 -527
rect -501 -595 -489 -561
rect -455 -595 -443 -561
rect -501 -629 -443 -595
rect -501 -663 -489 -629
rect -455 -663 -443 -629
rect -501 -697 -443 -663
rect -501 -731 -489 -697
rect -455 -731 -443 -697
rect -501 -765 -443 -731
rect -501 -799 -489 -765
rect -455 -799 -443 -765
rect -501 -833 -443 -799
rect -501 -867 -489 -833
rect -455 -867 -443 -833
rect -501 -901 -443 -867
rect -501 -935 -489 -901
rect -455 -935 -443 -901
rect -501 -969 -443 -935
rect -501 -1003 -489 -969
rect -455 -1003 -443 -969
rect -501 -1037 -443 -1003
rect -501 -1071 -489 -1037
rect -455 -1071 -443 -1037
rect -501 -1105 -443 -1071
rect -501 -1139 -489 -1105
rect -455 -1139 -443 -1105
rect -501 -1173 -443 -1139
rect -501 -1207 -489 -1173
rect -455 -1207 -443 -1173
rect -501 -1241 -443 -1207
rect -501 -1275 -489 -1241
rect -455 -1275 -443 -1241
rect -501 -1309 -443 -1275
rect -501 -1343 -489 -1309
rect -455 -1343 -443 -1309
rect -501 -1377 -443 -1343
rect -501 -1411 -489 -1377
rect -455 -1411 -443 -1377
rect -501 -1445 -443 -1411
rect -501 -1479 -489 -1445
rect -455 -1479 -443 -1445
rect -501 -1513 -443 -1479
rect -501 -1547 -489 -1513
rect -455 -1547 -443 -1513
rect -501 -1581 -443 -1547
rect -501 -1615 -489 -1581
rect -455 -1615 -443 -1581
rect -501 -1649 -443 -1615
rect -501 -1683 -489 -1649
rect -455 -1683 -443 -1649
rect -501 -1717 -443 -1683
rect -501 -1751 -489 -1717
rect -455 -1751 -443 -1717
rect -501 -1785 -443 -1751
rect -501 -1819 -489 -1785
rect -455 -1819 -443 -1785
rect -501 -1853 -443 -1819
rect -501 -1887 -489 -1853
rect -455 -1887 -443 -1853
rect -501 -1921 -443 -1887
rect -501 -1955 -489 -1921
rect -455 -1955 -443 -1921
rect -501 -1989 -443 -1955
rect -501 -2023 -489 -1989
rect -455 -2023 -443 -1989
rect -501 -2057 -443 -2023
rect -501 -2091 -489 -2057
rect -455 -2091 -443 -2057
rect -501 -2125 -443 -2091
rect -501 -2159 -489 -2125
rect -455 -2159 -443 -2125
rect -501 -2193 -443 -2159
rect -501 -2227 -489 -2193
rect -455 -2227 -443 -2193
rect -501 -2261 -443 -2227
rect -501 -2295 -489 -2261
rect -455 -2295 -443 -2261
rect -501 -2329 -443 -2295
rect -501 -2363 -489 -2329
rect -455 -2363 -443 -2329
rect -501 -2397 -443 -2363
rect -501 -2431 -489 -2397
rect -455 -2431 -443 -2397
rect -501 -2465 -443 -2431
rect -501 -2499 -489 -2465
rect -455 -2499 -443 -2465
rect -501 -2533 -443 -2499
rect -501 -2567 -489 -2533
rect -455 -2567 -443 -2533
rect -501 -2601 -443 -2567
rect -501 -2635 -489 -2601
rect -455 -2635 -443 -2601
rect -501 -2669 -443 -2635
rect -501 -2703 -489 -2669
rect -455 -2703 -443 -2669
rect -501 -2737 -443 -2703
rect -501 -2771 -489 -2737
rect -455 -2771 -443 -2737
rect -501 -2805 -443 -2771
rect -501 -2839 -489 -2805
rect -455 -2839 -443 -2805
rect -501 -2873 -443 -2839
rect -501 -2907 -489 -2873
rect -455 -2907 -443 -2873
rect -501 -2941 -443 -2907
rect -501 -2975 -489 -2941
rect -455 -2975 -443 -2941
rect -501 -3009 -443 -2975
rect -501 -3043 -489 -3009
rect -455 -3043 -443 -3009
rect -501 -3077 -443 -3043
rect -501 -3111 -489 -3077
rect -455 -3111 -443 -3077
rect -501 -3145 -443 -3111
rect -501 -3179 -489 -3145
rect -455 -3179 -443 -3145
rect -501 -3213 -443 -3179
rect -501 -3247 -489 -3213
rect -455 -3247 -443 -3213
rect -501 -3281 -443 -3247
rect -501 -3315 -489 -3281
rect -455 -3315 -443 -3281
rect -501 -3349 -443 -3315
rect -501 -3383 -489 -3349
rect -455 -3383 -443 -3349
rect -501 -3417 -443 -3383
rect -501 -3451 -489 -3417
rect -455 -3451 -443 -3417
rect -501 -3485 -443 -3451
rect -501 -3519 -489 -3485
rect -455 -3519 -443 -3485
rect -501 -3553 -443 -3519
rect -501 -3587 -489 -3553
rect -455 -3587 -443 -3553
rect -501 -3621 -443 -3587
rect -501 -3655 -489 -3621
rect -455 -3655 -443 -3621
rect -501 -3689 -443 -3655
rect -501 -3723 -489 -3689
rect -455 -3723 -443 -3689
rect -501 -3757 -443 -3723
rect -501 -3791 -489 -3757
rect -455 -3791 -443 -3757
rect -501 -3825 -443 -3791
rect -501 -3859 -489 -3825
rect -455 -3859 -443 -3825
rect -501 -3893 -443 -3859
rect -501 -3927 -489 -3893
rect -455 -3927 -443 -3893
rect -501 -3961 -443 -3927
rect -501 -3995 -489 -3961
rect -455 -3995 -443 -3961
rect -501 -4029 -443 -3995
rect -501 -4063 -489 -4029
rect -455 -4063 -443 -4029
rect -501 -4097 -443 -4063
rect -501 -4131 -489 -4097
rect -455 -4131 -443 -4097
rect -501 -4165 -443 -4131
rect -501 -4199 -489 -4165
rect -455 -4199 -443 -4165
rect -501 -4233 -443 -4199
rect -501 -4267 -489 -4233
rect -455 -4267 -443 -4233
rect -501 -4301 -443 -4267
rect -501 -4335 -489 -4301
rect -455 -4335 -443 -4301
rect -501 -4369 -443 -4335
rect -501 -4403 -489 -4369
rect -455 -4403 -443 -4369
rect -501 -4437 -443 -4403
rect -501 -4471 -489 -4437
rect -455 -4471 -443 -4437
rect -501 -4505 -443 -4471
rect -501 -4539 -489 -4505
rect -455 -4539 -443 -4505
rect -501 -4573 -443 -4539
rect -501 -4607 -489 -4573
rect -455 -4607 -443 -4573
rect -501 -4641 -443 -4607
rect -501 -4675 -489 -4641
rect -455 -4675 -443 -4641
rect -501 -4709 -443 -4675
rect -501 -4743 -489 -4709
rect -455 -4743 -443 -4709
rect -501 -4777 -443 -4743
rect -501 -4811 -489 -4777
rect -455 -4811 -443 -4777
rect -501 -4845 -443 -4811
rect -501 -4879 -489 -4845
rect -455 -4879 -443 -4845
rect -501 -4913 -443 -4879
rect -501 -4947 -489 -4913
rect -455 -4947 -443 -4913
rect -501 -4981 -443 -4947
rect -501 -5015 -489 -4981
rect -455 -5015 -443 -4981
rect -501 -5049 -443 -5015
rect -501 -5083 -489 -5049
rect -455 -5083 -443 -5049
rect -501 -5117 -443 -5083
rect -501 -5151 -489 -5117
rect -455 -5151 -443 -5117
rect -501 -5185 -443 -5151
rect -501 -5219 -489 -5185
rect -455 -5219 -443 -5185
rect -501 -5253 -443 -5219
rect -501 -5287 -489 -5253
rect -455 -5287 -443 -5253
rect -501 -5321 -443 -5287
rect -501 -5355 -489 -5321
rect -455 -5355 -443 -5321
rect -501 -5389 -443 -5355
rect -501 -5423 -489 -5389
rect -455 -5423 -443 -5389
rect -501 -5457 -443 -5423
rect -501 -5491 -489 -5457
rect -455 -5491 -443 -5457
rect -501 -5525 -443 -5491
rect -501 -5559 -489 -5525
rect -455 -5559 -443 -5525
rect -501 -5593 -443 -5559
rect -501 -5627 -489 -5593
rect -455 -5627 -443 -5593
rect -501 -5661 -443 -5627
rect -501 -5695 -489 -5661
rect -455 -5695 -443 -5661
rect -501 -5729 -443 -5695
rect -501 -5763 -489 -5729
rect -455 -5763 -443 -5729
rect -501 -5797 -443 -5763
rect -501 -5831 -489 -5797
rect -455 -5831 -443 -5797
rect -501 -5865 -443 -5831
rect -501 -5899 -489 -5865
rect -455 -5899 -443 -5865
rect -501 -5933 -443 -5899
rect -501 -5967 -489 -5933
rect -455 -5967 -443 -5933
rect -501 -6000 -443 -5967
rect -383 5967 -325 6000
rect -383 5933 -371 5967
rect -337 5933 -325 5967
rect -383 5899 -325 5933
rect -383 5865 -371 5899
rect -337 5865 -325 5899
rect -383 5831 -325 5865
rect -383 5797 -371 5831
rect -337 5797 -325 5831
rect -383 5763 -325 5797
rect -383 5729 -371 5763
rect -337 5729 -325 5763
rect -383 5695 -325 5729
rect -383 5661 -371 5695
rect -337 5661 -325 5695
rect -383 5627 -325 5661
rect -383 5593 -371 5627
rect -337 5593 -325 5627
rect -383 5559 -325 5593
rect -383 5525 -371 5559
rect -337 5525 -325 5559
rect -383 5491 -325 5525
rect -383 5457 -371 5491
rect -337 5457 -325 5491
rect -383 5423 -325 5457
rect -383 5389 -371 5423
rect -337 5389 -325 5423
rect -383 5355 -325 5389
rect -383 5321 -371 5355
rect -337 5321 -325 5355
rect -383 5287 -325 5321
rect -383 5253 -371 5287
rect -337 5253 -325 5287
rect -383 5219 -325 5253
rect -383 5185 -371 5219
rect -337 5185 -325 5219
rect -383 5151 -325 5185
rect -383 5117 -371 5151
rect -337 5117 -325 5151
rect -383 5083 -325 5117
rect -383 5049 -371 5083
rect -337 5049 -325 5083
rect -383 5015 -325 5049
rect -383 4981 -371 5015
rect -337 4981 -325 5015
rect -383 4947 -325 4981
rect -383 4913 -371 4947
rect -337 4913 -325 4947
rect -383 4879 -325 4913
rect -383 4845 -371 4879
rect -337 4845 -325 4879
rect -383 4811 -325 4845
rect -383 4777 -371 4811
rect -337 4777 -325 4811
rect -383 4743 -325 4777
rect -383 4709 -371 4743
rect -337 4709 -325 4743
rect -383 4675 -325 4709
rect -383 4641 -371 4675
rect -337 4641 -325 4675
rect -383 4607 -325 4641
rect -383 4573 -371 4607
rect -337 4573 -325 4607
rect -383 4539 -325 4573
rect -383 4505 -371 4539
rect -337 4505 -325 4539
rect -383 4471 -325 4505
rect -383 4437 -371 4471
rect -337 4437 -325 4471
rect -383 4403 -325 4437
rect -383 4369 -371 4403
rect -337 4369 -325 4403
rect -383 4335 -325 4369
rect -383 4301 -371 4335
rect -337 4301 -325 4335
rect -383 4267 -325 4301
rect -383 4233 -371 4267
rect -337 4233 -325 4267
rect -383 4199 -325 4233
rect -383 4165 -371 4199
rect -337 4165 -325 4199
rect -383 4131 -325 4165
rect -383 4097 -371 4131
rect -337 4097 -325 4131
rect -383 4063 -325 4097
rect -383 4029 -371 4063
rect -337 4029 -325 4063
rect -383 3995 -325 4029
rect -383 3961 -371 3995
rect -337 3961 -325 3995
rect -383 3927 -325 3961
rect -383 3893 -371 3927
rect -337 3893 -325 3927
rect -383 3859 -325 3893
rect -383 3825 -371 3859
rect -337 3825 -325 3859
rect -383 3791 -325 3825
rect -383 3757 -371 3791
rect -337 3757 -325 3791
rect -383 3723 -325 3757
rect -383 3689 -371 3723
rect -337 3689 -325 3723
rect -383 3655 -325 3689
rect -383 3621 -371 3655
rect -337 3621 -325 3655
rect -383 3587 -325 3621
rect -383 3553 -371 3587
rect -337 3553 -325 3587
rect -383 3519 -325 3553
rect -383 3485 -371 3519
rect -337 3485 -325 3519
rect -383 3451 -325 3485
rect -383 3417 -371 3451
rect -337 3417 -325 3451
rect -383 3383 -325 3417
rect -383 3349 -371 3383
rect -337 3349 -325 3383
rect -383 3315 -325 3349
rect -383 3281 -371 3315
rect -337 3281 -325 3315
rect -383 3247 -325 3281
rect -383 3213 -371 3247
rect -337 3213 -325 3247
rect -383 3179 -325 3213
rect -383 3145 -371 3179
rect -337 3145 -325 3179
rect -383 3111 -325 3145
rect -383 3077 -371 3111
rect -337 3077 -325 3111
rect -383 3043 -325 3077
rect -383 3009 -371 3043
rect -337 3009 -325 3043
rect -383 2975 -325 3009
rect -383 2941 -371 2975
rect -337 2941 -325 2975
rect -383 2907 -325 2941
rect -383 2873 -371 2907
rect -337 2873 -325 2907
rect -383 2839 -325 2873
rect -383 2805 -371 2839
rect -337 2805 -325 2839
rect -383 2771 -325 2805
rect -383 2737 -371 2771
rect -337 2737 -325 2771
rect -383 2703 -325 2737
rect -383 2669 -371 2703
rect -337 2669 -325 2703
rect -383 2635 -325 2669
rect -383 2601 -371 2635
rect -337 2601 -325 2635
rect -383 2567 -325 2601
rect -383 2533 -371 2567
rect -337 2533 -325 2567
rect -383 2499 -325 2533
rect -383 2465 -371 2499
rect -337 2465 -325 2499
rect -383 2431 -325 2465
rect -383 2397 -371 2431
rect -337 2397 -325 2431
rect -383 2363 -325 2397
rect -383 2329 -371 2363
rect -337 2329 -325 2363
rect -383 2295 -325 2329
rect -383 2261 -371 2295
rect -337 2261 -325 2295
rect -383 2227 -325 2261
rect -383 2193 -371 2227
rect -337 2193 -325 2227
rect -383 2159 -325 2193
rect -383 2125 -371 2159
rect -337 2125 -325 2159
rect -383 2091 -325 2125
rect -383 2057 -371 2091
rect -337 2057 -325 2091
rect -383 2023 -325 2057
rect -383 1989 -371 2023
rect -337 1989 -325 2023
rect -383 1955 -325 1989
rect -383 1921 -371 1955
rect -337 1921 -325 1955
rect -383 1887 -325 1921
rect -383 1853 -371 1887
rect -337 1853 -325 1887
rect -383 1819 -325 1853
rect -383 1785 -371 1819
rect -337 1785 -325 1819
rect -383 1751 -325 1785
rect -383 1717 -371 1751
rect -337 1717 -325 1751
rect -383 1683 -325 1717
rect -383 1649 -371 1683
rect -337 1649 -325 1683
rect -383 1615 -325 1649
rect -383 1581 -371 1615
rect -337 1581 -325 1615
rect -383 1547 -325 1581
rect -383 1513 -371 1547
rect -337 1513 -325 1547
rect -383 1479 -325 1513
rect -383 1445 -371 1479
rect -337 1445 -325 1479
rect -383 1411 -325 1445
rect -383 1377 -371 1411
rect -337 1377 -325 1411
rect -383 1343 -325 1377
rect -383 1309 -371 1343
rect -337 1309 -325 1343
rect -383 1275 -325 1309
rect -383 1241 -371 1275
rect -337 1241 -325 1275
rect -383 1207 -325 1241
rect -383 1173 -371 1207
rect -337 1173 -325 1207
rect -383 1139 -325 1173
rect -383 1105 -371 1139
rect -337 1105 -325 1139
rect -383 1071 -325 1105
rect -383 1037 -371 1071
rect -337 1037 -325 1071
rect -383 1003 -325 1037
rect -383 969 -371 1003
rect -337 969 -325 1003
rect -383 935 -325 969
rect -383 901 -371 935
rect -337 901 -325 935
rect -383 867 -325 901
rect -383 833 -371 867
rect -337 833 -325 867
rect -383 799 -325 833
rect -383 765 -371 799
rect -337 765 -325 799
rect -383 731 -325 765
rect -383 697 -371 731
rect -337 697 -325 731
rect -383 663 -325 697
rect -383 629 -371 663
rect -337 629 -325 663
rect -383 595 -325 629
rect -383 561 -371 595
rect -337 561 -325 595
rect -383 527 -325 561
rect -383 493 -371 527
rect -337 493 -325 527
rect -383 459 -325 493
rect -383 425 -371 459
rect -337 425 -325 459
rect -383 391 -325 425
rect -383 357 -371 391
rect -337 357 -325 391
rect -383 323 -325 357
rect -383 289 -371 323
rect -337 289 -325 323
rect -383 255 -325 289
rect -383 221 -371 255
rect -337 221 -325 255
rect -383 187 -325 221
rect -383 153 -371 187
rect -337 153 -325 187
rect -383 119 -325 153
rect -383 85 -371 119
rect -337 85 -325 119
rect -383 51 -325 85
rect -383 17 -371 51
rect -337 17 -325 51
rect -383 -17 -325 17
rect -383 -51 -371 -17
rect -337 -51 -325 -17
rect -383 -85 -325 -51
rect -383 -119 -371 -85
rect -337 -119 -325 -85
rect -383 -153 -325 -119
rect -383 -187 -371 -153
rect -337 -187 -325 -153
rect -383 -221 -325 -187
rect -383 -255 -371 -221
rect -337 -255 -325 -221
rect -383 -289 -325 -255
rect -383 -323 -371 -289
rect -337 -323 -325 -289
rect -383 -357 -325 -323
rect -383 -391 -371 -357
rect -337 -391 -325 -357
rect -383 -425 -325 -391
rect -383 -459 -371 -425
rect -337 -459 -325 -425
rect -383 -493 -325 -459
rect -383 -527 -371 -493
rect -337 -527 -325 -493
rect -383 -561 -325 -527
rect -383 -595 -371 -561
rect -337 -595 -325 -561
rect -383 -629 -325 -595
rect -383 -663 -371 -629
rect -337 -663 -325 -629
rect -383 -697 -325 -663
rect -383 -731 -371 -697
rect -337 -731 -325 -697
rect -383 -765 -325 -731
rect -383 -799 -371 -765
rect -337 -799 -325 -765
rect -383 -833 -325 -799
rect -383 -867 -371 -833
rect -337 -867 -325 -833
rect -383 -901 -325 -867
rect -383 -935 -371 -901
rect -337 -935 -325 -901
rect -383 -969 -325 -935
rect -383 -1003 -371 -969
rect -337 -1003 -325 -969
rect -383 -1037 -325 -1003
rect -383 -1071 -371 -1037
rect -337 -1071 -325 -1037
rect -383 -1105 -325 -1071
rect -383 -1139 -371 -1105
rect -337 -1139 -325 -1105
rect -383 -1173 -325 -1139
rect -383 -1207 -371 -1173
rect -337 -1207 -325 -1173
rect -383 -1241 -325 -1207
rect -383 -1275 -371 -1241
rect -337 -1275 -325 -1241
rect -383 -1309 -325 -1275
rect -383 -1343 -371 -1309
rect -337 -1343 -325 -1309
rect -383 -1377 -325 -1343
rect -383 -1411 -371 -1377
rect -337 -1411 -325 -1377
rect -383 -1445 -325 -1411
rect -383 -1479 -371 -1445
rect -337 -1479 -325 -1445
rect -383 -1513 -325 -1479
rect -383 -1547 -371 -1513
rect -337 -1547 -325 -1513
rect -383 -1581 -325 -1547
rect -383 -1615 -371 -1581
rect -337 -1615 -325 -1581
rect -383 -1649 -325 -1615
rect -383 -1683 -371 -1649
rect -337 -1683 -325 -1649
rect -383 -1717 -325 -1683
rect -383 -1751 -371 -1717
rect -337 -1751 -325 -1717
rect -383 -1785 -325 -1751
rect -383 -1819 -371 -1785
rect -337 -1819 -325 -1785
rect -383 -1853 -325 -1819
rect -383 -1887 -371 -1853
rect -337 -1887 -325 -1853
rect -383 -1921 -325 -1887
rect -383 -1955 -371 -1921
rect -337 -1955 -325 -1921
rect -383 -1989 -325 -1955
rect -383 -2023 -371 -1989
rect -337 -2023 -325 -1989
rect -383 -2057 -325 -2023
rect -383 -2091 -371 -2057
rect -337 -2091 -325 -2057
rect -383 -2125 -325 -2091
rect -383 -2159 -371 -2125
rect -337 -2159 -325 -2125
rect -383 -2193 -325 -2159
rect -383 -2227 -371 -2193
rect -337 -2227 -325 -2193
rect -383 -2261 -325 -2227
rect -383 -2295 -371 -2261
rect -337 -2295 -325 -2261
rect -383 -2329 -325 -2295
rect -383 -2363 -371 -2329
rect -337 -2363 -325 -2329
rect -383 -2397 -325 -2363
rect -383 -2431 -371 -2397
rect -337 -2431 -325 -2397
rect -383 -2465 -325 -2431
rect -383 -2499 -371 -2465
rect -337 -2499 -325 -2465
rect -383 -2533 -325 -2499
rect -383 -2567 -371 -2533
rect -337 -2567 -325 -2533
rect -383 -2601 -325 -2567
rect -383 -2635 -371 -2601
rect -337 -2635 -325 -2601
rect -383 -2669 -325 -2635
rect -383 -2703 -371 -2669
rect -337 -2703 -325 -2669
rect -383 -2737 -325 -2703
rect -383 -2771 -371 -2737
rect -337 -2771 -325 -2737
rect -383 -2805 -325 -2771
rect -383 -2839 -371 -2805
rect -337 -2839 -325 -2805
rect -383 -2873 -325 -2839
rect -383 -2907 -371 -2873
rect -337 -2907 -325 -2873
rect -383 -2941 -325 -2907
rect -383 -2975 -371 -2941
rect -337 -2975 -325 -2941
rect -383 -3009 -325 -2975
rect -383 -3043 -371 -3009
rect -337 -3043 -325 -3009
rect -383 -3077 -325 -3043
rect -383 -3111 -371 -3077
rect -337 -3111 -325 -3077
rect -383 -3145 -325 -3111
rect -383 -3179 -371 -3145
rect -337 -3179 -325 -3145
rect -383 -3213 -325 -3179
rect -383 -3247 -371 -3213
rect -337 -3247 -325 -3213
rect -383 -3281 -325 -3247
rect -383 -3315 -371 -3281
rect -337 -3315 -325 -3281
rect -383 -3349 -325 -3315
rect -383 -3383 -371 -3349
rect -337 -3383 -325 -3349
rect -383 -3417 -325 -3383
rect -383 -3451 -371 -3417
rect -337 -3451 -325 -3417
rect -383 -3485 -325 -3451
rect -383 -3519 -371 -3485
rect -337 -3519 -325 -3485
rect -383 -3553 -325 -3519
rect -383 -3587 -371 -3553
rect -337 -3587 -325 -3553
rect -383 -3621 -325 -3587
rect -383 -3655 -371 -3621
rect -337 -3655 -325 -3621
rect -383 -3689 -325 -3655
rect -383 -3723 -371 -3689
rect -337 -3723 -325 -3689
rect -383 -3757 -325 -3723
rect -383 -3791 -371 -3757
rect -337 -3791 -325 -3757
rect -383 -3825 -325 -3791
rect -383 -3859 -371 -3825
rect -337 -3859 -325 -3825
rect -383 -3893 -325 -3859
rect -383 -3927 -371 -3893
rect -337 -3927 -325 -3893
rect -383 -3961 -325 -3927
rect -383 -3995 -371 -3961
rect -337 -3995 -325 -3961
rect -383 -4029 -325 -3995
rect -383 -4063 -371 -4029
rect -337 -4063 -325 -4029
rect -383 -4097 -325 -4063
rect -383 -4131 -371 -4097
rect -337 -4131 -325 -4097
rect -383 -4165 -325 -4131
rect -383 -4199 -371 -4165
rect -337 -4199 -325 -4165
rect -383 -4233 -325 -4199
rect -383 -4267 -371 -4233
rect -337 -4267 -325 -4233
rect -383 -4301 -325 -4267
rect -383 -4335 -371 -4301
rect -337 -4335 -325 -4301
rect -383 -4369 -325 -4335
rect -383 -4403 -371 -4369
rect -337 -4403 -325 -4369
rect -383 -4437 -325 -4403
rect -383 -4471 -371 -4437
rect -337 -4471 -325 -4437
rect -383 -4505 -325 -4471
rect -383 -4539 -371 -4505
rect -337 -4539 -325 -4505
rect -383 -4573 -325 -4539
rect -383 -4607 -371 -4573
rect -337 -4607 -325 -4573
rect -383 -4641 -325 -4607
rect -383 -4675 -371 -4641
rect -337 -4675 -325 -4641
rect -383 -4709 -325 -4675
rect -383 -4743 -371 -4709
rect -337 -4743 -325 -4709
rect -383 -4777 -325 -4743
rect -383 -4811 -371 -4777
rect -337 -4811 -325 -4777
rect -383 -4845 -325 -4811
rect -383 -4879 -371 -4845
rect -337 -4879 -325 -4845
rect -383 -4913 -325 -4879
rect -383 -4947 -371 -4913
rect -337 -4947 -325 -4913
rect -383 -4981 -325 -4947
rect -383 -5015 -371 -4981
rect -337 -5015 -325 -4981
rect -383 -5049 -325 -5015
rect -383 -5083 -371 -5049
rect -337 -5083 -325 -5049
rect -383 -5117 -325 -5083
rect -383 -5151 -371 -5117
rect -337 -5151 -325 -5117
rect -383 -5185 -325 -5151
rect -383 -5219 -371 -5185
rect -337 -5219 -325 -5185
rect -383 -5253 -325 -5219
rect -383 -5287 -371 -5253
rect -337 -5287 -325 -5253
rect -383 -5321 -325 -5287
rect -383 -5355 -371 -5321
rect -337 -5355 -325 -5321
rect -383 -5389 -325 -5355
rect -383 -5423 -371 -5389
rect -337 -5423 -325 -5389
rect -383 -5457 -325 -5423
rect -383 -5491 -371 -5457
rect -337 -5491 -325 -5457
rect -383 -5525 -325 -5491
rect -383 -5559 -371 -5525
rect -337 -5559 -325 -5525
rect -383 -5593 -325 -5559
rect -383 -5627 -371 -5593
rect -337 -5627 -325 -5593
rect -383 -5661 -325 -5627
rect -383 -5695 -371 -5661
rect -337 -5695 -325 -5661
rect -383 -5729 -325 -5695
rect -383 -5763 -371 -5729
rect -337 -5763 -325 -5729
rect -383 -5797 -325 -5763
rect -383 -5831 -371 -5797
rect -337 -5831 -325 -5797
rect -383 -5865 -325 -5831
rect -383 -5899 -371 -5865
rect -337 -5899 -325 -5865
rect -383 -5933 -325 -5899
rect -383 -5967 -371 -5933
rect -337 -5967 -325 -5933
rect -383 -6000 -325 -5967
rect -265 5967 -207 6000
rect -265 5933 -253 5967
rect -219 5933 -207 5967
rect -265 5899 -207 5933
rect -265 5865 -253 5899
rect -219 5865 -207 5899
rect -265 5831 -207 5865
rect -265 5797 -253 5831
rect -219 5797 -207 5831
rect -265 5763 -207 5797
rect -265 5729 -253 5763
rect -219 5729 -207 5763
rect -265 5695 -207 5729
rect -265 5661 -253 5695
rect -219 5661 -207 5695
rect -265 5627 -207 5661
rect -265 5593 -253 5627
rect -219 5593 -207 5627
rect -265 5559 -207 5593
rect -265 5525 -253 5559
rect -219 5525 -207 5559
rect -265 5491 -207 5525
rect -265 5457 -253 5491
rect -219 5457 -207 5491
rect -265 5423 -207 5457
rect -265 5389 -253 5423
rect -219 5389 -207 5423
rect -265 5355 -207 5389
rect -265 5321 -253 5355
rect -219 5321 -207 5355
rect -265 5287 -207 5321
rect -265 5253 -253 5287
rect -219 5253 -207 5287
rect -265 5219 -207 5253
rect -265 5185 -253 5219
rect -219 5185 -207 5219
rect -265 5151 -207 5185
rect -265 5117 -253 5151
rect -219 5117 -207 5151
rect -265 5083 -207 5117
rect -265 5049 -253 5083
rect -219 5049 -207 5083
rect -265 5015 -207 5049
rect -265 4981 -253 5015
rect -219 4981 -207 5015
rect -265 4947 -207 4981
rect -265 4913 -253 4947
rect -219 4913 -207 4947
rect -265 4879 -207 4913
rect -265 4845 -253 4879
rect -219 4845 -207 4879
rect -265 4811 -207 4845
rect -265 4777 -253 4811
rect -219 4777 -207 4811
rect -265 4743 -207 4777
rect -265 4709 -253 4743
rect -219 4709 -207 4743
rect -265 4675 -207 4709
rect -265 4641 -253 4675
rect -219 4641 -207 4675
rect -265 4607 -207 4641
rect -265 4573 -253 4607
rect -219 4573 -207 4607
rect -265 4539 -207 4573
rect -265 4505 -253 4539
rect -219 4505 -207 4539
rect -265 4471 -207 4505
rect -265 4437 -253 4471
rect -219 4437 -207 4471
rect -265 4403 -207 4437
rect -265 4369 -253 4403
rect -219 4369 -207 4403
rect -265 4335 -207 4369
rect -265 4301 -253 4335
rect -219 4301 -207 4335
rect -265 4267 -207 4301
rect -265 4233 -253 4267
rect -219 4233 -207 4267
rect -265 4199 -207 4233
rect -265 4165 -253 4199
rect -219 4165 -207 4199
rect -265 4131 -207 4165
rect -265 4097 -253 4131
rect -219 4097 -207 4131
rect -265 4063 -207 4097
rect -265 4029 -253 4063
rect -219 4029 -207 4063
rect -265 3995 -207 4029
rect -265 3961 -253 3995
rect -219 3961 -207 3995
rect -265 3927 -207 3961
rect -265 3893 -253 3927
rect -219 3893 -207 3927
rect -265 3859 -207 3893
rect -265 3825 -253 3859
rect -219 3825 -207 3859
rect -265 3791 -207 3825
rect -265 3757 -253 3791
rect -219 3757 -207 3791
rect -265 3723 -207 3757
rect -265 3689 -253 3723
rect -219 3689 -207 3723
rect -265 3655 -207 3689
rect -265 3621 -253 3655
rect -219 3621 -207 3655
rect -265 3587 -207 3621
rect -265 3553 -253 3587
rect -219 3553 -207 3587
rect -265 3519 -207 3553
rect -265 3485 -253 3519
rect -219 3485 -207 3519
rect -265 3451 -207 3485
rect -265 3417 -253 3451
rect -219 3417 -207 3451
rect -265 3383 -207 3417
rect -265 3349 -253 3383
rect -219 3349 -207 3383
rect -265 3315 -207 3349
rect -265 3281 -253 3315
rect -219 3281 -207 3315
rect -265 3247 -207 3281
rect -265 3213 -253 3247
rect -219 3213 -207 3247
rect -265 3179 -207 3213
rect -265 3145 -253 3179
rect -219 3145 -207 3179
rect -265 3111 -207 3145
rect -265 3077 -253 3111
rect -219 3077 -207 3111
rect -265 3043 -207 3077
rect -265 3009 -253 3043
rect -219 3009 -207 3043
rect -265 2975 -207 3009
rect -265 2941 -253 2975
rect -219 2941 -207 2975
rect -265 2907 -207 2941
rect -265 2873 -253 2907
rect -219 2873 -207 2907
rect -265 2839 -207 2873
rect -265 2805 -253 2839
rect -219 2805 -207 2839
rect -265 2771 -207 2805
rect -265 2737 -253 2771
rect -219 2737 -207 2771
rect -265 2703 -207 2737
rect -265 2669 -253 2703
rect -219 2669 -207 2703
rect -265 2635 -207 2669
rect -265 2601 -253 2635
rect -219 2601 -207 2635
rect -265 2567 -207 2601
rect -265 2533 -253 2567
rect -219 2533 -207 2567
rect -265 2499 -207 2533
rect -265 2465 -253 2499
rect -219 2465 -207 2499
rect -265 2431 -207 2465
rect -265 2397 -253 2431
rect -219 2397 -207 2431
rect -265 2363 -207 2397
rect -265 2329 -253 2363
rect -219 2329 -207 2363
rect -265 2295 -207 2329
rect -265 2261 -253 2295
rect -219 2261 -207 2295
rect -265 2227 -207 2261
rect -265 2193 -253 2227
rect -219 2193 -207 2227
rect -265 2159 -207 2193
rect -265 2125 -253 2159
rect -219 2125 -207 2159
rect -265 2091 -207 2125
rect -265 2057 -253 2091
rect -219 2057 -207 2091
rect -265 2023 -207 2057
rect -265 1989 -253 2023
rect -219 1989 -207 2023
rect -265 1955 -207 1989
rect -265 1921 -253 1955
rect -219 1921 -207 1955
rect -265 1887 -207 1921
rect -265 1853 -253 1887
rect -219 1853 -207 1887
rect -265 1819 -207 1853
rect -265 1785 -253 1819
rect -219 1785 -207 1819
rect -265 1751 -207 1785
rect -265 1717 -253 1751
rect -219 1717 -207 1751
rect -265 1683 -207 1717
rect -265 1649 -253 1683
rect -219 1649 -207 1683
rect -265 1615 -207 1649
rect -265 1581 -253 1615
rect -219 1581 -207 1615
rect -265 1547 -207 1581
rect -265 1513 -253 1547
rect -219 1513 -207 1547
rect -265 1479 -207 1513
rect -265 1445 -253 1479
rect -219 1445 -207 1479
rect -265 1411 -207 1445
rect -265 1377 -253 1411
rect -219 1377 -207 1411
rect -265 1343 -207 1377
rect -265 1309 -253 1343
rect -219 1309 -207 1343
rect -265 1275 -207 1309
rect -265 1241 -253 1275
rect -219 1241 -207 1275
rect -265 1207 -207 1241
rect -265 1173 -253 1207
rect -219 1173 -207 1207
rect -265 1139 -207 1173
rect -265 1105 -253 1139
rect -219 1105 -207 1139
rect -265 1071 -207 1105
rect -265 1037 -253 1071
rect -219 1037 -207 1071
rect -265 1003 -207 1037
rect -265 969 -253 1003
rect -219 969 -207 1003
rect -265 935 -207 969
rect -265 901 -253 935
rect -219 901 -207 935
rect -265 867 -207 901
rect -265 833 -253 867
rect -219 833 -207 867
rect -265 799 -207 833
rect -265 765 -253 799
rect -219 765 -207 799
rect -265 731 -207 765
rect -265 697 -253 731
rect -219 697 -207 731
rect -265 663 -207 697
rect -265 629 -253 663
rect -219 629 -207 663
rect -265 595 -207 629
rect -265 561 -253 595
rect -219 561 -207 595
rect -265 527 -207 561
rect -265 493 -253 527
rect -219 493 -207 527
rect -265 459 -207 493
rect -265 425 -253 459
rect -219 425 -207 459
rect -265 391 -207 425
rect -265 357 -253 391
rect -219 357 -207 391
rect -265 323 -207 357
rect -265 289 -253 323
rect -219 289 -207 323
rect -265 255 -207 289
rect -265 221 -253 255
rect -219 221 -207 255
rect -265 187 -207 221
rect -265 153 -253 187
rect -219 153 -207 187
rect -265 119 -207 153
rect -265 85 -253 119
rect -219 85 -207 119
rect -265 51 -207 85
rect -265 17 -253 51
rect -219 17 -207 51
rect -265 -17 -207 17
rect -265 -51 -253 -17
rect -219 -51 -207 -17
rect -265 -85 -207 -51
rect -265 -119 -253 -85
rect -219 -119 -207 -85
rect -265 -153 -207 -119
rect -265 -187 -253 -153
rect -219 -187 -207 -153
rect -265 -221 -207 -187
rect -265 -255 -253 -221
rect -219 -255 -207 -221
rect -265 -289 -207 -255
rect -265 -323 -253 -289
rect -219 -323 -207 -289
rect -265 -357 -207 -323
rect -265 -391 -253 -357
rect -219 -391 -207 -357
rect -265 -425 -207 -391
rect -265 -459 -253 -425
rect -219 -459 -207 -425
rect -265 -493 -207 -459
rect -265 -527 -253 -493
rect -219 -527 -207 -493
rect -265 -561 -207 -527
rect -265 -595 -253 -561
rect -219 -595 -207 -561
rect -265 -629 -207 -595
rect -265 -663 -253 -629
rect -219 -663 -207 -629
rect -265 -697 -207 -663
rect -265 -731 -253 -697
rect -219 -731 -207 -697
rect -265 -765 -207 -731
rect -265 -799 -253 -765
rect -219 -799 -207 -765
rect -265 -833 -207 -799
rect -265 -867 -253 -833
rect -219 -867 -207 -833
rect -265 -901 -207 -867
rect -265 -935 -253 -901
rect -219 -935 -207 -901
rect -265 -969 -207 -935
rect -265 -1003 -253 -969
rect -219 -1003 -207 -969
rect -265 -1037 -207 -1003
rect -265 -1071 -253 -1037
rect -219 -1071 -207 -1037
rect -265 -1105 -207 -1071
rect -265 -1139 -253 -1105
rect -219 -1139 -207 -1105
rect -265 -1173 -207 -1139
rect -265 -1207 -253 -1173
rect -219 -1207 -207 -1173
rect -265 -1241 -207 -1207
rect -265 -1275 -253 -1241
rect -219 -1275 -207 -1241
rect -265 -1309 -207 -1275
rect -265 -1343 -253 -1309
rect -219 -1343 -207 -1309
rect -265 -1377 -207 -1343
rect -265 -1411 -253 -1377
rect -219 -1411 -207 -1377
rect -265 -1445 -207 -1411
rect -265 -1479 -253 -1445
rect -219 -1479 -207 -1445
rect -265 -1513 -207 -1479
rect -265 -1547 -253 -1513
rect -219 -1547 -207 -1513
rect -265 -1581 -207 -1547
rect -265 -1615 -253 -1581
rect -219 -1615 -207 -1581
rect -265 -1649 -207 -1615
rect -265 -1683 -253 -1649
rect -219 -1683 -207 -1649
rect -265 -1717 -207 -1683
rect -265 -1751 -253 -1717
rect -219 -1751 -207 -1717
rect -265 -1785 -207 -1751
rect -265 -1819 -253 -1785
rect -219 -1819 -207 -1785
rect -265 -1853 -207 -1819
rect -265 -1887 -253 -1853
rect -219 -1887 -207 -1853
rect -265 -1921 -207 -1887
rect -265 -1955 -253 -1921
rect -219 -1955 -207 -1921
rect -265 -1989 -207 -1955
rect -265 -2023 -253 -1989
rect -219 -2023 -207 -1989
rect -265 -2057 -207 -2023
rect -265 -2091 -253 -2057
rect -219 -2091 -207 -2057
rect -265 -2125 -207 -2091
rect -265 -2159 -253 -2125
rect -219 -2159 -207 -2125
rect -265 -2193 -207 -2159
rect -265 -2227 -253 -2193
rect -219 -2227 -207 -2193
rect -265 -2261 -207 -2227
rect -265 -2295 -253 -2261
rect -219 -2295 -207 -2261
rect -265 -2329 -207 -2295
rect -265 -2363 -253 -2329
rect -219 -2363 -207 -2329
rect -265 -2397 -207 -2363
rect -265 -2431 -253 -2397
rect -219 -2431 -207 -2397
rect -265 -2465 -207 -2431
rect -265 -2499 -253 -2465
rect -219 -2499 -207 -2465
rect -265 -2533 -207 -2499
rect -265 -2567 -253 -2533
rect -219 -2567 -207 -2533
rect -265 -2601 -207 -2567
rect -265 -2635 -253 -2601
rect -219 -2635 -207 -2601
rect -265 -2669 -207 -2635
rect -265 -2703 -253 -2669
rect -219 -2703 -207 -2669
rect -265 -2737 -207 -2703
rect -265 -2771 -253 -2737
rect -219 -2771 -207 -2737
rect -265 -2805 -207 -2771
rect -265 -2839 -253 -2805
rect -219 -2839 -207 -2805
rect -265 -2873 -207 -2839
rect -265 -2907 -253 -2873
rect -219 -2907 -207 -2873
rect -265 -2941 -207 -2907
rect -265 -2975 -253 -2941
rect -219 -2975 -207 -2941
rect -265 -3009 -207 -2975
rect -265 -3043 -253 -3009
rect -219 -3043 -207 -3009
rect -265 -3077 -207 -3043
rect -265 -3111 -253 -3077
rect -219 -3111 -207 -3077
rect -265 -3145 -207 -3111
rect -265 -3179 -253 -3145
rect -219 -3179 -207 -3145
rect -265 -3213 -207 -3179
rect -265 -3247 -253 -3213
rect -219 -3247 -207 -3213
rect -265 -3281 -207 -3247
rect -265 -3315 -253 -3281
rect -219 -3315 -207 -3281
rect -265 -3349 -207 -3315
rect -265 -3383 -253 -3349
rect -219 -3383 -207 -3349
rect -265 -3417 -207 -3383
rect -265 -3451 -253 -3417
rect -219 -3451 -207 -3417
rect -265 -3485 -207 -3451
rect -265 -3519 -253 -3485
rect -219 -3519 -207 -3485
rect -265 -3553 -207 -3519
rect -265 -3587 -253 -3553
rect -219 -3587 -207 -3553
rect -265 -3621 -207 -3587
rect -265 -3655 -253 -3621
rect -219 -3655 -207 -3621
rect -265 -3689 -207 -3655
rect -265 -3723 -253 -3689
rect -219 -3723 -207 -3689
rect -265 -3757 -207 -3723
rect -265 -3791 -253 -3757
rect -219 -3791 -207 -3757
rect -265 -3825 -207 -3791
rect -265 -3859 -253 -3825
rect -219 -3859 -207 -3825
rect -265 -3893 -207 -3859
rect -265 -3927 -253 -3893
rect -219 -3927 -207 -3893
rect -265 -3961 -207 -3927
rect -265 -3995 -253 -3961
rect -219 -3995 -207 -3961
rect -265 -4029 -207 -3995
rect -265 -4063 -253 -4029
rect -219 -4063 -207 -4029
rect -265 -4097 -207 -4063
rect -265 -4131 -253 -4097
rect -219 -4131 -207 -4097
rect -265 -4165 -207 -4131
rect -265 -4199 -253 -4165
rect -219 -4199 -207 -4165
rect -265 -4233 -207 -4199
rect -265 -4267 -253 -4233
rect -219 -4267 -207 -4233
rect -265 -4301 -207 -4267
rect -265 -4335 -253 -4301
rect -219 -4335 -207 -4301
rect -265 -4369 -207 -4335
rect -265 -4403 -253 -4369
rect -219 -4403 -207 -4369
rect -265 -4437 -207 -4403
rect -265 -4471 -253 -4437
rect -219 -4471 -207 -4437
rect -265 -4505 -207 -4471
rect -265 -4539 -253 -4505
rect -219 -4539 -207 -4505
rect -265 -4573 -207 -4539
rect -265 -4607 -253 -4573
rect -219 -4607 -207 -4573
rect -265 -4641 -207 -4607
rect -265 -4675 -253 -4641
rect -219 -4675 -207 -4641
rect -265 -4709 -207 -4675
rect -265 -4743 -253 -4709
rect -219 -4743 -207 -4709
rect -265 -4777 -207 -4743
rect -265 -4811 -253 -4777
rect -219 -4811 -207 -4777
rect -265 -4845 -207 -4811
rect -265 -4879 -253 -4845
rect -219 -4879 -207 -4845
rect -265 -4913 -207 -4879
rect -265 -4947 -253 -4913
rect -219 -4947 -207 -4913
rect -265 -4981 -207 -4947
rect -265 -5015 -253 -4981
rect -219 -5015 -207 -4981
rect -265 -5049 -207 -5015
rect -265 -5083 -253 -5049
rect -219 -5083 -207 -5049
rect -265 -5117 -207 -5083
rect -265 -5151 -253 -5117
rect -219 -5151 -207 -5117
rect -265 -5185 -207 -5151
rect -265 -5219 -253 -5185
rect -219 -5219 -207 -5185
rect -265 -5253 -207 -5219
rect -265 -5287 -253 -5253
rect -219 -5287 -207 -5253
rect -265 -5321 -207 -5287
rect -265 -5355 -253 -5321
rect -219 -5355 -207 -5321
rect -265 -5389 -207 -5355
rect -265 -5423 -253 -5389
rect -219 -5423 -207 -5389
rect -265 -5457 -207 -5423
rect -265 -5491 -253 -5457
rect -219 -5491 -207 -5457
rect -265 -5525 -207 -5491
rect -265 -5559 -253 -5525
rect -219 -5559 -207 -5525
rect -265 -5593 -207 -5559
rect -265 -5627 -253 -5593
rect -219 -5627 -207 -5593
rect -265 -5661 -207 -5627
rect -265 -5695 -253 -5661
rect -219 -5695 -207 -5661
rect -265 -5729 -207 -5695
rect -265 -5763 -253 -5729
rect -219 -5763 -207 -5729
rect -265 -5797 -207 -5763
rect -265 -5831 -253 -5797
rect -219 -5831 -207 -5797
rect -265 -5865 -207 -5831
rect -265 -5899 -253 -5865
rect -219 -5899 -207 -5865
rect -265 -5933 -207 -5899
rect -265 -5967 -253 -5933
rect -219 -5967 -207 -5933
rect -265 -6000 -207 -5967
rect -147 5967 -89 6000
rect -147 5933 -135 5967
rect -101 5933 -89 5967
rect -147 5899 -89 5933
rect -147 5865 -135 5899
rect -101 5865 -89 5899
rect -147 5831 -89 5865
rect -147 5797 -135 5831
rect -101 5797 -89 5831
rect -147 5763 -89 5797
rect -147 5729 -135 5763
rect -101 5729 -89 5763
rect -147 5695 -89 5729
rect -147 5661 -135 5695
rect -101 5661 -89 5695
rect -147 5627 -89 5661
rect -147 5593 -135 5627
rect -101 5593 -89 5627
rect -147 5559 -89 5593
rect -147 5525 -135 5559
rect -101 5525 -89 5559
rect -147 5491 -89 5525
rect -147 5457 -135 5491
rect -101 5457 -89 5491
rect -147 5423 -89 5457
rect -147 5389 -135 5423
rect -101 5389 -89 5423
rect -147 5355 -89 5389
rect -147 5321 -135 5355
rect -101 5321 -89 5355
rect -147 5287 -89 5321
rect -147 5253 -135 5287
rect -101 5253 -89 5287
rect -147 5219 -89 5253
rect -147 5185 -135 5219
rect -101 5185 -89 5219
rect -147 5151 -89 5185
rect -147 5117 -135 5151
rect -101 5117 -89 5151
rect -147 5083 -89 5117
rect -147 5049 -135 5083
rect -101 5049 -89 5083
rect -147 5015 -89 5049
rect -147 4981 -135 5015
rect -101 4981 -89 5015
rect -147 4947 -89 4981
rect -147 4913 -135 4947
rect -101 4913 -89 4947
rect -147 4879 -89 4913
rect -147 4845 -135 4879
rect -101 4845 -89 4879
rect -147 4811 -89 4845
rect -147 4777 -135 4811
rect -101 4777 -89 4811
rect -147 4743 -89 4777
rect -147 4709 -135 4743
rect -101 4709 -89 4743
rect -147 4675 -89 4709
rect -147 4641 -135 4675
rect -101 4641 -89 4675
rect -147 4607 -89 4641
rect -147 4573 -135 4607
rect -101 4573 -89 4607
rect -147 4539 -89 4573
rect -147 4505 -135 4539
rect -101 4505 -89 4539
rect -147 4471 -89 4505
rect -147 4437 -135 4471
rect -101 4437 -89 4471
rect -147 4403 -89 4437
rect -147 4369 -135 4403
rect -101 4369 -89 4403
rect -147 4335 -89 4369
rect -147 4301 -135 4335
rect -101 4301 -89 4335
rect -147 4267 -89 4301
rect -147 4233 -135 4267
rect -101 4233 -89 4267
rect -147 4199 -89 4233
rect -147 4165 -135 4199
rect -101 4165 -89 4199
rect -147 4131 -89 4165
rect -147 4097 -135 4131
rect -101 4097 -89 4131
rect -147 4063 -89 4097
rect -147 4029 -135 4063
rect -101 4029 -89 4063
rect -147 3995 -89 4029
rect -147 3961 -135 3995
rect -101 3961 -89 3995
rect -147 3927 -89 3961
rect -147 3893 -135 3927
rect -101 3893 -89 3927
rect -147 3859 -89 3893
rect -147 3825 -135 3859
rect -101 3825 -89 3859
rect -147 3791 -89 3825
rect -147 3757 -135 3791
rect -101 3757 -89 3791
rect -147 3723 -89 3757
rect -147 3689 -135 3723
rect -101 3689 -89 3723
rect -147 3655 -89 3689
rect -147 3621 -135 3655
rect -101 3621 -89 3655
rect -147 3587 -89 3621
rect -147 3553 -135 3587
rect -101 3553 -89 3587
rect -147 3519 -89 3553
rect -147 3485 -135 3519
rect -101 3485 -89 3519
rect -147 3451 -89 3485
rect -147 3417 -135 3451
rect -101 3417 -89 3451
rect -147 3383 -89 3417
rect -147 3349 -135 3383
rect -101 3349 -89 3383
rect -147 3315 -89 3349
rect -147 3281 -135 3315
rect -101 3281 -89 3315
rect -147 3247 -89 3281
rect -147 3213 -135 3247
rect -101 3213 -89 3247
rect -147 3179 -89 3213
rect -147 3145 -135 3179
rect -101 3145 -89 3179
rect -147 3111 -89 3145
rect -147 3077 -135 3111
rect -101 3077 -89 3111
rect -147 3043 -89 3077
rect -147 3009 -135 3043
rect -101 3009 -89 3043
rect -147 2975 -89 3009
rect -147 2941 -135 2975
rect -101 2941 -89 2975
rect -147 2907 -89 2941
rect -147 2873 -135 2907
rect -101 2873 -89 2907
rect -147 2839 -89 2873
rect -147 2805 -135 2839
rect -101 2805 -89 2839
rect -147 2771 -89 2805
rect -147 2737 -135 2771
rect -101 2737 -89 2771
rect -147 2703 -89 2737
rect -147 2669 -135 2703
rect -101 2669 -89 2703
rect -147 2635 -89 2669
rect -147 2601 -135 2635
rect -101 2601 -89 2635
rect -147 2567 -89 2601
rect -147 2533 -135 2567
rect -101 2533 -89 2567
rect -147 2499 -89 2533
rect -147 2465 -135 2499
rect -101 2465 -89 2499
rect -147 2431 -89 2465
rect -147 2397 -135 2431
rect -101 2397 -89 2431
rect -147 2363 -89 2397
rect -147 2329 -135 2363
rect -101 2329 -89 2363
rect -147 2295 -89 2329
rect -147 2261 -135 2295
rect -101 2261 -89 2295
rect -147 2227 -89 2261
rect -147 2193 -135 2227
rect -101 2193 -89 2227
rect -147 2159 -89 2193
rect -147 2125 -135 2159
rect -101 2125 -89 2159
rect -147 2091 -89 2125
rect -147 2057 -135 2091
rect -101 2057 -89 2091
rect -147 2023 -89 2057
rect -147 1989 -135 2023
rect -101 1989 -89 2023
rect -147 1955 -89 1989
rect -147 1921 -135 1955
rect -101 1921 -89 1955
rect -147 1887 -89 1921
rect -147 1853 -135 1887
rect -101 1853 -89 1887
rect -147 1819 -89 1853
rect -147 1785 -135 1819
rect -101 1785 -89 1819
rect -147 1751 -89 1785
rect -147 1717 -135 1751
rect -101 1717 -89 1751
rect -147 1683 -89 1717
rect -147 1649 -135 1683
rect -101 1649 -89 1683
rect -147 1615 -89 1649
rect -147 1581 -135 1615
rect -101 1581 -89 1615
rect -147 1547 -89 1581
rect -147 1513 -135 1547
rect -101 1513 -89 1547
rect -147 1479 -89 1513
rect -147 1445 -135 1479
rect -101 1445 -89 1479
rect -147 1411 -89 1445
rect -147 1377 -135 1411
rect -101 1377 -89 1411
rect -147 1343 -89 1377
rect -147 1309 -135 1343
rect -101 1309 -89 1343
rect -147 1275 -89 1309
rect -147 1241 -135 1275
rect -101 1241 -89 1275
rect -147 1207 -89 1241
rect -147 1173 -135 1207
rect -101 1173 -89 1207
rect -147 1139 -89 1173
rect -147 1105 -135 1139
rect -101 1105 -89 1139
rect -147 1071 -89 1105
rect -147 1037 -135 1071
rect -101 1037 -89 1071
rect -147 1003 -89 1037
rect -147 969 -135 1003
rect -101 969 -89 1003
rect -147 935 -89 969
rect -147 901 -135 935
rect -101 901 -89 935
rect -147 867 -89 901
rect -147 833 -135 867
rect -101 833 -89 867
rect -147 799 -89 833
rect -147 765 -135 799
rect -101 765 -89 799
rect -147 731 -89 765
rect -147 697 -135 731
rect -101 697 -89 731
rect -147 663 -89 697
rect -147 629 -135 663
rect -101 629 -89 663
rect -147 595 -89 629
rect -147 561 -135 595
rect -101 561 -89 595
rect -147 527 -89 561
rect -147 493 -135 527
rect -101 493 -89 527
rect -147 459 -89 493
rect -147 425 -135 459
rect -101 425 -89 459
rect -147 391 -89 425
rect -147 357 -135 391
rect -101 357 -89 391
rect -147 323 -89 357
rect -147 289 -135 323
rect -101 289 -89 323
rect -147 255 -89 289
rect -147 221 -135 255
rect -101 221 -89 255
rect -147 187 -89 221
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -221 -89 -187
rect -147 -255 -135 -221
rect -101 -255 -89 -221
rect -147 -289 -89 -255
rect -147 -323 -135 -289
rect -101 -323 -89 -289
rect -147 -357 -89 -323
rect -147 -391 -135 -357
rect -101 -391 -89 -357
rect -147 -425 -89 -391
rect -147 -459 -135 -425
rect -101 -459 -89 -425
rect -147 -493 -89 -459
rect -147 -527 -135 -493
rect -101 -527 -89 -493
rect -147 -561 -89 -527
rect -147 -595 -135 -561
rect -101 -595 -89 -561
rect -147 -629 -89 -595
rect -147 -663 -135 -629
rect -101 -663 -89 -629
rect -147 -697 -89 -663
rect -147 -731 -135 -697
rect -101 -731 -89 -697
rect -147 -765 -89 -731
rect -147 -799 -135 -765
rect -101 -799 -89 -765
rect -147 -833 -89 -799
rect -147 -867 -135 -833
rect -101 -867 -89 -833
rect -147 -901 -89 -867
rect -147 -935 -135 -901
rect -101 -935 -89 -901
rect -147 -969 -89 -935
rect -147 -1003 -135 -969
rect -101 -1003 -89 -969
rect -147 -1037 -89 -1003
rect -147 -1071 -135 -1037
rect -101 -1071 -89 -1037
rect -147 -1105 -89 -1071
rect -147 -1139 -135 -1105
rect -101 -1139 -89 -1105
rect -147 -1173 -89 -1139
rect -147 -1207 -135 -1173
rect -101 -1207 -89 -1173
rect -147 -1241 -89 -1207
rect -147 -1275 -135 -1241
rect -101 -1275 -89 -1241
rect -147 -1309 -89 -1275
rect -147 -1343 -135 -1309
rect -101 -1343 -89 -1309
rect -147 -1377 -89 -1343
rect -147 -1411 -135 -1377
rect -101 -1411 -89 -1377
rect -147 -1445 -89 -1411
rect -147 -1479 -135 -1445
rect -101 -1479 -89 -1445
rect -147 -1513 -89 -1479
rect -147 -1547 -135 -1513
rect -101 -1547 -89 -1513
rect -147 -1581 -89 -1547
rect -147 -1615 -135 -1581
rect -101 -1615 -89 -1581
rect -147 -1649 -89 -1615
rect -147 -1683 -135 -1649
rect -101 -1683 -89 -1649
rect -147 -1717 -89 -1683
rect -147 -1751 -135 -1717
rect -101 -1751 -89 -1717
rect -147 -1785 -89 -1751
rect -147 -1819 -135 -1785
rect -101 -1819 -89 -1785
rect -147 -1853 -89 -1819
rect -147 -1887 -135 -1853
rect -101 -1887 -89 -1853
rect -147 -1921 -89 -1887
rect -147 -1955 -135 -1921
rect -101 -1955 -89 -1921
rect -147 -1989 -89 -1955
rect -147 -2023 -135 -1989
rect -101 -2023 -89 -1989
rect -147 -2057 -89 -2023
rect -147 -2091 -135 -2057
rect -101 -2091 -89 -2057
rect -147 -2125 -89 -2091
rect -147 -2159 -135 -2125
rect -101 -2159 -89 -2125
rect -147 -2193 -89 -2159
rect -147 -2227 -135 -2193
rect -101 -2227 -89 -2193
rect -147 -2261 -89 -2227
rect -147 -2295 -135 -2261
rect -101 -2295 -89 -2261
rect -147 -2329 -89 -2295
rect -147 -2363 -135 -2329
rect -101 -2363 -89 -2329
rect -147 -2397 -89 -2363
rect -147 -2431 -135 -2397
rect -101 -2431 -89 -2397
rect -147 -2465 -89 -2431
rect -147 -2499 -135 -2465
rect -101 -2499 -89 -2465
rect -147 -2533 -89 -2499
rect -147 -2567 -135 -2533
rect -101 -2567 -89 -2533
rect -147 -2601 -89 -2567
rect -147 -2635 -135 -2601
rect -101 -2635 -89 -2601
rect -147 -2669 -89 -2635
rect -147 -2703 -135 -2669
rect -101 -2703 -89 -2669
rect -147 -2737 -89 -2703
rect -147 -2771 -135 -2737
rect -101 -2771 -89 -2737
rect -147 -2805 -89 -2771
rect -147 -2839 -135 -2805
rect -101 -2839 -89 -2805
rect -147 -2873 -89 -2839
rect -147 -2907 -135 -2873
rect -101 -2907 -89 -2873
rect -147 -2941 -89 -2907
rect -147 -2975 -135 -2941
rect -101 -2975 -89 -2941
rect -147 -3009 -89 -2975
rect -147 -3043 -135 -3009
rect -101 -3043 -89 -3009
rect -147 -3077 -89 -3043
rect -147 -3111 -135 -3077
rect -101 -3111 -89 -3077
rect -147 -3145 -89 -3111
rect -147 -3179 -135 -3145
rect -101 -3179 -89 -3145
rect -147 -3213 -89 -3179
rect -147 -3247 -135 -3213
rect -101 -3247 -89 -3213
rect -147 -3281 -89 -3247
rect -147 -3315 -135 -3281
rect -101 -3315 -89 -3281
rect -147 -3349 -89 -3315
rect -147 -3383 -135 -3349
rect -101 -3383 -89 -3349
rect -147 -3417 -89 -3383
rect -147 -3451 -135 -3417
rect -101 -3451 -89 -3417
rect -147 -3485 -89 -3451
rect -147 -3519 -135 -3485
rect -101 -3519 -89 -3485
rect -147 -3553 -89 -3519
rect -147 -3587 -135 -3553
rect -101 -3587 -89 -3553
rect -147 -3621 -89 -3587
rect -147 -3655 -135 -3621
rect -101 -3655 -89 -3621
rect -147 -3689 -89 -3655
rect -147 -3723 -135 -3689
rect -101 -3723 -89 -3689
rect -147 -3757 -89 -3723
rect -147 -3791 -135 -3757
rect -101 -3791 -89 -3757
rect -147 -3825 -89 -3791
rect -147 -3859 -135 -3825
rect -101 -3859 -89 -3825
rect -147 -3893 -89 -3859
rect -147 -3927 -135 -3893
rect -101 -3927 -89 -3893
rect -147 -3961 -89 -3927
rect -147 -3995 -135 -3961
rect -101 -3995 -89 -3961
rect -147 -4029 -89 -3995
rect -147 -4063 -135 -4029
rect -101 -4063 -89 -4029
rect -147 -4097 -89 -4063
rect -147 -4131 -135 -4097
rect -101 -4131 -89 -4097
rect -147 -4165 -89 -4131
rect -147 -4199 -135 -4165
rect -101 -4199 -89 -4165
rect -147 -4233 -89 -4199
rect -147 -4267 -135 -4233
rect -101 -4267 -89 -4233
rect -147 -4301 -89 -4267
rect -147 -4335 -135 -4301
rect -101 -4335 -89 -4301
rect -147 -4369 -89 -4335
rect -147 -4403 -135 -4369
rect -101 -4403 -89 -4369
rect -147 -4437 -89 -4403
rect -147 -4471 -135 -4437
rect -101 -4471 -89 -4437
rect -147 -4505 -89 -4471
rect -147 -4539 -135 -4505
rect -101 -4539 -89 -4505
rect -147 -4573 -89 -4539
rect -147 -4607 -135 -4573
rect -101 -4607 -89 -4573
rect -147 -4641 -89 -4607
rect -147 -4675 -135 -4641
rect -101 -4675 -89 -4641
rect -147 -4709 -89 -4675
rect -147 -4743 -135 -4709
rect -101 -4743 -89 -4709
rect -147 -4777 -89 -4743
rect -147 -4811 -135 -4777
rect -101 -4811 -89 -4777
rect -147 -4845 -89 -4811
rect -147 -4879 -135 -4845
rect -101 -4879 -89 -4845
rect -147 -4913 -89 -4879
rect -147 -4947 -135 -4913
rect -101 -4947 -89 -4913
rect -147 -4981 -89 -4947
rect -147 -5015 -135 -4981
rect -101 -5015 -89 -4981
rect -147 -5049 -89 -5015
rect -147 -5083 -135 -5049
rect -101 -5083 -89 -5049
rect -147 -5117 -89 -5083
rect -147 -5151 -135 -5117
rect -101 -5151 -89 -5117
rect -147 -5185 -89 -5151
rect -147 -5219 -135 -5185
rect -101 -5219 -89 -5185
rect -147 -5253 -89 -5219
rect -147 -5287 -135 -5253
rect -101 -5287 -89 -5253
rect -147 -5321 -89 -5287
rect -147 -5355 -135 -5321
rect -101 -5355 -89 -5321
rect -147 -5389 -89 -5355
rect -147 -5423 -135 -5389
rect -101 -5423 -89 -5389
rect -147 -5457 -89 -5423
rect -147 -5491 -135 -5457
rect -101 -5491 -89 -5457
rect -147 -5525 -89 -5491
rect -147 -5559 -135 -5525
rect -101 -5559 -89 -5525
rect -147 -5593 -89 -5559
rect -147 -5627 -135 -5593
rect -101 -5627 -89 -5593
rect -147 -5661 -89 -5627
rect -147 -5695 -135 -5661
rect -101 -5695 -89 -5661
rect -147 -5729 -89 -5695
rect -147 -5763 -135 -5729
rect -101 -5763 -89 -5729
rect -147 -5797 -89 -5763
rect -147 -5831 -135 -5797
rect -101 -5831 -89 -5797
rect -147 -5865 -89 -5831
rect -147 -5899 -135 -5865
rect -101 -5899 -89 -5865
rect -147 -5933 -89 -5899
rect -147 -5967 -135 -5933
rect -101 -5967 -89 -5933
rect -147 -6000 -89 -5967
rect -29 5967 29 6000
rect -29 5933 -17 5967
rect 17 5933 29 5967
rect -29 5899 29 5933
rect -29 5865 -17 5899
rect 17 5865 29 5899
rect -29 5831 29 5865
rect -29 5797 -17 5831
rect 17 5797 29 5831
rect -29 5763 29 5797
rect -29 5729 -17 5763
rect 17 5729 29 5763
rect -29 5695 29 5729
rect -29 5661 -17 5695
rect 17 5661 29 5695
rect -29 5627 29 5661
rect -29 5593 -17 5627
rect 17 5593 29 5627
rect -29 5559 29 5593
rect -29 5525 -17 5559
rect 17 5525 29 5559
rect -29 5491 29 5525
rect -29 5457 -17 5491
rect 17 5457 29 5491
rect -29 5423 29 5457
rect -29 5389 -17 5423
rect 17 5389 29 5423
rect -29 5355 29 5389
rect -29 5321 -17 5355
rect 17 5321 29 5355
rect -29 5287 29 5321
rect -29 5253 -17 5287
rect 17 5253 29 5287
rect -29 5219 29 5253
rect -29 5185 -17 5219
rect 17 5185 29 5219
rect -29 5151 29 5185
rect -29 5117 -17 5151
rect 17 5117 29 5151
rect -29 5083 29 5117
rect -29 5049 -17 5083
rect 17 5049 29 5083
rect -29 5015 29 5049
rect -29 4981 -17 5015
rect 17 4981 29 5015
rect -29 4947 29 4981
rect -29 4913 -17 4947
rect 17 4913 29 4947
rect -29 4879 29 4913
rect -29 4845 -17 4879
rect 17 4845 29 4879
rect -29 4811 29 4845
rect -29 4777 -17 4811
rect 17 4777 29 4811
rect -29 4743 29 4777
rect -29 4709 -17 4743
rect 17 4709 29 4743
rect -29 4675 29 4709
rect -29 4641 -17 4675
rect 17 4641 29 4675
rect -29 4607 29 4641
rect -29 4573 -17 4607
rect 17 4573 29 4607
rect -29 4539 29 4573
rect -29 4505 -17 4539
rect 17 4505 29 4539
rect -29 4471 29 4505
rect -29 4437 -17 4471
rect 17 4437 29 4471
rect -29 4403 29 4437
rect -29 4369 -17 4403
rect 17 4369 29 4403
rect -29 4335 29 4369
rect -29 4301 -17 4335
rect 17 4301 29 4335
rect -29 4267 29 4301
rect -29 4233 -17 4267
rect 17 4233 29 4267
rect -29 4199 29 4233
rect -29 4165 -17 4199
rect 17 4165 29 4199
rect -29 4131 29 4165
rect -29 4097 -17 4131
rect 17 4097 29 4131
rect -29 4063 29 4097
rect -29 4029 -17 4063
rect 17 4029 29 4063
rect -29 3995 29 4029
rect -29 3961 -17 3995
rect 17 3961 29 3995
rect -29 3927 29 3961
rect -29 3893 -17 3927
rect 17 3893 29 3927
rect -29 3859 29 3893
rect -29 3825 -17 3859
rect 17 3825 29 3859
rect -29 3791 29 3825
rect -29 3757 -17 3791
rect 17 3757 29 3791
rect -29 3723 29 3757
rect -29 3689 -17 3723
rect 17 3689 29 3723
rect -29 3655 29 3689
rect -29 3621 -17 3655
rect 17 3621 29 3655
rect -29 3587 29 3621
rect -29 3553 -17 3587
rect 17 3553 29 3587
rect -29 3519 29 3553
rect -29 3485 -17 3519
rect 17 3485 29 3519
rect -29 3451 29 3485
rect -29 3417 -17 3451
rect 17 3417 29 3451
rect -29 3383 29 3417
rect -29 3349 -17 3383
rect 17 3349 29 3383
rect -29 3315 29 3349
rect -29 3281 -17 3315
rect 17 3281 29 3315
rect -29 3247 29 3281
rect -29 3213 -17 3247
rect 17 3213 29 3247
rect -29 3179 29 3213
rect -29 3145 -17 3179
rect 17 3145 29 3179
rect -29 3111 29 3145
rect -29 3077 -17 3111
rect 17 3077 29 3111
rect -29 3043 29 3077
rect -29 3009 -17 3043
rect 17 3009 29 3043
rect -29 2975 29 3009
rect -29 2941 -17 2975
rect 17 2941 29 2975
rect -29 2907 29 2941
rect -29 2873 -17 2907
rect 17 2873 29 2907
rect -29 2839 29 2873
rect -29 2805 -17 2839
rect 17 2805 29 2839
rect -29 2771 29 2805
rect -29 2737 -17 2771
rect 17 2737 29 2771
rect -29 2703 29 2737
rect -29 2669 -17 2703
rect 17 2669 29 2703
rect -29 2635 29 2669
rect -29 2601 -17 2635
rect 17 2601 29 2635
rect -29 2567 29 2601
rect -29 2533 -17 2567
rect 17 2533 29 2567
rect -29 2499 29 2533
rect -29 2465 -17 2499
rect 17 2465 29 2499
rect -29 2431 29 2465
rect -29 2397 -17 2431
rect 17 2397 29 2431
rect -29 2363 29 2397
rect -29 2329 -17 2363
rect 17 2329 29 2363
rect -29 2295 29 2329
rect -29 2261 -17 2295
rect 17 2261 29 2295
rect -29 2227 29 2261
rect -29 2193 -17 2227
rect 17 2193 29 2227
rect -29 2159 29 2193
rect -29 2125 -17 2159
rect 17 2125 29 2159
rect -29 2091 29 2125
rect -29 2057 -17 2091
rect 17 2057 29 2091
rect -29 2023 29 2057
rect -29 1989 -17 2023
rect 17 1989 29 2023
rect -29 1955 29 1989
rect -29 1921 -17 1955
rect 17 1921 29 1955
rect -29 1887 29 1921
rect -29 1853 -17 1887
rect 17 1853 29 1887
rect -29 1819 29 1853
rect -29 1785 -17 1819
rect 17 1785 29 1819
rect -29 1751 29 1785
rect -29 1717 -17 1751
rect 17 1717 29 1751
rect -29 1683 29 1717
rect -29 1649 -17 1683
rect 17 1649 29 1683
rect -29 1615 29 1649
rect -29 1581 -17 1615
rect 17 1581 29 1615
rect -29 1547 29 1581
rect -29 1513 -17 1547
rect 17 1513 29 1547
rect -29 1479 29 1513
rect -29 1445 -17 1479
rect 17 1445 29 1479
rect -29 1411 29 1445
rect -29 1377 -17 1411
rect 17 1377 29 1411
rect -29 1343 29 1377
rect -29 1309 -17 1343
rect 17 1309 29 1343
rect -29 1275 29 1309
rect -29 1241 -17 1275
rect 17 1241 29 1275
rect -29 1207 29 1241
rect -29 1173 -17 1207
rect 17 1173 29 1207
rect -29 1139 29 1173
rect -29 1105 -17 1139
rect 17 1105 29 1139
rect -29 1071 29 1105
rect -29 1037 -17 1071
rect 17 1037 29 1071
rect -29 1003 29 1037
rect -29 969 -17 1003
rect 17 969 29 1003
rect -29 935 29 969
rect -29 901 -17 935
rect 17 901 29 935
rect -29 867 29 901
rect -29 833 -17 867
rect 17 833 29 867
rect -29 799 29 833
rect -29 765 -17 799
rect 17 765 29 799
rect -29 731 29 765
rect -29 697 -17 731
rect 17 697 29 731
rect -29 663 29 697
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -697 29 -663
rect -29 -731 -17 -697
rect 17 -731 29 -697
rect -29 -765 29 -731
rect -29 -799 -17 -765
rect 17 -799 29 -765
rect -29 -833 29 -799
rect -29 -867 -17 -833
rect 17 -867 29 -833
rect -29 -901 29 -867
rect -29 -935 -17 -901
rect 17 -935 29 -901
rect -29 -969 29 -935
rect -29 -1003 -17 -969
rect 17 -1003 29 -969
rect -29 -1037 29 -1003
rect -29 -1071 -17 -1037
rect 17 -1071 29 -1037
rect -29 -1105 29 -1071
rect -29 -1139 -17 -1105
rect 17 -1139 29 -1105
rect -29 -1173 29 -1139
rect -29 -1207 -17 -1173
rect 17 -1207 29 -1173
rect -29 -1241 29 -1207
rect -29 -1275 -17 -1241
rect 17 -1275 29 -1241
rect -29 -1309 29 -1275
rect -29 -1343 -17 -1309
rect 17 -1343 29 -1309
rect -29 -1377 29 -1343
rect -29 -1411 -17 -1377
rect 17 -1411 29 -1377
rect -29 -1445 29 -1411
rect -29 -1479 -17 -1445
rect 17 -1479 29 -1445
rect -29 -1513 29 -1479
rect -29 -1547 -17 -1513
rect 17 -1547 29 -1513
rect -29 -1581 29 -1547
rect -29 -1615 -17 -1581
rect 17 -1615 29 -1581
rect -29 -1649 29 -1615
rect -29 -1683 -17 -1649
rect 17 -1683 29 -1649
rect -29 -1717 29 -1683
rect -29 -1751 -17 -1717
rect 17 -1751 29 -1717
rect -29 -1785 29 -1751
rect -29 -1819 -17 -1785
rect 17 -1819 29 -1785
rect -29 -1853 29 -1819
rect -29 -1887 -17 -1853
rect 17 -1887 29 -1853
rect -29 -1921 29 -1887
rect -29 -1955 -17 -1921
rect 17 -1955 29 -1921
rect -29 -1989 29 -1955
rect -29 -2023 -17 -1989
rect 17 -2023 29 -1989
rect -29 -2057 29 -2023
rect -29 -2091 -17 -2057
rect 17 -2091 29 -2057
rect -29 -2125 29 -2091
rect -29 -2159 -17 -2125
rect 17 -2159 29 -2125
rect -29 -2193 29 -2159
rect -29 -2227 -17 -2193
rect 17 -2227 29 -2193
rect -29 -2261 29 -2227
rect -29 -2295 -17 -2261
rect 17 -2295 29 -2261
rect -29 -2329 29 -2295
rect -29 -2363 -17 -2329
rect 17 -2363 29 -2329
rect -29 -2397 29 -2363
rect -29 -2431 -17 -2397
rect 17 -2431 29 -2397
rect -29 -2465 29 -2431
rect -29 -2499 -17 -2465
rect 17 -2499 29 -2465
rect -29 -2533 29 -2499
rect -29 -2567 -17 -2533
rect 17 -2567 29 -2533
rect -29 -2601 29 -2567
rect -29 -2635 -17 -2601
rect 17 -2635 29 -2601
rect -29 -2669 29 -2635
rect -29 -2703 -17 -2669
rect 17 -2703 29 -2669
rect -29 -2737 29 -2703
rect -29 -2771 -17 -2737
rect 17 -2771 29 -2737
rect -29 -2805 29 -2771
rect -29 -2839 -17 -2805
rect 17 -2839 29 -2805
rect -29 -2873 29 -2839
rect -29 -2907 -17 -2873
rect 17 -2907 29 -2873
rect -29 -2941 29 -2907
rect -29 -2975 -17 -2941
rect 17 -2975 29 -2941
rect -29 -3009 29 -2975
rect -29 -3043 -17 -3009
rect 17 -3043 29 -3009
rect -29 -3077 29 -3043
rect -29 -3111 -17 -3077
rect 17 -3111 29 -3077
rect -29 -3145 29 -3111
rect -29 -3179 -17 -3145
rect 17 -3179 29 -3145
rect -29 -3213 29 -3179
rect -29 -3247 -17 -3213
rect 17 -3247 29 -3213
rect -29 -3281 29 -3247
rect -29 -3315 -17 -3281
rect 17 -3315 29 -3281
rect -29 -3349 29 -3315
rect -29 -3383 -17 -3349
rect 17 -3383 29 -3349
rect -29 -3417 29 -3383
rect -29 -3451 -17 -3417
rect 17 -3451 29 -3417
rect -29 -3485 29 -3451
rect -29 -3519 -17 -3485
rect 17 -3519 29 -3485
rect -29 -3553 29 -3519
rect -29 -3587 -17 -3553
rect 17 -3587 29 -3553
rect -29 -3621 29 -3587
rect -29 -3655 -17 -3621
rect 17 -3655 29 -3621
rect -29 -3689 29 -3655
rect -29 -3723 -17 -3689
rect 17 -3723 29 -3689
rect -29 -3757 29 -3723
rect -29 -3791 -17 -3757
rect 17 -3791 29 -3757
rect -29 -3825 29 -3791
rect -29 -3859 -17 -3825
rect 17 -3859 29 -3825
rect -29 -3893 29 -3859
rect -29 -3927 -17 -3893
rect 17 -3927 29 -3893
rect -29 -3961 29 -3927
rect -29 -3995 -17 -3961
rect 17 -3995 29 -3961
rect -29 -4029 29 -3995
rect -29 -4063 -17 -4029
rect 17 -4063 29 -4029
rect -29 -4097 29 -4063
rect -29 -4131 -17 -4097
rect 17 -4131 29 -4097
rect -29 -4165 29 -4131
rect -29 -4199 -17 -4165
rect 17 -4199 29 -4165
rect -29 -4233 29 -4199
rect -29 -4267 -17 -4233
rect 17 -4267 29 -4233
rect -29 -4301 29 -4267
rect -29 -4335 -17 -4301
rect 17 -4335 29 -4301
rect -29 -4369 29 -4335
rect -29 -4403 -17 -4369
rect 17 -4403 29 -4369
rect -29 -4437 29 -4403
rect -29 -4471 -17 -4437
rect 17 -4471 29 -4437
rect -29 -4505 29 -4471
rect -29 -4539 -17 -4505
rect 17 -4539 29 -4505
rect -29 -4573 29 -4539
rect -29 -4607 -17 -4573
rect 17 -4607 29 -4573
rect -29 -4641 29 -4607
rect -29 -4675 -17 -4641
rect 17 -4675 29 -4641
rect -29 -4709 29 -4675
rect -29 -4743 -17 -4709
rect 17 -4743 29 -4709
rect -29 -4777 29 -4743
rect -29 -4811 -17 -4777
rect 17 -4811 29 -4777
rect -29 -4845 29 -4811
rect -29 -4879 -17 -4845
rect 17 -4879 29 -4845
rect -29 -4913 29 -4879
rect -29 -4947 -17 -4913
rect 17 -4947 29 -4913
rect -29 -4981 29 -4947
rect -29 -5015 -17 -4981
rect 17 -5015 29 -4981
rect -29 -5049 29 -5015
rect -29 -5083 -17 -5049
rect 17 -5083 29 -5049
rect -29 -5117 29 -5083
rect -29 -5151 -17 -5117
rect 17 -5151 29 -5117
rect -29 -5185 29 -5151
rect -29 -5219 -17 -5185
rect 17 -5219 29 -5185
rect -29 -5253 29 -5219
rect -29 -5287 -17 -5253
rect 17 -5287 29 -5253
rect -29 -5321 29 -5287
rect -29 -5355 -17 -5321
rect 17 -5355 29 -5321
rect -29 -5389 29 -5355
rect -29 -5423 -17 -5389
rect 17 -5423 29 -5389
rect -29 -5457 29 -5423
rect -29 -5491 -17 -5457
rect 17 -5491 29 -5457
rect -29 -5525 29 -5491
rect -29 -5559 -17 -5525
rect 17 -5559 29 -5525
rect -29 -5593 29 -5559
rect -29 -5627 -17 -5593
rect 17 -5627 29 -5593
rect -29 -5661 29 -5627
rect -29 -5695 -17 -5661
rect 17 -5695 29 -5661
rect -29 -5729 29 -5695
rect -29 -5763 -17 -5729
rect 17 -5763 29 -5729
rect -29 -5797 29 -5763
rect -29 -5831 -17 -5797
rect 17 -5831 29 -5797
rect -29 -5865 29 -5831
rect -29 -5899 -17 -5865
rect 17 -5899 29 -5865
rect -29 -5933 29 -5899
rect -29 -5967 -17 -5933
rect 17 -5967 29 -5933
rect -29 -6000 29 -5967
rect 89 5967 147 6000
rect 89 5933 101 5967
rect 135 5933 147 5967
rect 89 5899 147 5933
rect 89 5865 101 5899
rect 135 5865 147 5899
rect 89 5831 147 5865
rect 89 5797 101 5831
rect 135 5797 147 5831
rect 89 5763 147 5797
rect 89 5729 101 5763
rect 135 5729 147 5763
rect 89 5695 147 5729
rect 89 5661 101 5695
rect 135 5661 147 5695
rect 89 5627 147 5661
rect 89 5593 101 5627
rect 135 5593 147 5627
rect 89 5559 147 5593
rect 89 5525 101 5559
rect 135 5525 147 5559
rect 89 5491 147 5525
rect 89 5457 101 5491
rect 135 5457 147 5491
rect 89 5423 147 5457
rect 89 5389 101 5423
rect 135 5389 147 5423
rect 89 5355 147 5389
rect 89 5321 101 5355
rect 135 5321 147 5355
rect 89 5287 147 5321
rect 89 5253 101 5287
rect 135 5253 147 5287
rect 89 5219 147 5253
rect 89 5185 101 5219
rect 135 5185 147 5219
rect 89 5151 147 5185
rect 89 5117 101 5151
rect 135 5117 147 5151
rect 89 5083 147 5117
rect 89 5049 101 5083
rect 135 5049 147 5083
rect 89 5015 147 5049
rect 89 4981 101 5015
rect 135 4981 147 5015
rect 89 4947 147 4981
rect 89 4913 101 4947
rect 135 4913 147 4947
rect 89 4879 147 4913
rect 89 4845 101 4879
rect 135 4845 147 4879
rect 89 4811 147 4845
rect 89 4777 101 4811
rect 135 4777 147 4811
rect 89 4743 147 4777
rect 89 4709 101 4743
rect 135 4709 147 4743
rect 89 4675 147 4709
rect 89 4641 101 4675
rect 135 4641 147 4675
rect 89 4607 147 4641
rect 89 4573 101 4607
rect 135 4573 147 4607
rect 89 4539 147 4573
rect 89 4505 101 4539
rect 135 4505 147 4539
rect 89 4471 147 4505
rect 89 4437 101 4471
rect 135 4437 147 4471
rect 89 4403 147 4437
rect 89 4369 101 4403
rect 135 4369 147 4403
rect 89 4335 147 4369
rect 89 4301 101 4335
rect 135 4301 147 4335
rect 89 4267 147 4301
rect 89 4233 101 4267
rect 135 4233 147 4267
rect 89 4199 147 4233
rect 89 4165 101 4199
rect 135 4165 147 4199
rect 89 4131 147 4165
rect 89 4097 101 4131
rect 135 4097 147 4131
rect 89 4063 147 4097
rect 89 4029 101 4063
rect 135 4029 147 4063
rect 89 3995 147 4029
rect 89 3961 101 3995
rect 135 3961 147 3995
rect 89 3927 147 3961
rect 89 3893 101 3927
rect 135 3893 147 3927
rect 89 3859 147 3893
rect 89 3825 101 3859
rect 135 3825 147 3859
rect 89 3791 147 3825
rect 89 3757 101 3791
rect 135 3757 147 3791
rect 89 3723 147 3757
rect 89 3689 101 3723
rect 135 3689 147 3723
rect 89 3655 147 3689
rect 89 3621 101 3655
rect 135 3621 147 3655
rect 89 3587 147 3621
rect 89 3553 101 3587
rect 135 3553 147 3587
rect 89 3519 147 3553
rect 89 3485 101 3519
rect 135 3485 147 3519
rect 89 3451 147 3485
rect 89 3417 101 3451
rect 135 3417 147 3451
rect 89 3383 147 3417
rect 89 3349 101 3383
rect 135 3349 147 3383
rect 89 3315 147 3349
rect 89 3281 101 3315
rect 135 3281 147 3315
rect 89 3247 147 3281
rect 89 3213 101 3247
rect 135 3213 147 3247
rect 89 3179 147 3213
rect 89 3145 101 3179
rect 135 3145 147 3179
rect 89 3111 147 3145
rect 89 3077 101 3111
rect 135 3077 147 3111
rect 89 3043 147 3077
rect 89 3009 101 3043
rect 135 3009 147 3043
rect 89 2975 147 3009
rect 89 2941 101 2975
rect 135 2941 147 2975
rect 89 2907 147 2941
rect 89 2873 101 2907
rect 135 2873 147 2907
rect 89 2839 147 2873
rect 89 2805 101 2839
rect 135 2805 147 2839
rect 89 2771 147 2805
rect 89 2737 101 2771
rect 135 2737 147 2771
rect 89 2703 147 2737
rect 89 2669 101 2703
rect 135 2669 147 2703
rect 89 2635 147 2669
rect 89 2601 101 2635
rect 135 2601 147 2635
rect 89 2567 147 2601
rect 89 2533 101 2567
rect 135 2533 147 2567
rect 89 2499 147 2533
rect 89 2465 101 2499
rect 135 2465 147 2499
rect 89 2431 147 2465
rect 89 2397 101 2431
rect 135 2397 147 2431
rect 89 2363 147 2397
rect 89 2329 101 2363
rect 135 2329 147 2363
rect 89 2295 147 2329
rect 89 2261 101 2295
rect 135 2261 147 2295
rect 89 2227 147 2261
rect 89 2193 101 2227
rect 135 2193 147 2227
rect 89 2159 147 2193
rect 89 2125 101 2159
rect 135 2125 147 2159
rect 89 2091 147 2125
rect 89 2057 101 2091
rect 135 2057 147 2091
rect 89 2023 147 2057
rect 89 1989 101 2023
rect 135 1989 147 2023
rect 89 1955 147 1989
rect 89 1921 101 1955
rect 135 1921 147 1955
rect 89 1887 147 1921
rect 89 1853 101 1887
rect 135 1853 147 1887
rect 89 1819 147 1853
rect 89 1785 101 1819
rect 135 1785 147 1819
rect 89 1751 147 1785
rect 89 1717 101 1751
rect 135 1717 147 1751
rect 89 1683 147 1717
rect 89 1649 101 1683
rect 135 1649 147 1683
rect 89 1615 147 1649
rect 89 1581 101 1615
rect 135 1581 147 1615
rect 89 1547 147 1581
rect 89 1513 101 1547
rect 135 1513 147 1547
rect 89 1479 147 1513
rect 89 1445 101 1479
rect 135 1445 147 1479
rect 89 1411 147 1445
rect 89 1377 101 1411
rect 135 1377 147 1411
rect 89 1343 147 1377
rect 89 1309 101 1343
rect 135 1309 147 1343
rect 89 1275 147 1309
rect 89 1241 101 1275
rect 135 1241 147 1275
rect 89 1207 147 1241
rect 89 1173 101 1207
rect 135 1173 147 1207
rect 89 1139 147 1173
rect 89 1105 101 1139
rect 135 1105 147 1139
rect 89 1071 147 1105
rect 89 1037 101 1071
rect 135 1037 147 1071
rect 89 1003 147 1037
rect 89 969 101 1003
rect 135 969 147 1003
rect 89 935 147 969
rect 89 901 101 935
rect 135 901 147 935
rect 89 867 147 901
rect 89 833 101 867
rect 135 833 147 867
rect 89 799 147 833
rect 89 765 101 799
rect 135 765 147 799
rect 89 731 147 765
rect 89 697 101 731
rect 135 697 147 731
rect 89 663 147 697
rect 89 629 101 663
rect 135 629 147 663
rect 89 595 147 629
rect 89 561 101 595
rect 135 561 147 595
rect 89 527 147 561
rect 89 493 101 527
rect 135 493 147 527
rect 89 459 147 493
rect 89 425 101 459
rect 135 425 147 459
rect 89 391 147 425
rect 89 357 101 391
rect 135 357 147 391
rect 89 323 147 357
rect 89 289 101 323
rect 135 289 147 323
rect 89 255 147 289
rect 89 221 101 255
rect 135 221 147 255
rect 89 187 147 221
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -221 147 -187
rect 89 -255 101 -221
rect 135 -255 147 -221
rect 89 -289 147 -255
rect 89 -323 101 -289
rect 135 -323 147 -289
rect 89 -357 147 -323
rect 89 -391 101 -357
rect 135 -391 147 -357
rect 89 -425 147 -391
rect 89 -459 101 -425
rect 135 -459 147 -425
rect 89 -493 147 -459
rect 89 -527 101 -493
rect 135 -527 147 -493
rect 89 -561 147 -527
rect 89 -595 101 -561
rect 135 -595 147 -561
rect 89 -629 147 -595
rect 89 -663 101 -629
rect 135 -663 147 -629
rect 89 -697 147 -663
rect 89 -731 101 -697
rect 135 -731 147 -697
rect 89 -765 147 -731
rect 89 -799 101 -765
rect 135 -799 147 -765
rect 89 -833 147 -799
rect 89 -867 101 -833
rect 135 -867 147 -833
rect 89 -901 147 -867
rect 89 -935 101 -901
rect 135 -935 147 -901
rect 89 -969 147 -935
rect 89 -1003 101 -969
rect 135 -1003 147 -969
rect 89 -1037 147 -1003
rect 89 -1071 101 -1037
rect 135 -1071 147 -1037
rect 89 -1105 147 -1071
rect 89 -1139 101 -1105
rect 135 -1139 147 -1105
rect 89 -1173 147 -1139
rect 89 -1207 101 -1173
rect 135 -1207 147 -1173
rect 89 -1241 147 -1207
rect 89 -1275 101 -1241
rect 135 -1275 147 -1241
rect 89 -1309 147 -1275
rect 89 -1343 101 -1309
rect 135 -1343 147 -1309
rect 89 -1377 147 -1343
rect 89 -1411 101 -1377
rect 135 -1411 147 -1377
rect 89 -1445 147 -1411
rect 89 -1479 101 -1445
rect 135 -1479 147 -1445
rect 89 -1513 147 -1479
rect 89 -1547 101 -1513
rect 135 -1547 147 -1513
rect 89 -1581 147 -1547
rect 89 -1615 101 -1581
rect 135 -1615 147 -1581
rect 89 -1649 147 -1615
rect 89 -1683 101 -1649
rect 135 -1683 147 -1649
rect 89 -1717 147 -1683
rect 89 -1751 101 -1717
rect 135 -1751 147 -1717
rect 89 -1785 147 -1751
rect 89 -1819 101 -1785
rect 135 -1819 147 -1785
rect 89 -1853 147 -1819
rect 89 -1887 101 -1853
rect 135 -1887 147 -1853
rect 89 -1921 147 -1887
rect 89 -1955 101 -1921
rect 135 -1955 147 -1921
rect 89 -1989 147 -1955
rect 89 -2023 101 -1989
rect 135 -2023 147 -1989
rect 89 -2057 147 -2023
rect 89 -2091 101 -2057
rect 135 -2091 147 -2057
rect 89 -2125 147 -2091
rect 89 -2159 101 -2125
rect 135 -2159 147 -2125
rect 89 -2193 147 -2159
rect 89 -2227 101 -2193
rect 135 -2227 147 -2193
rect 89 -2261 147 -2227
rect 89 -2295 101 -2261
rect 135 -2295 147 -2261
rect 89 -2329 147 -2295
rect 89 -2363 101 -2329
rect 135 -2363 147 -2329
rect 89 -2397 147 -2363
rect 89 -2431 101 -2397
rect 135 -2431 147 -2397
rect 89 -2465 147 -2431
rect 89 -2499 101 -2465
rect 135 -2499 147 -2465
rect 89 -2533 147 -2499
rect 89 -2567 101 -2533
rect 135 -2567 147 -2533
rect 89 -2601 147 -2567
rect 89 -2635 101 -2601
rect 135 -2635 147 -2601
rect 89 -2669 147 -2635
rect 89 -2703 101 -2669
rect 135 -2703 147 -2669
rect 89 -2737 147 -2703
rect 89 -2771 101 -2737
rect 135 -2771 147 -2737
rect 89 -2805 147 -2771
rect 89 -2839 101 -2805
rect 135 -2839 147 -2805
rect 89 -2873 147 -2839
rect 89 -2907 101 -2873
rect 135 -2907 147 -2873
rect 89 -2941 147 -2907
rect 89 -2975 101 -2941
rect 135 -2975 147 -2941
rect 89 -3009 147 -2975
rect 89 -3043 101 -3009
rect 135 -3043 147 -3009
rect 89 -3077 147 -3043
rect 89 -3111 101 -3077
rect 135 -3111 147 -3077
rect 89 -3145 147 -3111
rect 89 -3179 101 -3145
rect 135 -3179 147 -3145
rect 89 -3213 147 -3179
rect 89 -3247 101 -3213
rect 135 -3247 147 -3213
rect 89 -3281 147 -3247
rect 89 -3315 101 -3281
rect 135 -3315 147 -3281
rect 89 -3349 147 -3315
rect 89 -3383 101 -3349
rect 135 -3383 147 -3349
rect 89 -3417 147 -3383
rect 89 -3451 101 -3417
rect 135 -3451 147 -3417
rect 89 -3485 147 -3451
rect 89 -3519 101 -3485
rect 135 -3519 147 -3485
rect 89 -3553 147 -3519
rect 89 -3587 101 -3553
rect 135 -3587 147 -3553
rect 89 -3621 147 -3587
rect 89 -3655 101 -3621
rect 135 -3655 147 -3621
rect 89 -3689 147 -3655
rect 89 -3723 101 -3689
rect 135 -3723 147 -3689
rect 89 -3757 147 -3723
rect 89 -3791 101 -3757
rect 135 -3791 147 -3757
rect 89 -3825 147 -3791
rect 89 -3859 101 -3825
rect 135 -3859 147 -3825
rect 89 -3893 147 -3859
rect 89 -3927 101 -3893
rect 135 -3927 147 -3893
rect 89 -3961 147 -3927
rect 89 -3995 101 -3961
rect 135 -3995 147 -3961
rect 89 -4029 147 -3995
rect 89 -4063 101 -4029
rect 135 -4063 147 -4029
rect 89 -4097 147 -4063
rect 89 -4131 101 -4097
rect 135 -4131 147 -4097
rect 89 -4165 147 -4131
rect 89 -4199 101 -4165
rect 135 -4199 147 -4165
rect 89 -4233 147 -4199
rect 89 -4267 101 -4233
rect 135 -4267 147 -4233
rect 89 -4301 147 -4267
rect 89 -4335 101 -4301
rect 135 -4335 147 -4301
rect 89 -4369 147 -4335
rect 89 -4403 101 -4369
rect 135 -4403 147 -4369
rect 89 -4437 147 -4403
rect 89 -4471 101 -4437
rect 135 -4471 147 -4437
rect 89 -4505 147 -4471
rect 89 -4539 101 -4505
rect 135 -4539 147 -4505
rect 89 -4573 147 -4539
rect 89 -4607 101 -4573
rect 135 -4607 147 -4573
rect 89 -4641 147 -4607
rect 89 -4675 101 -4641
rect 135 -4675 147 -4641
rect 89 -4709 147 -4675
rect 89 -4743 101 -4709
rect 135 -4743 147 -4709
rect 89 -4777 147 -4743
rect 89 -4811 101 -4777
rect 135 -4811 147 -4777
rect 89 -4845 147 -4811
rect 89 -4879 101 -4845
rect 135 -4879 147 -4845
rect 89 -4913 147 -4879
rect 89 -4947 101 -4913
rect 135 -4947 147 -4913
rect 89 -4981 147 -4947
rect 89 -5015 101 -4981
rect 135 -5015 147 -4981
rect 89 -5049 147 -5015
rect 89 -5083 101 -5049
rect 135 -5083 147 -5049
rect 89 -5117 147 -5083
rect 89 -5151 101 -5117
rect 135 -5151 147 -5117
rect 89 -5185 147 -5151
rect 89 -5219 101 -5185
rect 135 -5219 147 -5185
rect 89 -5253 147 -5219
rect 89 -5287 101 -5253
rect 135 -5287 147 -5253
rect 89 -5321 147 -5287
rect 89 -5355 101 -5321
rect 135 -5355 147 -5321
rect 89 -5389 147 -5355
rect 89 -5423 101 -5389
rect 135 -5423 147 -5389
rect 89 -5457 147 -5423
rect 89 -5491 101 -5457
rect 135 -5491 147 -5457
rect 89 -5525 147 -5491
rect 89 -5559 101 -5525
rect 135 -5559 147 -5525
rect 89 -5593 147 -5559
rect 89 -5627 101 -5593
rect 135 -5627 147 -5593
rect 89 -5661 147 -5627
rect 89 -5695 101 -5661
rect 135 -5695 147 -5661
rect 89 -5729 147 -5695
rect 89 -5763 101 -5729
rect 135 -5763 147 -5729
rect 89 -5797 147 -5763
rect 89 -5831 101 -5797
rect 135 -5831 147 -5797
rect 89 -5865 147 -5831
rect 89 -5899 101 -5865
rect 135 -5899 147 -5865
rect 89 -5933 147 -5899
rect 89 -5967 101 -5933
rect 135 -5967 147 -5933
rect 89 -6000 147 -5967
rect 207 5967 265 6000
rect 207 5933 219 5967
rect 253 5933 265 5967
rect 207 5899 265 5933
rect 207 5865 219 5899
rect 253 5865 265 5899
rect 207 5831 265 5865
rect 207 5797 219 5831
rect 253 5797 265 5831
rect 207 5763 265 5797
rect 207 5729 219 5763
rect 253 5729 265 5763
rect 207 5695 265 5729
rect 207 5661 219 5695
rect 253 5661 265 5695
rect 207 5627 265 5661
rect 207 5593 219 5627
rect 253 5593 265 5627
rect 207 5559 265 5593
rect 207 5525 219 5559
rect 253 5525 265 5559
rect 207 5491 265 5525
rect 207 5457 219 5491
rect 253 5457 265 5491
rect 207 5423 265 5457
rect 207 5389 219 5423
rect 253 5389 265 5423
rect 207 5355 265 5389
rect 207 5321 219 5355
rect 253 5321 265 5355
rect 207 5287 265 5321
rect 207 5253 219 5287
rect 253 5253 265 5287
rect 207 5219 265 5253
rect 207 5185 219 5219
rect 253 5185 265 5219
rect 207 5151 265 5185
rect 207 5117 219 5151
rect 253 5117 265 5151
rect 207 5083 265 5117
rect 207 5049 219 5083
rect 253 5049 265 5083
rect 207 5015 265 5049
rect 207 4981 219 5015
rect 253 4981 265 5015
rect 207 4947 265 4981
rect 207 4913 219 4947
rect 253 4913 265 4947
rect 207 4879 265 4913
rect 207 4845 219 4879
rect 253 4845 265 4879
rect 207 4811 265 4845
rect 207 4777 219 4811
rect 253 4777 265 4811
rect 207 4743 265 4777
rect 207 4709 219 4743
rect 253 4709 265 4743
rect 207 4675 265 4709
rect 207 4641 219 4675
rect 253 4641 265 4675
rect 207 4607 265 4641
rect 207 4573 219 4607
rect 253 4573 265 4607
rect 207 4539 265 4573
rect 207 4505 219 4539
rect 253 4505 265 4539
rect 207 4471 265 4505
rect 207 4437 219 4471
rect 253 4437 265 4471
rect 207 4403 265 4437
rect 207 4369 219 4403
rect 253 4369 265 4403
rect 207 4335 265 4369
rect 207 4301 219 4335
rect 253 4301 265 4335
rect 207 4267 265 4301
rect 207 4233 219 4267
rect 253 4233 265 4267
rect 207 4199 265 4233
rect 207 4165 219 4199
rect 253 4165 265 4199
rect 207 4131 265 4165
rect 207 4097 219 4131
rect 253 4097 265 4131
rect 207 4063 265 4097
rect 207 4029 219 4063
rect 253 4029 265 4063
rect 207 3995 265 4029
rect 207 3961 219 3995
rect 253 3961 265 3995
rect 207 3927 265 3961
rect 207 3893 219 3927
rect 253 3893 265 3927
rect 207 3859 265 3893
rect 207 3825 219 3859
rect 253 3825 265 3859
rect 207 3791 265 3825
rect 207 3757 219 3791
rect 253 3757 265 3791
rect 207 3723 265 3757
rect 207 3689 219 3723
rect 253 3689 265 3723
rect 207 3655 265 3689
rect 207 3621 219 3655
rect 253 3621 265 3655
rect 207 3587 265 3621
rect 207 3553 219 3587
rect 253 3553 265 3587
rect 207 3519 265 3553
rect 207 3485 219 3519
rect 253 3485 265 3519
rect 207 3451 265 3485
rect 207 3417 219 3451
rect 253 3417 265 3451
rect 207 3383 265 3417
rect 207 3349 219 3383
rect 253 3349 265 3383
rect 207 3315 265 3349
rect 207 3281 219 3315
rect 253 3281 265 3315
rect 207 3247 265 3281
rect 207 3213 219 3247
rect 253 3213 265 3247
rect 207 3179 265 3213
rect 207 3145 219 3179
rect 253 3145 265 3179
rect 207 3111 265 3145
rect 207 3077 219 3111
rect 253 3077 265 3111
rect 207 3043 265 3077
rect 207 3009 219 3043
rect 253 3009 265 3043
rect 207 2975 265 3009
rect 207 2941 219 2975
rect 253 2941 265 2975
rect 207 2907 265 2941
rect 207 2873 219 2907
rect 253 2873 265 2907
rect 207 2839 265 2873
rect 207 2805 219 2839
rect 253 2805 265 2839
rect 207 2771 265 2805
rect 207 2737 219 2771
rect 253 2737 265 2771
rect 207 2703 265 2737
rect 207 2669 219 2703
rect 253 2669 265 2703
rect 207 2635 265 2669
rect 207 2601 219 2635
rect 253 2601 265 2635
rect 207 2567 265 2601
rect 207 2533 219 2567
rect 253 2533 265 2567
rect 207 2499 265 2533
rect 207 2465 219 2499
rect 253 2465 265 2499
rect 207 2431 265 2465
rect 207 2397 219 2431
rect 253 2397 265 2431
rect 207 2363 265 2397
rect 207 2329 219 2363
rect 253 2329 265 2363
rect 207 2295 265 2329
rect 207 2261 219 2295
rect 253 2261 265 2295
rect 207 2227 265 2261
rect 207 2193 219 2227
rect 253 2193 265 2227
rect 207 2159 265 2193
rect 207 2125 219 2159
rect 253 2125 265 2159
rect 207 2091 265 2125
rect 207 2057 219 2091
rect 253 2057 265 2091
rect 207 2023 265 2057
rect 207 1989 219 2023
rect 253 1989 265 2023
rect 207 1955 265 1989
rect 207 1921 219 1955
rect 253 1921 265 1955
rect 207 1887 265 1921
rect 207 1853 219 1887
rect 253 1853 265 1887
rect 207 1819 265 1853
rect 207 1785 219 1819
rect 253 1785 265 1819
rect 207 1751 265 1785
rect 207 1717 219 1751
rect 253 1717 265 1751
rect 207 1683 265 1717
rect 207 1649 219 1683
rect 253 1649 265 1683
rect 207 1615 265 1649
rect 207 1581 219 1615
rect 253 1581 265 1615
rect 207 1547 265 1581
rect 207 1513 219 1547
rect 253 1513 265 1547
rect 207 1479 265 1513
rect 207 1445 219 1479
rect 253 1445 265 1479
rect 207 1411 265 1445
rect 207 1377 219 1411
rect 253 1377 265 1411
rect 207 1343 265 1377
rect 207 1309 219 1343
rect 253 1309 265 1343
rect 207 1275 265 1309
rect 207 1241 219 1275
rect 253 1241 265 1275
rect 207 1207 265 1241
rect 207 1173 219 1207
rect 253 1173 265 1207
rect 207 1139 265 1173
rect 207 1105 219 1139
rect 253 1105 265 1139
rect 207 1071 265 1105
rect 207 1037 219 1071
rect 253 1037 265 1071
rect 207 1003 265 1037
rect 207 969 219 1003
rect 253 969 265 1003
rect 207 935 265 969
rect 207 901 219 935
rect 253 901 265 935
rect 207 867 265 901
rect 207 833 219 867
rect 253 833 265 867
rect 207 799 265 833
rect 207 765 219 799
rect 253 765 265 799
rect 207 731 265 765
rect 207 697 219 731
rect 253 697 265 731
rect 207 663 265 697
rect 207 629 219 663
rect 253 629 265 663
rect 207 595 265 629
rect 207 561 219 595
rect 253 561 265 595
rect 207 527 265 561
rect 207 493 219 527
rect 253 493 265 527
rect 207 459 265 493
rect 207 425 219 459
rect 253 425 265 459
rect 207 391 265 425
rect 207 357 219 391
rect 253 357 265 391
rect 207 323 265 357
rect 207 289 219 323
rect 253 289 265 323
rect 207 255 265 289
rect 207 221 219 255
rect 253 221 265 255
rect 207 187 265 221
rect 207 153 219 187
rect 253 153 265 187
rect 207 119 265 153
rect 207 85 219 119
rect 253 85 265 119
rect 207 51 265 85
rect 207 17 219 51
rect 253 17 265 51
rect 207 -17 265 17
rect 207 -51 219 -17
rect 253 -51 265 -17
rect 207 -85 265 -51
rect 207 -119 219 -85
rect 253 -119 265 -85
rect 207 -153 265 -119
rect 207 -187 219 -153
rect 253 -187 265 -153
rect 207 -221 265 -187
rect 207 -255 219 -221
rect 253 -255 265 -221
rect 207 -289 265 -255
rect 207 -323 219 -289
rect 253 -323 265 -289
rect 207 -357 265 -323
rect 207 -391 219 -357
rect 253 -391 265 -357
rect 207 -425 265 -391
rect 207 -459 219 -425
rect 253 -459 265 -425
rect 207 -493 265 -459
rect 207 -527 219 -493
rect 253 -527 265 -493
rect 207 -561 265 -527
rect 207 -595 219 -561
rect 253 -595 265 -561
rect 207 -629 265 -595
rect 207 -663 219 -629
rect 253 -663 265 -629
rect 207 -697 265 -663
rect 207 -731 219 -697
rect 253 -731 265 -697
rect 207 -765 265 -731
rect 207 -799 219 -765
rect 253 -799 265 -765
rect 207 -833 265 -799
rect 207 -867 219 -833
rect 253 -867 265 -833
rect 207 -901 265 -867
rect 207 -935 219 -901
rect 253 -935 265 -901
rect 207 -969 265 -935
rect 207 -1003 219 -969
rect 253 -1003 265 -969
rect 207 -1037 265 -1003
rect 207 -1071 219 -1037
rect 253 -1071 265 -1037
rect 207 -1105 265 -1071
rect 207 -1139 219 -1105
rect 253 -1139 265 -1105
rect 207 -1173 265 -1139
rect 207 -1207 219 -1173
rect 253 -1207 265 -1173
rect 207 -1241 265 -1207
rect 207 -1275 219 -1241
rect 253 -1275 265 -1241
rect 207 -1309 265 -1275
rect 207 -1343 219 -1309
rect 253 -1343 265 -1309
rect 207 -1377 265 -1343
rect 207 -1411 219 -1377
rect 253 -1411 265 -1377
rect 207 -1445 265 -1411
rect 207 -1479 219 -1445
rect 253 -1479 265 -1445
rect 207 -1513 265 -1479
rect 207 -1547 219 -1513
rect 253 -1547 265 -1513
rect 207 -1581 265 -1547
rect 207 -1615 219 -1581
rect 253 -1615 265 -1581
rect 207 -1649 265 -1615
rect 207 -1683 219 -1649
rect 253 -1683 265 -1649
rect 207 -1717 265 -1683
rect 207 -1751 219 -1717
rect 253 -1751 265 -1717
rect 207 -1785 265 -1751
rect 207 -1819 219 -1785
rect 253 -1819 265 -1785
rect 207 -1853 265 -1819
rect 207 -1887 219 -1853
rect 253 -1887 265 -1853
rect 207 -1921 265 -1887
rect 207 -1955 219 -1921
rect 253 -1955 265 -1921
rect 207 -1989 265 -1955
rect 207 -2023 219 -1989
rect 253 -2023 265 -1989
rect 207 -2057 265 -2023
rect 207 -2091 219 -2057
rect 253 -2091 265 -2057
rect 207 -2125 265 -2091
rect 207 -2159 219 -2125
rect 253 -2159 265 -2125
rect 207 -2193 265 -2159
rect 207 -2227 219 -2193
rect 253 -2227 265 -2193
rect 207 -2261 265 -2227
rect 207 -2295 219 -2261
rect 253 -2295 265 -2261
rect 207 -2329 265 -2295
rect 207 -2363 219 -2329
rect 253 -2363 265 -2329
rect 207 -2397 265 -2363
rect 207 -2431 219 -2397
rect 253 -2431 265 -2397
rect 207 -2465 265 -2431
rect 207 -2499 219 -2465
rect 253 -2499 265 -2465
rect 207 -2533 265 -2499
rect 207 -2567 219 -2533
rect 253 -2567 265 -2533
rect 207 -2601 265 -2567
rect 207 -2635 219 -2601
rect 253 -2635 265 -2601
rect 207 -2669 265 -2635
rect 207 -2703 219 -2669
rect 253 -2703 265 -2669
rect 207 -2737 265 -2703
rect 207 -2771 219 -2737
rect 253 -2771 265 -2737
rect 207 -2805 265 -2771
rect 207 -2839 219 -2805
rect 253 -2839 265 -2805
rect 207 -2873 265 -2839
rect 207 -2907 219 -2873
rect 253 -2907 265 -2873
rect 207 -2941 265 -2907
rect 207 -2975 219 -2941
rect 253 -2975 265 -2941
rect 207 -3009 265 -2975
rect 207 -3043 219 -3009
rect 253 -3043 265 -3009
rect 207 -3077 265 -3043
rect 207 -3111 219 -3077
rect 253 -3111 265 -3077
rect 207 -3145 265 -3111
rect 207 -3179 219 -3145
rect 253 -3179 265 -3145
rect 207 -3213 265 -3179
rect 207 -3247 219 -3213
rect 253 -3247 265 -3213
rect 207 -3281 265 -3247
rect 207 -3315 219 -3281
rect 253 -3315 265 -3281
rect 207 -3349 265 -3315
rect 207 -3383 219 -3349
rect 253 -3383 265 -3349
rect 207 -3417 265 -3383
rect 207 -3451 219 -3417
rect 253 -3451 265 -3417
rect 207 -3485 265 -3451
rect 207 -3519 219 -3485
rect 253 -3519 265 -3485
rect 207 -3553 265 -3519
rect 207 -3587 219 -3553
rect 253 -3587 265 -3553
rect 207 -3621 265 -3587
rect 207 -3655 219 -3621
rect 253 -3655 265 -3621
rect 207 -3689 265 -3655
rect 207 -3723 219 -3689
rect 253 -3723 265 -3689
rect 207 -3757 265 -3723
rect 207 -3791 219 -3757
rect 253 -3791 265 -3757
rect 207 -3825 265 -3791
rect 207 -3859 219 -3825
rect 253 -3859 265 -3825
rect 207 -3893 265 -3859
rect 207 -3927 219 -3893
rect 253 -3927 265 -3893
rect 207 -3961 265 -3927
rect 207 -3995 219 -3961
rect 253 -3995 265 -3961
rect 207 -4029 265 -3995
rect 207 -4063 219 -4029
rect 253 -4063 265 -4029
rect 207 -4097 265 -4063
rect 207 -4131 219 -4097
rect 253 -4131 265 -4097
rect 207 -4165 265 -4131
rect 207 -4199 219 -4165
rect 253 -4199 265 -4165
rect 207 -4233 265 -4199
rect 207 -4267 219 -4233
rect 253 -4267 265 -4233
rect 207 -4301 265 -4267
rect 207 -4335 219 -4301
rect 253 -4335 265 -4301
rect 207 -4369 265 -4335
rect 207 -4403 219 -4369
rect 253 -4403 265 -4369
rect 207 -4437 265 -4403
rect 207 -4471 219 -4437
rect 253 -4471 265 -4437
rect 207 -4505 265 -4471
rect 207 -4539 219 -4505
rect 253 -4539 265 -4505
rect 207 -4573 265 -4539
rect 207 -4607 219 -4573
rect 253 -4607 265 -4573
rect 207 -4641 265 -4607
rect 207 -4675 219 -4641
rect 253 -4675 265 -4641
rect 207 -4709 265 -4675
rect 207 -4743 219 -4709
rect 253 -4743 265 -4709
rect 207 -4777 265 -4743
rect 207 -4811 219 -4777
rect 253 -4811 265 -4777
rect 207 -4845 265 -4811
rect 207 -4879 219 -4845
rect 253 -4879 265 -4845
rect 207 -4913 265 -4879
rect 207 -4947 219 -4913
rect 253 -4947 265 -4913
rect 207 -4981 265 -4947
rect 207 -5015 219 -4981
rect 253 -5015 265 -4981
rect 207 -5049 265 -5015
rect 207 -5083 219 -5049
rect 253 -5083 265 -5049
rect 207 -5117 265 -5083
rect 207 -5151 219 -5117
rect 253 -5151 265 -5117
rect 207 -5185 265 -5151
rect 207 -5219 219 -5185
rect 253 -5219 265 -5185
rect 207 -5253 265 -5219
rect 207 -5287 219 -5253
rect 253 -5287 265 -5253
rect 207 -5321 265 -5287
rect 207 -5355 219 -5321
rect 253 -5355 265 -5321
rect 207 -5389 265 -5355
rect 207 -5423 219 -5389
rect 253 -5423 265 -5389
rect 207 -5457 265 -5423
rect 207 -5491 219 -5457
rect 253 -5491 265 -5457
rect 207 -5525 265 -5491
rect 207 -5559 219 -5525
rect 253 -5559 265 -5525
rect 207 -5593 265 -5559
rect 207 -5627 219 -5593
rect 253 -5627 265 -5593
rect 207 -5661 265 -5627
rect 207 -5695 219 -5661
rect 253 -5695 265 -5661
rect 207 -5729 265 -5695
rect 207 -5763 219 -5729
rect 253 -5763 265 -5729
rect 207 -5797 265 -5763
rect 207 -5831 219 -5797
rect 253 -5831 265 -5797
rect 207 -5865 265 -5831
rect 207 -5899 219 -5865
rect 253 -5899 265 -5865
rect 207 -5933 265 -5899
rect 207 -5967 219 -5933
rect 253 -5967 265 -5933
rect 207 -6000 265 -5967
rect 325 5967 383 6000
rect 325 5933 337 5967
rect 371 5933 383 5967
rect 325 5899 383 5933
rect 325 5865 337 5899
rect 371 5865 383 5899
rect 325 5831 383 5865
rect 325 5797 337 5831
rect 371 5797 383 5831
rect 325 5763 383 5797
rect 325 5729 337 5763
rect 371 5729 383 5763
rect 325 5695 383 5729
rect 325 5661 337 5695
rect 371 5661 383 5695
rect 325 5627 383 5661
rect 325 5593 337 5627
rect 371 5593 383 5627
rect 325 5559 383 5593
rect 325 5525 337 5559
rect 371 5525 383 5559
rect 325 5491 383 5525
rect 325 5457 337 5491
rect 371 5457 383 5491
rect 325 5423 383 5457
rect 325 5389 337 5423
rect 371 5389 383 5423
rect 325 5355 383 5389
rect 325 5321 337 5355
rect 371 5321 383 5355
rect 325 5287 383 5321
rect 325 5253 337 5287
rect 371 5253 383 5287
rect 325 5219 383 5253
rect 325 5185 337 5219
rect 371 5185 383 5219
rect 325 5151 383 5185
rect 325 5117 337 5151
rect 371 5117 383 5151
rect 325 5083 383 5117
rect 325 5049 337 5083
rect 371 5049 383 5083
rect 325 5015 383 5049
rect 325 4981 337 5015
rect 371 4981 383 5015
rect 325 4947 383 4981
rect 325 4913 337 4947
rect 371 4913 383 4947
rect 325 4879 383 4913
rect 325 4845 337 4879
rect 371 4845 383 4879
rect 325 4811 383 4845
rect 325 4777 337 4811
rect 371 4777 383 4811
rect 325 4743 383 4777
rect 325 4709 337 4743
rect 371 4709 383 4743
rect 325 4675 383 4709
rect 325 4641 337 4675
rect 371 4641 383 4675
rect 325 4607 383 4641
rect 325 4573 337 4607
rect 371 4573 383 4607
rect 325 4539 383 4573
rect 325 4505 337 4539
rect 371 4505 383 4539
rect 325 4471 383 4505
rect 325 4437 337 4471
rect 371 4437 383 4471
rect 325 4403 383 4437
rect 325 4369 337 4403
rect 371 4369 383 4403
rect 325 4335 383 4369
rect 325 4301 337 4335
rect 371 4301 383 4335
rect 325 4267 383 4301
rect 325 4233 337 4267
rect 371 4233 383 4267
rect 325 4199 383 4233
rect 325 4165 337 4199
rect 371 4165 383 4199
rect 325 4131 383 4165
rect 325 4097 337 4131
rect 371 4097 383 4131
rect 325 4063 383 4097
rect 325 4029 337 4063
rect 371 4029 383 4063
rect 325 3995 383 4029
rect 325 3961 337 3995
rect 371 3961 383 3995
rect 325 3927 383 3961
rect 325 3893 337 3927
rect 371 3893 383 3927
rect 325 3859 383 3893
rect 325 3825 337 3859
rect 371 3825 383 3859
rect 325 3791 383 3825
rect 325 3757 337 3791
rect 371 3757 383 3791
rect 325 3723 383 3757
rect 325 3689 337 3723
rect 371 3689 383 3723
rect 325 3655 383 3689
rect 325 3621 337 3655
rect 371 3621 383 3655
rect 325 3587 383 3621
rect 325 3553 337 3587
rect 371 3553 383 3587
rect 325 3519 383 3553
rect 325 3485 337 3519
rect 371 3485 383 3519
rect 325 3451 383 3485
rect 325 3417 337 3451
rect 371 3417 383 3451
rect 325 3383 383 3417
rect 325 3349 337 3383
rect 371 3349 383 3383
rect 325 3315 383 3349
rect 325 3281 337 3315
rect 371 3281 383 3315
rect 325 3247 383 3281
rect 325 3213 337 3247
rect 371 3213 383 3247
rect 325 3179 383 3213
rect 325 3145 337 3179
rect 371 3145 383 3179
rect 325 3111 383 3145
rect 325 3077 337 3111
rect 371 3077 383 3111
rect 325 3043 383 3077
rect 325 3009 337 3043
rect 371 3009 383 3043
rect 325 2975 383 3009
rect 325 2941 337 2975
rect 371 2941 383 2975
rect 325 2907 383 2941
rect 325 2873 337 2907
rect 371 2873 383 2907
rect 325 2839 383 2873
rect 325 2805 337 2839
rect 371 2805 383 2839
rect 325 2771 383 2805
rect 325 2737 337 2771
rect 371 2737 383 2771
rect 325 2703 383 2737
rect 325 2669 337 2703
rect 371 2669 383 2703
rect 325 2635 383 2669
rect 325 2601 337 2635
rect 371 2601 383 2635
rect 325 2567 383 2601
rect 325 2533 337 2567
rect 371 2533 383 2567
rect 325 2499 383 2533
rect 325 2465 337 2499
rect 371 2465 383 2499
rect 325 2431 383 2465
rect 325 2397 337 2431
rect 371 2397 383 2431
rect 325 2363 383 2397
rect 325 2329 337 2363
rect 371 2329 383 2363
rect 325 2295 383 2329
rect 325 2261 337 2295
rect 371 2261 383 2295
rect 325 2227 383 2261
rect 325 2193 337 2227
rect 371 2193 383 2227
rect 325 2159 383 2193
rect 325 2125 337 2159
rect 371 2125 383 2159
rect 325 2091 383 2125
rect 325 2057 337 2091
rect 371 2057 383 2091
rect 325 2023 383 2057
rect 325 1989 337 2023
rect 371 1989 383 2023
rect 325 1955 383 1989
rect 325 1921 337 1955
rect 371 1921 383 1955
rect 325 1887 383 1921
rect 325 1853 337 1887
rect 371 1853 383 1887
rect 325 1819 383 1853
rect 325 1785 337 1819
rect 371 1785 383 1819
rect 325 1751 383 1785
rect 325 1717 337 1751
rect 371 1717 383 1751
rect 325 1683 383 1717
rect 325 1649 337 1683
rect 371 1649 383 1683
rect 325 1615 383 1649
rect 325 1581 337 1615
rect 371 1581 383 1615
rect 325 1547 383 1581
rect 325 1513 337 1547
rect 371 1513 383 1547
rect 325 1479 383 1513
rect 325 1445 337 1479
rect 371 1445 383 1479
rect 325 1411 383 1445
rect 325 1377 337 1411
rect 371 1377 383 1411
rect 325 1343 383 1377
rect 325 1309 337 1343
rect 371 1309 383 1343
rect 325 1275 383 1309
rect 325 1241 337 1275
rect 371 1241 383 1275
rect 325 1207 383 1241
rect 325 1173 337 1207
rect 371 1173 383 1207
rect 325 1139 383 1173
rect 325 1105 337 1139
rect 371 1105 383 1139
rect 325 1071 383 1105
rect 325 1037 337 1071
rect 371 1037 383 1071
rect 325 1003 383 1037
rect 325 969 337 1003
rect 371 969 383 1003
rect 325 935 383 969
rect 325 901 337 935
rect 371 901 383 935
rect 325 867 383 901
rect 325 833 337 867
rect 371 833 383 867
rect 325 799 383 833
rect 325 765 337 799
rect 371 765 383 799
rect 325 731 383 765
rect 325 697 337 731
rect 371 697 383 731
rect 325 663 383 697
rect 325 629 337 663
rect 371 629 383 663
rect 325 595 383 629
rect 325 561 337 595
rect 371 561 383 595
rect 325 527 383 561
rect 325 493 337 527
rect 371 493 383 527
rect 325 459 383 493
rect 325 425 337 459
rect 371 425 383 459
rect 325 391 383 425
rect 325 357 337 391
rect 371 357 383 391
rect 325 323 383 357
rect 325 289 337 323
rect 371 289 383 323
rect 325 255 383 289
rect 325 221 337 255
rect 371 221 383 255
rect 325 187 383 221
rect 325 153 337 187
rect 371 153 383 187
rect 325 119 383 153
rect 325 85 337 119
rect 371 85 383 119
rect 325 51 383 85
rect 325 17 337 51
rect 371 17 383 51
rect 325 -17 383 17
rect 325 -51 337 -17
rect 371 -51 383 -17
rect 325 -85 383 -51
rect 325 -119 337 -85
rect 371 -119 383 -85
rect 325 -153 383 -119
rect 325 -187 337 -153
rect 371 -187 383 -153
rect 325 -221 383 -187
rect 325 -255 337 -221
rect 371 -255 383 -221
rect 325 -289 383 -255
rect 325 -323 337 -289
rect 371 -323 383 -289
rect 325 -357 383 -323
rect 325 -391 337 -357
rect 371 -391 383 -357
rect 325 -425 383 -391
rect 325 -459 337 -425
rect 371 -459 383 -425
rect 325 -493 383 -459
rect 325 -527 337 -493
rect 371 -527 383 -493
rect 325 -561 383 -527
rect 325 -595 337 -561
rect 371 -595 383 -561
rect 325 -629 383 -595
rect 325 -663 337 -629
rect 371 -663 383 -629
rect 325 -697 383 -663
rect 325 -731 337 -697
rect 371 -731 383 -697
rect 325 -765 383 -731
rect 325 -799 337 -765
rect 371 -799 383 -765
rect 325 -833 383 -799
rect 325 -867 337 -833
rect 371 -867 383 -833
rect 325 -901 383 -867
rect 325 -935 337 -901
rect 371 -935 383 -901
rect 325 -969 383 -935
rect 325 -1003 337 -969
rect 371 -1003 383 -969
rect 325 -1037 383 -1003
rect 325 -1071 337 -1037
rect 371 -1071 383 -1037
rect 325 -1105 383 -1071
rect 325 -1139 337 -1105
rect 371 -1139 383 -1105
rect 325 -1173 383 -1139
rect 325 -1207 337 -1173
rect 371 -1207 383 -1173
rect 325 -1241 383 -1207
rect 325 -1275 337 -1241
rect 371 -1275 383 -1241
rect 325 -1309 383 -1275
rect 325 -1343 337 -1309
rect 371 -1343 383 -1309
rect 325 -1377 383 -1343
rect 325 -1411 337 -1377
rect 371 -1411 383 -1377
rect 325 -1445 383 -1411
rect 325 -1479 337 -1445
rect 371 -1479 383 -1445
rect 325 -1513 383 -1479
rect 325 -1547 337 -1513
rect 371 -1547 383 -1513
rect 325 -1581 383 -1547
rect 325 -1615 337 -1581
rect 371 -1615 383 -1581
rect 325 -1649 383 -1615
rect 325 -1683 337 -1649
rect 371 -1683 383 -1649
rect 325 -1717 383 -1683
rect 325 -1751 337 -1717
rect 371 -1751 383 -1717
rect 325 -1785 383 -1751
rect 325 -1819 337 -1785
rect 371 -1819 383 -1785
rect 325 -1853 383 -1819
rect 325 -1887 337 -1853
rect 371 -1887 383 -1853
rect 325 -1921 383 -1887
rect 325 -1955 337 -1921
rect 371 -1955 383 -1921
rect 325 -1989 383 -1955
rect 325 -2023 337 -1989
rect 371 -2023 383 -1989
rect 325 -2057 383 -2023
rect 325 -2091 337 -2057
rect 371 -2091 383 -2057
rect 325 -2125 383 -2091
rect 325 -2159 337 -2125
rect 371 -2159 383 -2125
rect 325 -2193 383 -2159
rect 325 -2227 337 -2193
rect 371 -2227 383 -2193
rect 325 -2261 383 -2227
rect 325 -2295 337 -2261
rect 371 -2295 383 -2261
rect 325 -2329 383 -2295
rect 325 -2363 337 -2329
rect 371 -2363 383 -2329
rect 325 -2397 383 -2363
rect 325 -2431 337 -2397
rect 371 -2431 383 -2397
rect 325 -2465 383 -2431
rect 325 -2499 337 -2465
rect 371 -2499 383 -2465
rect 325 -2533 383 -2499
rect 325 -2567 337 -2533
rect 371 -2567 383 -2533
rect 325 -2601 383 -2567
rect 325 -2635 337 -2601
rect 371 -2635 383 -2601
rect 325 -2669 383 -2635
rect 325 -2703 337 -2669
rect 371 -2703 383 -2669
rect 325 -2737 383 -2703
rect 325 -2771 337 -2737
rect 371 -2771 383 -2737
rect 325 -2805 383 -2771
rect 325 -2839 337 -2805
rect 371 -2839 383 -2805
rect 325 -2873 383 -2839
rect 325 -2907 337 -2873
rect 371 -2907 383 -2873
rect 325 -2941 383 -2907
rect 325 -2975 337 -2941
rect 371 -2975 383 -2941
rect 325 -3009 383 -2975
rect 325 -3043 337 -3009
rect 371 -3043 383 -3009
rect 325 -3077 383 -3043
rect 325 -3111 337 -3077
rect 371 -3111 383 -3077
rect 325 -3145 383 -3111
rect 325 -3179 337 -3145
rect 371 -3179 383 -3145
rect 325 -3213 383 -3179
rect 325 -3247 337 -3213
rect 371 -3247 383 -3213
rect 325 -3281 383 -3247
rect 325 -3315 337 -3281
rect 371 -3315 383 -3281
rect 325 -3349 383 -3315
rect 325 -3383 337 -3349
rect 371 -3383 383 -3349
rect 325 -3417 383 -3383
rect 325 -3451 337 -3417
rect 371 -3451 383 -3417
rect 325 -3485 383 -3451
rect 325 -3519 337 -3485
rect 371 -3519 383 -3485
rect 325 -3553 383 -3519
rect 325 -3587 337 -3553
rect 371 -3587 383 -3553
rect 325 -3621 383 -3587
rect 325 -3655 337 -3621
rect 371 -3655 383 -3621
rect 325 -3689 383 -3655
rect 325 -3723 337 -3689
rect 371 -3723 383 -3689
rect 325 -3757 383 -3723
rect 325 -3791 337 -3757
rect 371 -3791 383 -3757
rect 325 -3825 383 -3791
rect 325 -3859 337 -3825
rect 371 -3859 383 -3825
rect 325 -3893 383 -3859
rect 325 -3927 337 -3893
rect 371 -3927 383 -3893
rect 325 -3961 383 -3927
rect 325 -3995 337 -3961
rect 371 -3995 383 -3961
rect 325 -4029 383 -3995
rect 325 -4063 337 -4029
rect 371 -4063 383 -4029
rect 325 -4097 383 -4063
rect 325 -4131 337 -4097
rect 371 -4131 383 -4097
rect 325 -4165 383 -4131
rect 325 -4199 337 -4165
rect 371 -4199 383 -4165
rect 325 -4233 383 -4199
rect 325 -4267 337 -4233
rect 371 -4267 383 -4233
rect 325 -4301 383 -4267
rect 325 -4335 337 -4301
rect 371 -4335 383 -4301
rect 325 -4369 383 -4335
rect 325 -4403 337 -4369
rect 371 -4403 383 -4369
rect 325 -4437 383 -4403
rect 325 -4471 337 -4437
rect 371 -4471 383 -4437
rect 325 -4505 383 -4471
rect 325 -4539 337 -4505
rect 371 -4539 383 -4505
rect 325 -4573 383 -4539
rect 325 -4607 337 -4573
rect 371 -4607 383 -4573
rect 325 -4641 383 -4607
rect 325 -4675 337 -4641
rect 371 -4675 383 -4641
rect 325 -4709 383 -4675
rect 325 -4743 337 -4709
rect 371 -4743 383 -4709
rect 325 -4777 383 -4743
rect 325 -4811 337 -4777
rect 371 -4811 383 -4777
rect 325 -4845 383 -4811
rect 325 -4879 337 -4845
rect 371 -4879 383 -4845
rect 325 -4913 383 -4879
rect 325 -4947 337 -4913
rect 371 -4947 383 -4913
rect 325 -4981 383 -4947
rect 325 -5015 337 -4981
rect 371 -5015 383 -4981
rect 325 -5049 383 -5015
rect 325 -5083 337 -5049
rect 371 -5083 383 -5049
rect 325 -5117 383 -5083
rect 325 -5151 337 -5117
rect 371 -5151 383 -5117
rect 325 -5185 383 -5151
rect 325 -5219 337 -5185
rect 371 -5219 383 -5185
rect 325 -5253 383 -5219
rect 325 -5287 337 -5253
rect 371 -5287 383 -5253
rect 325 -5321 383 -5287
rect 325 -5355 337 -5321
rect 371 -5355 383 -5321
rect 325 -5389 383 -5355
rect 325 -5423 337 -5389
rect 371 -5423 383 -5389
rect 325 -5457 383 -5423
rect 325 -5491 337 -5457
rect 371 -5491 383 -5457
rect 325 -5525 383 -5491
rect 325 -5559 337 -5525
rect 371 -5559 383 -5525
rect 325 -5593 383 -5559
rect 325 -5627 337 -5593
rect 371 -5627 383 -5593
rect 325 -5661 383 -5627
rect 325 -5695 337 -5661
rect 371 -5695 383 -5661
rect 325 -5729 383 -5695
rect 325 -5763 337 -5729
rect 371 -5763 383 -5729
rect 325 -5797 383 -5763
rect 325 -5831 337 -5797
rect 371 -5831 383 -5797
rect 325 -5865 383 -5831
rect 325 -5899 337 -5865
rect 371 -5899 383 -5865
rect 325 -5933 383 -5899
rect 325 -5967 337 -5933
rect 371 -5967 383 -5933
rect 325 -6000 383 -5967
rect 443 5967 501 6000
rect 443 5933 455 5967
rect 489 5933 501 5967
rect 443 5899 501 5933
rect 443 5865 455 5899
rect 489 5865 501 5899
rect 443 5831 501 5865
rect 443 5797 455 5831
rect 489 5797 501 5831
rect 443 5763 501 5797
rect 443 5729 455 5763
rect 489 5729 501 5763
rect 443 5695 501 5729
rect 443 5661 455 5695
rect 489 5661 501 5695
rect 443 5627 501 5661
rect 443 5593 455 5627
rect 489 5593 501 5627
rect 443 5559 501 5593
rect 443 5525 455 5559
rect 489 5525 501 5559
rect 443 5491 501 5525
rect 443 5457 455 5491
rect 489 5457 501 5491
rect 443 5423 501 5457
rect 443 5389 455 5423
rect 489 5389 501 5423
rect 443 5355 501 5389
rect 443 5321 455 5355
rect 489 5321 501 5355
rect 443 5287 501 5321
rect 443 5253 455 5287
rect 489 5253 501 5287
rect 443 5219 501 5253
rect 443 5185 455 5219
rect 489 5185 501 5219
rect 443 5151 501 5185
rect 443 5117 455 5151
rect 489 5117 501 5151
rect 443 5083 501 5117
rect 443 5049 455 5083
rect 489 5049 501 5083
rect 443 5015 501 5049
rect 443 4981 455 5015
rect 489 4981 501 5015
rect 443 4947 501 4981
rect 443 4913 455 4947
rect 489 4913 501 4947
rect 443 4879 501 4913
rect 443 4845 455 4879
rect 489 4845 501 4879
rect 443 4811 501 4845
rect 443 4777 455 4811
rect 489 4777 501 4811
rect 443 4743 501 4777
rect 443 4709 455 4743
rect 489 4709 501 4743
rect 443 4675 501 4709
rect 443 4641 455 4675
rect 489 4641 501 4675
rect 443 4607 501 4641
rect 443 4573 455 4607
rect 489 4573 501 4607
rect 443 4539 501 4573
rect 443 4505 455 4539
rect 489 4505 501 4539
rect 443 4471 501 4505
rect 443 4437 455 4471
rect 489 4437 501 4471
rect 443 4403 501 4437
rect 443 4369 455 4403
rect 489 4369 501 4403
rect 443 4335 501 4369
rect 443 4301 455 4335
rect 489 4301 501 4335
rect 443 4267 501 4301
rect 443 4233 455 4267
rect 489 4233 501 4267
rect 443 4199 501 4233
rect 443 4165 455 4199
rect 489 4165 501 4199
rect 443 4131 501 4165
rect 443 4097 455 4131
rect 489 4097 501 4131
rect 443 4063 501 4097
rect 443 4029 455 4063
rect 489 4029 501 4063
rect 443 3995 501 4029
rect 443 3961 455 3995
rect 489 3961 501 3995
rect 443 3927 501 3961
rect 443 3893 455 3927
rect 489 3893 501 3927
rect 443 3859 501 3893
rect 443 3825 455 3859
rect 489 3825 501 3859
rect 443 3791 501 3825
rect 443 3757 455 3791
rect 489 3757 501 3791
rect 443 3723 501 3757
rect 443 3689 455 3723
rect 489 3689 501 3723
rect 443 3655 501 3689
rect 443 3621 455 3655
rect 489 3621 501 3655
rect 443 3587 501 3621
rect 443 3553 455 3587
rect 489 3553 501 3587
rect 443 3519 501 3553
rect 443 3485 455 3519
rect 489 3485 501 3519
rect 443 3451 501 3485
rect 443 3417 455 3451
rect 489 3417 501 3451
rect 443 3383 501 3417
rect 443 3349 455 3383
rect 489 3349 501 3383
rect 443 3315 501 3349
rect 443 3281 455 3315
rect 489 3281 501 3315
rect 443 3247 501 3281
rect 443 3213 455 3247
rect 489 3213 501 3247
rect 443 3179 501 3213
rect 443 3145 455 3179
rect 489 3145 501 3179
rect 443 3111 501 3145
rect 443 3077 455 3111
rect 489 3077 501 3111
rect 443 3043 501 3077
rect 443 3009 455 3043
rect 489 3009 501 3043
rect 443 2975 501 3009
rect 443 2941 455 2975
rect 489 2941 501 2975
rect 443 2907 501 2941
rect 443 2873 455 2907
rect 489 2873 501 2907
rect 443 2839 501 2873
rect 443 2805 455 2839
rect 489 2805 501 2839
rect 443 2771 501 2805
rect 443 2737 455 2771
rect 489 2737 501 2771
rect 443 2703 501 2737
rect 443 2669 455 2703
rect 489 2669 501 2703
rect 443 2635 501 2669
rect 443 2601 455 2635
rect 489 2601 501 2635
rect 443 2567 501 2601
rect 443 2533 455 2567
rect 489 2533 501 2567
rect 443 2499 501 2533
rect 443 2465 455 2499
rect 489 2465 501 2499
rect 443 2431 501 2465
rect 443 2397 455 2431
rect 489 2397 501 2431
rect 443 2363 501 2397
rect 443 2329 455 2363
rect 489 2329 501 2363
rect 443 2295 501 2329
rect 443 2261 455 2295
rect 489 2261 501 2295
rect 443 2227 501 2261
rect 443 2193 455 2227
rect 489 2193 501 2227
rect 443 2159 501 2193
rect 443 2125 455 2159
rect 489 2125 501 2159
rect 443 2091 501 2125
rect 443 2057 455 2091
rect 489 2057 501 2091
rect 443 2023 501 2057
rect 443 1989 455 2023
rect 489 1989 501 2023
rect 443 1955 501 1989
rect 443 1921 455 1955
rect 489 1921 501 1955
rect 443 1887 501 1921
rect 443 1853 455 1887
rect 489 1853 501 1887
rect 443 1819 501 1853
rect 443 1785 455 1819
rect 489 1785 501 1819
rect 443 1751 501 1785
rect 443 1717 455 1751
rect 489 1717 501 1751
rect 443 1683 501 1717
rect 443 1649 455 1683
rect 489 1649 501 1683
rect 443 1615 501 1649
rect 443 1581 455 1615
rect 489 1581 501 1615
rect 443 1547 501 1581
rect 443 1513 455 1547
rect 489 1513 501 1547
rect 443 1479 501 1513
rect 443 1445 455 1479
rect 489 1445 501 1479
rect 443 1411 501 1445
rect 443 1377 455 1411
rect 489 1377 501 1411
rect 443 1343 501 1377
rect 443 1309 455 1343
rect 489 1309 501 1343
rect 443 1275 501 1309
rect 443 1241 455 1275
rect 489 1241 501 1275
rect 443 1207 501 1241
rect 443 1173 455 1207
rect 489 1173 501 1207
rect 443 1139 501 1173
rect 443 1105 455 1139
rect 489 1105 501 1139
rect 443 1071 501 1105
rect 443 1037 455 1071
rect 489 1037 501 1071
rect 443 1003 501 1037
rect 443 969 455 1003
rect 489 969 501 1003
rect 443 935 501 969
rect 443 901 455 935
rect 489 901 501 935
rect 443 867 501 901
rect 443 833 455 867
rect 489 833 501 867
rect 443 799 501 833
rect 443 765 455 799
rect 489 765 501 799
rect 443 731 501 765
rect 443 697 455 731
rect 489 697 501 731
rect 443 663 501 697
rect 443 629 455 663
rect 489 629 501 663
rect 443 595 501 629
rect 443 561 455 595
rect 489 561 501 595
rect 443 527 501 561
rect 443 493 455 527
rect 489 493 501 527
rect 443 459 501 493
rect 443 425 455 459
rect 489 425 501 459
rect 443 391 501 425
rect 443 357 455 391
rect 489 357 501 391
rect 443 323 501 357
rect 443 289 455 323
rect 489 289 501 323
rect 443 255 501 289
rect 443 221 455 255
rect 489 221 501 255
rect 443 187 501 221
rect 443 153 455 187
rect 489 153 501 187
rect 443 119 501 153
rect 443 85 455 119
rect 489 85 501 119
rect 443 51 501 85
rect 443 17 455 51
rect 489 17 501 51
rect 443 -17 501 17
rect 443 -51 455 -17
rect 489 -51 501 -17
rect 443 -85 501 -51
rect 443 -119 455 -85
rect 489 -119 501 -85
rect 443 -153 501 -119
rect 443 -187 455 -153
rect 489 -187 501 -153
rect 443 -221 501 -187
rect 443 -255 455 -221
rect 489 -255 501 -221
rect 443 -289 501 -255
rect 443 -323 455 -289
rect 489 -323 501 -289
rect 443 -357 501 -323
rect 443 -391 455 -357
rect 489 -391 501 -357
rect 443 -425 501 -391
rect 443 -459 455 -425
rect 489 -459 501 -425
rect 443 -493 501 -459
rect 443 -527 455 -493
rect 489 -527 501 -493
rect 443 -561 501 -527
rect 443 -595 455 -561
rect 489 -595 501 -561
rect 443 -629 501 -595
rect 443 -663 455 -629
rect 489 -663 501 -629
rect 443 -697 501 -663
rect 443 -731 455 -697
rect 489 -731 501 -697
rect 443 -765 501 -731
rect 443 -799 455 -765
rect 489 -799 501 -765
rect 443 -833 501 -799
rect 443 -867 455 -833
rect 489 -867 501 -833
rect 443 -901 501 -867
rect 443 -935 455 -901
rect 489 -935 501 -901
rect 443 -969 501 -935
rect 443 -1003 455 -969
rect 489 -1003 501 -969
rect 443 -1037 501 -1003
rect 443 -1071 455 -1037
rect 489 -1071 501 -1037
rect 443 -1105 501 -1071
rect 443 -1139 455 -1105
rect 489 -1139 501 -1105
rect 443 -1173 501 -1139
rect 443 -1207 455 -1173
rect 489 -1207 501 -1173
rect 443 -1241 501 -1207
rect 443 -1275 455 -1241
rect 489 -1275 501 -1241
rect 443 -1309 501 -1275
rect 443 -1343 455 -1309
rect 489 -1343 501 -1309
rect 443 -1377 501 -1343
rect 443 -1411 455 -1377
rect 489 -1411 501 -1377
rect 443 -1445 501 -1411
rect 443 -1479 455 -1445
rect 489 -1479 501 -1445
rect 443 -1513 501 -1479
rect 443 -1547 455 -1513
rect 489 -1547 501 -1513
rect 443 -1581 501 -1547
rect 443 -1615 455 -1581
rect 489 -1615 501 -1581
rect 443 -1649 501 -1615
rect 443 -1683 455 -1649
rect 489 -1683 501 -1649
rect 443 -1717 501 -1683
rect 443 -1751 455 -1717
rect 489 -1751 501 -1717
rect 443 -1785 501 -1751
rect 443 -1819 455 -1785
rect 489 -1819 501 -1785
rect 443 -1853 501 -1819
rect 443 -1887 455 -1853
rect 489 -1887 501 -1853
rect 443 -1921 501 -1887
rect 443 -1955 455 -1921
rect 489 -1955 501 -1921
rect 443 -1989 501 -1955
rect 443 -2023 455 -1989
rect 489 -2023 501 -1989
rect 443 -2057 501 -2023
rect 443 -2091 455 -2057
rect 489 -2091 501 -2057
rect 443 -2125 501 -2091
rect 443 -2159 455 -2125
rect 489 -2159 501 -2125
rect 443 -2193 501 -2159
rect 443 -2227 455 -2193
rect 489 -2227 501 -2193
rect 443 -2261 501 -2227
rect 443 -2295 455 -2261
rect 489 -2295 501 -2261
rect 443 -2329 501 -2295
rect 443 -2363 455 -2329
rect 489 -2363 501 -2329
rect 443 -2397 501 -2363
rect 443 -2431 455 -2397
rect 489 -2431 501 -2397
rect 443 -2465 501 -2431
rect 443 -2499 455 -2465
rect 489 -2499 501 -2465
rect 443 -2533 501 -2499
rect 443 -2567 455 -2533
rect 489 -2567 501 -2533
rect 443 -2601 501 -2567
rect 443 -2635 455 -2601
rect 489 -2635 501 -2601
rect 443 -2669 501 -2635
rect 443 -2703 455 -2669
rect 489 -2703 501 -2669
rect 443 -2737 501 -2703
rect 443 -2771 455 -2737
rect 489 -2771 501 -2737
rect 443 -2805 501 -2771
rect 443 -2839 455 -2805
rect 489 -2839 501 -2805
rect 443 -2873 501 -2839
rect 443 -2907 455 -2873
rect 489 -2907 501 -2873
rect 443 -2941 501 -2907
rect 443 -2975 455 -2941
rect 489 -2975 501 -2941
rect 443 -3009 501 -2975
rect 443 -3043 455 -3009
rect 489 -3043 501 -3009
rect 443 -3077 501 -3043
rect 443 -3111 455 -3077
rect 489 -3111 501 -3077
rect 443 -3145 501 -3111
rect 443 -3179 455 -3145
rect 489 -3179 501 -3145
rect 443 -3213 501 -3179
rect 443 -3247 455 -3213
rect 489 -3247 501 -3213
rect 443 -3281 501 -3247
rect 443 -3315 455 -3281
rect 489 -3315 501 -3281
rect 443 -3349 501 -3315
rect 443 -3383 455 -3349
rect 489 -3383 501 -3349
rect 443 -3417 501 -3383
rect 443 -3451 455 -3417
rect 489 -3451 501 -3417
rect 443 -3485 501 -3451
rect 443 -3519 455 -3485
rect 489 -3519 501 -3485
rect 443 -3553 501 -3519
rect 443 -3587 455 -3553
rect 489 -3587 501 -3553
rect 443 -3621 501 -3587
rect 443 -3655 455 -3621
rect 489 -3655 501 -3621
rect 443 -3689 501 -3655
rect 443 -3723 455 -3689
rect 489 -3723 501 -3689
rect 443 -3757 501 -3723
rect 443 -3791 455 -3757
rect 489 -3791 501 -3757
rect 443 -3825 501 -3791
rect 443 -3859 455 -3825
rect 489 -3859 501 -3825
rect 443 -3893 501 -3859
rect 443 -3927 455 -3893
rect 489 -3927 501 -3893
rect 443 -3961 501 -3927
rect 443 -3995 455 -3961
rect 489 -3995 501 -3961
rect 443 -4029 501 -3995
rect 443 -4063 455 -4029
rect 489 -4063 501 -4029
rect 443 -4097 501 -4063
rect 443 -4131 455 -4097
rect 489 -4131 501 -4097
rect 443 -4165 501 -4131
rect 443 -4199 455 -4165
rect 489 -4199 501 -4165
rect 443 -4233 501 -4199
rect 443 -4267 455 -4233
rect 489 -4267 501 -4233
rect 443 -4301 501 -4267
rect 443 -4335 455 -4301
rect 489 -4335 501 -4301
rect 443 -4369 501 -4335
rect 443 -4403 455 -4369
rect 489 -4403 501 -4369
rect 443 -4437 501 -4403
rect 443 -4471 455 -4437
rect 489 -4471 501 -4437
rect 443 -4505 501 -4471
rect 443 -4539 455 -4505
rect 489 -4539 501 -4505
rect 443 -4573 501 -4539
rect 443 -4607 455 -4573
rect 489 -4607 501 -4573
rect 443 -4641 501 -4607
rect 443 -4675 455 -4641
rect 489 -4675 501 -4641
rect 443 -4709 501 -4675
rect 443 -4743 455 -4709
rect 489 -4743 501 -4709
rect 443 -4777 501 -4743
rect 443 -4811 455 -4777
rect 489 -4811 501 -4777
rect 443 -4845 501 -4811
rect 443 -4879 455 -4845
rect 489 -4879 501 -4845
rect 443 -4913 501 -4879
rect 443 -4947 455 -4913
rect 489 -4947 501 -4913
rect 443 -4981 501 -4947
rect 443 -5015 455 -4981
rect 489 -5015 501 -4981
rect 443 -5049 501 -5015
rect 443 -5083 455 -5049
rect 489 -5083 501 -5049
rect 443 -5117 501 -5083
rect 443 -5151 455 -5117
rect 489 -5151 501 -5117
rect 443 -5185 501 -5151
rect 443 -5219 455 -5185
rect 489 -5219 501 -5185
rect 443 -5253 501 -5219
rect 443 -5287 455 -5253
rect 489 -5287 501 -5253
rect 443 -5321 501 -5287
rect 443 -5355 455 -5321
rect 489 -5355 501 -5321
rect 443 -5389 501 -5355
rect 443 -5423 455 -5389
rect 489 -5423 501 -5389
rect 443 -5457 501 -5423
rect 443 -5491 455 -5457
rect 489 -5491 501 -5457
rect 443 -5525 501 -5491
rect 443 -5559 455 -5525
rect 489 -5559 501 -5525
rect 443 -5593 501 -5559
rect 443 -5627 455 -5593
rect 489 -5627 501 -5593
rect 443 -5661 501 -5627
rect 443 -5695 455 -5661
rect 489 -5695 501 -5661
rect 443 -5729 501 -5695
rect 443 -5763 455 -5729
rect 489 -5763 501 -5729
rect 443 -5797 501 -5763
rect 443 -5831 455 -5797
rect 489 -5831 501 -5797
rect 443 -5865 501 -5831
rect 443 -5899 455 -5865
rect 489 -5899 501 -5865
rect 443 -5933 501 -5899
rect 443 -5967 455 -5933
rect 489 -5967 501 -5933
rect 443 -6000 501 -5967
rect 561 5967 619 6000
rect 561 5933 573 5967
rect 607 5933 619 5967
rect 561 5899 619 5933
rect 561 5865 573 5899
rect 607 5865 619 5899
rect 561 5831 619 5865
rect 561 5797 573 5831
rect 607 5797 619 5831
rect 561 5763 619 5797
rect 561 5729 573 5763
rect 607 5729 619 5763
rect 561 5695 619 5729
rect 561 5661 573 5695
rect 607 5661 619 5695
rect 561 5627 619 5661
rect 561 5593 573 5627
rect 607 5593 619 5627
rect 561 5559 619 5593
rect 561 5525 573 5559
rect 607 5525 619 5559
rect 561 5491 619 5525
rect 561 5457 573 5491
rect 607 5457 619 5491
rect 561 5423 619 5457
rect 561 5389 573 5423
rect 607 5389 619 5423
rect 561 5355 619 5389
rect 561 5321 573 5355
rect 607 5321 619 5355
rect 561 5287 619 5321
rect 561 5253 573 5287
rect 607 5253 619 5287
rect 561 5219 619 5253
rect 561 5185 573 5219
rect 607 5185 619 5219
rect 561 5151 619 5185
rect 561 5117 573 5151
rect 607 5117 619 5151
rect 561 5083 619 5117
rect 561 5049 573 5083
rect 607 5049 619 5083
rect 561 5015 619 5049
rect 561 4981 573 5015
rect 607 4981 619 5015
rect 561 4947 619 4981
rect 561 4913 573 4947
rect 607 4913 619 4947
rect 561 4879 619 4913
rect 561 4845 573 4879
rect 607 4845 619 4879
rect 561 4811 619 4845
rect 561 4777 573 4811
rect 607 4777 619 4811
rect 561 4743 619 4777
rect 561 4709 573 4743
rect 607 4709 619 4743
rect 561 4675 619 4709
rect 561 4641 573 4675
rect 607 4641 619 4675
rect 561 4607 619 4641
rect 561 4573 573 4607
rect 607 4573 619 4607
rect 561 4539 619 4573
rect 561 4505 573 4539
rect 607 4505 619 4539
rect 561 4471 619 4505
rect 561 4437 573 4471
rect 607 4437 619 4471
rect 561 4403 619 4437
rect 561 4369 573 4403
rect 607 4369 619 4403
rect 561 4335 619 4369
rect 561 4301 573 4335
rect 607 4301 619 4335
rect 561 4267 619 4301
rect 561 4233 573 4267
rect 607 4233 619 4267
rect 561 4199 619 4233
rect 561 4165 573 4199
rect 607 4165 619 4199
rect 561 4131 619 4165
rect 561 4097 573 4131
rect 607 4097 619 4131
rect 561 4063 619 4097
rect 561 4029 573 4063
rect 607 4029 619 4063
rect 561 3995 619 4029
rect 561 3961 573 3995
rect 607 3961 619 3995
rect 561 3927 619 3961
rect 561 3893 573 3927
rect 607 3893 619 3927
rect 561 3859 619 3893
rect 561 3825 573 3859
rect 607 3825 619 3859
rect 561 3791 619 3825
rect 561 3757 573 3791
rect 607 3757 619 3791
rect 561 3723 619 3757
rect 561 3689 573 3723
rect 607 3689 619 3723
rect 561 3655 619 3689
rect 561 3621 573 3655
rect 607 3621 619 3655
rect 561 3587 619 3621
rect 561 3553 573 3587
rect 607 3553 619 3587
rect 561 3519 619 3553
rect 561 3485 573 3519
rect 607 3485 619 3519
rect 561 3451 619 3485
rect 561 3417 573 3451
rect 607 3417 619 3451
rect 561 3383 619 3417
rect 561 3349 573 3383
rect 607 3349 619 3383
rect 561 3315 619 3349
rect 561 3281 573 3315
rect 607 3281 619 3315
rect 561 3247 619 3281
rect 561 3213 573 3247
rect 607 3213 619 3247
rect 561 3179 619 3213
rect 561 3145 573 3179
rect 607 3145 619 3179
rect 561 3111 619 3145
rect 561 3077 573 3111
rect 607 3077 619 3111
rect 561 3043 619 3077
rect 561 3009 573 3043
rect 607 3009 619 3043
rect 561 2975 619 3009
rect 561 2941 573 2975
rect 607 2941 619 2975
rect 561 2907 619 2941
rect 561 2873 573 2907
rect 607 2873 619 2907
rect 561 2839 619 2873
rect 561 2805 573 2839
rect 607 2805 619 2839
rect 561 2771 619 2805
rect 561 2737 573 2771
rect 607 2737 619 2771
rect 561 2703 619 2737
rect 561 2669 573 2703
rect 607 2669 619 2703
rect 561 2635 619 2669
rect 561 2601 573 2635
rect 607 2601 619 2635
rect 561 2567 619 2601
rect 561 2533 573 2567
rect 607 2533 619 2567
rect 561 2499 619 2533
rect 561 2465 573 2499
rect 607 2465 619 2499
rect 561 2431 619 2465
rect 561 2397 573 2431
rect 607 2397 619 2431
rect 561 2363 619 2397
rect 561 2329 573 2363
rect 607 2329 619 2363
rect 561 2295 619 2329
rect 561 2261 573 2295
rect 607 2261 619 2295
rect 561 2227 619 2261
rect 561 2193 573 2227
rect 607 2193 619 2227
rect 561 2159 619 2193
rect 561 2125 573 2159
rect 607 2125 619 2159
rect 561 2091 619 2125
rect 561 2057 573 2091
rect 607 2057 619 2091
rect 561 2023 619 2057
rect 561 1989 573 2023
rect 607 1989 619 2023
rect 561 1955 619 1989
rect 561 1921 573 1955
rect 607 1921 619 1955
rect 561 1887 619 1921
rect 561 1853 573 1887
rect 607 1853 619 1887
rect 561 1819 619 1853
rect 561 1785 573 1819
rect 607 1785 619 1819
rect 561 1751 619 1785
rect 561 1717 573 1751
rect 607 1717 619 1751
rect 561 1683 619 1717
rect 561 1649 573 1683
rect 607 1649 619 1683
rect 561 1615 619 1649
rect 561 1581 573 1615
rect 607 1581 619 1615
rect 561 1547 619 1581
rect 561 1513 573 1547
rect 607 1513 619 1547
rect 561 1479 619 1513
rect 561 1445 573 1479
rect 607 1445 619 1479
rect 561 1411 619 1445
rect 561 1377 573 1411
rect 607 1377 619 1411
rect 561 1343 619 1377
rect 561 1309 573 1343
rect 607 1309 619 1343
rect 561 1275 619 1309
rect 561 1241 573 1275
rect 607 1241 619 1275
rect 561 1207 619 1241
rect 561 1173 573 1207
rect 607 1173 619 1207
rect 561 1139 619 1173
rect 561 1105 573 1139
rect 607 1105 619 1139
rect 561 1071 619 1105
rect 561 1037 573 1071
rect 607 1037 619 1071
rect 561 1003 619 1037
rect 561 969 573 1003
rect 607 969 619 1003
rect 561 935 619 969
rect 561 901 573 935
rect 607 901 619 935
rect 561 867 619 901
rect 561 833 573 867
rect 607 833 619 867
rect 561 799 619 833
rect 561 765 573 799
rect 607 765 619 799
rect 561 731 619 765
rect 561 697 573 731
rect 607 697 619 731
rect 561 663 619 697
rect 561 629 573 663
rect 607 629 619 663
rect 561 595 619 629
rect 561 561 573 595
rect 607 561 619 595
rect 561 527 619 561
rect 561 493 573 527
rect 607 493 619 527
rect 561 459 619 493
rect 561 425 573 459
rect 607 425 619 459
rect 561 391 619 425
rect 561 357 573 391
rect 607 357 619 391
rect 561 323 619 357
rect 561 289 573 323
rect 607 289 619 323
rect 561 255 619 289
rect 561 221 573 255
rect 607 221 619 255
rect 561 187 619 221
rect 561 153 573 187
rect 607 153 619 187
rect 561 119 619 153
rect 561 85 573 119
rect 607 85 619 119
rect 561 51 619 85
rect 561 17 573 51
rect 607 17 619 51
rect 561 -17 619 17
rect 561 -51 573 -17
rect 607 -51 619 -17
rect 561 -85 619 -51
rect 561 -119 573 -85
rect 607 -119 619 -85
rect 561 -153 619 -119
rect 561 -187 573 -153
rect 607 -187 619 -153
rect 561 -221 619 -187
rect 561 -255 573 -221
rect 607 -255 619 -221
rect 561 -289 619 -255
rect 561 -323 573 -289
rect 607 -323 619 -289
rect 561 -357 619 -323
rect 561 -391 573 -357
rect 607 -391 619 -357
rect 561 -425 619 -391
rect 561 -459 573 -425
rect 607 -459 619 -425
rect 561 -493 619 -459
rect 561 -527 573 -493
rect 607 -527 619 -493
rect 561 -561 619 -527
rect 561 -595 573 -561
rect 607 -595 619 -561
rect 561 -629 619 -595
rect 561 -663 573 -629
rect 607 -663 619 -629
rect 561 -697 619 -663
rect 561 -731 573 -697
rect 607 -731 619 -697
rect 561 -765 619 -731
rect 561 -799 573 -765
rect 607 -799 619 -765
rect 561 -833 619 -799
rect 561 -867 573 -833
rect 607 -867 619 -833
rect 561 -901 619 -867
rect 561 -935 573 -901
rect 607 -935 619 -901
rect 561 -969 619 -935
rect 561 -1003 573 -969
rect 607 -1003 619 -969
rect 561 -1037 619 -1003
rect 561 -1071 573 -1037
rect 607 -1071 619 -1037
rect 561 -1105 619 -1071
rect 561 -1139 573 -1105
rect 607 -1139 619 -1105
rect 561 -1173 619 -1139
rect 561 -1207 573 -1173
rect 607 -1207 619 -1173
rect 561 -1241 619 -1207
rect 561 -1275 573 -1241
rect 607 -1275 619 -1241
rect 561 -1309 619 -1275
rect 561 -1343 573 -1309
rect 607 -1343 619 -1309
rect 561 -1377 619 -1343
rect 561 -1411 573 -1377
rect 607 -1411 619 -1377
rect 561 -1445 619 -1411
rect 561 -1479 573 -1445
rect 607 -1479 619 -1445
rect 561 -1513 619 -1479
rect 561 -1547 573 -1513
rect 607 -1547 619 -1513
rect 561 -1581 619 -1547
rect 561 -1615 573 -1581
rect 607 -1615 619 -1581
rect 561 -1649 619 -1615
rect 561 -1683 573 -1649
rect 607 -1683 619 -1649
rect 561 -1717 619 -1683
rect 561 -1751 573 -1717
rect 607 -1751 619 -1717
rect 561 -1785 619 -1751
rect 561 -1819 573 -1785
rect 607 -1819 619 -1785
rect 561 -1853 619 -1819
rect 561 -1887 573 -1853
rect 607 -1887 619 -1853
rect 561 -1921 619 -1887
rect 561 -1955 573 -1921
rect 607 -1955 619 -1921
rect 561 -1989 619 -1955
rect 561 -2023 573 -1989
rect 607 -2023 619 -1989
rect 561 -2057 619 -2023
rect 561 -2091 573 -2057
rect 607 -2091 619 -2057
rect 561 -2125 619 -2091
rect 561 -2159 573 -2125
rect 607 -2159 619 -2125
rect 561 -2193 619 -2159
rect 561 -2227 573 -2193
rect 607 -2227 619 -2193
rect 561 -2261 619 -2227
rect 561 -2295 573 -2261
rect 607 -2295 619 -2261
rect 561 -2329 619 -2295
rect 561 -2363 573 -2329
rect 607 -2363 619 -2329
rect 561 -2397 619 -2363
rect 561 -2431 573 -2397
rect 607 -2431 619 -2397
rect 561 -2465 619 -2431
rect 561 -2499 573 -2465
rect 607 -2499 619 -2465
rect 561 -2533 619 -2499
rect 561 -2567 573 -2533
rect 607 -2567 619 -2533
rect 561 -2601 619 -2567
rect 561 -2635 573 -2601
rect 607 -2635 619 -2601
rect 561 -2669 619 -2635
rect 561 -2703 573 -2669
rect 607 -2703 619 -2669
rect 561 -2737 619 -2703
rect 561 -2771 573 -2737
rect 607 -2771 619 -2737
rect 561 -2805 619 -2771
rect 561 -2839 573 -2805
rect 607 -2839 619 -2805
rect 561 -2873 619 -2839
rect 561 -2907 573 -2873
rect 607 -2907 619 -2873
rect 561 -2941 619 -2907
rect 561 -2975 573 -2941
rect 607 -2975 619 -2941
rect 561 -3009 619 -2975
rect 561 -3043 573 -3009
rect 607 -3043 619 -3009
rect 561 -3077 619 -3043
rect 561 -3111 573 -3077
rect 607 -3111 619 -3077
rect 561 -3145 619 -3111
rect 561 -3179 573 -3145
rect 607 -3179 619 -3145
rect 561 -3213 619 -3179
rect 561 -3247 573 -3213
rect 607 -3247 619 -3213
rect 561 -3281 619 -3247
rect 561 -3315 573 -3281
rect 607 -3315 619 -3281
rect 561 -3349 619 -3315
rect 561 -3383 573 -3349
rect 607 -3383 619 -3349
rect 561 -3417 619 -3383
rect 561 -3451 573 -3417
rect 607 -3451 619 -3417
rect 561 -3485 619 -3451
rect 561 -3519 573 -3485
rect 607 -3519 619 -3485
rect 561 -3553 619 -3519
rect 561 -3587 573 -3553
rect 607 -3587 619 -3553
rect 561 -3621 619 -3587
rect 561 -3655 573 -3621
rect 607 -3655 619 -3621
rect 561 -3689 619 -3655
rect 561 -3723 573 -3689
rect 607 -3723 619 -3689
rect 561 -3757 619 -3723
rect 561 -3791 573 -3757
rect 607 -3791 619 -3757
rect 561 -3825 619 -3791
rect 561 -3859 573 -3825
rect 607 -3859 619 -3825
rect 561 -3893 619 -3859
rect 561 -3927 573 -3893
rect 607 -3927 619 -3893
rect 561 -3961 619 -3927
rect 561 -3995 573 -3961
rect 607 -3995 619 -3961
rect 561 -4029 619 -3995
rect 561 -4063 573 -4029
rect 607 -4063 619 -4029
rect 561 -4097 619 -4063
rect 561 -4131 573 -4097
rect 607 -4131 619 -4097
rect 561 -4165 619 -4131
rect 561 -4199 573 -4165
rect 607 -4199 619 -4165
rect 561 -4233 619 -4199
rect 561 -4267 573 -4233
rect 607 -4267 619 -4233
rect 561 -4301 619 -4267
rect 561 -4335 573 -4301
rect 607 -4335 619 -4301
rect 561 -4369 619 -4335
rect 561 -4403 573 -4369
rect 607 -4403 619 -4369
rect 561 -4437 619 -4403
rect 561 -4471 573 -4437
rect 607 -4471 619 -4437
rect 561 -4505 619 -4471
rect 561 -4539 573 -4505
rect 607 -4539 619 -4505
rect 561 -4573 619 -4539
rect 561 -4607 573 -4573
rect 607 -4607 619 -4573
rect 561 -4641 619 -4607
rect 561 -4675 573 -4641
rect 607 -4675 619 -4641
rect 561 -4709 619 -4675
rect 561 -4743 573 -4709
rect 607 -4743 619 -4709
rect 561 -4777 619 -4743
rect 561 -4811 573 -4777
rect 607 -4811 619 -4777
rect 561 -4845 619 -4811
rect 561 -4879 573 -4845
rect 607 -4879 619 -4845
rect 561 -4913 619 -4879
rect 561 -4947 573 -4913
rect 607 -4947 619 -4913
rect 561 -4981 619 -4947
rect 561 -5015 573 -4981
rect 607 -5015 619 -4981
rect 561 -5049 619 -5015
rect 561 -5083 573 -5049
rect 607 -5083 619 -5049
rect 561 -5117 619 -5083
rect 561 -5151 573 -5117
rect 607 -5151 619 -5117
rect 561 -5185 619 -5151
rect 561 -5219 573 -5185
rect 607 -5219 619 -5185
rect 561 -5253 619 -5219
rect 561 -5287 573 -5253
rect 607 -5287 619 -5253
rect 561 -5321 619 -5287
rect 561 -5355 573 -5321
rect 607 -5355 619 -5321
rect 561 -5389 619 -5355
rect 561 -5423 573 -5389
rect 607 -5423 619 -5389
rect 561 -5457 619 -5423
rect 561 -5491 573 -5457
rect 607 -5491 619 -5457
rect 561 -5525 619 -5491
rect 561 -5559 573 -5525
rect 607 -5559 619 -5525
rect 561 -5593 619 -5559
rect 561 -5627 573 -5593
rect 607 -5627 619 -5593
rect 561 -5661 619 -5627
rect 561 -5695 573 -5661
rect 607 -5695 619 -5661
rect 561 -5729 619 -5695
rect 561 -5763 573 -5729
rect 607 -5763 619 -5729
rect 561 -5797 619 -5763
rect 561 -5831 573 -5797
rect 607 -5831 619 -5797
rect 561 -5865 619 -5831
rect 561 -5899 573 -5865
rect 607 -5899 619 -5865
rect 561 -5933 619 -5899
rect 561 -5967 573 -5933
rect 607 -5967 619 -5933
rect 561 -6000 619 -5967
<< ndiffc >>
rect -607 5933 -573 5967
rect -607 5865 -573 5899
rect -607 5797 -573 5831
rect -607 5729 -573 5763
rect -607 5661 -573 5695
rect -607 5593 -573 5627
rect -607 5525 -573 5559
rect -607 5457 -573 5491
rect -607 5389 -573 5423
rect -607 5321 -573 5355
rect -607 5253 -573 5287
rect -607 5185 -573 5219
rect -607 5117 -573 5151
rect -607 5049 -573 5083
rect -607 4981 -573 5015
rect -607 4913 -573 4947
rect -607 4845 -573 4879
rect -607 4777 -573 4811
rect -607 4709 -573 4743
rect -607 4641 -573 4675
rect -607 4573 -573 4607
rect -607 4505 -573 4539
rect -607 4437 -573 4471
rect -607 4369 -573 4403
rect -607 4301 -573 4335
rect -607 4233 -573 4267
rect -607 4165 -573 4199
rect -607 4097 -573 4131
rect -607 4029 -573 4063
rect -607 3961 -573 3995
rect -607 3893 -573 3927
rect -607 3825 -573 3859
rect -607 3757 -573 3791
rect -607 3689 -573 3723
rect -607 3621 -573 3655
rect -607 3553 -573 3587
rect -607 3485 -573 3519
rect -607 3417 -573 3451
rect -607 3349 -573 3383
rect -607 3281 -573 3315
rect -607 3213 -573 3247
rect -607 3145 -573 3179
rect -607 3077 -573 3111
rect -607 3009 -573 3043
rect -607 2941 -573 2975
rect -607 2873 -573 2907
rect -607 2805 -573 2839
rect -607 2737 -573 2771
rect -607 2669 -573 2703
rect -607 2601 -573 2635
rect -607 2533 -573 2567
rect -607 2465 -573 2499
rect -607 2397 -573 2431
rect -607 2329 -573 2363
rect -607 2261 -573 2295
rect -607 2193 -573 2227
rect -607 2125 -573 2159
rect -607 2057 -573 2091
rect -607 1989 -573 2023
rect -607 1921 -573 1955
rect -607 1853 -573 1887
rect -607 1785 -573 1819
rect -607 1717 -573 1751
rect -607 1649 -573 1683
rect -607 1581 -573 1615
rect -607 1513 -573 1547
rect -607 1445 -573 1479
rect -607 1377 -573 1411
rect -607 1309 -573 1343
rect -607 1241 -573 1275
rect -607 1173 -573 1207
rect -607 1105 -573 1139
rect -607 1037 -573 1071
rect -607 969 -573 1003
rect -607 901 -573 935
rect -607 833 -573 867
rect -607 765 -573 799
rect -607 697 -573 731
rect -607 629 -573 663
rect -607 561 -573 595
rect -607 493 -573 527
rect -607 425 -573 459
rect -607 357 -573 391
rect -607 289 -573 323
rect -607 221 -573 255
rect -607 153 -573 187
rect -607 85 -573 119
rect -607 17 -573 51
rect -607 -51 -573 -17
rect -607 -119 -573 -85
rect -607 -187 -573 -153
rect -607 -255 -573 -221
rect -607 -323 -573 -289
rect -607 -391 -573 -357
rect -607 -459 -573 -425
rect -607 -527 -573 -493
rect -607 -595 -573 -561
rect -607 -663 -573 -629
rect -607 -731 -573 -697
rect -607 -799 -573 -765
rect -607 -867 -573 -833
rect -607 -935 -573 -901
rect -607 -1003 -573 -969
rect -607 -1071 -573 -1037
rect -607 -1139 -573 -1105
rect -607 -1207 -573 -1173
rect -607 -1275 -573 -1241
rect -607 -1343 -573 -1309
rect -607 -1411 -573 -1377
rect -607 -1479 -573 -1445
rect -607 -1547 -573 -1513
rect -607 -1615 -573 -1581
rect -607 -1683 -573 -1649
rect -607 -1751 -573 -1717
rect -607 -1819 -573 -1785
rect -607 -1887 -573 -1853
rect -607 -1955 -573 -1921
rect -607 -2023 -573 -1989
rect -607 -2091 -573 -2057
rect -607 -2159 -573 -2125
rect -607 -2227 -573 -2193
rect -607 -2295 -573 -2261
rect -607 -2363 -573 -2329
rect -607 -2431 -573 -2397
rect -607 -2499 -573 -2465
rect -607 -2567 -573 -2533
rect -607 -2635 -573 -2601
rect -607 -2703 -573 -2669
rect -607 -2771 -573 -2737
rect -607 -2839 -573 -2805
rect -607 -2907 -573 -2873
rect -607 -2975 -573 -2941
rect -607 -3043 -573 -3009
rect -607 -3111 -573 -3077
rect -607 -3179 -573 -3145
rect -607 -3247 -573 -3213
rect -607 -3315 -573 -3281
rect -607 -3383 -573 -3349
rect -607 -3451 -573 -3417
rect -607 -3519 -573 -3485
rect -607 -3587 -573 -3553
rect -607 -3655 -573 -3621
rect -607 -3723 -573 -3689
rect -607 -3791 -573 -3757
rect -607 -3859 -573 -3825
rect -607 -3927 -573 -3893
rect -607 -3995 -573 -3961
rect -607 -4063 -573 -4029
rect -607 -4131 -573 -4097
rect -607 -4199 -573 -4165
rect -607 -4267 -573 -4233
rect -607 -4335 -573 -4301
rect -607 -4403 -573 -4369
rect -607 -4471 -573 -4437
rect -607 -4539 -573 -4505
rect -607 -4607 -573 -4573
rect -607 -4675 -573 -4641
rect -607 -4743 -573 -4709
rect -607 -4811 -573 -4777
rect -607 -4879 -573 -4845
rect -607 -4947 -573 -4913
rect -607 -5015 -573 -4981
rect -607 -5083 -573 -5049
rect -607 -5151 -573 -5117
rect -607 -5219 -573 -5185
rect -607 -5287 -573 -5253
rect -607 -5355 -573 -5321
rect -607 -5423 -573 -5389
rect -607 -5491 -573 -5457
rect -607 -5559 -573 -5525
rect -607 -5627 -573 -5593
rect -607 -5695 -573 -5661
rect -607 -5763 -573 -5729
rect -607 -5831 -573 -5797
rect -607 -5899 -573 -5865
rect -607 -5967 -573 -5933
rect -489 5933 -455 5967
rect -489 5865 -455 5899
rect -489 5797 -455 5831
rect -489 5729 -455 5763
rect -489 5661 -455 5695
rect -489 5593 -455 5627
rect -489 5525 -455 5559
rect -489 5457 -455 5491
rect -489 5389 -455 5423
rect -489 5321 -455 5355
rect -489 5253 -455 5287
rect -489 5185 -455 5219
rect -489 5117 -455 5151
rect -489 5049 -455 5083
rect -489 4981 -455 5015
rect -489 4913 -455 4947
rect -489 4845 -455 4879
rect -489 4777 -455 4811
rect -489 4709 -455 4743
rect -489 4641 -455 4675
rect -489 4573 -455 4607
rect -489 4505 -455 4539
rect -489 4437 -455 4471
rect -489 4369 -455 4403
rect -489 4301 -455 4335
rect -489 4233 -455 4267
rect -489 4165 -455 4199
rect -489 4097 -455 4131
rect -489 4029 -455 4063
rect -489 3961 -455 3995
rect -489 3893 -455 3927
rect -489 3825 -455 3859
rect -489 3757 -455 3791
rect -489 3689 -455 3723
rect -489 3621 -455 3655
rect -489 3553 -455 3587
rect -489 3485 -455 3519
rect -489 3417 -455 3451
rect -489 3349 -455 3383
rect -489 3281 -455 3315
rect -489 3213 -455 3247
rect -489 3145 -455 3179
rect -489 3077 -455 3111
rect -489 3009 -455 3043
rect -489 2941 -455 2975
rect -489 2873 -455 2907
rect -489 2805 -455 2839
rect -489 2737 -455 2771
rect -489 2669 -455 2703
rect -489 2601 -455 2635
rect -489 2533 -455 2567
rect -489 2465 -455 2499
rect -489 2397 -455 2431
rect -489 2329 -455 2363
rect -489 2261 -455 2295
rect -489 2193 -455 2227
rect -489 2125 -455 2159
rect -489 2057 -455 2091
rect -489 1989 -455 2023
rect -489 1921 -455 1955
rect -489 1853 -455 1887
rect -489 1785 -455 1819
rect -489 1717 -455 1751
rect -489 1649 -455 1683
rect -489 1581 -455 1615
rect -489 1513 -455 1547
rect -489 1445 -455 1479
rect -489 1377 -455 1411
rect -489 1309 -455 1343
rect -489 1241 -455 1275
rect -489 1173 -455 1207
rect -489 1105 -455 1139
rect -489 1037 -455 1071
rect -489 969 -455 1003
rect -489 901 -455 935
rect -489 833 -455 867
rect -489 765 -455 799
rect -489 697 -455 731
rect -489 629 -455 663
rect -489 561 -455 595
rect -489 493 -455 527
rect -489 425 -455 459
rect -489 357 -455 391
rect -489 289 -455 323
rect -489 221 -455 255
rect -489 153 -455 187
rect -489 85 -455 119
rect -489 17 -455 51
rect -489 -51 -455 -17
rect -489 -119 -455 -85
rect -489 -187 -455 -153
rect -489 -255 -455 -221
rect -489 -323 -455 -289
rect -489 -391 -455 -357
rect -489 -459 -455 -425
rect -489 -527 -455 -493
rect -489 -595 -455 -561
rect -489 -663 -455 -629
rect -489 -731 -455 -697
rect -489 -799 -455 -765
rect -489 -867 -455 -833
rect -489 -935 -455 -901
rect -489 -1003 -455 -969
rect -489 -1071 -455 -1037
rect -489 -1139 -455 -1105
rect -489 -1207 -455 -1173
rect -489 -1275 -455 -1241
rect -489 -1343 -455 -1309
rect -489 -1411 -455 -1377
rect -489 -1479 -455 -1445
rect -489 -1547 -455 -1513
rect -489 -1615 -455 -1581
rect -489 -1683 -455 -1649
rect -489 -1751 -455 -1717
rect -489 -1819 -455 -1785
rect -489 -1887 -455 -1853
rect -489 -1955 -455 -1921
rect -489 -2023 -455 -1989
rect -489 -2091 -455 -2057
rect -489 -2159 -455 -2125
rect -489 -2227 -455 -2193
rect -489 -2295 -455 -2261
rect -489 -2363 -455 -2329
rect -489 -2431 -455 -2397
rect -489 -2499 -455 -2465
rect -489 -2567 -455 -2533
rect -489 -2635 -455 -2601
rect -489 -2703 -455 -2669
rect -489 -2771 -455 -2737
rect -489 -2839 -455 -2805
rect -489 -2907 -455 -2873
rect -489 -2975 -455 -2941
rect -489 -3043 -455 -3009
rect -489 -3111 -455 -3077
rect -489 -3179 -455 -3145
rect -489 -3247 -455 -3213
rect -489 -3315 -455 -3281
rect -489 -3383 -455 -3349
rect -489 -3451 -455 -3417
rect -489 -3519 -455 -3485
rect -489 -3587 -455 -3553
rect -489 -3655 -455 -3621
rect -489 -3723 -455 -3689
rect -489 -3791 -455 -3757
rect -489 -3859 -455 -3825
rect -489 -3927 -455 -3893
rect -489 -3995 -455 -3961
rect -489 -4063 -455 -4029
rect -489 -4131 -455 -4097
rect -489 -4199 -455 -4165
rect -489 -4267 -455 -4233
rect -489 -4335 -455 -4301
rect -489 -4403 -455 -4369
rect -489 -4471 -455 -4437
rect -489 -4539 -455 -4505
rect -489 -4607 -455 -4573
rect -489 -4675 -455 -4641
rect -489 -4743 -455 -4709
rect -489 -4811 -455 -4777
rect -489 -4879 -455 -4845
rect -489 -4947 -455 -4913
rect -489 -5015 -455 -4981
rect -489 -5083 -455 -5049
rect -489 -5151 -455 -5117
rect -489 -5219 -455 -5185
rect -489 -5287 -455 -5253
rect -489 -5355 -455 -5321
rect -489 -5423 -455 -5389
rect -489 -5491 -455 -5457
rect -489 -5559 -455 -5525
rect -489 -5627 -455 -5593
rect -489 -5695 -455 -5661
rect -489 -5763 -455 -5729
rect -489 -5831 -455 -5797
rect -489 -5899 -455 -5865
rect -489 -5967 -455 -5933
rect -371 5933 -337 5967
rect -371 5865 -337 5899
rect -371 5797 -337 5831
rect -371 5729 -337 5763
rect -371 5661 -337 5695
rect -371 5593 -337 5627
rect -371 5525 -337 5559
rect -371 5457 -337 5491
rect -371 5389 -337 5423
rect -371 5321 -337 5355
rect -371 5253 -337 5287
rect -371 5185 -337 5219
rect -371 5117 -337 5151
rect -371 5049 -337 5083
rect -371 4981 -337 5015
rect -371 4913 -337 4947
rect -371 4845 -337 4879
rect -371 4777 -337 4811
rect -371 4709 -337 4743
rect -371 4641 -337 4675
rect -371 4573 -337 4607
rect -371 4505 -337 4539
rect -371 4437 -337 4471
rect -371 4369 -337 4403
rect -371 4301 -337 4335
rect -371 4233 -337 4267
rect -371 4165 -337 4199
rect -371 4097 -337 4131
rect -371 4029 -337 4063
rect -371 3961 -337 3995
rect -371 3893 -337 3927
rect -371 3825 -337 3859
rect -371 3757 -337 3791
rect -371 3689 -337 3723
rect -371 3621 -337 3655
rect -371 3553 -337 3587
rect -371 3485 -337 3519
rect -371 3417 -337 3451
rect -371 3349 -337 3383
rect -371 3281 -337 3315
rect -371 3213 -337 3247
rect -371 3145 -337 3179
rect -371 3077 -337 3111
rect -371 3009 -337 3043
rect -371 2941 -337 2975
rect -371 2873 -337 2907
rect -371 2805 -337 2839
rect -371 2737 -337 2771
rect -371 2669 -337 2703
rect -371 2601 -337 2635
rect -371 2533 -337 2567
rect -371 2465 -337 2499
rect -371 2397 -337 2431
rect -371 2329 -337 2363
rect -371 2261 -337 2295
rect -371 2193 -337 2227
rect -371 2125 -337 2159
rect -371 2057 -337 2091
rect -371 1989 -337 2023
rect -371 1921 -337 1955
rect -371 1853 -337 1887
rect -371 1785 -337 1819
rect -371 1717 -337 1751
rect -371 1649 -337 1683
rect -371 1581 -337 1615
rect -371 1513 -337 1547
rect -371 1445 -337 1479
rect -371 1377 -337 1411
rect -371 1309 -337 1343
rect -371 1241 -337 1275
rect -371 1173 -337 1207
rect -371 1105 -337 1139
rect -371 1037 -337 1071
rect -371 969 -337 1003
rect -371 901 -337 935
rect -371 833 -337 867
rect -371 765 -337 799
rect -371 697 -337 731
rect -371 629 -337 663
rect -371 561 -337 595
rect -371 493 -337 527
rect -371 425 -337 459
rect -371 357 -337 391
rect -371 289 -337 323
rect -371 221 -337 255
rect -371 153 -337 187
rect -371 85 -337 119
rect -371 17 -337 51
rect -371 -51 -337 -17
rect -371 -119 -337 -85
rect -371 -187 -337 -153
rect -371 -255 -337 -221
rect -371 -323 -337 -289
rect -371 -391 -337 -357
rect -371 -459 -337 -425
rect -371 -527 -337 -493
rect -371 -595 -337 -561
rect -371 -663 -337 -629
rect -371 -731 -337 -697
rect -371 -799 -337 -765
rect -371 -867 -337 -833
rect -371 -935 -337 -901
rect -371 -1003 -337 -969
rect -371 -1071 -337 -1037
rect -371 -1139 -337 -1105
rect -371 -1207 -337 -1173
rect -371 -1275 -337 -1241
rect -371 -1343 -337 -1309
rect -371 -1411 -337 -1377
rect -371 -1479 -337 -1445
rect -371 -1547 -337 -1513
rect -371 -1615 -337 -1581
rect -371 -1683 -337 -1649
rect -371 -1751 -337 -1717
rect -371 -1819 -337 -1785
rect -371 -1887 -337 -1853
rect -371 -1955 -337 -1921
rect -371 -2023 -337 -1989
rect -371 -2091 -337 -2057
rect -371 -2159 -337 -2125
rect -371 -2227 -337 -2193
rect -371 -2295 -337 -2261
rect -371 -2363 -337 -2329
rect -371 -2431 -337 -2397
rect -371 -2499 -337 -2465
rect -371 -2567 -337 -2533
rect -371 -2635 -337 -2601
rect -371 -2703 -337 -2669
rect -371 -2771 -337 -2737
rect -371 -2839 -337 -2805
rect -371 -2907 -337 -2873
rect -371 -2975 -337 -2941
rect -371 -3043 -337 -3009
rect -371 -3111 -337 -3077
rect -371 -3179 -337 -3145
rect -371 -3247 -337 -3213
rect -371 -3315 -337 -3281
rect -371 -3383 -337 -3349
rect -371 -3451 -337 -3417
rect -371 -3519 -337 -3485
rect -371 -3587 -337 -3553
rect -371 -3655 -337 -3621
rect -371 -3723 -337 -3689
rect -371 -3791 -337 -3757
rect -371 -3859 -337 -3825
rect -371 -3927 -337 -3893
rect -371 -3995 -337 -3961
rect -371 -4063 -337 -4029
rect -371 -4131 -337 -4097
rect -371 -4199 -337 -4165
rect -371 -4267 -337 -4233
rect -371 -4335 -337 -4301
rect -371 -4403 -337 -4369
rect -371 -4471 -337 -4437
rect -371 -4539 -337 -4505
rect -371 -4607 -337 -4573
rect -371 -4675 -337 -4641
rect -371 -4743 -337 -4709
rect -371 -4811 -337 -4777
rect -371 -4879 -337 -4845
rect -371 -4947 -337 -4913
rect -371 -5015 -337 -4981
rect -371 -5083 -337 -5049
rect -371 -5151 -337 -5117
rect -371 -5219 -337 -5185
rect -371 -5287 -337 -5253
rect -371 -5355 -337 -5321
rect -371 -5423 -337 -5389
rect -371 -5491 -337 -5457
rect -371 -5559 -337 -5525
rect -371 -5627 -337 -5593
rect -371 -5695 -337 -5661
rect -371 -5763 -337 -5729
rect -371 -5831 -337 -5797
rect -371 -5899 -337 -5865
rect -371 -5967 -337 -5933
rect -253 5933 -219 5967
rect -253 5865 -219 5899
rect -253 5797 -219 5831
rect -253 5729 -219 5763
rect -253 5661 -219 5695
rect -253 5593 -219 5627
rect -253 5525 -219 5559
rect -253 5457 -219 5491
rect -253 5389 -219 5423
rect -253 5321 -219 5355
rect -253 5253 -219 5287
rect -253 5185 -219 5219
rect -253 5117 -219 5151
rect -253 5049 -219 5083
rect -253 4981 -219 5015
rect -253 4913 -219 4947
rect -253 4845 -219 4879
rect -253 4777 -219 4811
rect -253 4709 -219 4743
rect -253 4641 -219 4675
rect -253 4573 -219 4607
rect -253 4505 -219 4539
rect -253 4437 -219 4471
rect -253 4369 -219 4403
rect -253 4301 -219 4335
rect -253 4233 -219 4267
rect -253 4165 -219 4199
rect -253 4097 -219 4131
rect -253 4029 -219 4063
rect -253 3961 -219 3995
rect -253 3893 -219 3927
rect -253 3825 -219 3859
rect -253 3757 -219 3791
rect -253 3689 -219 3723
rect -253 3621 -219 3655
rect -253 3553 -219 3587
rect -253 3485 -219 3519
rect -253 3417 -219 3451
rect -253 3349 -219 3383
rect -253 3281 -219 3315
rect -253 3213 -219 3247
rect -253 3145 -219 3179
rect -253 3077 -219 3111
rect -253 3009 -219 3043
rect -253 2941 -219 2975
rect -253 2873 -219 2907
rect -253 2805 -219 2839
rect -253 2737 -219 2771
rect -253 2669 -219 2703
rect -253 2601 -219 2635
rect -253 2533 -219 2567
rect -253 2465 -219 2499
rect -253 2397 -219 2431
rect -253 2329 -219 2363
rect -253 2261 -219 2295
rect -253 2193 -219 2227
rect -253 2125 -219 2159
rect -253 2057 -219 2091
rect -253 1989 -219 2023
rect -253 1921 -219 1955
rect -253 1853 -219 1887
rect -253 1785 -219 1819
rect -253 1717 -219 1751
rect -253 1649 -219 1683
rect -253 1581 -219 1615
rect -253 1513 -219 1547
rect -253 1445 -219 1479
rect -253 1377 -219 1411
rect -253 1309 -219 1343
rect -253 1241 -219 1275
rect -253 1173 -219 1207
rect -253 1105 -219 1139
rect -253 1037 -219 1071
rect -253 969 -219 1003
rect -253 901 -219 935
rect -253 833 -219 867
rect -253 765 -219 799
rect -253 697 -219 731
rect -253 629 -219 663
rect -253 561 -219 595
rect -253 493 -219 527
rect -253 425 -219 459
rect -253 357 -219 391
rect -253 289 -219 323
rect -253 221 -219 255
rect -253 153 -219 187
rect -253 85 -219 119
rect -253 17 -219 51
rect -253 -51 -219 -17
rect -253 -119 -219 -85
rect -253 -187 -219 -153
rect -253 -255 -219 -221
rect -253 -323 -219 -289
rect -253 -391 -219 -357
rect -253 -459 -219 -425
rect -253 -527 -219 -493
rect -253 -595 -219 -561
rect -253 -663 -219 -629
rect -253 -731 -219 -697
rect -253 -799 -219 -765
rect -253 -867 -219 -833
rect -253 -935 -219 -901
rect -253 -1003 -219 -969
rect -253 -1071 -219 -1037
rect -253 -1139 -219 -1105
rect -253 -1207 -219 -1173
rect -253 -1275 -219 -1241
rect -253 -1343 -219 -1309
rect -253 -1411 -219 -1377
rect -253 -1479 -219 -1445
rect -253 -1547 -219 -1513
rect -253 -1615 -219 -1581
rect -253 -1683 -219 -1649
rect -253 -1751 -219 -1717
rect -253 -1819 -219 -1785
rect -253 -1887 -219 -1853
rect -253 -1955 -219 -1921
rect -253 -2023 -219 -1989
rect -253 -2091 -219 -2057
rect -253 -2159 -219 -2125
rect -253 -2227 -219 -2193
rect -253 -2295 -219 -2261
rect -253 -2363 -219 -2329
rect -253 -2431 -219 -2397
rect -253 -2499 -219 -2465
rect -253 -2567 -219 -2533
rect -253 -2635 -219 -2601
rect -253 -2703 -219 -2669
rect -253 -2771 -219 -2737
rect -253 -2839 -219 -2805
rect -253 -2907 -219 -2873
rect -253 -2975 -219 -2941
rect -253 -3043 -219 -3009
rect -253 -3111 -219 -3077
rect -253 -3179 -219 -3145
rect -253 -3247 -219 -3213
rect -253 -3315 -219 -3281
rect -253 -3383 -219 -3349
rect -253 -3451 -219 -3417
rect -253 -3519 -219 -3485
rect -253 -3587 -219 -3553
rect -253 -3655 -219 -3621
rect -253 -3723 -219 -3689
rect -253 -3791 -219 -3757
rect -253 -3859 -219 -3825
rect -253 -3927 -219 -3893
rect -253 -3995 -219 -3961
rect -253 -4063 -219 -4029
rect -253 -4131 -219 -4097
rect -253 -4199 -219 -4165
rect -253 -4267 -219 -4233
rect -253 -4335 -219 -4301
rect -253 -4403 -219 -4369
rect -253 -4471 -219 -4437
rect -253 -4539 -219 -4505
rect -253 -4607 -219 -4573
rect -253 -4675 -219 -4641
rect -253 -4743 -219 -4709
rect -253 -4811 -219 -4777
rect -253 -4879 -219 -4845
rect -253 -4947 -219 -4913
rect -253 -5015 -219 -4981
rect -253 -5083 -219 -5049
rect -253 -5151 -219 -5117
rect -253 -5219 -219 -5185
rect -253 -5287 -219 -5253
rect -253 -5355 -219 -5321
rect -253 -5423 -219 -5389
rect -253 -5491 -219 -5457
rect -253 -5559 -219 -5525
rect -253 -5627 -219 -5593
rect -253 -5695 -219 -5661
rect -253 -5763 -219 -5729
rect -253 -5831 -219 -5797
rect -253 -5899 -219 -5865
rect -253 -5967 -219 -5933
rect -135 5933 -101 5967
rect -135 5865 -101 5899
rect -135 5797 -101 5831
rect -135 5729 -101 5763
rect -135 5661 -101 5695
rect -135 5593 -101 5627
rect -135 5525 -101 5559
rect -135 5457 -101 5491
rect -135 5389 -101 5423
rect -135 5321 -101 5355
rect -135 5253 -101 5287
rect -135 5185 -101 5219
rect -135 5117 -101 5151
rect -135 5049 -101 5083
rect -135 4981 -101 5015
rect -135 4913 -101 4947
rect -135 4845 -101 4879
rect -135 4777 -101 4811
rect -135 4709 -101 4743
rect -135 4641 -101 4675
rect -135 4573 -101 4607
rect -135 4505 -101 4539
rect -135 4437 -101 4471
rect -135 4369 -101 4403
rect -135 4301 -101 4335
rect -135 4233 -101 4267
rect -135 4165 -101 4199
rect -135 4097 -101 4131
rect -135 4029 -101 4063
rect -135 3961 -101 3995
rect -135 3893 -101 3927
rect -135 3825 -101 3859
rect -135 3757 -101 3791
rect -135 3689 -101 3723
rect -135 3621 -101 3655
rect -135 3553 -101 3587
rect -135 3485 -101 3519
rect -135 3417 -101 3451
rect -135 3349 -101 3383
rect -135 3281 -101 3315
rect -135 3213 -101 3247
rect -135 3145 -101 3179
rect -135 3077 -101 3111
rect -135 3009 -101 3043
rect -135 2941 -101 2975
rect -135 2873 -101 2907
rect -135 2805 -101 2839
rect -135 2737 -101 2771
rect -135 2669 -101 2703
rect -135 2601 -101 2635
rect -135 2533 -101 2567
rect -135 2465 -101 2499
rect -135 2397 -101 2431
rect -135 2329 -101 2363
rect -135 2261 -101 2295
rect -135 2193 -101 2227
rect -135 2125 -101 2159
rect -135 2057 -101 2091
rect -135 1989 -101 2023
rect -135 1921 -101 1955
rect -135 1853 -101 1887
rect -135 1785 -101 1819
rect -135 1717 -101 1751
rect -135 1649 -101 1683
rect -135 1581 -101 1615
rect -135 1513 -101 1547
rect -135 1445 -101 1479
rect -135 1377 -101 1411
rect -135 1309 -101 1343
rect -135 1241 -101 1275
rect -135 1173 -101 1207
rect -135 1105 -101 1139
rect -135 1037 -101 1071
rect -135 969 -101 1003
rect -135 901 -101 935
rect -135 833 -101 867
rect -135 765 -101 799
rect -135 697 -101 731
rect -135 629 -101 663
rect -135 561 -101 595
rect -135 493 -101 527
rect -135 425 -101 459
rect -135 357 -101 391
rect -135 289 -101 323
rect -135 221 -101 255
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -135 -255 -101 -221
rect -135 -323 -101 -289
rect -135 -391 -101 -357
rect -135 -459 -101 -425
rect -135 -527 -101 -493
rect -135 -595 -101 -561
rect -135 -663 -101 -629
rect -135 -731 -101 -697
rect -135 -799 -101 -765
rect -135 -867 -101 -833
rect -135 -935 -101 -901
rect -135 -1003 -101 -969
rect -135 -1071 -101 -1037
rect -135 -1139 -101 -1105
rect -135 -1207 -101 -1173
rect -135 -1275 -101 -1241
rect -135 -1343 -101 -1309
rect -135 -1411 -101 -1377
rect -135 -1479 -101 -1445
rect -135 -1547 -101 -1513
rect -135 -1615 -101 -1581
rect -135 -1683 -101 -1649
rect -135 -1751 -101 -1717
rect -135 -1819 -101 -1785
rect -135 -1887 -101 -1853
rect -135 -1955 -101 -1921
rect -135 -2023 -101 -1989
rect -135 -2091 -101 -2057
rect -135 -2159 -101 -2125
rect -135 -2227 -101 -2193
rect -135 -2295 -101 -2261
rect -135 -2363 -101 -2329
rect -135 -2431 -101 -2397
rect -135 -2499 -101 -2465
rect -135 -2567 -101 -2533
rect -135 -2635 -101 -2601
rect -135 -2703 -101 -2669
rect -135 -2771 -101 -2737
rect -135 -2839 -101 -2805
rect -135 -2907 -101 -2873
rect -135 -2975 -101 -2941
rect -135 -3043 -101 -3009
rect -135 -3111 -101 -3077
rect -135 -3179 -101 -3145
rect -135 -3247 -101 -3213
rect -135 -3315 -101 -3281
rect -135 -3383 -101 -3349
rect -135 -3451 -101 -3417
rect -135 -3519 -101 -3485
rect -135 -3587 -101 -3553
rect -135 -3655 -101 -3621
rect -135 -3723 -101 -3689
rect -135 -3791 -101 -3757
rect -135 -3859 -101 -3825
rect -135 -3927 -101 -3893
rect -135 -3995 -101 -3961
rect -135 -4063 -101 -4029
rect -135 -4131 -101 -4097
rect -135 -4199 -101 -4165
rect -135 -4267 -101 -4233
rect -135 -4335 -101 -4301
rect -135 -4403 -101 -4369
rect -135 -4471 -101 -4437
rect -135 -4539 -101 -4505
rect -135 -4607 -101 -4573
rect -135 -4675 -101 -4641
rect -135 -4743 -101 -4709
rect -135 -4811 -101 -4777
rect -135 -4879 -101 -4845
rect -135 -4947 -101 -4913
rect -135 -5015 -101 -4981
rect -135 -5083 -101 -5049
rect -135 -5151 -101 -5117
rect -135 -5219 -101 -5185
rect -135 -5287 -101 -5253
rect -135 -5355 -101 -5321
rect -135 -5423 -101 -5389
rect -135 -5491 -101 -5457
rect -135 -5559 -101 -5525
rect -135 -5627 -101 -5593
rect -135 -5695 -101 -5661
rect -135 -5763 -101 -5729
rect -135 -5831 -101 -5797
rect -135 -5899 -101 -5865
rect -135 -5967 -101 -5933
rect -17 5933 17 5967
rect -17 5865 17 5899
rect -17 5797 17 5831
rect -17 5729 17 5763
rect -17 5661 17 5695
rect -17 5593 17 5627
rect -17 5525 17 5559
rect -17 5457 17 5491
rect -17 5389 17 5423
rect -17 5321 17 5355
rect -17 5253 17 5287
rect -17 5185 17 5219
rect -17 5117 17 5151
rect -17 5049 17 5083
rect -17 4981 17 5015
rect -17 4913 17 4947
rect -17 4845 17 4879
rect -17 4777 17 4811
rect -17 4709 17 4743
rect -17 4641 17 4675
rect -17 4573 17 4607
rect -17 4505 17 4539
rect -17 4437 17 4471
rect -17 4369 17 4403
rect -17 4301 17 4335
rect -17 4233 17 4267
rect -17 4165 17 4199
rect -17 4097 17 4131
rect -17 4029 17 4063
rect -17 3961 17 3995
rect -17 3893 17 3927
rect -17 3825 17 3859
rect -17 3757 17 3791
rect -17 3689 17 3723
rect -17 3621 17 3655
rect -17 3553 17 3587
rect -17 3485 17 3519
rect -17 3417 17 3451
rect -17 3349 17 3383
rect -17 3281 17 3315
rect -17 3213 17 3247
rect -17 3145 17 3179
rect -17 3077 17 3111
rect -17 3009 17 3043
rect -17 2941 17 2975
rect -17 2873 17 2907
rect -17 2805 17 2839
rect -17 2737 17 2771
rect -17 2669 17 2703
rect -17 2601 17 2635
rect -17 2533 17 2567
rect -17 2465 17 2499
rect -17 2397 17 2431
rect -17 2329 17 2363
rect -17 2261 17 2295
rect -17 2193 17 2227
rect -17 2125 17 2159
rect -17 2057 17 2091
rect -17 1989 17 2023
rect -17 1921 17 1955
rect -17 1853 17 1887
rect -17 1785 17 1819
rect -17 1717 17 1751
rect -17 1649 17 1683
rect -17 1581 17 1615
rect -17 1513 17 1547
rect -17 1445 17 1479
rect -17 1377 17 1411
rect -17 1309 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1139
rect -17 1037 17 1071
rect -17 969 17 1003
rect -17 901 17 935
rect -17 833 17 867
rect -17 765 17 799
rect -17 697 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -697
rect -17 -799 17 -765
rect -17 -867 17 -833
rect -17 -935 17 -901
rect -17 -1003 17 -969
rect -17 -1071 17 -1037
rect -17 -1139 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1309
rect -17 -1411 17 -1377
rect -17 -1479 17 -1445
rect -17 -1547 17 -1513
rect -17 -1615 17 -1581
rect -17 -1683 17 -1649
rect -17 -1751 17 -1717
rect -17 -1819 17 -1785
rect -17 -1887 17 -1853
rect -17 -1955 17 -1921
rect -17 -2023 17 -1989
rect -17 -2091 17 -2057
rect -17 -2159 17 -2125
rect -17 -2227 17 -2193
rect -17 -2295 17 -2261
rect -17 -2363 17 -2329
rect -17 -2431 17 -2397
rect -17 -2499 17 -2465
rect -17 -2567 17 -2533
rect -17 -2635 17 -2601
rect -17 -2703 17 -2669
rect -17 -2771 17 -2737
rect -17 -2839 17 -2805
rect -17 -2907 17 -2873
rect -17 -2975 17 -2941
rect -17 -3043 17 -3009
rect -17 -3111 17 -3077
rect -17 -3179 17 -3145
rect -17 -3247 17 -3213
rect -17 -3315 17 -3281
rect -17 -3383 17 -3349
rect -17 -3451 17 -3417
rect -17 -3519 17 -3485
rect -17 -3587 17 -3553
rect -17 -3655 17 -3621
rect -17 -3723 17 -3689
rect -17 -3791 17 -3757
rect -17 -3859 17 -3825
rect -17 -3927 17 -3893
rect -17 -3995 17 -3961
rect -17 -4063 17 -4029
rect -17 -4131 17 -4097
rect -17 -4199 17 -4165
rect -17 -4267 17 -4233
rect -17 -4335 17 -4301
rect -17 -4403 17 -4369
rect -17 -4471 17 -4437
rect -17 -4539 17 -4505
rect -17 -4607 17 -4573
rect -17 -4675 17 -4641
rect -17 -4743 17 -4709
rect -17 -4811 17 -4777
rect -17 -4879 17 -4845
rect -17 -4947 17 -4913
rect -17 -5015 17 -4981
rect -17 -5083 17 -5049
rect -17 -5151 17 -5117
rect -17 -5219 17 -5185
rect -17 -5287 17 -5253
rect -17 -5355 17 -5321
rect -17 -5423 17 -5389
rect -17 -5491 17 -5457
rect -17 -5559 17 -5525
rect -17 -5627 17 -5593
rect -17 -5695 17 -5661
rect -17 -5763 17 -5729
rect -17 -5831 17 -5797
rect -17 -5899 17 -5865
rect -17 -5967 17 -5933
rect 101 5933 135 5967
rect 101 5865 135 5899
rect 101 5797 135 5831
rect 101 5729 135 5763
rect 101 5661 135 5695
rect 101 5593 135 5627
rect 101 5525 135 5559
rect 101 5457 135 5491
rect 101 5389 135 5423
rect 101 5321 135 5355
rect 101 5253 135 5287
rect 101 5185 135 5219
rect 101 5117 135 5151
rect 101 5049 135 5083
rect 101 4981 135 5015
rect 101 4913 135 4947
rect 101 4845 135 4879
rect 101 4777 135 4811
rect 101 4709 135 4743
rect 101 4641 135 4675
rect 101 4573 135 4607
rect 101 4505 135 4539
rect 101 4437 135 4471
rect 101 4369 135 4403
rect 101 4301 135 4335
rect 101 4233 135 4267
rect 101 4165 135 4199
rect 101 4097 135 4131
rect 101 4029 135 4063
rect 101 3961 135 3995
rect 101 3893 135 3927
rect 101 3825 135 3859
rect 101 3757 135 3791
rect 101 3689 135 3723
rect 101 3621 135 3655
rect 101 3553 135 3587
rect 101 3485 135 3519
rect 101 3417 135 3451
rect 101 3349 135 3383
rect 101 3281 135 3315
rect 101 3213 135 3247
rect 101 3145 135 3179
rect 101 3077 135 3111
rect 101 3009 135 3043
rect 101 2941 135 2975
rect 101 2873 135 2907
rect 101 2805 135 2839
rect 101 2737 135 2771
rect 101 2669 135 2703
rect 101 2601 135 2635
rect 101 2533 135 2567
rect 101 2465 135 2499
rect 101 2397 135 2431
rect 101 2329 135 2363
rect 101 2261 135 2295
rect 101 2193 135 2227
rect 101 2125 135 2159
rect 101 2057 135 2091
rect 101 1989 135 2023
rect 101 1921 135 1955
rect 101 1853 135 1887
rect 101 1785 135 1819
rect 101 1717 135 1751
rect 101 1649 135 1683
rect 101 1581 135 1615
rect 101 1513 135 1547
rect 101 1445 135 1479
rect 101 1377 135 1411
rect 101 1309 135 1343
rect 101 1241 135 1275
rect 101 1173 135 1207
rect 101 1105 135 1139
rect 101 1037 135 1071
rect 101 969 135 1003
rect 101 901 135 935
rect 101 833 135 867
rect 101 765 135 799
rect 101 697 135 731
rect 101 629 135 663
rect 101 561 135 595
rect 101 493 135 527
rect 101 425 135 459
rect 101 357 135 391
rect 101 289 135 323
rect 101 221 135 255
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 101 -255 135 -221
rect 101 -323 135 -289
rect 101 -391 135 -357
rect 101 -459 135 -425
rect 101 -527 135 -493
rect 101 -595 135 -561
rect 101 -663 135 -629
rect 101 -731 135 -697
rect 101 -799 135 -765
rect 101 -867 135 -833
rect 101 -935 135 -901
rect 101 -1003 135 -969
rect 101 -1071 135 -1037
rect 101 -1139 135 -1105
rect 101 -1207 135 -1173
rect 101 -1275 135 -1241
rect 101 -1343 135 -1309
rect 101 -1411 135 -1377
rect 101 -1479 135 -1445
rect 101 -1547 135 -1513
rect 101 -1615 135 -1581
rect 101 -1683 135 -1649
rect 101 -1751 135 -1717
rect 101 -1819 135 -1785
rect 101 -1887 135 -1853
rect 101 -1955 135 -1921
rect 101 -2023 135 -1989
rect 101 -2091 135 -2057
rect 101 -2159 135 -2125
rect 101 -2227 135 -2193
rect 101 -2295 135 -2261
rect 101 -2363 135 -2329
rect 101 -2431 135 -2397
rect 101 -2499 135 -2465
rect 101 -2567 135 -2533
rect 101 -2635 135 -2601
rect 101 -2703 135 -2669
rect 101 -2771 135 -2737
rect 101 -2839 135 -2805
rect 101 -2907 135 -2873
rect 101 -2975 135 -2941
rect 101 -3043 135 -3009
rect 101 -3111 135 -3077
rect 101 -3179 135 -3145
rect 101 -3247 135 -3213
rect 101 -3315 135 -3281
rect 101 -3383 135 -3349
rect 101 -3451 135 -3417
rect 101 -3519 135 -3485
rect 101 -3587 135 -3553
rect 101 -3655 135 -3621
rect 101 -3723 135 -3689
rect 101 -3791 135 -3757
rect 101 -3859 135 -3825
rect 101 -3927 135 -3893
rect 101 -3995 135 -3961
rect 101 -4063 135 -4029
rect 101 -4131 135 -4097
rect 101 -4199 135 -4165
rect 101 -4267 135 -4233
rect 101 -4335 135 -4301
rect 101 -4403 135 -4369
rect 101 -4471 135 -4437
rect 101 -4539 135 -4505
rect 101 -4607 135 -4573
rect 101 -4675 135 -4641
rect 101 -4743 135 -4709
rect 101 -4811 135 -4777
rect 101 -4879 135 -4845
rect 101 -4947 135 -4913
rect 101 -5015 135 -4981
rect 101 -5083 135 -5049
rect 101 -5151 135 -5117
rect 101 -5219 135 -5185
rect 101 -5287 135 -5253
rect 101 -5355 135 -5321
rect 101 -5423 135 -5389
rect 101 -5491 135 -5457
rect 101 -5559 135 -5525
rect 101 -5627 135 -5593
rect 101 -5695 135 -5661
rect 101 -5763 135 -5729
rect 101 -5831 135 -5797
rect 101 -5899 135 -5865
rect 101 -5967 135 -5933
rect 219 5933 253 5967
rect 219 5865 253 5899
rect 219 5797 253 5831
rect 219 5729 253 5763
rect 219 5661 253 5695
rect 219 5593 253 5627
rect 219 5525 253 5559
rect 219 5457 253 5491
rect 219 5389 253 5423
rect 219 5321 253 5355
rect 219 5253 253 5287
rect 219 5185 253 5219
rect 219 5117 253 5151
rect 219 5049 253 5083
rect 219 4981 253 5015
rect 219 4913 253 4947
rect 219 4845 253 4879
rect 219 4777 253 4811
rect 219 4709 253 4743
rect 219 4641 253 4675
rect 219 4573 253 4607
rect 219 4505 253 4539
rect 219 4437 253 4471
rect 219 4369 253 4403
rect 219 4301 253 4335
rect 219 4233 253 4267
rect 219 4165 253 4199
rect 219 4097 253 4131
rect 219 4029 253 4063
rect 219 3961 253 3995
rect 219 3893 253 3927
rect 219 3825 253 3859
rect 219 3757 253 3791
rect 219 3689 253 3723
rect 219 3621 253 3655
rect 219 3553 253 3587
rect 219 3485 253 3519
rect 219 3417 253 3451
rect 219 3349 253 3383
rect 219 3281 253 3315
rect 219 3213 253 3247
rect 219 3145 253 3179
rect 219 3077 253 3111
rect 219 3009 253 3043
rect 219 2941 253 2975
rect 219 2873 253 2907
rect 219 2805 253 2839
rect 219 2737 253 2771
rect 219 2669 253 2703
rect 219 2601 253 2635
rect 219 2533 253 2567
rect 219 2465 253 2499
rect 219 2397 253 2431
rect 219 2329 253 2363
rect 219 2261 253 2295
rect 219 2193 253 2227
rect 219 2125 253 2159
rect 219 2057 253 2091
rect 219 1989 253 2023
rect 219 1921 253 1955
rect 219 1853 253 1887
rect 219 1785 253 1819
rect 219 1717 253 1751
rect 219 1649 253 1683
rect 219 1581 253 1615
rect 219 1513 253 1547
rect 219 1445 253 1479
rect 219 1377 253 1411
rect 219 1309 253 1343
rect 219 1241 253 1275
rect 219 1173 253 1207
rect 219 1105 253 1139
rect 219 1037 253 1071
rect 219 969 253 1003
rect 219 901 253 935
rect 219 833 253 867
rect 219 765 253 799
rect 219 697 253 731
rect 219 629 253 663
rect 219 561 253 595
rect 219 493 253 527
rect 219 425 253 459
rect 219 357 253 391
rect 219 289 253 323
rect 219 221 253 255
rect 219 153 253 187
rect 219 85 253 119
rect 219 17 253 51
rect 219 -51 253 -17
rect 219 -119 253 -85
rect 219 -187 253 -153
rect 219 -255 253 -221
rect 219 -323 253 -289
rect 219 -391 253 -357
rect 219 -459 253 -425
rect 219 -527 253 -493
rect 219 -595 253 -561
rect 219 -663 253 -629
rect 219 -731 253 -697
rect 219 -799 253 -765
rect 219 -867 253 -833
rect 219 -935 253 -901
rect 219 -1003 253 -969
rect 219 -1071 253 -1037
rect 219 -1139 253 -1105
rect 219 -1207 253 -1173
rect 219 -1275 253 -1241
rect 219 -1343 253 -1309
rect 219 -1411 253 -1377
rect 219 -1479 253 -1445
rect 219 -1547 253 -1513
rect 219 -1615 253 -1581
rect 219 -1683 253 -1649
rect 219 -1751 253 -1717
rect 219 -1819 253 -1785
rect 219 -1887 253 -1853
rect 219 -1955 253 -1921
rect 219 -2023 253 -1989
rect 219 -2091 253 -2057
rect 219 -2159 253 -2125
rect 219 -2227 253 -2193
rect 219 -2295 253 -2261
rect 219 -2363 253 -2329
rect 219 -2431 253 -2397
rect 219 -2499 253 -2465
rect 219 -2567 253 -2533
rect 219 -2635 253 -2601
rect 219 -2703 253 -2669
rect 219 -2771 253 -2737
rect 219 -2839 253 -2805
rect 219 -2907 253 -2873
rect 219 -2975 253 -2941
rect 219 -3043 253 -3009
rect 219 -3111 253 -3077
rect 219 -3179 253 -3145
rect 219 -3247 253 -3213
rect 219 -3315 253 -3281
rect 219 -3383 253 -3349
rect 219 -3451 253 -3417
rect 219 -3519 253 -3485
rect 219 -3587 253 -3553
rect 219 -3655 253 -3621
rect 219 -3723 253 -3689
rect 219 -3791 253 -3757
rect 219 -3859 253 -3825
rect 219 -3927 253 -3893
rect 219 -3995 253 -3961
rect 219 -4063 253 -4029
rect 219 -4131 253 -4097
rect 219 -4199 253 -4165
rect 219 -4267 253 -4233
rect 219 -4335 253 -4301
rect 219 -4403 253 -4369
rect 219 -4471 253 -4437
rect 219 -4539 253 -4505
rect 219 -4607 253 -4573
rect 219 -4675 253 -4641
rect 219 -4743 253 -4709
rect 219 -4811 253 -4777
rect 219 -4879 253 -4845
rect 219 -4947 253 -4913
rect 219 -5015 253 -4981
rect 219 -5083 253 -5049
rect 219 -5151 253 -5117
rect 219 -5219 253 -5185
rect 219 -5287 253 -5253
rect 219 -5355 253 -5321
rect 219 -5423 253 -5389
rect 219 -5491 253 -5457
rect 219 -5559 253 -5525
rect 219 -5627 253 -5593
rect 219 -5695 253 -5661
rect 219 -5763 253 -5729
rect 219 -5831 253 -5797
rect 219 -5899 253 -5865
rect 219 -5967 253 -5933
rect 337 5933 371 5967
rect 337 5865 371 5899
rect 337 5797 371 5831
rect 337 5729 371 5763
rect 337 5661 371 5695
rect 337 5593 371 5627
rect 337 5525 371 5559
rect 337 5457 371 5491
rect 337 5389 371 5423
rect 337 5321 371 5355
rect 337 5253 371 5287
rect 337 5185 371 5219
rect 337 5117 371 5151
rect 337 5049 371 5083
rect 337 4981 371 5015
rect 337 4913 371 4947
rect 337 4845 371 4879
rect 337 4777 371 4811
rect 337 4709 371 4743
rect 337 4641 371 4675
rect 337 4573 371 4607
rect 337 4505 371 4539
rect 337 4437 371 4471
rect 337 4369 371 4403
rect 337 4301 371 4335
rect 337 4233 371 4267
rect 337 4165 371 4199
rect 337 4097 371 4131
rect 337 4029 371 4063
rect 337 3961 371 3995
rect 337 3893 371 3927
rect 337 3825 371 3859
rect 337 3757 371 3791
rect 337 3689 371 3723
rect 337 3621 371 3655
rect 337 3553 371 3587
rect 337 3485 371 3519
rect 337 3417 371 3451
rect 337 3349 371 3383
rect 337 3281 371 3315
rect 337 3213 371 3247
rect 337 3145 371 3179
rect 337 3077 371 3111
rect 337 3009 371 3043
rect 337 2941 371 2975
rect 337 2873 371 2907
rect 337 2805 371 2839
rect 337 2737 371 2771
rect 337 2669 371 2703
rect 337 2601 371 2635
rect 337 2533 371 2567
rect 337 2465 371 2499
rect 337 2397 371 2431
rect 337 2329 371 2363
rect 337 2261 371 2295
rect 337 2193 371 2227
rect 337 2125 371 2159
rect 337 2057 371 2091
rect 337 1989 371 2023
rect 337 1921 371 1955
rect 337 1853 371 1887
rect 337 1785 371 1819
rect 337 1717 371 1751
rect 337 1649 371 1683
rect 337 1581 371 1615
rect 337 1513 371 1547
rect 337 1445 371 1479
rect 337 1377 371 1411
rect 337 1309 371 1343
rect 337 1241 371 1275
rect 337 1173 371 1207
rect 337 1105 371 1139
rect 337 1037 371 1071
rect 337 969 371 1003
rect 337 901 371 935
rect 337 833 371 867
rect 337 765 371 799
rect 337 697 371 731
rect 337 629 371 663
rect 337 561 371 595
rect 337 493 371 527
rect 337 425 371 459
rect 337 357 371 391
rect 337 289 371 323
rect 337 221 371 255
rect 337 153 371 187
rect 337 85 371 119
rect 337 17 371 51
rect 337 -51 371 -17
rect 337 -119 371 -85
rect 337 -187 371 -153
rect 337 -255 371 -221
rect 337 -323 371 -289
rect 337 -391 371 -357
rect 337 -459 371 -425
rect 337 -527 371 -493
rect 337 -595 371 -561
rect 337 -663 371 -629
rect 337 -731 371 -697
rect 337 -799 371 -765
rect 337 -867 371 -833
rect 337 -935 371 -901
rect 337 -1003 371 -969
rect 337 -1071 371 -1037
rect 337 -1139 371 -1105
rect 337 -1207 371 -1173
rect 337 -1275 371 -1241
rect 337 -1343 371 -1309
rect 337 -1411 371 -1377
rect 337 -1479 371 -1445
rect 337 -1547 371 -1513
rect 337 -1615 371 -1581
rect 337 -1683 371 -1649
rect 337 -1751 371 -1717
rect 337 -1819 371 -1785
rect 337 -1887 371 -1853
rect 337 -1955 371 -1921
rect 337 -2023 371 -1989
rect 337 -2091 371 -2057
rect 337 -2159 371 -2125
rect 337 -2227 371 -2193
rect 337 -2295 371 -2261
rect 337 -2363 371 -2329
rect 337 -2431 371 -2397
rect 337 -2499 371 -2465
rect 337 -2567 371 -2533
rect 337 -2635 371 -2601
rect 337 -2703 371 -2669
rect 337 -2771 371 -2737
rect 337 -2839 371 -2805
rect 337 -2907 371 -2873
rect 337 -2975 371 -2941
rect 337 -3043 371 -3009
rect 337 -3111 371 -3077
rect 337 -3179 371 -3145
rect 337 -3247 371 -3213
rect 337 -3315 371 -3281
rect 337 -3383 371 -3349
rect 337 -3451 371 -3417
rect 337 -3519 371 -3485
rect 337 -3587 371 -3553
rect 337 -3655 371 -3621
rect 337 -3723 371 -3689
rect 337 -3791 371 -3757
rect 337 -3859 371 -3825
rect 337 -3927 371 -3893
rect 337 -3995 371 -3961
rect 337 -4063 371 -4029
rect 337 -4131 371 -4097
rect 337 -4199 371 -4165
rect 337 -4267 371 -4233
rect 337 -4335 371 -4301
rect 337 -4403 371 -4369
rect 337 -4471 371 -4437
rect 337 -4539 371 -4505
rect 337 -4607 371 -4573
rect 337 -4675 371 -4641
rect 337 -4743 371 -4709
rect 337 -4811 371 -4777
rect 337 -4879 371 -4845
rect 337 -4947 371 -4913
rect 337 -5015 371 -4981
rect 337 -5083 371 -5049
rect 337 -5151 371 -5117
rect 337 -5219 371 -5185
rect 337 -5287 371 -5253
rect 337 -5355 371 -5321
rect 337 -5423 371 -5389
rect 337 -5491 371 -5457
rect 337 -5559 371 -5525
rect 337 -5627 371 -5593
rect 337 -5695 371 -5661
rect 337 -5763 371 -5729
rect 337 -5831 371 -5797
rect 337 -5899 371 -5865
rect 337 -5967 371 -5933
rect 455 5933 489 5967
rect 455 5865 489 5899
rect 455 5797 489 5831
rect 455 5729 489 5763
rect 455 5661 489 5695
rect 455 5593 489 5627
rect 455 5525 489 5559
rect 455 5457 489 5491
rect 455 5389 489 5423
rect 455 5321 489 5355
rect 455 5253 489 5287
rect 455 5185 489 5219
rect 455 5117 489 5151
rect 455 5049 489 5083
rect 455 4981 489 5015
rect 455 4913 489 4947
rect 455 4845 489 4879
rect 455 4777 489 4811
rect 455 4709 489 4743
rect 455 4641 489 4675
rect 455 4573 489 4607
rect 455 4505 489 4539
rect 455 4437 489 4471
rect 455 4369 489 4403
rect 455 4301 489 4335
rect 455 4233 489 4267
rect 455 4165 489 4199
rect 455 4097 489 4131
rect 455 4029 489 4063
rect 455 3961 489 3995
rect 455 3893 489 3927
rect 455 3825 489 3859
rect 455 3757 489 3791
rect 455 3689 489 3723
rect 455 3621 489 3655
rect 455 3553 489 3587
rect 455 3485 489 3519
rect 455 3417 489 3451
rect 455 3349 489 3383
rect 455 3281 489 3315
rect 455 3213 489 3247
rect 455 3145 489 3179
rect 455 3077 489 3111
rect 455 3009 489 3043
rect 455 2941 489 2975
rect 455 2873 489 2907
rect 455 2805 489 2839
rect 455 2737 489 2771
rect 455 2669 489 2703
rect 455 2601 489 2635
rect 455 2533 489 2567
rect 455 2465 489 2499
rect 455 2397 489 2431
rect 455 2329 489 2363
rect 455 2261 489 2295
rect 455 2193 489 2227
rect 455 2125 489 2159
rect 455 2057 489 2091
rect 455 1989 489 2023
rect 455 1921 489 1955
rect 455 1853 489 1887
rect 455 1785 489 1819
rect 455 1717 489 1751
rect 455 1649 489 1683
rect 455 1581 489 1615
rect 455 1513 489 1547
rect 455 1445 489 1479
rect 455 1377 489 1411
rect 455 1309 489 1343
rect 455 1241 489 1275
rect 455 1173 489 1207
rect 455 1105 489 1139
rect 455 1037 489 1071
rect 455 969 489 1003
rect 455 901 489 935
rect 455 833 489 867
rect 455 765 489 799
rect 455 697 489 731
rect 455 629 489 663
rect 455 561 489 595
rect 455 493 489 527
rect 455 425 489 459
rect 455 357 489 391
rect 455 289 489 323
rect 455 221 489 255
rect 455 153 489 187
rect 455 85 489 119
rect 455 17 489 51
rect 455 -51 489 -17
rect 455 -119 489 -85
rect 455 -187 489 -153
rect 455 -255 489 -221
rect 455 -323 489 -289
rect 455 -391 489 -357
rect 455 -459 489 -425
rect 455 -527 489 -493
rect 455 -595 489 -561
rect 455 -663 489 -629
rect 455 -731 489 -697
rect 455 -799 489 -765
rect 455 -867 489 -833
rect 455 -935 489 -901
rect 455 -1003 489 -969
rect 455 -1071 489 -1037
rect 455 -1139 489 -1105
rect 455 -1207 489 -1173
rect 455 -1275 489 -1241
rect 455 -1343 489 -1309
rect 455 -1411 489 -1377
rect 455 -1479 489 -1445
rect 455 -1547 489 -1513
rect 455 -1615 489 -1581
rect 455 -1683 489 -1649
rect 455 -1751 489 -1717
rect 455 -1819 489 -1785
rect 455 -1887 489 -1853
rect 455 -1955 489 -1921
rect 455 -2023 489 -1989
rect 455 -2091 489 -2057
rect 455 -2159 489 -2125
rect 455 -2227 489 -2193
rect 455 -2295 489 -2261
rect 455 -2363 489 -2329
rect 455 -2431 489 -2397
rect 455 -2499 489 -2465
rect 455 -2567 489 -2533
rect 455 -2635 489 -2601
rect 455 -2703 489 -2669
rect 455 -2771 489 -2737
rect 455 -2839 489 -2805
rect 455 -2907 489 -2873
rect 455 -2975 489 -2941
rect 455 -3043 489 -3009
rect 455 -3111 489 -3077
rect 455 -3179 489 -3145
rect 455 -3247 489 -3213
rect 455 -3315 489 -3281
rect 455 -3383 489 -3349
rect 455 -3451 489 -3417
rect 455 -3519 489 -3485
rect 455 -3587 489 -3553
rect 455 -3655 489 -3621
rect 455 -3723 489 -3689
rect 455 -3791 489 -3757
rect 455 -3859 489 -3825
rect 455 -3927 489 -3893
rect 455 -3995 489 -3961
rect 455 -4063 489 -4029
rect 455 -4131 489 -4097
rect 455 -4199 489 -4165
rect 455 -4267 489 -4233
rect 455 -4335 489 -4301
rect 455 -4403 489 -4369
rect 455 -4471 489 -4437
rect 455 -4539 489 -4505
rect 455 -4607 489 -4573
rect 455 -4675 489 -4641
rect 455 -4743 489 -4709
rect 455 -4811 489 -4777
rect 455 -4879 489 -4845
rect 455 -4947 489 -4913
rect 455 -5015 489 -4981
rect 455 -5083 489 -5049
rect 455 -5151 489 -5117
rect 455 -5219 489 -5185
rect 455 -5287 489 -5253
rect 455 -5355 489 -5321
rect 455 -5423 489 -5389
rect 455 -5491 489 -5457
rect 455 -5559 489 -5525
rect 455 -5627 489 -5593
rect 455 -5695 489 -5661
rect 455 -5763 489 -5729
rect 455 -5831 489 -5797
rect 455 -5899 489 -5865
rect 455 -5967 489 -5933
rect 573 5933 607 5967
rect 573 5865 607 5899
rect 573 5797 607 5831
rect 573 5729 607 5763
rect 573 5661 607 5695
rect 573 5593 607 5627
rect 573 5525 607 5559
rect 573 5457 607 5491
rect 573 5389 607 5423
rect 573 5321 607 5355
rect 573 5253 607 5287
rect 573 5185 607 5219
rect 573 5117 607 5151
rect 573 5049 607 5083
rect 573 4981 607 5015
rect 573 4913 607 4947
rect 573 4845 607 4879
rect 573 4777 607 4811
rect 573 4709 607 4743
rect 573 4641 607 4675
rect 573 4573 607 4607
rect 573 4505 607 4539
rect 573 4437 607 4471
rect 573 4369 607 4403
rect 573 4301 607 4335
rect 573 4233 607 4267
rect 573 4165 607 4199
rect 573 4097 607 4131
rect 573 4029 607 4063
rect 573 3961 607 3995
rect 573 3893 607 3927
rect 573 3825 607 3859
rect 573 3757 607 3791
rect 573 3689 607 3723
rect 573 3621 607 3655
rect 573 3553 607 3587
rect 573 3485 607 3519
rect 573 3417 607 3451
rect 573 3349 607 3383
rect 573 3281 607 3315
rect 573 3213 607 3247
rect 573 3145 607 3179
rect 573 3077 607 3111
rect 573 3009 607 3043
rect 573 2941 607 2975
rect 573 2873 607 2907
rect 573 2805 607 2839
rect 573 2737 607 2771
rect 573 2669 607 2703
rect 573 2601 607 2635
rect 573 2533 607 2567
rect 573 2465 607 2499
rect 573 2397 607 2431
rect 573 2329 607 2363
rect 573 2261 607 2295
rect 573 2193 607 2227
rect 573 2125 607 2159
rect 573 2057 607 2091
rect 573 1989 607 2023
rect 573 1921 607 1955
rect 573 1853 607 1887
rect 573 1785 607 1819
rect 573 1717 607 1751
rect 573 1649 607 1683
rect 573 1581 607 1615
rect 573 1513 607 1547
rect 573 1445 607 1479
rect 573 1377 607 1411
rect 573 1309 607 1343
rect 573 1241 607 1275
rect 573 1173 607 1207
rect 573 1105 607 1139
rect 573 1037 607 1071
rect 573 969 607 1003
rect 573 901 607 935
rect 573 833 607 867
rect 573 765 607 799
rect 573 697 607 731
rect 573 629 607 663
rect 573 561 607 595
rect 573 493 607 527
rect 573 425 607 459
rect 573 357 607 391
rect 573 289 607 323
rect 573 221 607 255
rect 573 153 607 187
rect 573 85 607 119
rect 573 17 607 51
rect 573 -51 607 -17
rect 573 -119 607 -85
rect 573 -187 607 -153
rect 573 -255 607 -221
rect 573 -323 607 -289
rect 573 -391 607 -357
rect 573 -459 607 -425
rect 573 -527 607 -493
rect 573 -595 607 -561
rect 573 -663 607 -629
rect 573 -731 607 -697
rect 573 -799 607 -765
rect 573 -867 607 -833
rect 573 -935 607 -901
rect 573 -1003 607 -969
rect 573 -1071 607 -1037
rect 573 -1139 607 -1105
rect 573 -1207 607 -1173
rect 573 -1275 607 -1241
rect 573 -1343 607 -1309
rect 573 -1411 607 -1377
rect 573 -1479 607 -1445
rect 573 -1547 607 -1513
rect 573 -1615 607 -1581
rect 573 -1683 607 -1649
rect 573 -1751 607 -1717
rect 573 -1819 607 -1785
rect 573 -1887 607 -1853
rect 573 -1955 607 -1921
rect 573 -2023 607 -1989
rect 573 -2091 607 -2057
rect 573 -2159 607 -2125
rect 573 -2227 607 -2193
rect 573 -2295 607 -2261
rect 573 -2363 607 -2329
rect 573 -2431 607 -2397
rect 573 -2499 607 -2465
rect 573 -2567 607 -2533
rect 573 -2635 607 -2601
rect 573 -2703 607 -2669
rect 573 -2771 607 -2737
rect 573 -2839 607 -2805
rect 573 -2907 607 -2873
rect 573 -2975 607 -2941
rect 573 -3043 607 -3009
rect 573 -3111 607 -3077
rect 573 -3179 607 -3145
rect 573 -3247 607 -3213
rect 573 -3315 607 -3281
rect 573 -3383 607 -3349
rect 573 -3451 607 -3417
rect 573 -3519 607 -3485
rect 573 -3587 607 -3553
rect 573 -3655 607 -3621
rect 573 -3723 607 -3689
rect 573 -3791 607 -3757
rect 573 -3859 607 -3825
rect 573 -3927 607 -3893
rect 573 -3995 607 -3961
rect 573 -4063 607 -4029
rect 573 -4131 607 -4097
rect 573 -4199 607 -4165
rect 573 -4267 607 -4233
rect 573 -4335 607 -4301
rect 573 -4403 607 -4369
rect 573 -4471 607 -4437
rect 573 -4539 607 -4505
rect 573 -4607 607 -4573
rect 573 -4675 607 -4641
rect 573 -4743 607 -4709
rect 573 -4811 607 -4777
rect 573 -4879 607 -4845
rect 573 -4947 607 -4913
rect 573 -5015 607 -4981
rect 573 -5083 607 -5049
rect 573 -5151 607 -5117
rect 573 -5219 607 -5185
rect 573 -5287 607 -5253
rect 573 -5355 607 -5321
rect 573 -5423 607 -5389
rect 573 -5491 607 -5457
rect 573 -5559 607 -5525
rect 573 -5627 607 -5593
rect 573 -5695 607 -5661
rect 573 -5763 607 -5729
rect 573 -5831 607 -5797
rect 573 -5899 607 -5865
rect 573 -5967 607 -5933
<< poly >>
rect -564 6072 -498 6088
rect -564 6038 -548 6072
rect -514 6038 -498 6072
rect -564 6022 -498 6038
rect -446 6078 -380 6088
rect -328 6078 -262 6088
rect -446 6032 -262 6078
rect -446 6022 -380 6032
rect -328 6022 -262 6032
rect -210 6078 -144 6088
rect -92 6078 -26 6088
rect -210 6032 -26 6078
rect -210 6022 -144 6032
rect -92 6022 -26 6032
rect 26 6078 92 6088
rect 144 6078 210 6088
rect 26 6032 210 6078
rect 26 6022 92 6032
rect 144 6022 210 6032
rect 262 6078 328 6088
rect 380 6078 446 6088
rect 498 6083 564 6088
rect 262 6032 446 6078
rect 262 6022 328 6032
rect 380 6022 446 6032
rect 497 6029 566 6083
rect 498 6022 564 6029
rect -561 6000 -501 6022
rect -443 6000 -383 6022
rect -325 6000 -265 6022
rect -207 6000 -147 6022
rect -89 6000 -29 6022
rect 29 6000 89 6022
rect 147 6000 207 6022
rect 265 6000 325 6022
rect 383 6000 443 6022
rect 501 6000 561 6022
rect -561 -6022 -501 -6000
rect -443 -6022 -383 -6000
rect -325 -6022 -265 -6000
rect -207 -6022 -147 -6000
rect -89 -6022 -29 -6000
rect 29 -6022 89 -6000
rect 147 -6022 207 -6000
rect 265 -6022 325 -6000
rect 383 -6022 443 -6000
rect 501 -6022 561 -6000
rect -564 -6032 -498 -6022
rect -446 -6032 -380 -6022
rect -564 -6078 -380 -6032
rect -564 -6088 -498 -6078
rect -446 -6088 -380 -6078
rect -328 -6032 -262 -6022
rect -210 -6032 -144 -6022
rect -328 -6078 -144 -6032
rect -328 -6088 -262 -6078
rect -210 -6088 -144 -6078
rect -92 -6032 -26 -6022
rect 26 -6032 92 -6022
rect -92 -6078 92 -6032
rect -92 -6088 -26 -6078
rect 26 -6088 92 -6078
rect 144 -6032 210 -6022
rect 262 -6032 328 -6022
rect 144 -6078 328 -6032
rect 144 -6088 210 -6078
rect 262 -6088 328 -6078
rect 380 -6032 446 -6022
rect 498 -6032 564 -6022
rect 380 -6078 564 -6032
rect 380 -6088 446 -6078
rect 498 -6088 564 -6078
<< polycont >>
rect -548 6038 -514 6072
<< locali >>
rect -564 6038 -548 6072
rect -514 6038 -498 6072
rect -607 5967 -573 6004
rect -607 5899 -573 5923
rect -607 5831 -573 5851
rect -607 5763 -573 5779
rect -607 5695 -573 5707
rect -607 5627 -573 5635
rect -607 5559 -573 5563
rect -607 5453 -573 5457
rect -607 5381 -573 5389
rect -607 5309 -573 5321
rect -607 5237 -573 5253
rect -607 5165 -573 5185
rect -607 5093 -573 5117
rect -607 5021 -573 5049
rect -607 4949 -573 4981
rect -607 4879 -573 4913
rect -607 4811 -573 4843
rect -607 4743 -573 4771
rect -607 4675 -573 4699
rect -607 4607 -573 4627
rect -607 4539 -573 4555
rect -607 4471 -573 4483
rect -607 4403 -573 4411
rect -607 4335 -573 4339
rect -607 4229 -573 4233
rect -607 4157 -573 4165
rect -607 4085 -573 4097
rect -607 4013 -573 4029
rect -607 3941 -573 3961
rect -607 3869 -573 3893
rect -607 3797 -573 3825
rect -607 3725 -573 3757
rect -607 3655 -573 3689
rect -607 3587 -573 3619
rect -607 3519 -573 3547
rect -607 3451 -573 3475
rect -607 3383 -573 3403
rect -607 3315 -573 3331
rect -607 3247 -573 3259
rect -607 3179 -573 3187
rect -607 3111 -573 3115
rect -607 3005 -573 3009
rect -607 2933 -573 2941
rect -607 2861 -573 2873
rect -607 2789 -573 2805
rect -607 2717 -573 2737
rect -607 2645 -573 2669
rect -607 2573 -573 2601
rect -607 2501 -573 2533
rect -607 2431 -573 2465
rect -607 2363 -573 2395
rect -607 2295 -573 2323
rect -607 2227 -573 2251
rect -607 2159 -573 2179
rect -607 2091 -573 2107
rect -607 2023 -573 2035
rect -607 1955 -573 1963
rect -607 1887 -573 1891
rect -607 1781 -573 1785
rect -607 1709 -573 1717
rect -607 1637 -573 1649
rect -607 1565 -573 1581
rect -607 1493 -573 1513
rect -607 1421 -573 1445
rect -607 1349 -573 1377
rect -607 1277 -573 1309
rect -607 1207 -573 1241
rect -607 1139 -573 1171
rect -607 1071 -573 1099
rect -607 1003 -573 1027
rect -607 935 -573 955
rect -607 867 -573 883
rect -607 799 -573 811
rect -607 731 -573 739
rect -607 663 -573 667
rect -607 557 -573 561
rect -607 485 -573 493
rect -607 413 -573 425
rect -607 341 -573 357
rect -607 269 -573 289
rect -607 197 -573 221
rect -607 125 -573 153
rect -607 53 -573 85
rect -607 -17 -573 17
rect -607 -85 -573 -53
rect -607 -153 -573 -125
rect -607 -221 -573 -197
rect -607 -289 -573 -269
rect -607 -357 -573 -341
rect -607 -425 -573 -413
rect -607 -493 -573 -485
rect -607 -561 -573 -557
rect -607 -667 -573 -663
rect -607 -739 -573 -731
rect -607 -811 -573 -799
rect -607 -883 -573 -867
rect -607 -955 -573 -935
rect -607 -1027 -573 -1003
rect -607 -1099 -573 -1071
rect -607 -1171 -573 -1139
rect -607 -1241 -573 -1207
rect -607 -1309 -573 -1277
rect -607 -1377 -573 -1349
rect -607 -1445 -573 -1421
rect -607 -1513 -573 -1493
rect -607 -1581 -573 -1565
rect -607 -1649 -573 -1637
rect -607 -1717 -573 -1709
rect -607 -1785 -573 -1781
rect -607 -1891 -573 -1887
rect -607 -1963 -573 -1955
rect -607 -2035 -573 -2023
rect -607 -2107 -573 -2091
rect -607 -2179 -573 -2159
rect -607 -2251 -573 -2227
rect -607 -2323 -573 -2295
rect -607 -2395 -573 -2363
rect -607 -2465 -573 -2431
rect -607 -2533 -573 -2501
rect -607 -2601 -573 -2573
rect -607 -2669 -573 -2645
rect -607 -2737 -573 -2717
rect -607 -2805 -573 -2789
rect -607 -2873 -573 -2861
rect -607 -2941 -573 -2933
rect -607 -3009 -573 -3005
rect -607 -3115 -573 -3111
rect -607 -3187 -573 -3179
rect -607 -3259 -573 -3247
rect -607 -3331 -573 -3315
rect -607 -3403 -573 -3383
rect -607 -3475 -573 -3451
rect -607 -3547 -573 -3519
rect -607 -3619 -573 -3587
rect -607 -3689 -573 -3655
rect -607 -3757 -573 -3725
rect -607 -3825 -573 -3797
rect -607 -3893 -573 -3869
rect -607 -3961 -573 -3941
rect -607 -4029 -573 -4013
rect -607 -4097 -573 -4085
rect -607 -4165 -573 -4157
rect -607 -4233 -573 -4229
rect -607 -4339 -573 -4335
rect -607 -4411 -573 -4403
rect -607 -4483 -573 -4471
rect -607 -4555 -573 -4539
rect -607 -4627 -573 -4607
rect -607 -4699 -573 -4675
rect -607 -4771 -573 -4743
rect -607 -4843 -573 -4811
rect -607 -4913 -573 -4879
rect -607 -4981 -573 -4949
rect -607 -5049 -573 -5021
rect -607 -5117 -573 -5093
rect -607 -5185 -573 -5165
rect -607 -5253 -573 -5237
rect -607 -5321 -573 -5309
rect -607 -5389 -573 -5381
rect -607 -5457 -573 -5453
rect -607 -5563 -573 -5559
rect -607 -5635 -573 -5627
rect -607 -5707 -573 -5695
rect -607 -5779 -573 -5763
rect -607 -5851 -573 -5831
rect -607 -5923 -573 -5899
rect -607 -6004 -573 -5967
rect -489 5967 -455 6004
rect -489 5899 -455 5923
rect -489 5831 -455 5851
rect -489 5763 -455 5779
rect -489 5695 -455 5707
rect -489 5627 -455 5635
rect -489 5559 -455 5563
rect -489 5453 -455 5457
rect -489 5381 -455 5389
rect -489 5309 -455 5321
rect -489 5237 -455 5253
rect -489 5165 -455 5185
rect -489 5093 -455 5117
rect -489 5021 -455 5049
rect -489 4949 -455 4981
rect -489 4879 -455 4913
rect -489 4811 -455 4843
rect -489 4743 -455 4771
rect -489 4675 -455 4699
rect -489 4607 -455 4627
rect -489 4539 -455 4555
rect -489 4471 -455 4483
rect -489 4403 -455 4411
rect -489 4335 -455 4339
rect -489 4229 -455 4233
rect -489 4157 -455 4165
rect -489 4085 -455 4097
rect -489 4013 -455 4029
rect -489 3941 -455 3961
rect -489 3869 -455 3893
rect -489 3797 -455 3825
rect -489 3725 -455 3757
rect -489 3655 -455 3689
rect -489 3587 -455 3619
rect -489 3519 -455 3547
rect -489 3451 -455 3475
rect -489 3383 -455 3403
rect -489 3315 -455 3331
rect -489 3247 -455 3259
rect -489 3179 -455 3187
rect -489 3111 -455 3115
rect -489 3005 -455 3009
rect -489 2933 -455 2941
rect -489 2861 -455 2873
rect -489 2789 -455 2805
rect -489 2717 -455 2737
rect -489 2645 -455 2669
rect -489 2573 -455 2601
rect -489 2501 -455 2533
rect -489 2431 -455 2465
rect -489 2363 -455 2395
rect -489 2295 -455 2323
rect -489 2227 -455 2251
rect -489 2159 -455 2179
rect -489 2091 -455 2107
rect -489 2023 -455 2035
rect -489 1955 -455 1963
rect -489 1887 -455 1891
rect -489 1781 -455 1785
rect -489 1709 -455 1717
rect -489 1637 -455 1649
rect -489 1565 -455 1581
rect -489 1493 -455 1513
rect -489 1421 -455 1445
rect -489 1349 -455 1377
rect -489 1277 -455 1309
rect -489 1207 -455 1241
rect -489 1139 -455 1171
rect -489 1071 -455 1099
rect -489 1003 -455 1027
rect -489 935 -455 955
rect -489 867 -455 883
rect -489 799 -455 811
rect -489 731 -455 739
rect -489 663 -455 667
rect -489 557 -455 561
rect -489 485 -455 493
rect -489 413 -455 425
rect -489 341 -455 357
rect -489 269 -455 289
rect -489 197 -455 221
rect -489 125 -455 153
rect -489 53 -455 85
rect -489 -17 -455 17
rect -489 -85 -455 -53
rect -489 -153 -455 -125
rect -489 -221 -455 -197
rect -489 -289 -455 -269
rect -489 -357 -455 -341
rect -489 -425 -455 -413
rect -489 -493 -455 -485
rect -489 -561 -455 -557
rect -489 -667 -455 -663
rect -489 -739 -455 -731
rect -489 -811 -455 -799
rect -489 -883 -455 -867
rect -489 -955 -455 -935
rect -489 -1027 -455 -1003
rect -489 -1099 -455 -1071
rect -489 -1171 -455 -1139
rect -489 -1241 -455 -1207
rect -489 -1309 -455 -1277
rect -489 -1377 -455 -1349
rect -489 -1445 -455 -1421
rect -489 -1513 -455 -1493
rect -489 -1581 -455 -1565
rect -489 -1649 -455 -1637
rect -489 -1717 -455 -1709
rect -489 -1785 -455 -1781
rect -489 -1891 -455 -1887
rect -489 -1963 -455 -1955
rect -489 -2035 -455 -2023
rect -489 -2107 -455 -2091
rect -489 -2179 -455 -2159
rect -489 -2251 -455 -2227
rect -489 -2323 -455 -2295
rect -489 -2395 -455 -2363
rect -489 -2465 -455 -2431
rect -489 -2533 -455 -2501
rect -489 -2601 -455 -2573
rect -489 -2669 -455 -2645
rect -489 -2737 -455 -2717
rect -489 -2805 -455 -2789
rect -489 -2873 -455 -2861
rect -489 -2941 -455 -2933
rect -489 -3009 -455 -3005
rect -489 -3115 -455 -3111
rect -489 -3187 -455 -3179
rect -489 -3259 -455 -3247
rect -489 -3331 -455 -3315
rect -489 -3403 -455 -3383
rect -489 -3475 -455 -3451
rect -489 -3547 -455 -3519
rect -489 -3619 -455 -3587
rect -489 -3689 -455 -3655
rect -489 -3757 -455 -3725
rect -489 -3825 -455 -3797
rect -489 -3893 -455 -3869
rect -489 -3961 -455 -3941
rect -489 -4029 -455 -4013
rect -489 -4097 -455 -4085
rect -489 -4165 -455 -4157
rect -489 -4233 -455 -4229
rect -489 -4339 -455 -4335
rect -489 -4411 -455 -4403
rect -489 -4483 -455 -4471
rect -489 -4555 -455 -4539
rect -489 -4627 -455 -4607
rect -489 -4699 -455 -4675
rect -489 -4771 -455 -4743
rect -489 -4843 -455 -4811
rect -489 -4913 -455 -4879
rect -489 -4981 -455 -4949
rect -489 -5049 -455 -5021
rect -489 -5117 -455 -5093
rect -489 -5185 -455 -5165
rect -489 -5253 -455 -5237
rect -489 -5321 -455 -5309
rect -489 -5389 -455 -5381
rect -489 -5457 -455 -5453
rect -489 -5563 -455 -5559
rect -489 -5635 -455 -5627
rect -489 -5707 -455 -5695
rect -489 -5779 -455 -5763
rect -489 -5851 -455 -5831
rect -489 -5923 -455 -5899
rect -489 -6004 -455 -5967
rect -371 5967 -337 6004
rect -371 5899 -337 5923
rect -371 5831 -337 5851
rect -371 5763 -337 5779
rect -371 5695 -337 5707
rect -371 5627 -337 5635
rect -371 5559 -337 5563
rect -371 5453 -337 5457
rect -371 5381 -337 5389
rect -371 5309 -337 5321
rect -371 5237 -337 5253
rect -371 5165 -337 5185
rect -371 5093 -337 5117
rect -371 5021 -337 5049
rect -371 4949 -337 4981
rect -371 4879 -337 4913
rect -371 4811 -337 4843
rect -371 4743 -337 4771
rect -371 4675 -337 4699
rect -371 4607 -337 4627
rect -371 4539 -337 4555
rect -371 4471 -337 4483
rect -371 4403 -337 4411
rect -371 4335 -337 4339
rect -371 4229 -337 4233
rect -371 4157 -337 4165
rect -371 4085 -337 4097
rect -371 4013 -337 4029
rect -371 3941 -337 3961
rect -371 3869 -337 3893
rect -371 3797 -337 3825
rect -371 3725 -337 3757
rect -371 3655 -337 3689
rect -371 3587 -337 3619
rect -371 3519 -337 3547
rect -371 3451 -337 3475
rect -371 3383 -337 3403
rect -371 3315 -337 3331
rect -371 3247 -337 3259
rect -371 3179 -337 3187
rect -371 3111 -337 3115
rect -371 3005 -337 3009
rect -371 2933 -337 2941
rect -371 2861 -337 2873
rect -371 2789 -337 2805
rect -371 2717 -337 2737
rect -371 2645 -337 2669
rect -371 2573 -337 2601
rect -371 2501 -337 2533
rect -371 2431 -337 2465
rect -371 2363 -337 2395
rect -371 2295 -337 2323
rect -371 2227 -337 2251
rect -371 2159 -337 2179
rect -371 2091 -337 2107
rect -371 2023 -337 2035
rect -371 1955 -337 1963
rect -371 1887 -337 1891
rect -371 1781 -337 1785
rect -371 1709 -337 1717
rect -371 1637 -337 1649
rect -371 1565 -337 1581
rect -371 1493 -337 1513
rect -371 1421 -337 1445
rect -371 1349 -337 1377
rect -371 1277 -337 1309
rect -371 1207 -337 1241
rect -371 1139 -337 1171
rect -371 1071 -337 1099
rect -371 1003 -337 1027
rect -371 935 -337 955
rect -371 867 -337 883
rect -371 799 -337 811
rect -371 731 -337 739
rect -371 663 -337 667
rect -371 557 -337 561
rect -371 485 -337 493
rect -371 413 -337 425
rect -371 341 -337 357
rect -371 269 -337 289
rect -371 197 -337 221
rect -371 125 -337 153
rect -371 53 -337 85
rect -371 -17 -337 17
rect -371 -85 -337 -53
rect -371 -153 -337 -125
rect -371 -221 -337 -197
rect -371 -289 -337 -269
rect -371 -357 -337 -341
rect -371 -425 -337 -413
rect -371 -493 -337 -485
rect -371 -561 -337 -557
rect -371 -667 -337 -663
rect -371 -739 -337 -731
rect -371 -811 -337 -799
rect -371 -883 -337 -867
rect -371 -955 -337 -935
rect -371 -1027 -337 -1003
rect -371 -1099 -337 -1071
rect -371 -1171 -337 -1139
rect -371 -1241 -337 -1207
rect -371 -1309 -337 -1277
rect -371 -1377 -337 -1349
rect -371 -1445 -337 -1421
rect -371 -1513 -337 -1493
rect -371 -1581 -337 -1565
rect -371 -1649 -337 -1637
rect -371 -1717 -337 -1709
rect -371 -1785 -337 -1781
rect -371 -1891 -337 -1887
rect -371 -1963 -337 -1955
rect -371 -2035 -337 -2023
rect -371 -2107 -337 -2091
rect -371 -2179 -337 -2159
rect -371 -2251 -337 -2227
rect -371 -2323 -337 -2295
rect -371 -2395 -337 -2363
rect -371 -2465 -337 -2431
rect -371 -2533 -337 -2501
rect -371 -2601 -337 -2573
rect -371 -2669 -337 -2645
rect -371 -2737 -337 -2717
rect -371 -2805 -337 -2789
rect -371 -2873 -337 -2861
rect -371 -2941 -337 -2933
rect -371 -3009 -337 -3005
rect -371 -3115 -337 -3111
rect -371 -3187 -337 -3179
rect -371 -3259 -337 -3247
rect -371 -3331 -337 -3315
rect -371 -3403 -337 -3383
rect -371 -3475 -337 -3451
rect -371 -3547 -337 -3519
rect -371 -3619 -337 -3587
rect -371 -3689 -337 -3655
rect -371 -3757 -337 -3725
rect -371 -3825 -337 -3797
rect -371 -3893 -337 -3869
rect -371 -3961 -337 -3941
rect -371 -4029 -337 -4013
rect -371 -4097 -337 -4085
rect -371 -4165 -337 -4157
rect -371 -4233 -337 -4229
rect -371 -4339 -337 -4335
rect -371 -4411 -337 -4403
rect -371 -4483 -337 -4471
rect -371 -4555 -337 -4539
rect -371 -4627 -337 -4607
rect -371 -4699 -337 -4675
rect -371 -4771 -337 -4743
rect -371 -4843 -337 -4811
rect -371 -4913 -337 -4879
rect -371 -4981 -337 -4949
rect -371 -5049 -337 -5021
rect -371 -5117 -337 -5093
rect -371 -5185 -337 -5165
rect -371 -5253 -337 -5237
rect -371 -5321 -337 -5309
rect -371 -5389 -337 -5381
rect -371 -5457 -337 -5453
rect -371 -5563 -337 -5559
rect -371 -5635 -337 -5627
rect -371 -5707 -337 -5695
rect -371 -5779 -337 -5763
rect -371 -5851 -337 -5831
rect -371 -5923 -337 -5899
rect -371 -6004 -337 -5967
rect -253 5967 -219 6004
rect -253 5899 -219 5923
rect -253 5831 -219 5851
rect -253 5763 -219 5779
rect -253 5695 -219 5707
rect -253 5627 -219 5635
rect -253 5559 -219 5563
rect -253 5453 -219 5457
rect -253 5381 -219 5389
rect -253 5309 -219 5321
rect -253 5237 -219 5253
rect -253 5165 -219 5185
rect -253 5093 -219 5117
rect -253 5021 -219 5049
rect -253 4949 -219 4981
rect -253 4879 -219 4913
rect -253 4811 -219 4843
rect -253 4743 -219 4771
rect -253 4675 -219 4699
rect -253 4607 -219 4627
rect -253 4539 -219 4555
rect -253 4471 -219 4483
rect -253 4403 -219 4411
rect -253 4335 -219 4339
rect -253 4229 -219 4233
rect -253 4157 -219 4165
rect -253 4085 -219 4097
rect -253 4013 -219 4029
rect -253 3941 -219 3961
rect -253 3869 -219 3893
rect -253 3797 -219 3825
rect -253 3725 -219 3757
rect -253 3655 -219 3689
rect -253 3587 -219 3619
rect -253 3519 -219 3547
rect -253 3451 -219 3475
rect -253 3383 -219 3403
rect -253 3315 -219 3331
rect -253 3247 -219 3259
rect -253 3179 -219 3187
rect -253 3111 -219 3115
rect -253 3005 -219 3009
rect -253 2933 -219 2941
rect -253 2861 -219 2873
rect -253 2789 -219 2805
rect -253 2717 -219 2737
rect -253 2645 -219 2669
rect -253 2573 -219 2601
rect -253 2501 -219 2533
rect -253 2431 -219 2465
rect -253 2363 -219 2395
rect -253 2295 -219 2323
rect -253 2227 -219 2251
rect -253 2159 -219 2179
rect -253 2091 -219 2107
rect -253 2023 -219 2035
rect -253 1955 -219 1963
rect -253 1887 -219 1891
rect -253 1781 -219 1785
rect -253 1709 -219 1717
rect -253 1637 -219 1649
rect -253 1565 -219 1581
rect -253 1493 -219 1513
rect -253 1421 -219 1445
rect -253 1349 -219 1377
rect -253 1277 -219 1309
rect -253 1207 -219 1241
rect -253 1139 -219 1171
rect -253 1071 -219 1099
rect -253 1003 -219 1027
rect -253 935 -219 955
rect -253 867 -219 883
rect -253 799 -219 811
rect -253 731 -219 739
rect -253 663 -219 667
rect -253 557 -219 561
rect -253 485 -219 493
rect -253 413 -219 425
rect -253 341 -219 357
rect -253 269 -219 289
rect -253 197 -219 221
rect -253 125 -219 153
rect -253 53 -219 85
rect -253 -17 -219 17
rect -253 -85 -219 -53
rect -253 -153 -219 -125
rect -253 -221 -219 -197
rect -253 -289 -219 -269
rect -253 -357 -219 -341
rect -253 -425 -219 -413
rect -253 -493 -219 -485
rect -253 -561 -219 -557
rect -253 -667 -219 -663
rect -253 -739 -219 -731
rect -253 -811 -219 -799
rect -253 -883 -219 -867
rect -253 -955 -219 -935
rect -253 -1027 -219 -1003
rect -253 -1099 -219 -1071
rect -253 -1171 -219 -1139
rect -253 -1241 -219 -1207
rect -253 -1309 -219 -1277
rect -253 -1377 -219 -1349
rect -253 -1445 -219 -1421
rect -253 -1513 -219 -1493
rect -253 -1581 -219 -1565
rect -253 -1649 -219 -1637
rect -253 -1717 -219 -1709
rect -253 -1785 -219 -1781
rect -253 -1891 -219 -1887
rect -253 -1963 -219 -1955
rect -253 -2035 -219 -2023
rect -253 -2107 -219 -2091
rect -253 -2179 -219 -2159
rect -253 -2251 -219 -2227
rect -253 -2323 -219 -2295
rect -253 -2395 -219 -2363
rect -253 -2465 -219 -2431
rect -253 -2533 -219 -2501
rect -253 -2601 -219 -2573
rect -253 -2669 -219 -2645
rect -253 -2737 -219 -2717
rect -253 -2805 -219 -2789
rect -253 -2873 -219 -2861
rect -253 -2941 -219 -2933
rect -253 -3009 -219 -3005
rect -253 -3115 -219 -3111
rect -253 -3187 -219 -3179
rect -253 -3259 -219 -3247
rect -253 -3331 -219 -3315
rect -253 -3403 -219 -3383
rect -253 -3475 -219 -3451
rect -253 -3547 -219 -3519
rect -253 -3619 -219 -3587
rect -253 -3689 -219 -3655
rect -253 -3757 -219 -3725
rect -253 -3825 -219 -3797
rect -253 -3893 -219 -3869
rect -253 -3961 -219 -3941
rect -253 -4029 -219 -4013
rect -253 -4097 -219 -4085
rect -253 -4165 -219 -4157
rect -253 -4233 -219 -4229
rect -253 -4339 -219 -4335
rect -253 -4411 -219 -4403
rect -253 -4483 -219 -4471
rect -253 -4555 -219 -4539
rect -253 -4627 -219 -4607
rect -253 -4699 -219 -4675
rect -253 -4771 -219 -4743
rect -253 -4843 -219 -4811
rect -253 -4913 -219 -4879
rect -253 -4981 -219 -4949
rect -253 -5049 -219 -5021
rect -253 -5117 -219 -5093
rect -253 -5185 -219 -5165
rect -253 -5253 -219 -5237
rect -253 -5321 -219 -5309
rect -253 -5389 -219 -5381
rect -253 -5457 -219 -5453
rect -253 -5563 -219 -5559
rect -253 -5635 -219 -5627
rect -253 -5707 -219 -5695
rect -253 -5779 -219 -5763
rect -253 -5851 -219 -5831
rect -253 -5923 -219 -5899
rect -253 -6004 -219 -5967
rect -135 5967 -101 6004
rect -135 5899 -101 5923
rect -135 5831 -101 5851
rect -135 5763 -101 5779
rect -135 5695 -101 5707
rect -135 5627 -101 5635
rect -135 5559 -101 5563
rect -135 5453 -101 5457
rect -135 5381 -101 5389
rect -135 5309 -101 5321
rect -135 5237 -101 5253
rect -135 5165 -101 5185
rect -135 5093 -101 5117
rect -135 5021 -101 5049
rect -135 4949 -101 4981
rect -135 4879 -101 4913
rect -135 4811 -101 4843
rect -135 4743 -101 4771
rect -135 4675 -101 4699
rect -135 4607 -101 4627
rect -135 4539 -101 4555
rect -135 4471 -101 4483
rect -135 4403 -101 4411
rect -135 4335 -101 4339
rect -135 4229 -101 4233
rect -135 4157 -101 4165
rect -135 4085 -101 4097
rect -135 4013 -101 4029
rect -135 3941 -101 3961
rect -135 3869 -101 3893
rect -135 3797 -101 3825
rect -135 3725 -101 3757
rect -135 3655 -101 3689
rect -135 3587 -101 3619
rect -135 3519 -101 3547
rect -135 3451 -101 3475
rect -135 3383 -101 3403
rect -135 3315 -101 3331
rect -135 3247 -101 3259
rect -135 3179 -101 3187
rect -135 3111 -101 3115
rect -135 3005 -101 3009
rect -135 2933 -101 2941
rect -135 2861 -101 2873
rect -135 2789 -101 2805
rect -135 2717 -101 2737
rect -135 2645 -101 2669
rect -135 2573 -101 2601
rect -135 2501 -101 2533
rect -135 2431 -101 2465
rect -135 2363 -101 2395
rect -135 2295 -101 2323
rect -135 2227 -101 2251
rect -135 2159 -101 2179
rect -135 2091 -101 2107
rect -135 2023 -101 2035
rect -135 1955 -101 1963
rect -135 1887 -101 1891
rect -135 1781 -101 1785
rect -135 1709 -101 1717
rect -135 1637 -101 1649
rect -135 1565 -101 1581
rect -135 1493 -101 1513
rect -135 1421 -101 1445
rect -135 1349 -101 1377
rect -135 1277 -101 1309
rect -135 1207 -101 1241
rect -135 1139 -101 1171
rect -135 1071 -101 1099
rect -135 1003 -101 1027
rect -135 935 -101 955
rect -135 867 -101 883
rect -135 799 -101 811
rect -135 731 -101 739
rect -135 663 -101 667
rect -135 557 -101 561
rect -135 485 -101 493
rect -135 413 -101 425
rect -135 341 -101 357
rect -135 269 -101 289
rect -135 197 -101 221
rect -135 125 -101 153
rect -135 53 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -53
rect -135 -153 -101 -125
rect -135 -221 -101 -197
rect -135 -289 -101 -269
rect -135 -357 -101 -341
rect -135 -425 -101 -413
rect -135 -493 -101 -485
rect -135 -561 -101 -557
rect -135 -667 -101 -663
rect -135 -739 -101 -731
rect -135 -811 -101 -799
rect -135 -883 -101 -867
rect -135 -955 -101 -935
rect -135 -1027 -101 -1003
rect -135 -1099 -101 -1071
rect -135 -1171 -101 -1139
rect -135 -1241 -101 -1207
rect -135 -1309 -101 -1277
rect -135 -1377 -101 -1349
rect -135 -1445 -101 -1421
rect -135 -1513 -101 -1493
rect -135 -1581 -101 -1565
rect -135 -1649 -101 -1637
rect -135 -1717 -101 -1709
rect -135 -1785 -101 -1781
rect -135 -1891 -101 -1887
rect -135 -1963 -101 -1955
rect -135 -2035 -101 -2023
rect -135 -2107 -101 -2091
rect -135 -2179 -101 -2159
rect -135 -2251 -101 -2227
rect -135 -2323 -101 -2295
rect -135 -2395 -101 -2363
rect -135 -2465 -101 -2431
rect -135 -2533 -101 -2501
rect -135 -2601 -101 -2573
rect -135 -2669 -101 -2645
rect -135 -2737 -101 -2717
rect -135 -2805 -101 -2789
rect -135 -2873 -101 -2861
rect -135 -2941 -101 -2933
rect -135 -3009 -101 -3005
rect -135 -3115 -101 -3111
rect -135 -3187 -101 -3179
rect -135 -3259 -101 -3247
rect -135 -3331 -101 -3315
rect -135 -3403 -101 -3383
rect -135 -3475 -101 -3451
rect -135 -3547 -101 -3519
rect -135 -3619 -101 -3587
rect -135 -3689 -101 -3655
rect -135 -3757 -101 -3725
rect -135 -3825 -101 -3797
rect -135 -3893 -101 -3869
rect -135 -3961 -101 -3941
rect -135 -4029 -101 -4013
rect -135 -4097 -101 -4085
rect -135 -4165 -101 -4157
rect -135 -4233 -101 -4229
rect -135 -4339 -101 -4335
rect -135 -4411 -101 -4403
rect -135 -4483 -101 -4471
rect -135 -4555 -101 -4539
rect -135 -4627 -101 -4607
rect -135 -4699 -101 -4675
rect -135 -4771 -101 -4743
rect -135 -4843 -101 -4811
rect -135 -4913 -101 -4879
rect -135 -4981 -101 -4949
rect -135 -5049 -101 -5021
rect -135 -5117 -101 -5093
rect -135 -5185 -101 -5165
rect -135 -5253 -101 -5237
rect -135 -5321 -101 -5309
rect -135 -5389 -101 -5381
rect -135 -5457 -101 -5453
rect -135 -5563 -101 -5559
rect -135 -5635 -101 -5627
rect -135 -5707 -101 -5695
rect -135 -5779 -101 -5763
rect -135 -5851 -101 -5831
rect -135 -5923 -101 -5899
rect -135 -6004 -101 -5967
rect -17 5967 17 6004
rect -17 5899 17 5923
rect -17 5831 17 5851
rect -17 5763 17 5779
rect -17 5695 17 5707
rect -17 5627 17 5635
rect -17 5559 17 5563
rect -17 5453 17 5457
rect -17 5381 17 5389
rect -17 5309 17 5321
rect -17 5237 17 5253
rect -17 5165 17 5185
rect -17 5093 17 5117
rect -17 5021 17 5049
rect -17 4949 17 4981
rect -17 4879 17 4913
rect -17 4811 17 4843
rect -17 4743 17 4771
rect -17 4675 17 4699
rect -17 4607 17 4627
rect -17 4539 17 4555
rect -17 4471 17 4483
rect -17 4403 17 4411
rect -17 4335 17 4339
rect -17 4229 17 4233
rect -17 4157 17 4165
rect -17 4085 17 4097
rect -17 4013 17 4029
rect -17 3941 17 3961
rect -17 3869 17 3893
rect -17 3797 17 3825
rect -17 3725 17 3757
rect -17 3655 17 3689
rect -17 3587 17 3619
rect -17 3519 17 3547
rect -17 3451 17 3475
rect -17 3383 17 3403
rect -17 3315 17 3331
rect -17 3247 17 3259
rect -17 3179 17 3187
rect -17 3111 17 3115
rect -17 3005 17 3009
rect -17 2933 17 2941
rect -17 2861 17 2873
rect -17 2789 17 2805
rect -17 2717 17 2737
rect -17 2645 17 2669
rect -17 2573 17 2601
rect -17 2501 17 2533
rect -17 2431 17 2465
rect -17 2363 17 2395
rect -17 2295 17 2323
rect -17 2227 17 2251
rect -17 2159 17 2179
rect -17 2091 17 2107
rect -17 2023 17 2035
rect -17 1955 17 1963
rect -17 1887 17 1891
rect -17 1781 17 1785
rect -17 1709 17 1717
rect -17 1637 17 1649
rect -17 1565 17 1581
rect -17 1493 17 1513
rect -17 1421 17 1445
rect -17 1349 17 1377
rect -17 1277 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1171
rect -17 1071 17 1099
rect -17 1003 17 1027
rect -17 935 17 955
rect -17 867 17 883
rect -17 799 17 811
rect -17 731 17 739
rect -17 663 17 667
rect -17 557 17 561
rect -17 485 17 493
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -493 17 -485
rect -17 -561 17 -557
rect -17 -667 17 -663
rect -17 -739 17 -731
rect -17 -811 17 -799
rect -17 -883 17 -867
rect -17 -955 17 -935
rect -17 -1027 17 -1003
rect -17 -1099 17 -1071
rect -17 -1171 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1277
rect -17 -1377 17 -1349
rect -17 -1445 17 -1421
rect -17 -1513 17 -1493
rect -17 -1581 17 -1565
rect -17 -1649 17 -1637
rect -17 -1717 17 -1709
rect -17 -1785 17 -1781
rect -17 -1891 17 -1887
rect -17 -1963 17 -1955
rect -17 -2035 17 -2023
rect -17 -2107 17 -2091
rect -17 -2179 17 -2159
rect -17 -2251 17 -2227
rect -17 -2323 17 -2295
rect -17 -2395 17 -2363
rect -17 -2465 17 -2431
rect -17 -2533 17 -2501
rect -17 -2601 17 -2573
rect -17 -2669 17 -2645
rect -17 -2737 17 -2717
rect -17 -2805 17 -2789
rect -17 -2873 17 -2861
rect -17 -2941 17 -2933
rect -17 -3009 17 -3005
rect -17 -3115 17 -3111
rect -17 -3187 17 -3179
rect -17 -3259 17 -3247
rect -17 -3331 17 -3315
rect -17 -3403 17 -3383
rect -17 -3475 17 -3451
rect -17 -3547 17 -3519
rect -17 -3619 17 -3587
rect -17 -3689 17 -3655
rect -17 -3757 17 -3725
rect -17 -3825 17 -3797
rect -17 -3893 17 -3869
rect -17 -3961 17 -3941
rect -17 -4029 17 -4013
rect -17 -4097 17 -4085
rect -17 -4165 17 -4157
rect -17 -4233 17 -4229
rect -17 -4339 17 -4335
rect -17 -4411 17 -4403
rect -17 -4483 17 -4471
rect -17 -4555 17 -4539
rect -17 -4627 17 -4607
rect -17 -4699 17 -4675
rect -17 -4771 17 -4743
rect -17 -4843 17 -4811
rect -17 -4913 17 -4879
rect -17 -4981 17 -4949
rect -17 -5049 17 -5021
rect -17 -5117 17 -5093
rect -17 -5185 17 -5165
rect -17 -5253 17 -5237
rect -17 -5321 17 -5309
rect -17 -5389 17 -5381
rect -17 -5457 17 -5453
rect -17 -5563 17 -5559
rect -17 -5635 17 -5627
rect -17 -5707 17 -5695
rect -17 -5779 17 -5763
rect -17 -5851 17 -5831
rect -17 -5923 17 -5899
rect -17 -6004 17 -5967
rect 101 5967 135 6004
rect 101 5899 135 5923
rect 101 5831 135 5851
rect 101 5763 135 5779
rect 101 5695 135 5707
rect 101 5627 135 5635
rect 101 5559 135 5563
rect 101 5453 135 5457
rect 101 5381 135 5389
rect 101 5309 135 5321
rect 101 5237 135 5253
rect 101 5165 135 5185
rect 101 5093 135 5117
rect 101 5021 135 5049
rect 101 4949 135 4981
rect 101 4879 135 4913
rect 101 4811 135 4843
rect 101 4743 135 4771
rect 101 4675 135 4699
rect 101 4607 135 4627
rect 101 4539 135 4555
rect 101 4471 135 4483
rect 101 4403 135 4411
rect 101 4335 135 4339
rect 101 4229 135 4233
rect 101 4157 135 4165
rect 101 4085 135 4097
rect 101 4013 135 4029
rect 101 3941 135 3961
rect 101 3869 135 3893
rect 101 3797 135 3825
rect 101 3725 135 3757
rect 101 3655 135 3689
rect 101 3587 135 3619
rect 101 3519 135 3547
rect 101 3451 135 3475
rect 101 3383 135 3403
rect 101 3315 135 3331
rect 101 3247 135 3259
rect 101 3179 135 3187
rect 101 3111 135 3115
rect 101 3005 135 3009
rect 101 2933 135 2941
rect 101 2861 135 2873
rect 101 2789 135 2805
rect 101 2717 135 2737
rect 101 2645 135 2669
rect 101 2573 135 2601
rect 101 2501 135 2533
rect 101 2431 135 2465
rect 101 2363 135 2395
rect 101 2295 135 2323
rect 101 2227 135 2251
rect 101 2159 135 2179
rect 101 2091 135 2107
rect 101 2023 135 2035
rect 101 1955 135 1963
rect 101 1887 135 1891
rect 101 1781 135 1785
rect 101 1709 135 1717
rect 101 1637 135 1649
rect 101 1565 135 1581
rect 101 1493 135 1513
rect 101 1421 135 1445
rect 101 1349 135 1377
rect 101 1277 135 1309
rect 101 1207 135 1241
rect 101 1139 135 1171
rect 101 1071 135 1099
rect 101 1003 135 1027
rect 101 935 135 955
rect 101 867 135 883
rect 101 799 135 811
rect 101 731 135 739
rect 101 663 135 667
rect 101 557 135 561
rect 101 485 135 493
rect 101 413 135 425
rect 101 341 135 357
rect 101 269 135 289
rect 101 197 135 221
rect 101 125 135 153
rect 101 53 135 85
rect 101 -17 135 17
rect 101 -85 135 -53
rect 101 -153 135 -125
rect 101 -221 135 -197
rect 101 -289 135 -269
rect 101 -357 135 -341
rect 101 -425 135 -413
rect 101 -493 135 -485
rect 101 -561 135 -557
rect 101 -667 135 -663
rect 101 -739 135 -731
rect 101 -811 135 -799
rect 101 -883 135 -867
rect 101 -955 135 -935
rect 101 -1027 135 -1003
rect 101 -1099 135 -1071
rect 101 -1171 135 -1139
rect 101 -1241 135 -1207
rect 101 -1309 135 -1277
rect 101 -1377 135 -1349
rect 101 -1445 135 -1421
rect 101 -1513 135 -1493
rect 101 -1581 135 -1565
rect 101 -1649 135 -1637
rect 101 -1717 135 -1709
rect 101 -1785 135 -1781
rect 101 -1891 135 -1887
rect 101 -1963 135 -1955
rect 101 -2035 135 -2023
rect 101 -2107 135 -2091
rect 101 -2179 135 -2159
rect 101 -2251 135 -2227
rect 101 -2323 135 -2295
rect 101 -2395 135 -2363
rect 101 -2465 135 -2431
rect 101 -2533 135 -2501
rect 101 -2601 135 -2573
rect 101 -2669 135 -2645
rect 101 -2737 135 -2717
rect 101 -2805 135 -2789
rect 101 -2873 135 -2861
rect 101 -2941 135 -2933
rect 101 -3009 135 -3005
rect 101 -3115 135 -3111
rect 101 -3187 135 -3179
rect 101 -3259 135 -3247
rect 101 -3331 135 -3315
rect 101 -3403 135 -3383
rect 101 -3475 135 -3451
rect 101 -3547 135 -3519
rect 101 -3619 135 -3587
rect 101 -3689 135 -3655
rect 101 -3757 135 -3725
rect 101 -3825 135 -3797
rect 101 -3893 135 -3869
rect 101 -3961 135 -3941
rect 101 -4029 135 -4013
rect 101 -4097 135 -4085
rect 101 -4165 135 -4157
rect 101 -4233 135 -4229
rect 101 -4339 135 -4335
rect 101 -4411 135 -4403
rect 101 -4483 135 -4471
rect 101 -4555 135 -4539
rect 101 -4627 135 -4607
rect 101 -4699 135 -4675
rect 101 -4771 135 -4743
rect 101 -4843 135 -4811
rect 101 -4913 135 -4879
rect 101 -4981 135 -4949
rect 101 -5049 135 -5021
rect 101 -5117 135 -5093
rect 101 -5185 135 -5165
rect 101 -5253 135 -5237
rect 101 -5321 135 -5309
rect 101 -5389 135 -5381
rect 101 -5457 135 -5453
rect 101 -5563 135 -5559
rect 101 -5635 135 -5627
rect 101 -5707 135 -5695
rect 101 -5779 135 -5763
rect 101 -5851 135 -5831
rect 101 -5923 135 -5899
rect 101 -6004 135 -5967
rect 219 5967 253 6004
rect 219 5899 253 5923
rect 219 5831 253 5851
rect 219 5763 253 5779
rect 219 5695 253 5707
rect 219 5627 253 5635
rect 219 5559 253 5563
rect 219 5453 253 5457
rect 219 5381 253 5389
rect 219 5309 253 5321
rect 219 5237 253 5253
rect 219 5165 253 5185
rect 219 5093 253 5117
rect 219 5021 253 5049
rect 219 4949 253 4981
rect 219 4879 253 4913
rect 219 4811 253 4843
rect 219 4743 253 4771
rect 219 4675 253 4699
rect 219 4607 253 4627
rect 219 4539 253 4555
rect 219 4471 253 4483
rect 219 4403 253 4411
rect 219 4335 253 4339
rect 219 4229 253 4233
rect 219 4157 253 4165
rect 219 4085 253 4097
rect 219 4013 253 4029
rect 219 3941 253 3961
rect 219 3869 253 3893
rect 219 3797 253 3825
rect 219 3725 253 3757
rect 219 3655 253 3689
rect 219 3587 253 3619
rect 219 3519 253 3547
rect 219 3451 253 3475
rect 219 3383 253 3403
rect 219 3315 253 3331
rect 219 3247 253 3259
rect 219 3179 253 3187
rect 219 3111 253 3115
rect 219 3005 253 3009
rect 219 2933 253 2941
rect 219 2861 253 2873
rect 219 2789 253 2805
rect 219 2717 253 2737
rect 219 2645 253 2669
rect 219 2573 253 2601
rect 219 2501 253 2533
rect 219 2431 253 2465
rect 219 2363 253 2395
rect 219 2295 253 2323
rect 219 2227 253 2251
rect 219 2159 253 2179
rect 219 2091 253 2107
rect 219 2023 253 2035
rect 219 1955 253 1963
rect 219 1887 253 1891
rect 219 1781 253 1785
rect 219 1709 253 1717
rect 219 1637 253 1649
rect 219 1565 253 1581
rect 219 1493 253 1513
rect 219 1421 253 1445
rect 219 1349 253 1377
rect 219 1277 253 1309
rect 219 1207 253 1241
rect 219 1139 253 1171
rect 219 1071 253 1099
rect 219 1003 253 1027
rect 219 935 253 955
rect 219 867 253 883
rect 219 799 253 811
rect 219 731 253 739
rect 219 663 253 667
rect 219 557 253 561
rect 219 485 253 493
rect 219 413 253 425
rect 219 341 253 357
rect 219 269 253 289
rect 219 197 253 221
rect 219 125 253 153
rect 219 53 253 85
rect 219 -17 253 17
rect 219 -85 253 -53
rect 219 -153 253 -125
rect 219 -221 253 -197
rect 219 -289 253 -269
rect 219 -357 253 -341
rect 219 -425 253 -413
rect 219 -493 253 -485
rect 219 -561 253 -557
rect 219 -667 253 -663
rect 219 -739 253 -731
rect 219 -811 253 -799
rect 219 -883 253 -867
rect 219 -955 253 -935
rect 219 -1027 253 -1003
rect 219 -1099 253 -1071
rect 219 -1171 253 -1139
rect 219 -1241 253 -1207
rect 219 -1309 253 -1277
rect 219 -1377 253 -1349
rect 219 -1445 253 -1421
rect 219 -1513 253 -1493
rect 219 -1581 253 -1565
rect 219 -1649 253 -1637
rect 219 -1717 253 -1709
rect 219 -1785 253 -1781
rect 219 -1891 253 -1887
rect 219 -1963 253 -1955
rect 219 -2035 253 -2023
rect 219 -2107 253 -2091
rect 219 -2179 253 -2159
rect 219 -2251 253 -2227
rect 219 -2323 253 -2295
rect 219 -2395 253 -2363
rect 219 -2465 253 -2431
rect 219 -2533 253 -2501
rect 219 -2601 253 -2573
rect 219 -2669 253 -2645
rect 219 -2737 253 -2717
rect 219 -2805 253 -2789
rect 219 -2873 253 -2861
rect 219 -2941 253 -2933
rect 219 -3009 253 -3005
rect 219 -3115 253 -3111
rect 219 -3187 253 -3179
rect 219 -3259 253 -3247
rect 219 -3331 253 -3315
rect 219 -3403 253 -3383
rect 219 -3475 253 -3451
rect 219 -3547 253 -3519
rect 219 -3619 253 -3587
rect 219 -3689 253 -3655
rect 219 -3757 253 -3725
rect 219 -3825 253 -3797
rect 219 -3893 253 -3869
rect 219 -3961 253 -3941
rect 219 -4029 253 -4013
rect 219 -4097 253 -4085
rect 219 -4165 253 -4157
rect 219 -4233 253 -4229
rect 219 -4339 253 -4335
rect 219 -4411 253 -4403
rect 219 -4483 253 -4471
rect 219 -4555 253 -4539
rect 219 -4627 253 -4607
rect 219 -4699 253 -4675
rect 219 -4771 253 -4743
rect 219 -4843 253 -4811
rect 219 -4913 253 -4879
rect 219 -4981 253 -4949
rect 219 -5049 253 -5021
rect 219 -5117 253 -5093
rect 219 -5185 253 -5165
rect 219 -5253 253 -5237
rect 219 -5321 253 -5309
rect 219 -5389 253 -5381
rect 219 -5457 253 -5453
rect 219 -5563 253 -5559
rect 219 -5635 253 -5627
rect 219 -5707 253 -5695
rect 219 -5779 253 -5763
rect 219 -5851 253 -5831
rect 219 -5923 253 -5899
rect 219 -6004 253 -5967
rect 337 5967 371 6004
rect 337 5899 371 5923
rect 337 5831 371 5851
rect 337 5763 371 5779
rect 337 5695 371 5707
rect 337 5627 371 5635
rect 337 5559 371 5563
rect 337 5453 371 5457
rect 337 5381 371 5389
rect 337 5309 371 5321
rect 337 5237 371 5253
rect 337 5165 371 5185
rect 337 5093 371 5117
rect 337 5021 371 5049
rect 337 4949 371 4981
rect 337 4879 371 4913
rect 337 4811 371 4843
rect 337 4743 371 4771
rect 337 4675 371 4699
rect 337 4607 371 4627
rect 337 4539 371 4555
rect 337 4471 371 4483
rect 337 4403 371 4411
rect 337 4335 371 4339
rect 337 4229 371 4233
rect 337 4157 371 4165
rect 337 4085 371 4097
rect 337 4013 371 4029
rect 337 3941 371 3961
rect 337 3869 371 3893
rect 337 3797 371 3825
rect 337 3725 371 3757
rect 337 3655 371 3689
rect 337 3587 371 3619
rect 337 3519 371 3547
rect 337 3451 371 3475
rect 337 3383 371 3403
rect 337 3315 371 3331
rect 337 3247 371 3259
rect 337 3179 371 3187
rect 337 3111 371 3115
rect 337 3005 371 3009
rect 337 2933 371 2941
rect 337 2861 371 2873
rect 337 2789 371 2805
rect 337 2717 371 2737
rect 337 2645 371 2669
rect 337 2573 371 2601
rect 337 2501 371 2533
rect 337 2431 371 2465
rect 337 2363 371 2395
rect 337 2295 371 2323
rect 337 2227 371 2251
rect 337 2159 371 2179
rect 337 2091 371 2107
rect 337 2023 371 2035
rect 337 1955 371 1963
rect 337 1887 371 1891
rect 337 1781 371 1785
rect 337 1709 371 1717
rect 337 1637 371 1649
rect 337 1565 371 1581
rect 337 1493 371 1513
rect 337 1421 371 1445
rect 337 1349 371 1377
rect 337 1277 371 1309
rect 337 1207 371 1241
rect 337 1139 371 1171
rect 337 1071 371 1099
rect 337 1003 371 1027
rect 337 935 371 955
rect 337 867 371 883
rect 337 799 371 811
rect 337 731 371 739
rect 337 663 371 667
rect 337 557 371 561
rect 337 485 371 493
rect 337 413 371 425
rect 337 341 371 357
rect 337 269 371 289
rect 337 197 371 221
rect 337 125 371 153
rect 337 53 371 85
rect 337 -17 371 17
rect 337 -85 371 -53
rect 337 -153 371 -125
rect 337 -221 371 -197
rect 337 -289 371 -269
rect 337 -357 371 -341
rect 337 -425 371 -413
rect 337 -493 371 -485
rect 337 -561 371 -557
rect 337 -667 371 -663
rect 337 -739 371 -731
rect 337 -811 371 -799
rect 337 -883 371 -867
rect 337 -955 371 -935
rect 337 -1027 371 -1003
rect 337 -1099 371 -1071
rect 337 -1171 371 -1139
rect 337 -1241 371 -1207
rect 337 -1309 371 -1277
rect 337 -1377 371 -1349
rect 337 -1445 371 -1421
rect 337 -1513 371 -1493
rect 337 -1581 371 -1565
rect 337 -1649 371 -1637
rect 337 -1717 371 -1709
rect 337 -1785 371 -1781
rect 337 -1891 371 -1887
rect 337 -1963 371 -1955
rect 337 -2035 371 -2023
rect 337 -2107 371 -2091
rect 337 -2179 371 -2159
rect 337 -2251 371 -2227
rect 337 -2323 371 -2295
rect 337 -2395 371 -2363
rect 337 -2465 371 -2431
rect 337 -2533 371 -2501
rect 337 -2601 371 -2573
rect 337 -2669 371 -2645
rect 337 -2737 371 -2717
rect 337 -2805 371 -2789
rect 337 -2873 371 -2861
rect 337 -2941 371 -2933
rect 337 -3009 371 -3005
rect 337 -3115 371 -3111
rect 337 -3187 371 -3179
rect 337 -3259 371 -3247
rect 337 -3331 371 -3315
rect 337 -3403 371 -3383
rect 337 -3475 371 -3451
rect 337 -3547 371 -3519
rect 337 -3619 371 -3587
rect 337 -3689 371 -3655
rect 337 -3757 371 -3725
rect 337 -3825 371 -3797
rect 337 -3893 371 -3869
rect 337 -3961 371 -3941
rect 337 -4029 371 -4013
rect 337 -4097 371 -4085
rect 337 -4165 371 -4157
rect 337 -4233 371 -4229
rect 337 -4339 371 -4335
rect 337 -4411 371 -4403
rect 337 -4483 371 -4471
rect 337 -4555 371 -4539
rect 337 -4627 371 -4607
rect 337 -4699 371 -4675
rect 337 -4771 371 -4743
rect 337 -4843 371 -4811
rect 337 -4913 371 -4879
rect 337 -4981 371 -4949
rect 337 -5049 371 -5021
rect 337 -5117 371 -5093
rect 337 -5185 371 -5165
rect 337 -5253 371 -5237
rect 337 -5321 371 -5309
rect 337 -5389 371 -5381
rect 337 -5457 371 -5453
rect 337 -5563 371 -5559
rect 337 -5635 371 -5627
rect 337 -5707 371 -5695
rect 337 -5779 371 -5763
rect 337 -5851 371 -5831
rect 337 -5923 371 -5899
rect 337 -6004 371 -5967
rect 455 5967 489 6004
rect 455 5899 489 5923
rect 455 5831 489 5851
rect 455 5763 489 5779
rect 455 5695 489 5707
rect 455 5627 489 5635
rect 455 5559 489 5563
rect 455 5453 489 5457
rect 455 5381 489 5389
rect 455 5309 489 5321
rect 455 5237 489 5253
rect 455 5165 489 5185
rect 455 5093 489 5117
rect 455 5021 489 5049
rect 455 4949 489 4981
rect 455 4879 489 4913
rect 455 4811 489 4843
rect 455 4743 489 4771
rect 455 4675 489 4699
rect 455 4607 489 4627
rect 455 4539 489 4555
rect 455 4471 489 4483
rect 455 4403 489 4411
rect 455 4335 489 4339
rect 455 4229 489 4233
rect 455 4157 489 4165
rect 455 4085 489 4097
rect 455 4013 489 4029
rect 455 3941 489 3961
rect 455 3869 489 3893
rect 455 3797 489 3825
rect 455 3725 489 3757
rect 455 3655 489 3689
rect 455 3587 489 3619
rect 455 3519 489 3547
rect 455 3451 489 3475
rect 455 3383 489 3403
rect 455 3315 489 3331
rect 455 3247 489 3259
rect 455 3179 489 3187
rect 455 3111 489 3115
rect 455 3005 489 3009
rect 455 2933 489 2941
rect 455 2861 489 2873
rect 455 2789 489 2805
rect 455 2717 489 2737
rect 455 2645 489 2669
rect 455 2573 489 2601
rect 455 2501 489 2533
rect 455 2431 489 2465
rect 455 2363 489 2395
rect 455 2295 489 2323
rect 455 2227 489 2251
rect 455 2159 489 2179
rect 455 2091 489 2107
rect 455 2023 489 2035
rect 455 1955 489 1963
rect 455 1887 489 1891
rect 455 1781 489 1785
rect 455 1709 489 1717
rect 455 1637 489 1649
rect 455 1565 489 1581
rect 455 1493 489 1513
rect 455 1421 489 1445
rect 455 1349 489 1377
rect 455 1277 489 1309
rect 455 1207 489 1241
rect 455 1139 489 1171
rect 455 1071 489 1099
rect 455 1003 489 1027
rect 455 935 489 955
rect 455 867 489 883
rect 455 799 489 811
rect 455 731 489 739
rect 455 663 489 667
rect 455 557 489 561
rect 455 485 489 493
rect 455 413 489 425
rect 455 341 489 357
rect 455 269 489 289
rect 455 197 489 221
rect 455 125 489 153
rect 455 53 489 85
rect 455 -17 489 17
rect 455 -85 489 -53
rect 455 -153 489 -125
rect 455 -221 489 -197
rect 455 -289 489 -269
rect 455 -357 489 -341
rect 455 -425 489 -413
rect 455 -493 489 -485
rect 455 -561 489 -557
rect 455 -667 489 -663
rect 455 -739 489 -731
rect 455 -811 489 -799
rect 455 -883 489 -867
rect 455 -955 489 -935
rect 455 -1027 489 -1003
rect 455 -1099 489 -1071
rect 455 -1171 489 -1139
rect 455 -1241 489 -1207
rect 455 -1309 489 -1277
rect 455 -1377 489 -1349
rect 455 -1445 489 -1421
rect 455 -1513 489 -1493
rect 455 -1581 489 -1565
rect 455 -1649 489 -1637
rect 455 -1717 489 -1709
rect 455 -1785 489 -1781
rect 455 -1891 489 -1887
rect 455 -1963 489 -1955
rect 455 -2035 489 -2023
rect 455 -2107 489 -2091
rect 455 -2179 489 -2159
rect 455 -2251 489 -2227
rect 455 -2323 489 -2295
rect 455 -2395 489 -2363
rect 455 -2465 489 -2431
rect 455 -2533 489 -2501
rect 455 -2601 489 -2573
rect 455 -2669 489 -2645
rect 455 -2737 489 -2717
rect 455 -2805 489 -2789
rect 455 -2873 489 -2861
rect 455 -2941 489 -2933
rect 455 -3009 489 -3005
rect 455 -3115 489 -3111
rect 455 -3187 489 -3179
rect 455 -3259 489 -3247
rect 455 -3331 489 -3315
rect 455 -3403 489 -3383
rect 455 -3475 489 -3451
rect 455 -3547 489 -3519
rect 455 -3619 489 -3587
rect 455 -3689 489 -3655
rect 455 -3757 489 -3725
rect 455 -3825 489 -3797
rect 455 -3893 489 -3869
rect 455 -3961 489 -3941
rect 455 -4029 489 -4013
rect 455 -4097 489 -4085
rect 455 -4165 489 -4157
rect 455 -4233 489 -4229
rect 455 -4339 489 -4335
rect 455 -4411 489 -4403
rect 455 -4483 489 -4471
rect 455 -4555 489 -4539
rect 455 -4627 489 -4607
rect 455 -4699 489 -4675
rect 455 -4771 489 -4743
rect 455 -4843 489 -4811
rect 455 -4913 489 -4879
rect 455 -4981 489 -4949
rect 455 -5049 489 -5021
rect 455 -5117 489 -5093
rect 455 -5185 489 -5165
rect 455 -5253 489 -5237
rect 455 -5321 489 -5309
rect 455 -5389 489 -5381
rect 455 -5457 489 -5453
rect 455 -5563 489 -5559
rect 455 -5635 489 -5627
rect 455 -5707 489 -5695
rect 455 -5779 489 -5763
rect 455 -5851 489 -5831
rect 455 -5923 489 -5899
rect 455 -6004 489 -5967
rect 573 5967 607 6004
rect 573 5899 607 5923
rect 573 5831 607 5851
rect 573 5763 607 5779
rect 573 5695 607 5707
rect 573 5627 607 5635
rect 573 5559 607 5563
rect 573 5453 607 5457
rect 573 5381 607 5389
rect 573 5309 607 5321
rect 573 5237 607 5253
rect 573 5165 607 5185
rect 573 5093 607 5117
rect 573 5021 607 5049
rect 573 4949 607 4981
rect 573 4879 607 4913
rect 573 4811 607 4843
rect 573 4743 607 4771
rect 573 4675 607 4699
rect 573 4607 607 4627
rect 573 4539 607 4555
rect 573 4471 607 4483
rect 573 4403 607 4411
rect 573 4335 607 4339
rect 573 4229 607 4233
rect 573 4157 607 4165
rect 573 4085 607 4097
rect 573 4013 607 4029
rect 573 3941 607 3961
rect 573 3869 607 3893
rect 573 3797 607 3825
rect 573 3725 607 3757
rect 573 3655 607 3689
rect 573 3587 607 3619
rect 573 3519 607 3547
rect 573 3451 607 3475
rect 573 3383 607 3403
rect 573 3315 607 3331
rect 573 3247 607 3259
rect 573 3179 607 3187
rect 573 3111 607 3115
rect 573 3005 607 3009
rect 573 2933 607 2941
rect 573 2861 607 2873
rect 573 2789 607 2805
rect 573 2717 607 2737
rect 573 2645 607 2669
rect 573 2573 607 2601
rect 573 2501 607 2533
rect 573 2431 607 2465
rect 573 2363 607 2395
rect 573 2295 607 2323
rect 573 2227 607 2251
rect 573 2159 607 2179
rect 573 2091 607 2107
rect 573 2023 607 2035
rect 573 1955 607 1963
rect 573 1887 607 1891
rect 573 1781 607 1785
rect 573 1709 607 1717
rect 573 1637 607 1649
rect 573 1565 607 1581
rect 573 1493 607 1513
rect 573 1421 607 1445
rect 573 1349 607 1377
rect 573 1277 607 1309
rect 573 1207 607 1241
rect 573 1139 607 1171
rect 573 1071 607 1099
rect 573 1003 607 1027
rect 573 935 607 955
rect 573 867 607 883
rect 573 799 607 811
rect 573 731 607 739
rect 573 663 607 667
rect 573 557 607 561
rect 573 485 607 493
rect 573 413 607 425
rect 573 341 607 357
rect 573 269 607 289
rect 573 197 607 221
rect 573 125 607 153
rect 573 53 607 85
rect 573 -17 607 17
rect 573 -85 607 -53
rect 573 -153 607 -125
rect 573 -221 607 -197
rect 573 -289 607 -269
rect 573 -357 607 -341
rect 573 -425 607 -413
rect 573 -493 607 -485
rect 573 -561 607 -557
rect 573 -667 607 -663
rect 573 -739 607 -731
rect 573 -811 607 -799
rect 573 -883 607 -867
rect 573 -955 607 -935
rect 573 -1027 607 -1003
rect 573 -1099 607 -1071
rect 573 -1171 607 -1139
rect 573 -1241 607 -1207
rect 573 -1309 607 -1277
rect 573 -1377 607 -1349
rect 573 -1445 607 -1421
rect 573 -1513 607 -1493
rect 573 -1581 607 -1565
rect 573 -1649 607 -1637
rect 573 -1717 607 -1709
rect 573 -1785 607 -1781
rect 573 -1891 607 -1887
rect 573 -1963 607 -1955
rect 573 -2035 607 -2023
rect 573 -2107 607 -2091
rect 573 -2179 607 -2159
rect 573 -2251 607 -2227
rect 573 -2323 607 -2295
rect 573 -2395 607 -2363
rect 573 -2465 607 -2431
rect 573 -2533 607 -2501
rect 573 -2601 607 -2573
rect 573 -2669 607 -2645
rect 573 -2737 607 -2717
rect 573 -2805 607 -2789
rect 573 -2873 607 -2861
rect 573 -2941 607 -2933
rect 573 -3009 607 -3005
rect 573 -3115 607 -3111
rect 573 -3187 607 -3179
rect 573 -3259 607 -3247
rect 573 -3331 607 -3315
rect 573 -3403 607 -3383
rect 573 -3475 607 -3451
rect 573 -3547 607 -3519
rect 573 -3619 607 -3587
rect 573 -3689 607 -3655
rect 573 -3757 607 -3725
rect 573 -3825 607 -3797
rect 573 -3893 607 -3869
rect 573 -3961 607 -3941
rect 573 -4029 607 -4013
rect 573 -4097 607 -4085
rect 573 -4165 607 -4157
rect 573 -4233 607 -4229
rect 573 -4339 607 -4335
rect 573 -4411 607 -4403
rect 573 -4483 607 -4471
rect 573 -4555 607 -4539
rect 573 -4627 607 -4607
rect 573 -4699 607 -4675
rect 573 -4771 607 -4743
rect 573 -4843 607 -4811
rect 573 -4913 607 -4879
rect 573 -4981 607 -4949
rect 573 -5049 607 -5021
rect 573 -5117 607 -5093
rect 573 -5185 607 -5165
rect 573 -5253 607 -5237
rect 573 -5321 607 -5309
rect 573 -5389 607 -5381
rect 573 -5457 607 -5453
rect 573 -5563 607 -5559
rect 573 -5635 607 -5627
rect 573 -5707 607 -5695
rect 573 -5779 607 -5763
rect 573 -5851 607 -5831
rect 573 -5923 607 -5899
rect 573 -6004 607 -5967
<< viali >>
rect -548 6038 -514 6072
rect -607 5933 -573 5957
rect -607 5923 -573 5933
rect -607 5865 -573 5885
rect -607 5851 -573 5865
rect -607 5797 -573 5813
rect -607 5779 -573 5797
rect -607 5729 -573 5741
rect -607 5707 -573 5729
rect -607 5661 -573 5669
rect -607 5635 -573 5661
rect -607 5593 -573 5597
rect -607 5563 -573 5593
rect -607 5491 -573 5525
rect -607 5423 -573 5453
rect -607 5419 -573 5423
rect -607 5355 -573 5381
rect -607 5347 -573 5355
rect -607 5287 -573 5309
rect -607 5275 -573 5287
rect -607 5219 -573 5237
rect -607 5203 -573 5219
rect -607 5151 -573 5165
rect -607 5131 -573 5151
rect -607 5083 -573 5093
rect -607 5059 -573 5083
rect -607 5015 -573 5021
rect -607 4987 -573 5015
rect -607 4947 -573 4949
rect -607 4915 -573 4947
rect -607 4845 -573 4877
rect -607 4843 -573 4845
rect -607 4777 -573 4805
rect -607 4771 -573 4777
rect -607 4709 -573 4733
rect -607 4699 -573 4709
rect -607 4641 -573 4661
rect -607 4627 -573 4641
rect -607 4573 -573 4589
rect -607 4555 -573 4573
rect -607 4505 -573 4517
rect -607 4483 -573 4505
rect -607 4437 -573 4445
rect -607 4411 -573 4437
rect -607 4369 -573 4373
rect -607 4339 -573 4369
rect -607 4267 -573 4301
rect -607 4199 -573 4229
rect -607 4195 -573 4199
rect -607 4131 -573 4157
rect -607 4123 -573 4131
rect -607 4063 -573 4085
rect -607 4051 -573 4063
rect -607 3995 -573 4013
rect -607 3979 -573 3995
rect -607 3927 -573 3941
rect -607 3907 -573 3927
rect -607 3859 -573 3869
rect -607 3835 -573 3859
rect -607 3791 -573 3797
rect -607 3763 -573 3791
rect -607 3723 -573 3725
rect -607 3691 -573 3723
rect -607 3621 -573 3653
rect -607 3619 -573 3621
rect -607 3553 -573 3581
rect -607 3547 -573 3553
rect -607 3485 -573 3509
rect -607 3475 -573 3485
rect -607 3417 -573 3437
rect -607 3403 -573 3417
rect -607 3349 -573 3365
rect -607 3331 -573 3349
rect -607 3281 -573 3293
rect -607 3259 -573 3281
rect -607 3213 -573 3221
rect -607 3187 -573 3213
rect -607 3145 -573 3149
rect -607 3115 -573 3145
rect -607 3043 -573 3077
rect -607 2975 -573 3005
rect -607 2971 -573 2975
rect -607 2907 -573 2933
rect -607 2899 -573 2907
rect -607 2839 -573 2861
rect -607 2827 -573 2839
rect -607 2771 -573 2789
rect -607 2755 -573 2771
rect -607 2703 -573 2717
rect -607 2683 -573 2703
rect -607 2635 -573 2645
rect -607 2611 -573 2635
rect -607 2567 -573 2573
rect -607 2539 -573 2567
rect -607 2499 -573 2501
rect -607 2467 -573 2499
rect -607 2397 -573 2429
rect -607 2395 -573 2397
rect -607 2329 -573 2357
rect -607 2323 -573 2329
rect -607 2261 -573 2285
rect -607 2251 -573 2261
rect -607 2193 -573 2213
rect -607 2179 -573 2193
rect -607 2125 -573 2141
rect -607 2107 -573 2125
rect -607 2057 -573 2069
rect -607 2035 -573 2057
rect -607 1989 -573 1997
rect -607 1963 -573 1989
rect -607 1921 -573 1925
rect -607 1891 -573 1921
rect -607 1819 -573 1853
rect -607 1751 -573 1781
rect -607 1747 -573 1751
rect -607 1683 -573 1709
rect -607 1675 -573 1683
rect -607 1615 -573 1637
rect -607 1603 -573 1615
rect -607 1547 -573 1565
rect -607 1531 -573 1547
rect -607 1479 -573 1493
rect -607 1459 -573 1479
rect -607 1411 -573 1421
rect -607 1387 -573 1411
rect -607 1343 -573 1349
rect -607 1315 -573 1343
rect -607 1275 -573 1277
rect -607 1243 -573 1275
rect -607 1173 -573 1205
rect -607 1171 -573 1173
rect -607 1105 -573 1133
rect -607 1099 -573 1105
rect -607 1037 -573 1061
rect -607 1027 -573 1037
rect -607 969 -573 989
rect -607 955 -573 969
rect -607 901 -573 917
rect -607 883 -573 901
rect -607 833 -573 845
rect -607 811 -573 833
rect -607 765 -573 773
rect -607 739 -573 765
rect -607 697 -573 701
rect -607 667 -573 697
rect -607 595 -573 629
rect -607 527 -573 557
rect -607 523 -573 527
rect -607 459 -573 485
rect -607 451 -573 459
rect -607 391 -573 413
rect -607 379 -573 391
rect -607 323 -573 341
rect -607 307 -573 323
rect -607 255 -573 269
rect -607 235 -573 255
rect -607 187 -573 197
rect -607 163 -573 187
rect -607 119 -573 125
rect -607 91 -573 119
rect -607 51 -573 53
rect -607 19 -573 51
rect -607 -51 -573 -19
rect -607 -53 -573 -51
rect -607 -119 -573 -91
rect -607 -125 -573 -119
rect -607 -187 -573 -163
rect -607 -197 -573 -187
rect -607 -255 -573 -235
rect -607 -269 -573 -255
rect -607 -323 -573 -307
rect -607 -341 -573 -323
rect -607 -391 -573 -379
rect -607 -413 -573 -391
rect -607 -459 -573 -451
rect -607 -485 -573 -459
rect -607 -527 -573 -523
rect -607 -557 -573 -527
rect -607 -629 -573 -595
rect -607 -697 -573 -667
rect -607 -701 -573 -697
rect -607 -765 -573 -739
rect -607 -773 -573 -765
rect -607 -833 -573 -811
rect -607 -845 -573 -833
rect -607 -901 -573 -883
rect -607 -917 -573 -901
rect -607 -969 -573 -955
rect -607 -989 -573 -969
rect -607 -1037 -573 -1027
rect -607 -1061 -573 -1037
rect -607 -1105 -573 -1099
rect -607 -1133 -573 -1105
rect -607 -1173 -573 -1171
rect -607 -1205 -573 -1173
rect -607 -1275 -573 -1243
rect -607 -1277 -573 -1275
rect -607 -1343 -573 -1315
rect -607 -1349 -573 -1343
rect -607 -1411 -573 -1387
rect -607 -1421 -573 -1411
rect -607 -1479 -573 -1459
rect -607 -1493 -573 -1479
rect -607 -1547 -573 -1531
rect -607 -1565 -573 -1547
rect -607 -1615 -573 -1603
rect -607 -1637 -573 -1615
rect -607 -1683 -573 -1675
rect -607 -1709 -573 -1683
rect -607 -1751 -573 -1747
rect -607 -1781 -573 -1751
rect -607 -1853 -573 -1819
rect -607 -1921 -573 -1891
rect -607 -1925 -573 -1921
rect -607 -1989 -573 -1963
rect -607 -1997 -573 -1989
rect -607 -2057 -573 -2035
rect -607 -2069 -573 -2057
rect -607 -2125 -573 -2107
rect -607 -2141 -573 -2125
rect -607 -2193 -573 -2179
rect -607 -2213 -573 -2193
rect -607 -2261 -573 -2251
rect -607 -2285 -573 -2261
rect -607 -2329 -573 -2323
rect -607 -2357 -573 -2329
rect -607 -2397 -573 -2395
rect -607 -2429 -573 -2397
rect -607 -2499 -573 -2467
rect -607 -2501 -573 -2499
rect -607 -2567 -573 -2539
rect -607 -2573 -573 -2567
rect -607 -2635 -573 -2611
rect -607 -2645 -573 -2635
rect -607 -2703 -573 -2683
rect -607 -2717 -573 -2703
rect -607 -2771 -573 -2755
rect -607 -2789 -573 -2771
rect -607 -2839 -573 -2827
rect -607 -2861 -573 -2839
rect -607 -2907 -573 -2899
rect -607 -2933 -573 -2907
rect -607 -2975 -573 -2971
rect -607 -3005 -573 -2975
rect -607 -3077 -573 -3043
rect -607 -3145 -573 -3115
rect -607 -3149 -573 -3145
rect -607 -3213 -573 -3187
rect -607 -3221 -573 -3213
rect -607 -3281 -573 -3259
rect -607 -3293 -573 -3281
rect -607 -3349 -573 -3331
rect -607 -3365 -573 -3349
rect -607 -3417 -573 -3403
rect -607 -3437 -573 -3417
rect -607 -3485 -573 -3475
rect -607 -3509 -573 -3485
rect -607 -3553 -573 -3547
rect -607 -3581 -573 -3553
rect -607 -3621 -573 -3619
rect -607 -3653 -573 -3621
rect -607 -3723 -573 -3691
rect -607 -3725 -573 -3723
rect -607 -3791 -573 -3763
rect -607 -3797 -573 -3791
rect -607 -3859 -573 -3835
rect -607 -3869 -573 -3859
rect -607 -3927 -573 -3907
rect -607 -3941 -573 -3927
rect -607 -3995 -573 -3979
rect -607 -4013 -573 -3995
rect -607 -4063 -573 -4051
rect -607 -4085 -573 -4063
rect -607 -4131 -573 -4123
rect -607 -4157 -573 -4131
rect -607 -4199 -573 -4195
rect -607 -4229 -573 -4199
rect -607 -4301 -573 -4267
rect -607 -4369 -573 -4339
rect -607 -4373 -573 -4369
rect -607 -4437 -573 -4411
rect -607 -4445 -573 -4437
rect -607 -4505 -573 -4483
rect -607 -4517 -573 -4505
rect -607 -4573 -573 -4555
rect -607 -4589 -573 -4573
rect -607 -4641 -573 -4627
rect -607 -4661 -573 -4641
rect -607 -4709 -573 -4699
rect -607 -4733 -573 -4709
rect -607 -4777 -573 -4771
rect -607 -4805 -573 -4777
rect -607 -4845 -573 -4843
rect -607 -4877 -573 -4845
rect -607 -4947 -573 -4915
rect -607 -4949 -573 -4947
rect -607 -5015 -573 -4987
rect -607 -5021 -573 -5015
rect -607 -5083 -573 -5059
rect -607 -5093 -573 -5083
rect -607 -5151 -573 -5131
rect -607 -5165 -573 -5151
rect -607 -5219 -573 -5203
rect -607 -5237 -573 -5219
rect -607 -5287 -573 -5275
rect -607 -5309 -573 -5287
rect -607 -5355 -573 -5347
rect -607 -5381 -573 -5355
rect -607 -5423 -573 -5419
rect -607 -5453 -573 -5423
rect -607 -5525 -573 -5491
rect -607 -5593 -573 -5563
rect -607 -5597 -573 -5593
rect -607 -5661 -573 -5635
rect -607 -5669 -573 -5661
rect -607 -5729 -573 -5707
rect -607 -5741 -573 -5729
rect -607 -5797 -573 -5779
rect -607 -5813 -573 -5797
rect -607 -5865 -573 -5851
rect -607 -5885 -573 -5865
rect -607 -5933 -573 -5923
rect -607 -5957 -573 -5933
rect -489 5933 -455 5957
rect -489 5923 -455 5933
rect -489 5865 -455 5885
rect -489 5851 -455 5865
rect -489 5797 -455 5813
rect -489 5779 -455 5797
rect -489 5729 -455 5741
rect -489 5707 -455 5729
rect -489 5661 -455 5669
rect -489 5635 -455 5661
rect -489 5593 -455 5597
rect -489 5563 -455 5593
rect -489 5491 -455 5525
rect -489 5423 -455 5453
rect -489 5419 -455 5423
rect -489 5355 -455 5381
rect -489 5347 -455 5355
rect -489 5287 -455 5309
rect -489 5275 -455 5287
rect -489 5219 -455 5237
rect -489 5203 -455 5219
rect -489 5151 -455 5165
rect -489 5131 -455 5151
rect -489 5083 -455 5093
rect -489 5059 -455 5083
rect -489 5015 -455 5021
rect -489 4987 -455 5015
rect -489 4947 -455 4949
rect -489 4915 -455 4947
rect -489 4845 -455 4877
rect -489 4843 -455 4845
rect -489 4777 -455 4805
rect -489 4771 -455 4777
rect -489 4709 -455 4733
rect -489 4699 -455 4709
rect -489 4641 -455 4661
rect -489 4627 -455 4641
rect -489 4573 -455 4589
rect -489 4555 -455 4573
rect -489 4505 -455 4517
rect -489 4483 -455 4505
rect -489 4437 -455 4445
rect -489 4411 -455 4437
rect -489 4369 -455 4373
rect -489 4339 -455 4369
rect -489 4267 -455 4301
rect -489 4199 -455 4229
rect -489 4195 -455 4199
rect -489 4131 -455 4157
rect -489 4123 -455 4131
rect -489 4063 -455 4085
rect -489 4051 -455 4063
rect -489 3995 -455 4013
rect -489 3979 -455 3995
rect -489 3927 -455 3941
rect -489 3907 -455 3927
rect -489 3859 -455 3869
rect -489 3835 -455 3859
rect -489 3791 -455 3797
rect -489 3763 -455 3791
rect -489 3723 -455 3725
rect -489 3691 -455 3723
rect -489 3621 -455 3653
rect -489 3619 -455 3621
rect -489 3553 -455 3581
rect -489 3547 -455 3553
rect -489 3485 -455 3509
rect -489 3475 -455 3485
rect -489 3417 -455 3437
rect -489 3403 -455 3417
rect -489 3349 -455 3365
rect -489 3331 -455 3349
rect -489 3281 -455 3293
rect -489 3259 -455 3281
rect -489 3213 -455 3221
rect -489 3187 -455 3213
rect -489 3145 -455 3149
rect -489 3115 -455 3145
rect -489 3043 -455 3077
rect -489 2975 -455 3005
rect -489 2971 -455 2975
rect -489 2907 -455 2933
rect -489 2899 -455 2907
rect -489 2839 -455 2861
rect -489 2827 -455 2839
rect -489 2771 -455 2789
rect -489 2755 -455 2771
rect -489 2703 -455 2717
rect -489 2683 -455 2703
rect -489 2635 -455 2645
rect -489 2611 -455 2635
rect -489 2567 -455 2573
rect -489 2539 -455 2567
rect -489 2499 -455 2501
rect -489 2467 -455 2499
rect -489 2397 -455 2429
rect -489 2395 -455 2397
rect -489 2329 -455 2357
rect -489 2323 -455 2329
rect -489 2261 -455 2285
rect -489 2251 -455 2261
rect -489 2193 -455 2213
rect -489 2179 -455 2193
rect -489 2125 -455 2141
rect -489 2107 -455 2125
rect -489 2057 -455 2069
rect -489 2035 -455 2057
rect -489 1989 -455 1997
rect -489 1963 -455 1989
rect -489 1921 -455 1925
rect -489 1891 -455 1921
rect -489 1819 -455 1853
rect -489 1751 -455 1781
rect -489 1747 -455 1751
rect -489 1683 -455 1709
rect -489 1675 -455 1683
rect -489 1615 -455 1637
rect -489 1603 -455 1615
rect -489 1547 -455 1565
rect -489 1531 -455 1547
rect -489 1479 -455 1493
rect -489 1459 -455 1479
rect -489 1411 -455 1421
rect -489 1387 -455 1411
rect -489 1343 -455 1349
rect -489 1315 -455 1343
rect -489 1275 -455 1277
rect -489 1243 -455 1275
rect -489 1173 -455 1205
rect -489 1171 -455 1173
rect -489 1105 -455 1133
rect -489 1099 -455 1105
rect -489 1037 -455 1061
rect -489 1027 -455 1037
rect -489 969 -455 989
rect -489 955 -455 969
rect -489 901 -455 917
rect -489 883 -455 901
rect -489 833 -455 845
rect -489 811 -455 833
rect -489 765 -455 773
rect -489 739 -455 765
rect -489 697 -455 701
rect -489 667 -455 697
rect -489 595 -455 629
rect -489 527 -455 557
rect -489 523 -455 527
rect -489 459 -455 485
rect -489 451 -455 459
rect -489 391 -455 413
rect -489 379 -455 391
rect -489 323 -455 341
rect -489 307 -455 323
rect -489 255 -455 269
rect -489 235 -455 255
rect -489 187 -455 197
rect -489 163 -455 187
rect -489 119 -455 125
rect -489 91 -455 119
rect -489 51 -455 53
rect -489 19 -455 51
rect -489 -51 -455 -19
rect -489 -53 -455 -51
rect -489 -119 -455 -91
rect -489 -125 -455 -119
rect -489 -187 -455 -163
rect -489 -197 -455 -187
rect -489 -255 -455 -235
rect -489 -269 -455 -255
rect -489 -323 -455 -307
rect -489 -341 -455 -323
rect -489 -391 -455 -379
rect -489 -413 -455 -391
rect -489 -459 -455 -451
rect -489 -485 -455 -459
rect -489 -527 -455 -523
rect -489 -557 -455 -527
rect -489 -629 -455 -595
rect -489 -697 -455 -667
rect -489 -701 -455 -697
rect -489 -765 -455 -739
rect -489 -773 -455 -765
rect -489 -833 -455 -811
rect -489 -845 -455 -833
rect -489 -901 -455 -883
rect -489 -917 -455 -901
rect -489 -969 -455 -955
rect -489 -989 -455 -969
rect -489 -1037 -455 -1027
rect -489 -1061 -455 -1037
rect -489 -1105 -455 -1099
rect -489 -1133 -455 -1105
rect -489 -1173 -455 -1171
rect -489 -1205 -455 -1173
rect -489 -1275 -455 -1243
rect -489 -1277 -455 -1275
rect -489 -1343 -455 -1315
rect -489 -1349 -455 -1343
rect -489 -1411 -455 -1387
rect -489 -1421 -455 -1411
rect -489 -1479 -455 -1459
rect -489 -1493 -455 -1479
rect -489 -1547 -455 -1531
rect -489 -1565 -455 -1547
rect -489 -1615 -455 -1603
rect -489 -1637 -455 -1615
rect -489 -1683 -455 -1675
rect -489 -1709 -455 -1683
rect -489 -1751 -455 -1747
rect -489 -1781 -455 -1751
rect -489 -1853 -455 -1819
rect -489 -1921 -455 -1891
rect -489 -1925 -455 -1921
rect -489 -1989 -455 -1963
rect -489 -1997 -455 -1989
rect -489 -2057 -455 -2035
rect -489 -2069 -455 -2057
rect -489 -2125 -455 -2107
rect -489 -2141 -455 -2125
rect -489 -2193 -455 -2179
rect -489 -2213 -455 -2193
rect -489 -2261 -455 -2251
rect -489 -2285 -455 -2261
rect -489 -2329 -455 -2323
rect -489 -2357 -455 -2329
rect -489 -2397 -455 -2395
rect -489 -2429 -455 -2397
rect -489 -2499 -455 -2467
rect -489 -2501 -455 -2499
rect -489 -2567 -455 -2539
rect -489 -2573 -455 -2567
rect -489 -2635 -455 -2611
rect -489 -2645 -455 -2635
rect -489 -2703 -455 -2683
rect -489 -2717 -455 -2703
rect -489 -2771 -455 -2755
rect -489 -2789 -455 -2771
rect -489 -2839 -455 -2827
rect -489 -2861 -455 -2839
rect -489 -2907 -455 -2899
rect -489 -2933 -455 -2907
rect -489 -2975 -455 -2971
rect -489 -3005 -455 -2975
rect -489 -3077 -455 -3043
rect -489 -3145 -455 -3115
rect -489 -3149 -455 -3145
rect -489 -3213 -455 -3187
rect -489 -3221 -455 -3213
rect -489 -3281 -455 -3259
rect -489 -3293 -455 -3281
rect -489 -3349 -455 -3331
rect -489 -3365 -455 -3349
rect -489 -3417 -455 -3403
rect -489 -3437 -455 -3417
rect -489 -3485 -455 -3475
rect -489 -3509 -455 -3485
rect -489 -3553 -455 -3547
rect -489 -3581 -455 -3553
rect -489 -3621 -455 -3619
rect -489 -3653 -455 -3621
rect -489 -3723 -455 -3691
rect -489 -3725 -455 -3723
rect -489 -3791 -455 -3763
rect -489 -3797 -455 -3791
rect -489 -3859 -455 -3835
rect -489 -3869 -455 -3859
rect -489 -3927 -455 -3907
rect -489 -3941 -455 -3927
rect -489 -3995 -455 -3979
rect -489 -4013 -455 -3995
rect -489 -4063 -455 -4051
rect -489 -4085 -455 -4063
rect -489 -4131 -455 -4123
rect -489 -4157 -455 -4131
rect -489 -4199 -455 -4195
rect -489 -4229 -455 -4199
rect -489 -4301 -455 -4267
rect -489 -4369 -455 -4339
rect -489 -4373 -455 -4369
rect -489 -4437 -455 -4411
rect -489 -4445 -455 -4437
rect -489 -4505 -455 -4483
rect -489 -4517 -455 -4505
rect -489 -4573 -455 -4555
rect -489 -4589 -455 -4573
rect -489 -4641 -455 -4627
rect -489 -4661 -455 -4641
rect -489 -4709 -455 -4699
rect -489 -4733 -455 -4709
rect -489 -4777 -455 -4771
rect -489 -4805 -455 -4777
rect -489 -4845 -455 -4843
rect -489 -4877 -455 -4845
rect -489 -4947 -455 -4915
rect -489 -4949 -455 -4947
rect -489 -5015 -455 -4987
rect -489 -5021 -455 -5015
rect -489 -5083 -455 -5059
rect -489 -5093 -455 -5083
rect -489 -5151 -455 -5131
rect -489 -5165 -455 -5151
rect -489 -5219 -455 -5203
rect -489 -5237 -455 -5219
rect -489 -5287 -455 -5275
rect -489 -5309 -455 -5287
rect -489 -5355 -455 -5347
rect -489 -5381 -455 -5355
rect -489 -5423 -455 -5419
rect -489 -5453 -455 -5423
rect -489 -5525 -455 -5491
rect -489 -5593 -455 -5563
rect -489 -5597 -455 -5593
rect -489 -5661 -455 -5635
rect -489 -5669 -455 -5661
rect -489 -5729 -455 -5707
rect -489 -5741 -455 -5729
rect -489 -5797 -455 -5779
rect -489 -5813 -455 -5797
rect -489 -5865 -455 -5851
rect -489 -5885 -455 -5865
rect -489 -5933 -455 -5923
rect -489 -5957 -455 -5933
rect -371 5933 -337 5957
rect -371 5923 -337 5933
rect -371 5865 -337 5885
rect -371 5851 -337 5865
rect -371 5797 -337 5813
rect -371 5779 -337 5797
rect -371 5729 -337 5741
rect -371 5707 -337 5729
rect -371 5661 -337 5669
rect -371 5635 -337 5661
rect -371 5593 -337 5597
rect -371 5563 -337 5593
rect -371 5491 -337 5525
rect -371 5423 -337 5453
rect -371 5419 -337 5423
rect -371 5355 -337 5381
rect -371 5347 -337 5355
rect -371 5287 -337 5309
rect -371 5275 -337 5287
rect -371 5219 -337 5237
rect -371 5203 -337 5219
rect -371 5151 -337 5165
rect -371 5131 -337 5151
rect -371 5083 -337 5093
rect -371 5059 -337 5083
rect -371 5015 -337 5021
rect -371 4987 -337 5015
rect -371 4947 -337 4949
rect -371 4915 -337 4947
rect -371 4845 -337 4877
rect -371 4843 -337 4845
rect -371 4777 -337 4805
rect -371 4771 -337 4777
rect -371 4709 -337 4733
rect -371 4699 -337 4709
rect -371 4641 -337 4661
rect -371 4627 -337 4641
rect -371 4573 -337 4589
rect -371 4555 -337 4573
rect -371 4505 -337 4517
rect -371 4483 -337 4505
rect -371 4437 -337 4445
rect -371 4411 -337 4437
rect -371 4369 -337 4373
rect -371 4339 -337 4369
rect -371 4267 -337 4301
rect -371 4199 -337 4229
rect -371 4195 -337 4199
rect -371 4131 -337 4157
rect -371 4123 -337 4131
rect -371 4063 -337 4085
rect -371 4051 -337 4063
rect -371 3995 -337 4013
rect -371 3979 -337 3995
rect -371 3927 -337 3941
rect -371 3907 -337 3927
rect -371 3859 -337 3869
rect -371 3835 -337 3859
rect -371 3791 -337 3797
rect -371 3763 -337 3791
rect -371 3723 -337 3725
rect -371 3691 -337 3723
rect -371 3621 -337 3653
rect -371 3619 -337 3621
rect -371 3553 -337 3581
rect -371 3547 -337 3553
rect -371 3485 -337 3509
rect -371 3475 -337 3485
rect -371 3417 -337 3437
rect -371 3403 -337 3417
rect -371 3349 -337 3365
rect -371 3331 -337 3349
rect -371 3281 -337 3293
rect -371 3259 -337 3281
rect -371 3213 -337 3221
rect -371 3187 -337 3213
rect -371 3145 -337 3149
rect -371 3115 -337 3145
rect -371 3043 -337 3077
rect -371 2975 -337 3005
rect -371 2971 -337 2975
rect -371 2907 -337 2933
rect -371 2899 -337 2907
rect -371 2839 -337 2861
rect -371 2827 -337 2839
rect -371 2771 -337 2789
rect -371 2755 -337 2771
rect -371 2703 -337 2717
rect -371 2683 -337 2703
rect -371 2635 -337 2645
rect -371 2611 -337 2635
rect -371 2567 -337 2573
rect -371 2539 -337 2567
rect -371 2499 -337 2501
rect -371 2467 -337 2499
rect -371 2397 -337 2429
rect -371 2395 -337 2397
rect -371 2329 -337 2357
rect -371 2323 -337 2329
rect -371 2261 -337 2285
rect -371 2251 -337 2261
rect -371 2193 -337 2213
rect -371 2179 -337 2193
rect -371 2125 -337 2141
rect -371 2107 -337 2125
rect -371 2057 -337 2069
rect -371 2035 -337 2057
rect -371 1989 -337 1997
rect -371 1963 -337 1989
rect -371 1921 -337 1925
rect -371 1891 -337 1921
rect -371 1819 -337 1853
rect -371 1751 -337 1781
rect -371 1747 -337 1751
rect -371 1683 -337 1709
rect -371 1675 -337 1683
rect -371 1615 -337 1637
rect -371 1603 -337 1615
rect -371 1547 -337 1565
rect -371 1531 -337 1547
rect -371 1479 -337 1493
rect -371 1459 -337 1479
rect -371 1411 -337 1421
rect -371 1387 -337 1411
rect -371 1343 -337 1349
rect -371 1315 -337 1343
rect -371 1275 -337 1277
rect -371 1243 -337 1275
rect -371 1173 -337 1205
rect -371 1171 -337 1173
rect -371 1105 -337 1133
rect -371 1099 -337 1105
rect -371 1037 -337 1061
rect -371 1027 -337 1037
rect -371 969 -337 989
rect -371 955 -337 969
rect -371 901 -337 917
rect -371 883 -337 901
rect -371 833 -337 845
rect -371 811 -337 833
rect -371 765 -337 773
rect -371 739 -337 765
rect -371 697 -337 701
rect -371 667 -337 697
rect -371 595 -337 629
rect -371 527 -337 557
rect -371 523 -337 527
rect -371 459 -337 485
rect -371 451 -337 459
rect -371 391 -337 413
rect -371 379 -337 391
rect -371 323 -337 341
rect -371 307 -337 323
rect -371 255 -337 269
rect -371 235 -337 255
rect -371 187 -337 197
rect -371 163 -337 187
rect -371 119 -337 125
rect -371 91 -337 119
rect -371 51 -337 53
rect -371 19 -337 51
rect -371 -51 -337 -19
rect -371 -53 -337 -51
rect -371 -119 -337 -91
rect -371 -125 -337 -119
rect -371 -187 -337 -163
rect -371 -197 -337 -187
rect -371 -255 -337 -235
rect -371 -269 -337 -255
rect -371 -323 -337 -307
rect -371 -341 -337 -323
rect -371 -391 -337 -379
rect -371 -413 -337 -391
rect -371 -459 -337 -451
rect -371 -485 -337 -459
rect -371 -527 -337 -523
rect -371 -557 -337 -527
rect -371 -629 -337 -595
rect -371 -697 -337 -667
rect -371 -701 -337 -697
rect -371 -765 -337 -739
rect -371 -773 -337 -765
rect -371 -833 -337 -811
rect -371 -845 -337 -833
rect -371 -901 -337 -883
rect -371 -917 -337 -901
rect -371 -969 -337 -955
rect -371 -989 -337 -969
rect -371 -1037 -337 -1027
rect -371 -1061 -337 -1037
rect -371 -1105 -337 -1099
rect -371 -1133 -337 -1105
rect -371 -1173 -337 -1171
rect -371 -1205 -337 -1173
rect -371 -1275 -337 -1243
rect -371 -1277 -337 -1275
rect -371 -1343 -337 -1315
rect -371 -1349 -337 -1343
rect -371 -1411 -337 -1387
rect -371 -1421 -337 -1411
rect -371 -1479 -337 -1459
rect -371 -1493 -337 -1479
rect -371 -1547 -337 -1531
rect -371 -1565 -337 -1547
rect -371 -1615 -337 -1603
rect -371 -1637 -337 -1615
rect -371 -1683 -337 -1675
rect -371 -1709 -337 -1683
rect -371 -1751 -337 -1747
rect -371 -1781 -337 -1751
rect -371 -1853 -337 -1819
rect -371 -1921 -337 -1891
rect -371 -1925 -337 -1921
rect -371 -1989 -337 -1963
rect -371 -1997 -337 -1989
rect -371 -2057 -337 -2035
rect -371 -2069 -337 -2057
rect -371 -2125 -337 -2107
rect -371 -2141 -337 -2125
rect -371 -2193 -337 -2179
rect -371 -2213 -337 -2193
rect -371 -2261 -337 -2251
rect -371 -2285 -337 -2261
rect -371 -2329 -337 -2323
rect -371 -2357 -337 -2329
rect -371 -2397 -337 -2395
rect -371 -2429 -337 -2397
rect -371 -2499 -337 -2467
rect -371 -2501 -337 -2499
rect -371 -2567 -337 -2539
rect -371 -2573 -337 -2567
rect -371 -2635 -337 -2611
rect -371 -2645 -337 -2635
rect -371 -2703 -337 -2683
rect -371 -2717 -337 -2703
rect -371 -2771 -337 -2755
rect -371 -2789 -337 -2771
rect -371 -2839 -337 -2827
rect -371 -2861 -337 -2839
rect -371 -2907 -337 -2899
rect -371 -2933 -337 -2907
rect -371 -2975 -337 -2971
rect -371 -3005 -337 -2975
rect -371 -3077 -337 -3043
rect -371 -3145 -337 -3115
rect -371 -3149 -337 -3145
rect -371 -3213 -337 -3187
rect -371 -3221 -337 -3213
rect -371 -3281 -337 -3259
rect -371 -3293 -337 -3281
rect -371 -3349 -337 -3331
rect -371 -3365 -337 -3349
rect -371 -3417 -337 -3403
rect -371 -3437 -337 -3417
rect -371 -3485 -337 -3475
rect -371 -3509 -337 -3485
rect -371 -3553 -337 -3547
rect -371 -3581 -337 -3553
rect -371 -3621 -337 -3619
rect -371 -3653 -337 -3621
rect -371 -3723 -337 -3691
rect -371 -3725 -337 -3723
rect -371 -3791 -337 -3763
rect -371 -3797 -337 -3791
rect -371 -3859 -337 -3835
rect -371 -3869 -337 -3859
rect -371 -3927 -337 -3907
rect -371 -3941 -337 -3927
rect -371 -3995 -337 -3979
rect -371 -4013 -337 -3995
rect -371 -4063 -337 -4051
rect -371 -4085 -337 -4063
rect -371 -4131 -337 -4123
rect -371 -4157 -337 -4131
rect -371 -4199 -337 -4195
rect -371 -4229 -337 -4199
rect -371 -4301 -337 -4267
rect -371 -4369 -337 -4339
rect -371 -4373 -337 -4369
rect -371 -4437 -337 -4411
rect -371 -4445 -337 -4437
rect -371 -4505 -337 -4483
rect -371 -4517 -337 -4505
rect -371 -4573 -337 -4555
rect -371 -4589 -337 -4573
rect -371 -4641 -337 -4627
rect -371 -4661 -337 -4641
rect -371 -4709 -337 -4699
rect -371 -4733 -337 -4709
rect -371 -4777 -337 -4771
rect -371 -4805 -337 -4777
rect -371 -4845 -337 -4843
rect -371 -4877 -337 -4845
rect -371 -4947 -337 -4915
rect -371 -4949 -337 -4947
rect -371 -5015 -337 -4987
rect -371 -5021 -337 -5015
rect -371 -5083 -337 -5059
rect -371 -5093 -337 -5083
rect -371 -5151 -337 -5131
rect -371 -5165 -337 -5151
rect -371 -5219 -337 -5203
rect -371 -5237 -337 -5219
rect -371 -5287 -337 -5275
rect -371 -5309 -337 -5287
rect -371 -5355 -337 -5347
rect -371 -5381 -337 -5355
rect -371 -5423 -337 -5419
rect -371 -5453 -337 -5423
rect -371 -5525 -337 -5491
rect -371 -5593 -337 -5563
rect -371 -5597 -337 -5593
rect -371 -5661 -337 -5635
rect -371 -5669 -337 -5661
rect -371 -5729 -337 -5707
rect -371 -5741 -337 -5729
rect -371 -5797 -337 -5779
rect -371 -5813 -337 -5797
rect -371 -5865 -337 -5851
rect -371 -5885 -337 -5865
rect -371 -5933 -337 -5923
rect -371 -5957 -337 -5933
rect -253 5933 -219 5957
rect -253 5923 -219 5933
rect -253 5865 -219 5885
rect -253 5851 -219 5865
rect -253 5797 -219 5813
rect -253 5779 -219 5797
rect -253 5729 -219 5741
rect -253 5707 -219 5729
rect -253 5661 -219 5669
rect -253 5635 -219 5661
rect -253 5593 -219 5597
rect -253 5563 -219 5593
rect -253 5491 -219 5525
rect -253 5423 -219 5453
rect -253 5419 -219 5423
rect -253 5355 -219 5381
rect -253 5347 -219 5355
rect -253 5287 -219 5309
rect -253 5275 -219 5287
rect -253 5219 -219 5237
rect -253 5203 -219 5219
rect -253 5151 -219 5165
rect -253 5131 -219 5151
rect -253 5083 -219 5093
rect -253 5059 -219 5083
rect -253 5015 -219 5021
rect -253 4987 -219 5015
rect -253 4947 -219 4949
rect -253 4915 -219 4947
rect -253 4845 -219 4877
rect -253 4843 -219 4845
rect -253 4777 -219 4805
rect -253 4771 -219 4777
rect -253 4709 -219 4733
rect -253 4699 -219 4709
rect -253 4641 -219 4661
rect -253 4627 -219 4641
rect -253 4573 -219 4589
rect -253 4555 -219 4573
rect -253 4505 -219 4517
rect -253 4483 -219 4505
rect -253 4437 -219 4445
rect -253 4411 -219 4437
rect -253 4369 -219 4373
rect -253 4339 -219 4369
rect -253 4267 -219 4301
rect -253 4199 -219 4229
rect -253 4195 -219 4199
rect -253 4131 -219 4157
rect -253 4123 -219 4131
rect -253 4063 -219 4085
rect -253 4051 -219 4063
rect -253 3995 -219 4013
rect -253 3979 -219 3995
rect -253 3927 -219 3941
rect -253 3907 -219 3927
rect -253 3859 -219 3869
rect -253 3835 -219 3859
rect -253 3791 -219 3797
rect -253 3763 -219 3791
rect -253 3723 -219 3725
rect -253 3691 -219 3723
rect -253 3621 -219 3653
rect -253 3619 -219 3621
rect -253 3553 -219 3581
rect -253 3547 -219 3553
rect -253 3485 -219 3509
rect -253 3475 -219 3485
rect -253 3417 -219 3437
rect -253 3403 -219 3417
rect -253 3349 -219 3365
rect -253 3331 -219 3349
rect -253 3281 -219 3293
rect -253 3259 -219 3281
rect -253 3213 -219 3221
rect -253 3187 -219 3213
rect -253 3145 -219 3149
rect -253 3115 -219 3145
rect -253 3043 -219 3077
rect -253 2975 -219 3005
rect -253 2971 -219 2975
rect -253 2907 -219 2933
rect -253 2899 -219 2907
rect -253 2839 -219 2861
rect -253 2827 -219 2839
rect -253 2771 -219 2789
rect -253 2755 -219 2771
rect -253 2703 -219 2717
rect -253 2683 -219 2703
rect -253 2635 -219 2645
rect -253 2611 -219 2635
rect -253 2567 -219 2573
rect -253 2539 -219 2567
rect -253 2499 -219 2501
rect -253 2467 -219 2499
rect -253 2397 -219 2429
rect -253 2395 -219 2397
rect -253 2329 -219 2357
rect -253 2323 -219 2329
rect -253 2261 -219 2285
rect -253 2251 -219 2261
rect -253 2193 -219 2213
rect -253 2179 -219 2193
rect -253 2125 -219 2141
rect -253 2107 -219 2125
rect -253 2057 -219 2069
rect -253 2035 -219 2057
rect -253 1989 -219 1997
rect -253 1963 -219 1989
rect -253 1921 -219 1925
rect -253 1891 -219 1921
rect -253 1819 -219 1853
rect -253 1751 -219 1781
rect -253 1747 -219 1751
rect -253 1683 -219 1709
rect -253 1675 -219 1683
rect -253 1615 -219 1637
rect -253 1603 -219 1615
rect -253 1547 -219 1565
rect -253 1531 -219 1547
rect -253 1479 -219 1493
rect -253 1459 -219 1479
rect -253 1411 -219 1421
rect -253 1387 -219 1411
rect -253 1343 -219 1349
rect -253 1315 -219 1343
rect -253 1275 -219 1277
rect -253 1243 -219 1275
rect -253 1173 -219 1205
rect -253 1171 -219 1173
rect -253 1105 -219 1133
rect -253 1099 -219 1105
rect -253 1037 -219 1061
rect -253 1027 -219 1037
rect -253 969 -219 989
rect -253 955 -219 969
rect -253 901 -219 917
rect -253 883 -219 901
rect -253 833 -219 845
rect -253 811 -219 833
rect -253 765 -219 773
rect -253 739 -219 765
rect -253 697 -219 701
rect -253 667 -219 697
rect -253 595 -219 629
rect -253 527 -219 557
rect -253 523 -219 527
rect -253 459 -219 485
rect -253 451 -219 459
rect -253 391 -219 413
rect -253 379 -219 391
rect -253 323 -219 341
rect -253 307 -219 323
rect -253 255 -219 269
rect -253 235 -219 255
rect -253 187 -219 197
rect -253 163 -219 187
rect -253 119 -219 125
rect -253 91 -219 119
rect -253 51 -219 53
rect -253 19 -219 51
rect -253 -51 -219 -19
rect -253 -53 -219 -51
rect -253 -119 -219 -91
rect -253 -125 -219 -119
rect -253 -187 -219 -163
rect -253 -197 -219 -187
rect -253 -255 -219 -235
rect -253 -269 -219 -255
rect -253 -323 -219 -307
rect -253 -341 -219 -323
rect -253 -391 -219 -379
rect -253 -413 -219 -391
rect -253 -459 -219 -451
rect -253 -485 -219 -459
rect -253 -527 -219 -523
rect -253 -557 -219 -527
rect -253 -629 -219 -595
rect -253 -697 -219 -667
rect -253 -701 -219 -697
rect -253 -765 -219 -739
rect -253 -773 -219 -765
rect -253 -833 -219 -811
rect -253 -845 -219 -833
rect -253 -901 -219 -883
rect -253 -917 -219 -901
rect -253 -969 -219 -955
rect -253 -989 -219 -969
rect -253 -1037 -219 -1027
rect -253 -1061 -219 -1037
rect -253 -1105 -219 -1099
rect -253 -1133 -219 -1105
rect -253 -1173 -219 -1171
rect -253 -1205 -219 -1173
rect -253 -1275 -219 -1243
rect -253 -1277 -219 -1275
rect -253 -1343 -219 -1315
rect -253 -1349 -219 -1343
rect -253 -1411 -219 -1387
rect -253 -1421 -219 -1411
rect -253 -1479 -219 -1459
rect -253 -1493 -219 -1479
rect -253 -1547 -219 -1531
rect -253 -1565 -219 -1547
rect -253 -1615 -219 -1603
rect -253 -1637 -219 -1615
rect -253 -1683 -219 -1675
rect -253 -1709 -219 -1683
rect -253 -1751 -219 -1747
rect -253 -1781 -219 -1751
rect -253 -1853 -219 -1819
rect -253 -1921 -219 -1891
rect -253 -1925 -219 -1921
rect -253 -1989 -219 -1963
rect -253 -1997 -219 -1989
rect -253 -2057 -219 -2035
rect -253 -2069 -219 -2057
rect -253 -2125 -219 -2107
rect -253 -2141 -219 -2125
rect -253 -2193 -219 -2179
rect -253 -2213 -219 -2193
rect -253 -2261 -219 -2251
rect -253 -2285 -219 -2261
rect -253 -2329 -219 -2323
rect -253 -2357 -219 -2329
rect -253 -2397 -219 -2395
rect -253 -2429 -219 -2397
rect -253 -2499 -219 -2467
rect -253 -2501 -219 -2499
rect -253 -2567 -219 -2539
rect -253 -2573 -219 -2567
rect -253 -2635 -219 -2611
rect -253 -2645 -219 -2635
rect -253 -2703 -219 -2683
rect -253 -2717 -219 -2703
rect -253 -2771 -219 -2755
rect -253 -2789 -219 -2771
rect -253 -2839 -219 -2827
rect -253 -2861 -219 -2839
rect -253 -2907 -219 -2899
rect -253 -2933 -219 -2907
rect -253 -2975 -219 -2971
rect -253 -3005 -219 -2975
rect -253 -3077 -219 -3043
rect -253 -3145 -219 -3115
rect -253 -3149 -219 -3145
rect -253 -3213 -219 -3187
rect -253 -3221 -219 -3213
rect -253 -3281 -219 -3259
rect -253 -3293 -219 -3281
rect -253 -3349 -219 -3331
rect -253 -3365 -219 -3349
rect -253 -3417 -219 -3403
rect -253 -3437 -219 -3417
rect -253 -3485 -219 -3475
rect -253 -3509 -219 -3485
rect -253 -3553 -219 -3547
rect -253 -3581 -219 -3553
rect -253 -3621 -219 -3619
rect -253 -3653 -219 -3621
rect -253 -3723 -219 -3691
rect -253 -3725 -219 -3723
rect -253 -3791 -219 -3763
rect -253 -3797 -219 -3791
rect -253 -3859 -219 -3835
rect -253 -3869 -219 -3859
rect -253 -3927 -219 -3907
rect -253 -3941 -219 -3927
rect -253 -3995 -219 -3979
rect -253 -4013 -219 -3995
rect -253 -4063 -219 -4051
rect -253 -4085 -219 -4063
rect -253 -4131 -219 -4123
rect -253 -4157 -219 -4131
rect -253 -4199 -219 -4195
rect -253 -4229 -219 -4199
rect -253 -4301 -219 -4267
rect -253 -4369 -219 -4339
rect -253 -4373 -219 -4369
rect -253 -4437 -219 -4411
rect -253 -4445 -219 -4437
rect -253 -4505 -219 -4483
rect -253 -4517 -219 -4505
rect -253 -4573 -219 -4555
rect -253 -4589 -219 -4573
rect -253 -4641 -219 -4627
rect -253 -4661 -219 -4641
rect -253 -4709 -219 -4699
rect -253 -4733 -219 -4709
rect -253 -4777 -219 -4771
rect -253 -4805 -219 -4777
rect -253 -4845 -219 -4843
rect -253 -4877 -219 -4845
rect -253 -4947 -219 -4915
rect -253 -4949 -219 -4947
rect -253 -5015 -219 -4987
rect -253 -5021 -219 -5015
rect -253 -5083 -219 -5059
rect -253 -5093 -219 -5083
rect -253 -5151 -219 -5131
rect -253 -5165 -219 -5151
rect -253 -5219 -219 -5203
rect -253 -5237 -219 -5219
rect -253 -5287 -219 -5275
rect -253 -5309 -219 -5287
rect -253 -5355 -219 -5347
rect -253 -5381 -219 -5355
rect -253 -5423 -219 -5419
rect -253 -5453 -219 -5423
rect -253 -5525 -219 -5491
rect -253 -5593 -219 -5563
rect -253 -5597 -219 -5593
rect -253 -5661 -219 -5635
rect -253 -5669 -219 -5661
rect -253 -5729 -219 -5707
rect -253 -5741 -219 -5729
rect -253 -5797 -219 -5779
rect -253 -5813 -219 -5797
rect -253 -5865 -219 -5851
rect -253 -5885 -219 -5865
rect -253 -5933 -219 -5923
rect -253 -5957 -219 -5933
rect -135 5933 -101 5957
rect -135 5923 -101 5933
rect -135 5865 -101 5885
rect -135 5851 -101 5865
rect -135 5797 -101 5813
rect -135 5779 -101 5797
rect -135 5729 -101 5741
rect -135 5707 -101 5729
rect -135 5661 -101 5669
rect -135 5635 -101 5661
rect -135 5593 -101 5597
rect -135 5563 -101 5593
rect -135 5491 -101 5525
rect -135 5423 -101 5453
rect -135 5419 -101 5423
rect -135 5355 -101 5381
rect -135 5347 -101 5355
rect -135 5287 -101 5309
rect -135 5275 -101 5287
rect -135 5219 -101 5237
rect -135 5203 -101 5219
rect -135 5151 -101 5165
rect -135 5131 -101 5151
rect -135 5083 -101 5093
rect -135 5059 -101 5083
rect -135 5015 -101 5021
rect -135 4987 -101 5015
rect -135 4947 -101 4949
rect -135 4915 -101 4947
rect -135 4845 -101 4877
rect -135 4843 -101 4845
rect -135 4777 -101 4805
rect -135 4771 -101 4777
rect -135 4709 -101 4733
rect -135 4699 -101 4709
rect -135 4641 -101 4661
rect -135 4627 -101 4641
rect -135 4573 -101 4589
rect -135 4555 -101 4573
rect -135 4505 -101 4517
rect -135 4483 -101 4505
rect -135 4437 -101 4445
rect -135 4411 -101 4437
rect -135 4369 -101 4373
rect -135 4339 -101 4369
rect -135 4267 -101 4301
rect -135 4199 -101 4229
rect -135 4195 -101 4199
rect -135 4131 -101 4157
rect -135 4123 -101 4131
rect -135 4063 -101 4085
rect -135 4051 -101 4063
rect -135 3995 -101 4013
rect -135 3979 -101 3995
rect -135 3927 -101 3941
rect -135 3907 -101 3927
rect -135 3859 -101 3869
rect -135 3835 -101 3859
rect -135 3791 -101 3797
rect -135 3763 -101 3791
rect -135 3723 -101 3725
rect -135 3691 -101 3723
rect -135 3621 -101 3653
rect -135 3619 -101 3621
rect -135 3553 -101 3581
rect -135 3547 -101 3553
rect -135 3485 -101 3509
rect -135 3475 -101 3485
rect -135 3417 -101 3437
rect -135 3403 -101 3417
rect -135 3349 -101 3365
rect -135 3331 -101 3349
rect -135 3281 -101 3293
rect -135 3259 -101 3281
rect -135 3213 -101 3221
rect -135 3187 -101 3213
rect -135 3145 -101 3149
rect -135 3115 -101 3145
rect -135 3043 -101 3077
rect -135 2975 -101 3005
rect -135 2971 -101 2975
rect -135 2907 -101 2933
rect -135 2899 -101 2907
rect -135 2839 -101 2861
rect -135 2827 -101 2839
rect -135 2771 -101 2789
rect -135 2755 -101 2771
rect -135 2703 -101 2717
rect -135 2683 -101 2703
rect -135 2635 -101 2645
rect -135 2611 -101 2635
rect -135 2567 -101 2573
rect -135 2539 -101 2567
rect -135 2499 -101 2501
rect -135 2467 -101 2499
rect -135 2397 -101 2429
rect -135 2395 -101 2397
rect -135 2329 -101 2357
rect -135 2323 -101 2329
rect -135 2261 -101 2285
rect -135 2251 -101 2261
rect -135 2193 -101 2213
rect -135 2179 -101 2193
rect -135 2125 -101 2141
rect -135 2107 -101 2125
rect -135 2057 -101 2069
rect -135 2035 -101 2057
rect -135 1989 -101 1997
rect -135 1963 -101 1989
rect -135 1921 -101 1925
rect -135 1891 -101 1921
rect -135 1819 -101 1853
rect -135 1751 -101 1781
rect -135 1747 -101 1751
rect -135 1683 -101 1709
rect -135 1675 -101 1683
rect -135 1615 -101 1637
rect -135 1603 -101 1615
rect -135 1547 -101 1565
rect -135 1531 -101 1547
rect -135 1479 -101 1493
rect -135 1459 -101 1479
rect -135 1411 -101 1421
rect -135 1387 -101 1411
rect -135 1343 -101 1349
rect -135 1315 -101 1343
rect -135 1275 -101 1277
rect -135 1243 -101 1275
rect -135 1173 -101 1205
rect -135 1171 -101 1173
rect -135 1105 -101 1133
rect -135 1099 -101 1105
rect -135 1037 -101 1061
rect -135 1027 -101 1037
rect -135 969 -101 989
rect -135 955 -101 969
rect -135 901 -101 917
rect -135 883 -101 901
rect -135 833 -101 845
rect -135 811 -101 833
rect -135 765 -101 773
rect -135 739 -101 765
rect -135 697 -101 701
rect -135 667 -101 697
rect -135 595 -101 629
rect -135 527 -101 557
rect -135 523 -101 527
rect -135 459 -101 485
rect -135 451 -101 459
rect -135 391 -101 413
rect -135 379 -101 391
rect -135 323 -101 341
rect -135 307 -101 323
rect -135 255 -101 269
rect -135 235 -101 255
rect -135 187 -101 197
rect -135 163 -101 187
rect -135 119 -101 125
rect -135 91 -101 119
rect -135 51 -101 53
rect -135 19 -101 51
rect -135 -51 -101 -19
rect -135 -53 -101 -51
rect -135 -119 -101 -91
rect -135 -125 -101 -119
rect -135 -187 -101 -163
rect -135 -197 -101 -187
rect -135 -255 -101 -235
rect -135 -269 -101 -255
rect -135 -323 -101 -307
rect -135 -341 -101 -323
rect -135 -391 -101 -379
rect -135 -413 -101 -391
rect -135 -459 -101 -451
rect -135 -485 -101 -459
rect -135 -527 -101 -523
rect -135 -557 -101 -527
rect -135 -629 -101 -595
rect -135 -697 -101 -667
rect -135 -701 -101 -697
rect -135 -765 -101 -739
rect -135 -773 -101 -765
rect -135 -833 -101 -811
rect -135 -845 -101 -833
rect -135 -901 -101 -883
rect -135 -917 -101 -901
rect -135 -969 -101 -955
rect -135 -989 -101 -969
rect -135 -1037 -101 -1027
rect -135 -1061 -101 -1037
rect -135 -1105 -101 -1099
rect -135 -1133 -101 -1105
rect -135 -1173 -101 -1171
rect -135 -1205 -101 -1173
rect -135 -1275 -101 -1243
rect -135 -1277 -101 -1275
rect -135 -1343 -101 -1315
rect -135 -1349 -101 -1343
rect -135 -1411 -101 -1387
rect -135 -1421 -101 -1411
rect -135 -1479 -101 -1459
rect -135 -1493 -101 -1479
rect -135 -1547 -101 -1531
rect -135 -1565 -101 -1547
rect -135 -1615 -101 -1603
rect -135 -1637 -101 -1615
rect -135 -1683 -101 -1675
rect -135 -1709 -101 -1683
rect -135 -1751 -101 -1747
rect -135 -1781 -101 -1751
rect -135 -1853 -101 -1819
rect -135 -1921 -101 -1891
rect -135 -1925 -101 -1921
rect -135 -1989 -101 -1963
rect -135 -1997 -101 -1989
rect -135 -2057 -101 -2035
rect -135 -2069 -101 -2057
rect -135 -2125 -101 -2107
rect -135 -2141 -101 -2125
rect -135 -2193 -101 -2179
rect -135 -2213 -101 -2193
rect -135 -2261 -101 -2251
rect -135 -2285 -101 -2261
rect -135 -2329 -101 -2323
rect -135 -2357 -101 -2329
rect -135 -2397 -101 -2395
rect -135 -2429 -101 -2397
rect -135 -2499 -101 -2467
rect -135 -2501 -101 -2499
rect -135 -2567 -101 -2539
rect -135 -2573 -101 -2567
rect -135 -2635 -101 -2611
rect -135 -2645 -101 -2635
rect -135 -2703 -101 -2683
rect -135 -2717 -101 -2703
rect -135 -2771 -101 -2755
rect -135 -2789 -101 -2771
rect -135 -2839 -101 -2827
rect -135 -2861 -101 -2839
rect -135 -2907 -101 -2899
rect -135 -2933 -101 -2907
rect -135 -2975 -101 -2971
rect -135 -3005 -101 -2975
rect -135 -3077 -101 -3043
rect -135 -3145 -101 -3115
rect -135 -3149 -101 -3145
rect -135 -3213 -101 -3187
rect -135 -3221 -101 -3213
rect -135 -3281 -101 -3259
rect -135 -3293 -101 -3281
rect -135 -3349 -101 -3331
rect -135 -3365 -101 -3349
rect -135 -3417 -101 -3403
rect -135 -3437 -101 -3417
rect -135 -3485 -101 -3475
rect -135 -3509 -101 -3485
rect -135 -3553 -101 -3547
rect -135 -3581 -101 -3553
rect -135 -3621 -101 -3619
rect -135 -3653 -101 -3621
rect -135 -3723 -101 -3691
rect -135 -3725 -101 -3723
rect -135 -3791 -101 -3763
rect -135 -3797 -101 -3791
rect -135 -3859 -101 -3835
rect -135 -3869 -101 -3859
rect -135 -3927 -101 -3907
rect -135 -3941 -101 -3927
rect -135 -3995 -101 -3979
rect -135 -4013 -101 -3995
rect -135 -4063 -101 -4051
rect -135 -4085 -101 -4063
rect -135 -4131 -101 -4123
rect -135 -4157 -101 -4131
rect -135 -4199 -101 -4195
rect -135 -4229 -101 -4199
rect -135 -4301 -101 -4267
rect -135 -4369 -101 -4339
rect -135 -4373 -101 -4369
rect -135 -4437 -101 -4411
rect -135 -4445 -101 -4437
rect -135 -4505 -101 -4483
rect -135 -4517 -101 -4505
rect -135 -4573 -101 -4555
rect -135 -4589 -101 -4573
rect -135 -4641 -101 -4627
rect -135 -4661 -101 -4641
rect -135 -4709 -101 -4699
rect -135 -4733 -101 -4709
rect -135 -4777 -101 -4771
rect -135 -4805 -101 -4777
rect -135 -4845 -101 -4843
rect -135 -4877 -101 -4845
rect -135 -4947 -101 -4915
rect -135 -4949 -101 -4947
rect -135 -5015 -101 -4987
rect -135 -5021 -101 -5015
rect -135 -5083 -101 -5059
rect -135 -5093 -101 -5083
rect -135 -5151 -101 -5131
rect -135 -5165 -101 -5151
rect -135 -5219 -101 -5203
rect -135 -5237 -101 -5219
rect -135 -5287 -101 -5275
rect -135 -5309 -101 -5287
rect -135 -5355 -101 -5347
rect -135 -5381 -101 -5355
rect -135 -5423 -101 -5419
rect -135 -5453 -101 -5423
rect -135 -5525 -101 -5491
rect -135 -5593 -101 -5563
rect -135 -5597 -101 -5593
rect -135 -5661 -101 -5635
rect -135 -5669 -101 -5661
rect -135 -5729 -101 -5707
rect -135 -5741 -101 -5729
rect -135 -5797 -101 -5779
rect -135 -5813 -101 -5797
rect -135 -5865 -101 -5851
rect -135 -5885 -101 -5865
rect -135 -5933 -101 -5923
rect -135 -5957 -101 -5933
rect -17 5933 17 5957
rect -17 5923 17 5933
rect -17 5865 17 5885
rect -17 5851 17 5865
rect -17 5797 17 5813
rect -17 5779 17 5797
rect -17 5729 17 5741
rect -17 5707 17 5729
rect -17 5661 17 5669
rect -17 5635 17 5661
rect -17 5593 17 5597
rect -17 5563 17 5593
rect -17 5491 17 5525
rect -17 5423 17 5453
rect -17 5419 17 5423
rect -17 5355 17 5381
rect -17 5347 17 5355
rect -17 5287 17 5309
rect -17 5275 17 5287
rect -17 5219 17 5237
rect -17 5203 17 5219
rect -17 5151 17 5165
rect -17 5131 17 5151
rect -17 5083 17 5093
rect -17 5059 17 5083
rect -17 5015 17 5021
rect -17 4987 17 5015
rect -17 4947 17 4949
rect -17 4915 17 4947
rect -17 4845 17 4877
rect -17 4843 17 4845
rect -17 4777 17 4805
rect -17 4771 17 4777
rect -17 4709 17 4733
rect -17 4699 17 4709
rect -17 4641 17 4661
rect -17 4627 17 4641
rect -17 4573 17 4589
rect -17 4555 17 4573
rect -17 4505 17 4517
rect -17 4483 17 4505
rect -17 4437 17 4445
rect -17 4411 17 4437
rect -17 4369 17 4373
rect -17 4339 17 4369
rect -17 4267 17 4301
rect -17 4199 17 4229
rect -17 4195 17 4199
rect -17 4131 17 4157
rect -17 4123 17 4131
rect -17 4063 17 4085
rect -17 4051 17 4063
rect -17 3995 17 4013
rect -17 3979 17 3995
rect -17 3927 17 3941
rect -17 3907 17 3927
rect -17 3859 17 3869
rect -17 3835 17 3859
rect -17 3791 17 3797
rect -17 3763 17 3791
rect -17 3723 17 3725
rect -17 3691 17 3723
rect -17 3621 17 3653
rect -17 3619 17 3621
rect -17 3553 17 3581
rect -17 3547 17 3553
rect -17 3485 17 3509
rect -17 3475 17 3485
rect -17 3417 17 3437
rect -17 3403 17 3417
rect -17 3349 17 3365
rect -17 3331 17 3349
rect -17 3281 17 3293
rect -17 3259 17 3281
rect -17 3213 17 3221
rect -17 3187 17 3213
rect -17 3145 17 3149
rect -17 3115 17 3145
rect -17 3043 17 3077
rect -17 2975 17 3005
rect -17 2971 17 2975
rect -17 2907 17 2933
rect -17 2899 17 2907
rect -17 2839 17 2861
rect -17 2827 17 2839
rect -17 2771 17 2789
rect -17 2755 17 2771
rect -17 2703 17 2717
rect -17 2683 17 2703
rect -17 2635 17 2645
rect -17 2611 17 2635
rect -17 2567 17 2573
rect -17 2539 17 2567
rect -17 2499 17 2501
rect -17 2467 17 2499
rect -17 2397 17 2429
rect -17 2395 17 2397
rect -17 2329 17 2357
rect -17 2323 17 2329
rect -17 2261 17 2285
rect -17 2251 17 2261
rect -17 2193 17 2213
rect -17 2179 17 2193
rect -17 2125 17 2141
rect -17 2107 17 2125
rect -17 2057 17 2069
rect -17 2035 17 2057
rect -17 1989 17 1997
rect -17 1963 17 1989
rect -17 1921 17 1925
rect -17 1891 17 1921
rect -17 1819 17 1853
rect -17 1751 17 1781
rect -17 1747 17 1751
rect -17 1683 17 1709
rect -17 1675 17 1683
rect -17 1615 17 1637
rect -17 1603 17 1615
rect -17 1547 17 1565
rect -17 1531 17 1547
rect -17 1479 17 1493
rect -17 1459 17 1479
rect -17 1411 17 1421
rect -17 1387 17 1411
rect -17 1343 17 1349
rect -17 1315 17 1343
rect -17 1275 17 1277
rect -17 1243 17 1275
rect -17 1173 17 1205
rect -17 1171 17 1173
rect -17 1105 17 1133
rect -17 1099 17 1105
rect -17 1037 17 1061
rect -17 1027 17 1037
rect -17 969 17 989
rect -17 955 17 969
rect -17 901 17 917
rect -17 883 17 901
rect -17 833 17 845
rect -17 811 17 833
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect -17 -833 17 -811
rect -17 -845 17 -833
rect -17 -901 17 -883
rect -17 -917 17 -901
rect -17 -969 17 -955
rect -17 -989 17 -969
rect -17 -1037 17 -1027
rect -17 -1061 17 -1037
rect -17 -1105 17 -1099
rect -17 -1133 17 -1105
rect -17 -1173 17 -1171
rect -17 -1205 17 -1173
rect -17 -1275 17 -1243
rect -17 -1277 17 -1275
rect -17 -1343 17 -1315
rect -17 -1349 17 -1343
rect -17 -1411 17 -1387
rect -17 -1421 17 -1411
rect -17 -1479 17 -1459
rect -17 -1493 17 -1479
rect -17 -1547 17 -1531
rect -17 -1565 17 -1547
rect -17 -1615 17 -1603
rect -17 -1637 17 -1615
rect -17 -1683 17 -1675
rect -17 -1709 17 -1683
rect -17 -1751 17 -1747
rect -17 -1781 17 -1751
rect -17 -1853 17 -1819
rect -17 -1921 17 -1891
rect -17 -1925 17 -1921
rect -17 -1989 17 -1963
rect -17 -1997 17 -1989
rect -17 -2057 17 -2035
rect -17 -2069 17 -2057
rect -17 -2125 17 -2107
rect -17 -2141 17 -2125
rect -17 -2193 17 -2179
rect -17 -2213 17 -2193
rect -17 -2261 17 -2251
rect -17 -2285 17 -2261
rect -17 -2329 17 -2323
rect -17 -2357 17 -2329
rect -17 -2397 17 -2395
rect -17 -2429 17 -2397
rect -17 -2499 17 -2467
rect -17 -2501 17 -2499
rect -17 -2567 17 -2539
rect -17 -2573 17 -2567
rect -17 -2635 17 -2611
rect -17 -2645 17 -2635
rect -17 -2703 17 -2683
rect -17 -2717 17 -2703
rect -17 -2771 17 -2755
rect -17 -2789 17 -2771
rect -17 -2839 17 -2827
rect -17 -2861 17 -2839
rect -17 -2907 17 -2899
rect -17 -2933 17 -2907
rect -17 -2975 17 -2971
rect -17 -3005 17 -2975
rect -17 -3077 17 -3043
rect -17 -3145 17 -3115
rect -17 -3149 17 -3145
rect -17 -3213 17 -3187
rect -17 -3221 17 -3213
rect -17 -3281 17 -3259
rect -17 -3293 17 -3281
rect -17 -3349 17 -3331
rect -17 -3365 17 -3349
rect -17 -3417 17 -3403
rect -17 -3437 17 -3417
rect -17 -3485 17 -3475
rect -17 -3509 17 -3485
rect -17 -3553 17 -3547
rect -17 -3581 17 -3553
rect -17 -3621 17 -3619
rect -17 -3653 17 -3621
rect -17 -3723 17 -3691
rect -17 -3725 17 -3723
rect -17 -3791 17 -3763
rect -17 -3797 17 -3791
rect -17 -3859 17 -3835
rect -17 -3869 17 -3859
rect -17 -3927 17 -3907
rect -17 -3941 17 -3927
rect -17 -3995 17 -3979
rect -17 -4013 17 -3995
rect -17 -4063 17 -4051
rect -17 -4085 17 -4063
rect -17 -4131 17 -4123
rect -17 -4157 17 -4131
rect -17 -4199 17 -4195
rect -17 -4229 17 -4199
rect -17 -4301 17 -4267
rect -17 -4369 17 -4339
rect -17 -4373 17 -4369
rect -17 -4437 17 -4411
rect -17 -4445 17 -4437
rect -17 -4505 17 -4483
rect -17 -4517 17 -4505
rect -17 -4573 17 -4555
rect -17 -4589 17 -4573
rect -17 -4641 17 -4627
rect -17 -4661 17 -4641
rect -17 -4709 17 -4699
rect -17 -4733 17 -4709
rect -17 -4777 17 -4771
rect -17 -4805 17 -4777
rect -17 -4845 17 -4843
rect -17 -4877 17 -4845
rect -17 -4947 17 -4915
rect -17 -4949 17 -4947
rect -17 -5015 17 -4987
rect -17 -5021 17 -5015
rect -17 -5083 17 -5059
rect -17 -5093 17 -5083
rect -17 -5151 17 -5131
rect -17 -5165 17 -5151
rect -17 -5219 17 -5203
rect -17 -5237 17 -5219
rect -17 -5287 17 -5275
rect -17 -5309 17 -5287
rect -17 -5355 17 -5347
rect -17 -5381 17 -5355
rect -17 -5423 17 -5419
rect -17 -5453 17 -5423
rect -17 -5525 17 -5491
rect -17 -5593 17 -5563
rect -17 -5597 17 -5593
rect -17 -5661 17 -5635
rect -17 -5669 17 -5661
rect -17 -5729 17 -5707
rect -17 -5741 17 -5729
rect -17 -5797 17 -5779
rect -17 -5813 17 -5797
rect -17 -5865 17 -5851
rect -17 -5885 17 -5865
rect -17 -5933 17 -5923
rect -17 -5957 17 -5933
rect 101 5933 135 5957
rect 101 5923 135 5933
rect 101 5865 135 5885
rect 101 5851 135 5865
rect 101 5797 135 5813
rect 101 5779 135 5797
rect 101 5729 135 5741
rect 101 5707 135 5729
rect 101 5661 135 5669
rect 101 5635 135 5661
rect 101 5593 135 5597
rect 101 5563 135 5593
rect 101 5491 135 5525
rect 101 5423 135 5453
rect 101 5419 135 5423
rect 101 5355 135 5381
rect 101 5347 135 5355
rect 101 5287 135 5309
rect 101 5275 135 5287
rect 101 5219 135 5237
rect 101 5203 135 5219
rect 101 5151 135 5165
rect 101 5131 135 5151
rect 101 5083 135 5093
rect 101 5059 135 5083
rect 101 5015 135 5021
rect 101 4987 135 5015
rect 101 4947 135 4949
rect 101 4915 135 4947
rect 101 4845 135 4877
rect 101 4843 135 4845
rect 101 4777 135 4805
rect 101 4771 135 4777
rect 101 4709 135 4733
rect 101 4699 135 4709
rect 101 4641 135 4661
rect 101 4627 135 4641
rect 101 4573 135 4589
rect 101 4555 135 4573
rect 101 4505 135 4517
rect 101 4483 135 4505
rect 101 4437 135 4445
rect 101 4411 135 4437
rect 101 4369 135 4373
rect 101 4339 135 4369
rect 101 4267 135 4301
rect 101 4199 135 4229
rect 101 4195 135 4199
rect 101 4131 135 4157
rect 101 4123 135 4131
rect 101 4063 135 4085
rect 101 4051 135 4063
rect 101 3995 135 4013
rect 101 3979 135 3995
rect 101 3927 135 3941
rect 101 3907 135 3927
rect 101 3859 135 3869
rect 101 3835 135 3859
rect 101 3791 135 3797
rect 101 3763 135 3791
rect 101 3723 135 3725
rect 101 3691 135 3723
rect 101 3621 135 3653
rect 101 3619 135 3621
rect 101 3553 135 3581
rect 101 3547 135 3553
rect 101 3485 135 3509
rect 101 3475 135 3485
rect 101 3417 135 3437
rect 101 3403 135 3417
rect 101 3349 135 3365
rect 101 3331 135 3349
rect 101 3281 135 3293
rect 101 3259 135 3281
rect 101 3213 135 3221
rect 101 3187 135 3213
rect 101 3145 135 3149
rect 101 3115 135 3145
rect 101 3043 135 3077
rect 101 2975 135 3005
rect 101 2971 135 2975
rect 101 2907 135 2933
rect 101 2899 135 2907
rect 101 2839 135 2861
rect 101 2827 135 2839
rect 101 2771 135 2789
rect 101 2755 135 2771
rect 101 2703 135 2717
rect 101 2683 135 2703
rect 101 2635 135 2645
rect 101 2611 135 2635
rect 101 2567 135 2573
rect 101 2539 135 2567
rect 101 2499 135 2501
rect 101 2467 135 2499
rect 101 2397 135 2429
rect 101 2395 135 2397
rect 101 2329 135 2357
rect 101 2323 135 2329
rect 101 2261 135 2285
rect 101 2251 135 2261
rect 101 2193 135 2213
rect 101 2179 135 2193
rect 101 2125 135 2141
rect 101 2107 135 2125
rect 101 2057 135 2069
rect 101 2035 135 2057
rect 101 1989 135 1997
rect 101 1963 135 1989
rect 101 1921 135 1925
rect 101 1891 135 1921
rect 101 1819 135 1853
rect 101 1751 135 1781
rect 101 1747 135 1751
rect 101 1683 135 1709
rect 101 1675 135 1683
rect 101 1615 135 1637
rect 101 1603 135 1615
rect 101 1547 135 1565
rect 101 1531 135 1547
rect 101 1479 135 1493
rect 101 1459 135 1479
rect 101 1411 135 1421
rect 101 1387 135 1411
rect 101 1343 135 1349
rect 101 1315 135 1343
rect 101 1275 135 1277
rect 101 1243 135 1275
rect 101 1173 135 1205
rect 101 1171 135 1173
rect 101 1105 135 1133
rect 101 1099 135 1105
rect 101 1037 135 1061
rect 101 1027 135 1037
rect 101 969 135 989
rect 101 955 135 969
rect 101 901 135 917
rect 101 883 135 901
rect 101 833 135 845
rect 101 811 135 833
rect 101 765 135 773
rect 101 739 135 765
rect 101 697 135 701
rect 101 667 135 697
rect 101 595 135 629
rect 101 527 135 557
rect 101 523 135 527
rect 101 459 135 485
rect 101 451 135 459
rect 101 391 135 413
rect 101 379 135 391
rect 101 323 135 341
rect 101 307 135 323
rect 101 255 135 269
rect 101 235 135 255
rect 101 187 135 197
rect 101 163 135 187
rect 101 119 135 125
rect 101 91 135 119
rect 101 51 135 53
rect 101 19 135 51
rect 101 -51 135 -19
rect 101 -53 135 -51
rect 101 -119 135 -91
rect 101 -125 135 -119
rect 101 -187 135 -163
rect 101 -197 135 -187
rect 101 -255 135 -235
rect 101 -269 135 -255
rect 101 -323 135 -307
rect 101 -341 135 -323
rect 101 -391 135 -379
rect 101 -413 135 -391
rect 101 -459 135 -451
rect 101 -485 135 -459
rect 101 -527 135 -523
rect 101 -557 135 -527
rect 101 -629 135 -595
rect 101 -697 135 -667
rect 101 -701 135 -697
rect 101 -765 135 -739
rect 101 -773 135 -765
rect 101 -833 135 -811
rect 101 -845 135 -833
rect 101 -901 135 -883
rect 101 -917 135 -901
rect 101 -969 135 -955
rect 101 -989 135 -969
rect 101 -1037 135 -1027
rect 101 -1061 135 -1037
rect 101 -1105 135 -1099
rect 101 -1133 135 -1105
rect 101 -1173 135 -1171
rect 101 -1205 135 -1173
rect 101 -1275 135 -1243
rect 101 -1277 135 -1275
rect 101 -1343 135 -1315
rect 101 -1349 135 -1343
rect 101 -1411 135 -1387
rect 101 -1421 135 -1411
rect 101 -1479 135 -1459
rect 101 -1493 135 -1479
rect 101 -1547 135 -1531
rect 101 -1565 135 -1547
rect 101 -1615 135 -1603
rect 101 -1637 135 -1615
rect 101 -1683 135 -1675
rect 101 -1709 135 -1683
rect 101 -1751 135 -1747
rect 101 -1781 135 -1751
rect 101 -1853 135 -1819
rect 101 -1921 135 -1891
rect 101 -1925 135 -1921
rect 101 -1989 135 -1963
rect 101 -1997 135 -1989
rect 101 -2057 135 -2035
rect 101 -2069 135 -2057
rect 101 -2125 135 -2107
rect 101 -2141 135 -2125
rect 101 -2193 135 -2179
rect 101 -2213 135 -2193
rect 101 -2261 135 -2251
rect 101 -2285 135 -2261
rect 101 -2329 135 -2323
rect 101 -2357 135 -2329
rect 101 -2397 135 -2395
rect 101 -2429 135 -2397
rect 101 -2499 135 -2467
rect 101 -2501 135 -2499
rect 101 -2567 135 -2539
rect 101 -2573 135 -2567
rect 101 -2635 135 -2611
rect 101 -2645 135 -2635
rect 101 -2703 135 -2683
rect 101 -2717 135 -2703
rect 101 -2771 135 -2755
rect 101 -2789 135 -2771
rect 101 -2839 135 -2827
rect 101 -2861 135 -2839
rect 101 -2907 135 -2899
rect 101 -2933 135 -2907
rect 101 -2975 135 -2971
rect 101 -3005 135 -2975
rect 101 -3077 135 -3043
rect 101 -3145 135 -3115
rect 101 -3149 135 -3145
rect 101 -3213 135 -3187
rect 101 -3221 135 -3213
rect 101 -3281 135 -3259
rect 101 -3293 135 -3281
rect 101 -3349 135 -3331
rect 101 -3365 135 -3349
rect 101 -3417 135 -3403
rect 101 -3437 135 -3417
rect 101 -3485 135 -3475
rect 101 -3509 135 -3485
rect 101 -3553 135 -3547
rect 101 -3581 135 -3553
rect 101 -3621 135 -3619
rect 101 -3653 135 -3621
rect 101 -3723 135 -3691
rect 101 -3725 135 -3723
rect 101 -3791 135 -3763
rect 101 -3797 135 -3791
rect 101 -3859 135 -3835
rect 101 -3869 135 -3859
rect 101 -3927 135 -3907
rect 101 -3941 135 -3927
rect 101 -3995 135 -3979
rect 101 -4013 135 -3995
rect 101 -4063 135 -4051
rect 101 -4085 135 -4063
rect 101 -4131 135 -4123
rect 101 -4157 135 -4131
rect 101 -4199 135 -4195
rect 101 -4229 135 -4199
rect 101 -4301 135 -4267
rect 101 -4369 135 -4339
rect 101 -4373 135 -4369
rect 101 -4437 135 -4411
rect 101 -4445 135 -4437
rect 101 -4505 135 -4483
rect 101 -4517 135 -4505
rect 101 -4573 135 -4555
rect 101 -4589 135 -4573
rect 101 -4641 135 -4627
rect 101 -4661 135 -4641
rect 101 -4709 135 -4699
rect 101 -4733 135 -4709
rect 101 -4777 135 -4771
rect 101 -4805 135 -4777
rect 101 -4845 135 -4843
rect 101 -4877 135 -4845
rect 101 -4947 135 -4915
rect 101 -4949 135 -4947
rect 101 -5015 135 -4987
rect 101 -5021 135 -5015
rect 101 -5083 135 -5059
rect 101 -5093 135 -5083
rect 101 -5151 135 -5131
rect 101 -5165 135 -5151
rect 101 -5219 135 -5203
rect 101 -5237 135 -5219
rect 101 -5287 135 -5275
rect 101 -5309 135 -5287
rect 101 -5355 135 -5347
rect 101 -5381 135 -5355
rect 101 -5423 135 -5419
rect 101 -5453 135 -5423
rect 101 -5525 135 -5491
rect 101 -5593 135 -5563
rect 101 -5597 135 -5593
rect 101 -5661 135 -5635
rect 101 -5669 135 -5661
rect 101 -5729 135 -5707
rect 101 -5741 135 -5729
rect 101 -5797 135 -5779
rect 101 -5813 135 -5797
rect 101 -5865 135 -5851
rect 101 -5885 135 -5865
rect 101 -5933 135 -5923
rect 101 -5957 135 -5933
rect 219 5933 253 5957
rect 219 5923 253 5933
rect 219 5865 253 5885
rect 219 5851 253 5865
rect 219 5797 253 5813
rect 219 5779 253 5797
rect 219 5729 253 5741
rect 219 5707 253 5729
rect 219 5661 253 5669
rect 219 5635 253 5661
rect 219 5593 253 5597
rect 219 5563 253 5593
rect 219 5491 253 5525
rect 219 5423 253 5453
rect 219 5419 253 5423
rect 219 5355 253 5381
rect 219 5347 253 5355
rect 219 5287 253 5309
rect 219 5275 253 5287
rect 219 5219 253 5237
rect 219 5203 253 5219
rect 219 5151 253 5165
rect 219 5131 253 5151
rect 219 5083 253 5093
rect 219 5059 253 5083
rect 219 5015 253 5021
rect 219 4987 253 5015
rect 219 4947 253 4949
rect 219 4915 253 4947
rect 219 4845 253 4877
rect 219 4843 253 4845
rect 219 4777 253 4805
rect 219 4771 253 4777
rect 219 4709 253 4733
rect 219 4699 253 4709
rect 219 4641 253 4661
rect 219 4627 253 4641
rect 219 4573 253 4589
rect 219 4555 253 4573
rect 219 4505 253 4517
rect 219 4483 253 4505
rect 219 4437 253 4445
rect 219 4411 253 4437
rect 219 4369 253 4373
rect 219 4339 253 4369
rect 219 4267 253 4301
rect 219 4199 253 4229
rect 219 4195 253 4199
rect 219 4131 253 4157
rect 219 4123 253 4131
rect 219 4063 253 4085
rect 219 4051 253 4063
rect 219 3995 253 4013
rect 219 3979 253 3995
rect 219 3927 253 3941
rect 219 3907 253 3927
rect 219 3859 253 3869
rect 219 3835 253 3859
rect 219 3791 253 3797
rect 219 3763 253 3791
rect 219 3723 253 3725
rect 219 3691 253 3723
rect 219 3621 253 3653
rect 219 3619 253 3621
rect 219 3553 253 3581
rect 219 3547 253 3553
rect 219 3485 253 3509
rect 219 3475 253 3485
rect 219 3417 253 3437
rect 219 3403 253 3417
rect 219 3349 253 3365
rect 219 3331 253 3349
rect 219 3281 253 3293
rect 219 3259 253 3281
rect 219 3213 253 3221
rect 219 3187 253 3213
rect 219 3145 253 3149
rect 219 3115 253 3145
rect 219 3043 253 3077
rect 219 2975 253 3005
rect 219 2971 253 2975
rect 219 2907 253 2933
rect 219 2899 253 2907
rect 219 2839 253 2861
rect 219 2827 253 2839
rect 219 2771 253 2789
rect 219 2755 253 2771
rect 219 2703 253 2717
rect 219 2683 253 2703
rect 219 2635 253 2645
rect 219 2611 253 2635
rect 219 2567 253 2573
rect 219 2539 253 2567
rect 219 2499 253 2501
rect 219 2467 253 2499
rect 219 2397 253 2429
rect 219 2395 253 2397
rect 219 2329 253 2357
rect 219 2323 253 2329
rect 219 2261 253 2285
rect 219 2251 253 2261
rect 219 2193 253 2213
rect 219 2179 253 2193
rect 219 2125 253 2141
rect 219 2107 253 2125
rect 219 2057 253 2069
rect 219 2035 253 2057
rect 219 1989 253 1997
rect 219 1963 253 1989
rect 219 1921 253 1925
rect 219 1891 253 1921
rect 219 1819 253 1853
rect 219 1751 253 1781
rect 219 1747 253 1751
rect 219 1683 253 1709
rect 219 1675 253 1683
rect 219 1615 253 1637
rect 219 1603 253 1615
rect 219 1547 253 1565
rect 219 1531 253 1547
rect 219 1479 253 1493
rect 219 1459 253 1479
rect 219 1411 253 1421
rect 219 1387 253 1411
rect 219 1343 253 1349
rect 219 1315 253 1343
rect 219 1275 253 1277
rect 219 1243 253 1275
rect 219 1173 253 1205
rect 219 1171 253 1173
rect 219 1105 253 1133
rect 219 1099 253 1105
rect 219 1037 253 1061
rect 219 1027 253 1037
rect 219 969 253 989
rect 219 955 253 969
rect 219 901 253 917
rect 219 883 253 901
rect 219 833 253 845
rect 219 811 253 833
rect 219 765 253 773
rect 219 739 253 765
rect 219 697 253 701
rect 219 667 253 697
rect 219 595 253 629
rect 219 527 253 557
rect 219 523 253 527
rect 219 459 253 485
rect 219 451 253 459
rect 219 391 253 413
rect 219 379 253 391
rect 219 323 253 341
rect 219 307 253 323
rect 219 255 253 269
rect 219 235 253 255
rect 219 187 253 197
rect 219 163 253 187
rect 219 119 253 125
rect 219 91 253 119
rect 219 51 253 53
rect 219 19 253 51
rect 219 -51 253 -19
rect 219 -53 253 -51
rect 219 -119 253 -91
rect 219 -125 253 -119
rect 219 -187 253 -163
rect 219 -197 253 -187
rect 219 -255 253 -235
rect 219 -269 253 -255
rect 219 -323 253 -307
rect 219 -341 253 -323
rect 219 -391 253 -379
rect 219 -413 253 -391
rect 219 -459 253 -451
rect 219 -485 253 -459
rect 219 -527 253 -523
rect 219 -557 253 -527
rect 219 -629 253 -595
rect 219 -697 253 -667
rect 219 -701 253 -697
rect 219 -765 253 -739
rect 219 -773 253 -765
rect 219 -833 253 -811
rect 219 -845 253 -833
rect 219 -901 253 -883
rect 219 -917 253 -901
rect 219 -969 253 -955
rect 219 -989 253 -969
rect 219 -1037 253 -1027
rect 219 -1061 253 -1037
rect 219 -1105 253 -1099
rect 219 -1133 253 -1105
rect 219 -1173 253 -1171
rect 219 -1205 253 -1173
rect 219 -1275 253 -1243
rect 219 -1277 253 -1275
rect 219 -1343 253 -1315
rect 219 -1349 253 -1343
rect 219 -1411 253 -1387
rect 219 -1421 253 -1411
rect 219 -1479 253 -1459
rect 219 -1493 253 -1479
rect 219 -1547 253 -1531
rect 219 -1565 253 -1547
rect 219 -1615 253 -1603
rect 219 -1637 253 -1615
rect 219 -1683 253 -1675
rect 219 -1709 253 -1683
rect 219 -1751 253 -1747
rect 219 -1781 253 -1751
rect 219 -1853 253 -1819
rect 219 -1921 253 -1891
rect 219 -1925 253 -1921
rect 219 -1989 253 -1963
rect 219 -1997 253 -1989
rect 219 -2057 253 -2035
rect 219 -2069 253 -2057
rect 219 -2125 253 -2107
rect 219 -2141 253 -2125
rect 219 -2193 253 -2179
rect 219 -2213 253 -2193
rect 219 -2261 253 -2251
rect 219 -2285 253 -2261
rect 219 -2329 253 -2323
rect 219 -2357 253 -2329
rect 219 -2397 253 -2395
rect 219 -2429 253 -2397
rect 219 -2499 253 -2467
rect 219 -2501 253 -2499
rect 219 -2567 253 -2539
rect 219 -2573 253 -2567
rect 219 -2635 253 -2611
rect 219 -2645 253 -2635
rect 219 -2703 253 -2683
rect 219 -2717 253 -2703
rect 219 -2771 253 -2755
rect 219 -2789 253 -2771
rect 219 -2839 253 -2827
rect 219 -2861 253 -2839
rect 219 -2907 253 -2899
rect 219 -2933 253 -2907
rect 219 -2975 253 -2971
rect 219 -3005 253 -2975
rect 219 -3077 253 -3043
rect 219 -3145 253 -3115
rect 219 -3149 253 -3145
rect 219 -3213 253 -3187
rect 219 -3221 253 -3213
rect 219 -3281 253 -3259
rect 219 -3293 253 -3281
rect 219 -3349 253 -3331
rect 219 -3365 253 -3349
rect 219 -3417 253 -3403
rect 219 -3437 253 -3417
rect 219 -3485 253 -3475
rect 219 -3509 253 -3485
rect 219 -3553 253 -3547
rect 219 -3581 253 -3553
rect 219 -3621 253 -3619
rect 219 -3653 253 -3621
rect 219 -3723 253 -3691
rect 219 -3725 253 -3723
rect 219 -3791 253 -3763
rect 219 -3797 253 -3791
rect 219 -3859 253 -3835
rect 219 -3869 253 -3859
rect 219 -3927 253 -3907
rect 219 -3941 253 -3927
rect 219 -3995 253 -3979
rect 219 -4013 253 -3995
rect 219 -4063 253 -4051
rect 219 -4085 253 -4063
rect 219 -4131 253 -4123
rect 219 -4157 253 -4131
rect 219 -4199 253 -4195
rect 219 -4229 253 -4199
rect 219 -4301 253 -4267
rect 219 -4369 253 -4339
rect 219 -4373 253 -4369
rect 219 -4437 253 -4411
rect 219 -4445 253 -4437
rect 219 -4505 253 -4483
rect 219 -4517 253 -4505
rect 219 -4573 253 -4555
rect 219 -4589 253 -4573
rect 219 -4641 253 -4627
rect 219 -4661 253 -4641
rect 219 -4709 253 -4699
rect 219 -4733 253 -4709
rect 219 -4777 253 -4771
rect 219 -4805 253 -4777
rect 219 -4845 253 -4843
rect 219 -4877 253 -4845
rect 219 -4947 253 -4915
rect 219 -4949 253 -4947
rect 219 -5015 253 -4987
rect 219 -5021 253 -5015
rect 219 -5083 253 -5059
rect 219 -5093 253 -5083
rect 219 -5151 253 -5131
rect 219 -5165 253 -5151
rect 219 -5219 253 -5203
rect 219 -5237 253 -5219
rect 219 -5287 253 -5275
rect 219 -5309 253 -5287
rect 219 -5355 253 -5347
rect 219 -5381 253 -5355
rect 219 -5423 253 -5419
rect 219 -5453 253 -5423
rect 219 -5525 253 -5491
rect 219 -5593 253 -5563
rect 219 -5597 253 -5593
rect 219 -5661 253 -5635
rect 219 -5669 253 -5661
rect 219 -5729 253 -5707
rect 219 -5741 253 -5729
rect 219 -5797 253 -5779
rect 219 -5813 253 -5797
rect 219 -5865 253 -5851
rect 219 -5885 253 -5865
rect 219 -5933 253 -5923
rect 219 -5957 253 -5933
rect 337 5933 371 5957
rect 337 5923 371 5933
rect 337 5865 371 5885
rect 337 5851 371 5865
rect 337 5797 371 5813
rect 337 5779 371 5797
rect 337 5729 371 5741
rect 337 5707 371 5729
rect 337 5661 371 5669
rect 337 5635 371 5661
rect 337 5593 371 5597
rect 337 5563 371 5593
rect 337 5491 371 5525
rect 337 5423 371 5453
rect 337 5419 371 5423
rect 337 5355 371 5381
rect 337 5347 371 5355
rect 337 5287 371 5309
rect 337 5275 371 5287
rect 337 5219 371 5237
rect 337 5203 371 5219
rect 337 5151 371 5165
rect 337 5131 371 5151
rect 337 5083 371 5093
rect 337 5059 371 5083
rect 337 5015 371 5021
rect 337 4987 371 5015
rect 337 4947 371 4949
rect 337 4915 371 4947
rect 337 4845 371 4877
rect 337 4843 371 4845
rect 337 4777 371 4805
rect 337 4771 371 4777
rect 337 4709 371 4733
rect 337 4699 371 4709
rect 337 4641 371 4661
rect 337 4627 371 4641
rect 337 4573 371 4589
rect 337 4555 371 4573
rect 337 4505 371 4517
rect 337 4483 371 4505
rect 337 4437 371 4445
rect 337 4411 371 4437
rect 337 4369 371 4373
rect 337 4339 371 4369
rect 337 4267 371 4301
rect 337 4199 371 4229
rect 337 4195 371 4199
rect 337 4131 371 4157
rect 337 4123 371 4131
rect 337 4063 371 4085
rect 337 4051 371 4063
rect 337 3995 371 4013
rect 337 3979 371 3995
rect 337 3927 371 3941
rect 337 3907 371 3927
rect 337 3859 371 3869
rect 337 3835 371 3859
rect 337 3791 371 3797
rect 337 3763 371 3791
rect 337 3723 371 3725
rect 337 3691 371 3723
rect 337 3621 371 3653
rect 337 3619 371 3621
rect 337 3553 371 3581
rect 337 3547 371 3553
rect 337 3485 371 3509
rect 337 3475 371 3485
rect 337 3417 371 3437
rect 337 3403 371 3417
rect 337 3349 371 3365
rect 337 3331 371 3349
rect 337 3281 371 3293
rect 337 3259 371 3281
rect 337 3213 371 3221
rect 337 3187 371 3213
rect 337 3145 371 3149
rect 337 3115 371 3145
rect 337 3043 371 3077
rect 337 2975 371 3005
rect 337 2971 371 2975
rect 337 2907 371 2933
rect 337 2899 371 2907
rect 337 2839 371 2861
rect 337 2827 371 2839
rect 337 2771 371 2789
rect 337 2755 371 2771
rect 337 2703 371 2717
rect 337 2683 371 2703
rect 337 2635 371 2645
rect 337 2611 371 2635
rect 337 2567 371 2573
rect 337 2539 371 2567
rect 337 2499 371 2501
rect 337 2467 371 2499
rect 337 2397 371 2429
rect 337 2395 371 2397
rect 337 2329 371 2357
rect 337 2323 371 2329
rect 337 2261 371 2285
rect 337 2251 371 2261
rect 337 2193 371 2213
rect 337 2179 371 2193
rect 337 2125 371 2141
rect 337 2107 371 2125
rect 337 2057 371 2069
rect 337 2035 371 2057
rect 337 1989 371 1997
rect 337 1963 371 1989
rect 337 1921 371 1925
rect 337 1891 371 1921
rect 337 1819 371 1853
rect 337 1751 371 1781
rect 337 1747 371 1751
rect 337 1683 371 1709
rect 337 1675 371 1683
rect 337 1615 371 1637
rect 337 1603 371 1615
rect 337 1547 371 1565
rect 337 1531 371 1547
rect 337 1479 371 1493
rect 337 1459 371 1479
rect 337 1411 371 1421
rect 337 1387 371 1411
rect 337 1343 371 1349
rect 337 1315 371 1343
rect 337 1275 371 1277
rect 337 1243 371 1275
rect 337 1173 371 1205
rect 337 1171 371 1173
rect 337 1105 371 1133
rect 337 1099 371 1105
rect 337 1037 371 1061
rect 337 1027 371 1037
rect 337 969 371 989
rect 337 955 371 969
rect 337 901 371 917
rect 337 883 371 901
rect 337 833 371 845
rect 337 811 371 833
rect 337 765 371 773
rect 337 739 371 765
rect 337 697 371 701
rect 337 667 371 697
rect 337 595 371 629
rect 337 527 371 557
rect 337 523 371 527
rect 337 459 371 485
rect 337 451 371 459
rect 337 391 371 413
rect 337 379 371 391
rect 337 323 371 341
rect 337 307 371 323
rect 337 255 371 269
rect 337 235 371 255
rect 337 187 371 197
rect 337 163 371 187
rect 337 119 371 125
rect 337 91 371 119
rect 337 51 371 53
rect 337 19 371 51
rect 337 -51 371 -19
rect 337 -53 371 -51
rect 337 -119 371 -91
rect 337 -125 371 -119
rect 337 -187 371 -163
rect 337 -197 371 -187
rect 337 -255 371 -235
rect 337 -269 371 -255
rect 337 -323 371 -307
rect 337 -341 371 -323
rect 337 -391 371 -379
rect 337 -413 371 -391
rect 337 -459 371 -451
rect 337 -485 371 -459
rect 337 -527 371 -523
rect 337 -557 371 -527
rect 337 -629 371 -595
rect 337 -697 371 -667
rect 337 -701 371 -697
rect 337 -765 371 -739
rect 337 -773 371 -765
rect 337 -833 371 -811
rect 337 -845 371 -833
rect 337 -901 371 -883
rect 337 -917 371 -901
rect 337 -969 371 -955
rect 337 -989 371 -969
rect 337 -1037 371 -1027
rect 337 -1061 371 -1037
rect 337 -1105 371 -1099
rect 337 -1133 371 -1105
rect 337 -1173 371 -1171
rect 337 -1205 371 -1173
rect 337 -1275 371 -1243
rect 337 -1277 371 -1275
rect 337 -1343 371 -1315
rect 337 -1349 371 -1343
rect 337 -1411 371 -1387
rect 337 -1421 371 -1411
rect 337 -1479 371 -1459
rect 337 -1493 371 -1479
rect 337 -1547 371 -1531
rect 337 -1565 371 -1547
rect 337 -1615 371 -1603
rect 337 -1637 371 -1615
rect 337 -1683 371 -1675
rect 337 -1709 371 -1683
rect 337 -1751 371 -1747
rect 337 -1781 371 -1751
rect 337 -1853 371 -1819
rect 337 -1921 371 -1891
rect 337 -1925 371 -1921
rect 337 -1989 371 -1963
rect 337 -1997 371 -1989
rect 337 -2057 371 -2035
rect 337 -2069 371 -2057
rect 337 -2125 371 -2107
rect 337 -2141 371 -2125
rect 337 -2193 371 -2179
rect 337 -2213 371 -2193
rect 337 -2261 371 -2251
rect 337 -2285 371 -2261
rect 337 -2329 371 -2323
rect 337 -2357 371 -2329
rect 337 -2397 371 -2395
rect 337 -2429 371 -2397
rect 337 -2499 371 -2467
rect 337 -2501 371 -2499
rect 337 -2567 371 -2539
rect 337 -2573 371 -2567
rect 337 -2635 371 -2611
rect 337 -2645 371 -2635
rect 337 -2703 371 -2683
rect 337 -2717 371 -2703
rect 337 -2771 371 -2755
rect 337 -2789 371 -2771
rect 337 -2839 371 -2827
rect 337 -2861 371 -2839
rect 337 -2907 371 -2899
rect 337 -2933 371 -2907
rect 337 -2975 371 -2971
rect 337 -3005 371 -2975
rect 337 -3077 371 -3043
rect 337 -3145 371 -3115
rect 337 -3149 371 -3145
rect 337 -3213 371 -3187
rect 337 -3221 371 -3213
rect 337 -3281 371 -3259
rect 337 -3293 371 -3281
rect 337 -3349 371 -3331
rect 337 -3365 371 -3349
rect 337 -3417 371 -3403
rect 337 -3437 371 -3417
rect 337 -3485 371 -3475
rect 337 -3509 371 -3485
rect 337 -3553 371 -3547
rect 337 -3581 371 -3553
rect 337 -3621 371 -3619
rect 337 -3653 371 -3621
rect 337 -3723 371 -3691
rect 337 -3725 371 -3723
rect 337 -3791 371 -3763
rect 337 -3797 371 -3791
rect 337 -3859 371 -3835
rect 337 -3869 371 -3859
rect 337 -3927 371 -3907
rect 337 -3941 371 -3927
rect 337 -3995 371 -3979
rect 337 -4013 371 -3995
rect 337 -4063 371 -4051
rect 337 -4085 371 -4063
rect 337 -4131 371 -4123
rect 337 -4157 371 -4131
rect 337 -4199 371 -4195
rect 337 -4229 371 -4199
rect 337 -4301 371 -4267
rect 337 -4369 371 -4339
rect 337 -4373 371 -4369
rect 337 -4437 371 -4411
rect 337 -4445 371 -4437
rect 337 -4505 371 -4483
rect 337 -4517 371 -4505
rect 337 -4573 371 -4555
rect 337 -4589 371 -4573
rect 337 -4641 371 -4627
rect 337 -4661 371 -4641
rect 337 -4709 371 -4699
rect 337 -4733 371 -4709
rect 337 -4777 371 -4771
rect 337 -4805 371 -4777
rect 337 -4845 371 -4843
rect 337 -4877 371 -4845
rect 337 -4947 371 -4915
rect 337 -4949 371 -4947
rect 337 -5015 371 -4987
rect 337 -5021 371 -5015
rect 337 -5083 371 -5059
rect 337 -5093 371 -5083
rect 337 -5151 371 -5131
rect 337 -5165 371 -5151
rect 337 -5219 371 -5203
rect 337 -5237 371 -5219
rect 337 -5287 371 -5275
rect 337 -5309 371 -5287
rect 337 -5355 371 -5347
rect 337 -5381 371 -5355
rect 337 -5423 371 -5419
rect 337 -5453 371 -5423
rect 337 -5525 371 -5491
rect 337 -5593 371 -5563
rect 337 -5597 371 -5593
rect 337 -5661 371 -5635
rect 337 -5669 371 -5661
rect 337 -5729 371 -5707
rect 337 -5741 371 -5729
rect 337 -5797 371 -5779
rect 337 -5813 371 -5797
rect 337 -5865 371 -5851
rect 337 -5885 371 -5865
rect 337 -5933 371 -5923
rect 337 -5957 371 -5933
rect 455 5933 489 5957
rect 455 5923 489 5933
rect 455 5865 489 5885
rect 455 5851 489 5865
rect 455 5797 489 5813
rect 455 5779 489 5797
rect 455 5729 489 5741
rect 455 5707 489 5729
rect 455 5661 489 5669
rect 455 5635 489 5661
rect 455 5593 489 5597
rect 455 5563 489 5593
rect 455 5491 489 5525
rect 455 5423 489 5453
rect 455 5419 489 5423
rect 455 5355 489 5381
rect 455 5347 489 5355
rect 455 5287 489 5309
rect 455 5275 489 5287
rect 455 5219 489 5237
rect 455 5203 489 5219
rect 455 5151 489 5165
rect 455 5131 489 5151
rect 455 5083 489 5093
rect 455 5059 489 5083
rect 455 5015 489 5021
rect 455 4987 489 5015
rect 455 4947 489 4949
rect 455 4915 489 4947
rect 455 4845 489 4877
rect 455 4843 489 4845
rect 455 4777 489 4805
rect 455 4771 489 4777
rect 455 4709 489 4733
rect 455 4699 489 4709
rect 455 4641 489 4661
rect 455 4627 489 4641
rect 455 4573 489 4589
rect 455 4555 489 4573
rect 455 4505 489 4517
rect 455 4483 489 4505
rect 455 4437 489 4445
rect 455 4411 489 4437
rect 455 4369 489 4373
rect 455 4339 489 4369
rect 455 4267 489 4301
rect 455 4199 489 4229
rect 455 4195 489 4199
rect 455 4131 489 4157
rect 455 4123 489 4131
rect 455 4063 489 4085
rect 455 4051 489 4063
rect 455 3995 489 4013
rect 455 3979 489 3995
rect 455 3927 489 3941
rect 455 3907 489 3927
rect 455 3859 489 3869
rect 455 3835 489 3859
rect 455 3791 489 3797
rect 455 3763 489 3791
rect 455 3723 489 3725
rect 455 3691 489 3723
rect 455 3621 489 3653
rect 455 3619 489 3621
rect 455 3553 489 3581
rect 455 3547 489 3553
rect 455 3485 489 3509
rect 455 3475 489 3485
rect 455 3417 489 3437
rect 455 3403 489 3417
rect 455 3349 489 3365
rect 455 3331 489 3349
rect 455 3281 489 3293
rect 455 3259 489 3281
rect 455 3213 489 3221
rect 455 3187 489 3213
rect 455 3145 489 3149
rect 455 3115 489 3145
rect 455 3043 489 3077
rect 455 2975 489 3005
rect 455 2971 489 2975
rect 455 2907 489 2933
rect 455 2899 489 2907
rect 455 2839 489 2861
rect 455 2827 489 2839
rect 455 2771 489 2789
rect 455 2755 489 2771
rect 455 2703 489 2717
rect 455 2683 489 2703
rect 455 2635 489 2645
rect 455 2611 489 2635
rect 455 2567 489 2573
rect 455 2539 489 2567
rect 455 2499 489 2501
rect 455 2467 489 2499
rect 455 2397 489 2429
rect 455 2395 489 2397
rect 455 2329 489 2357
rect 455 2323 489 2329
rect 455 2261 489 2285
rect 455 2251 489 2261
rect 455 2193 489 2213
rect 455 2179 489 2193
rect 455 2125 489 2141
rect 455 2107 489 2125
rect 455 2057 489 2069
rect 455 2035 489 2057
rect 455 1989 489 1997
rect 455 1963 489 1989
rect 455 1921 489 1925
rect 455 1891 489 1921
rect 455 1819 489 1853
rect 455 1751 489 1781
rect 455 1747 489 1751
rect 455 1683 489 1709
rect 455 1675 489 1683
rect 455 1615 489 1637
rect 455 1603 489 1615
rect 455 1547 489 1565
rect 455 1531 489 1547
rect 455 1479 489 1493
rect 455 1459 489 1479
rect 455 1411 489 1421
rect 455 1387 489 1411
rect 455 1343 489 1349
rect 455 1315 489 1343
rect 455 1275 489 1277
rect 455 1243 489 1275
rect 455 1173 489 1205
rect 455 1171 489 1173
rect 455 1105 489 1133
rect 455 1099 489 1105
rect 455 1037 489 1061
rect 455 1027 489 1037
rect 455 969 489 989
rect 455 955 489 969
rect 455 901 489 917
rect 455 883 489 901
rect 455 833 489 845
rect 455 811 489 833
rect 455 765 489 773
rect 455 739 489 765
rect 455 697 489 701
rect 455 667 489 697
rect 455 595 489 629
rect 455 527 489 557
rect 455 523 489 527
rect 455 459 489 485
rect 455 451 489 459
rect 455 391 489 413
rect 455 379 489 391
rect 455 323 489 341
rect 455 307 489 323
rect 455 255 489 269
rect 455 235 489 255
rect 455 187 489 197
rect 455 163 489 187
rect 455 119 489 125
rect 455 91 489 119
rect 455 51 489 53
rect 455 19 489 51
rect 455 -51 489 -19
rect 455 -53 489 -51
rect 455 -119 489 -91
rect 455 -125 489 -119
rect 455 -187 489 -163
rect 455 -197 489 -187
rect 455 -255 489 -235
rect 455 -269 489 -255
rect 455 -323 489 -307
rect 455 -341 489 -323
rect 455 -391 489 -379
rect 455 -413 489 -391
rect 455 -459 489 -451
rect 455 -485 489 -459
rect 455 -527 489 -523
rect 455 -557 489 -527
rect 455 -629 489 -595
rect 455 -697 489 -667
rect 455 -701 489 -697
rect 455 -765 489 -739
rect 455 -773 489 -765
rect 455 -833 489 -811
rect 455 -845 489 -833
rect 455 -901 489 -883
rect 455 -917 489 -901
rect 455 -969 489 -955
rect 455 -989 489 -969
rect 455 -1037 489 -1027
rect 455 -1061 489 -1037
rect 455 -1105 489 -1099
rect 455 -1133 489 -1105
rect 455 -1173 489 -1171
rect 455 -1205 489 -1173
rect 455 -1275 489 -1243
rect 455 -1277 489 -1275
rect 455 -1343 489 -1315
rect 455 -1349 489 -1343
rect 455 -1411 489 -1387
rect 455 -1421 489 -1411
rect 455 -1479 489 -1459
rect 455 -1493 489 -1479
rect 455 -1547 489 -1531
rect 455 -1565 489 -1547
rect 455 -1615 489 -1603
rect 455 -1637 489 -1615
rect 455 -1683 489 -1675
rect 455 -1709 489 -1683
rect 455 -1751 489 -1747
rect 455 -1781 489 -1751
rect 455 -1853 489 -1819
rect 455 -1921 489 -1891
rect 455 -1925 489 -1921
rect 455 -1989 489 -1963
rect 455 -1997 489 -1989
rect 455 -2057 489 -2035
rect 455 -2069 489 -2057
rect 455 -2125 489 -2107
rect 455 -2141 489 -2125
rect 455 -2193 489 -2179
rect 455 -2213 489 -2193
rect 455 -2261 489 -2251
rect 455 -2285 489 -2261
rect 455 -2329 489 -2323
rect 455 -2357 489 -2329
rect 455 -2397 489 -2395
rect 455 -2429 489 -2397
rect 455 -2499 489 -2467
rect 455 -2501 489 -2499
rect 455 -2567 489 -2539
rect 455 -2573 489 -2567
rect 455 -2635 489 -2611
rect 455 -2645 489 -2635
rect 455 -2703 489 -2683
rect 455 -2717 489 -2703
rect 455 -2771 489 -2755
rect 455 -2789 489 -2771
rect 455 -2839 489 -2827
rect 455 -2861 489 -2839
rect 455 -2907 489 -2899
rect 455 -2933 489 -2907
rect 455 -2975 489 -2971
rect 455 -3005 489 -2975
rect 455 -3077 489 -3043
rect 455 -3145 489 -3115
rect 455 -3149 489 -3145
rect 455 -3213 489 -3187
rect 455 -3221 489 -3213
rect 455 -3281 489 -3259
rect 455 -3293 489 -3281
rect 455 -3349 489 -3331
rect 455 -3365 489 -3349
rect 455 -3417 489 -3403
rect 455 -3437 489 -3417
rect 455 -3485 489 -3475
rect 455 -3509 489 -3485
rect 455 -3553 489 -3547
rect 455 -3581 489 -3553
rect 455 -3621 489 -3619
rect 455 -3653 489 -3621
rect 455 -3723 489 -3691
rect 455 -3725 489 -3723
rect 455 -3791 489 -3763
rect 455 -3797 489 -3791
rect 455 -3859 489 -3835
rect 455 -3869 489 -3859
rect 455 -3927 489 -3907
rect 455 -3941 489 -3927
rect 455 -3995 489 -3979
rect 455 -4013 489 -3995
rect 455 -4063 489 -4051
rect 455 -4085 489 -4063
rect 455 -4131 489 -4123
rect 455 -4157 489 -4131
rect 455 -4199 489 -4195
rect 455 -4229 489 -4199
rect 455 -4301 489 -4267
rect 455 -4369 489 -4339
rect 455 -4373 489 -4369
rect 455 -4437 489 -4411
rect 455 -4445 489 -4437
rect 455 -4505 489 -4483
rect 455 -4517 489 -4505
rect 455 -4573 489 -4555
rect 455 -4589 489 -4573
rect 455 -4641 489 -4627
rect 455 -4661 489 -4641
rect 455 -4709 489 -4699
rect 455 -4733 489 -4709
rect 455 -4777 489 -4771
rect 455 -4805 489 -4777
rect 455 -4845 489 -4843
rect 455 -4877 489 -4845
rect 455 -4947 489 -4915
rect 455 -4949 489 -4947
rect 455 -5015 489 -4987
rect 455 -5021 489 -5015
rect 455 -5083 489 -5059
rect 455 -5093 489 -5083
rect 455 -5151 489 -5131
rect 455 -5165 489 -5151
rect 455 -5219 489 -5203
rect 455 -5237 489 -5219
rect 455 -5287 489 -5275
rect 455 -5309 489 -5287
rect 455 -5355 489 -5347
rect 455 -5381 489 -5355
rect 455 -5423 489 -5419
rect 455 -5453 489 -5423
rect 455 -5525 489 -5491
rect 455 -5593 489 -5563
rect 455 -5597 489 -5593
rect 455 -5661 489 -5635
rect 455 -5669 489 -5661
rect 455 -5729 489 -5707
rect 455 -5741 489 -5729
rect 455 -5797 489 -5779
rect 455 -5813 489 -5797
rect 455 -5865 489 -5851
rect 455 -5885 489 -5865
rect 455 -5933 489 -5923
rect 455 -5957 489 -5933
rect 573 5933 607 5957
rect 573 5923 607 5933
rect 573 5865 607 5885
rect 573 5851 607 5865
rect 573 5797 607 5813
rect 573 5779 607 5797
rect 573 5729 607 5741
rect 573 5707 607 5729
rect 573 5661 607 5669
rect 573 5635 607 5661
rect 573 5593 607 5597
rect 573 5563 607 5593
rect 573 5491 607 5525
rect 573 5423 607 5453
rect 573 5419 607 5423
rect 573 5355 607 5381
rect 573 5347 607 5355
rect 573 5287 607 5309
rect 573 5275 607 5287
rect 573 5219 607 5237
rect 573 5203 607 5219
rect 573 5151 607 5165
rect 573 5131 607 5151
rect 573 5083 607 5093
rect 573 5059 607 5083
rect 573 5015 607 5021
rect 573 4987 607 5015
rect 573 4947 607 4949
rect 573 4915 607 4947
rect 573 4845 607 4877
rect 573 4843 607 4845
rect 573 4777 607 4805
rect 573 4771 607 4777
rect 573 4709 607 4733
rect 573 4699 607 4709
rect 573 4641 607 4661
rect 573 4627 607 4641
rect 573 4573 607 4589
rect 573 4555 607 4573
rect 573 4505 607 4517
rect 573 4483 607 4505
rect 573 4437 607 4445
rect 573 4411 607 4437
rect 573 4369 607 4373
rect 573 4339 607 4369
rect 573 4267 607 4301
rect 573 4199 607 4229
rect 573 4195 607 4199
rect 573 4131 607 4157
rect 573 4123 607 4131
rect 573 4063 607 4085
rect 573 4051 607 4063
rect 573 3995 607 4013
rect 573 3979 607 3995
rect 573 3927 607 3941
rect 573 3907 607 3927
rect 573 3859 607 3869
rect 573 3835 607 3859
rect 573 3791 607 3797
rect 573 3763 607 3791
rect 573 3723 607 3725
rect 573 3691 607 3723
rect 573 3621 607 3653
rect 573 3619 607 3621
rect 573 3553 607 3581
rect 573 3547 607 3553
rect 573 3485 607 3509
rect 573 3475 607 3485
rect 573 3417 607 3437
rect 573 3403 607 3417
rect 573 3349 607 3365
rect 573 3331 607 3349
rect 573 3281 607 3293
rect 573 3259 607 3281
rect 573 3213 607 3221
rect 573 3187 607 3213
rect 573 3145 607 3149
rect 573 3115 607 3145
rect 573 3043 607 3077
rect 573 2975 607 3005
rect 573 2971 607 2975
rect 573 2907 607 2933
rect 573 2899 607 2907
rect 573 2839 607 2861
rect 573 2827 607 2839
rect 573 2771 607 2789
rect 573 2755 607 2771
rect 573 2703 607 2717
rect 573 2683 607 2703
rect 573 2635 607 2645
rect 573 2611 607 2635
rect 573 2567 607 2573
rect 573 2539 607 2567
rect 573 2499 607 2501
rect 573 2467 607 2499
rect 573 2397 607 2429
rect 573 2395 607 2397
rect 573 2329 607 2357
rect 573 2323 607 2329
rect 573 2261 607 2285
rect 573 2251 607 2261
rect 573 2193 607 2213
rect 573 2179 607 2193
rect 573 2125 607 2141
rect 573 2107 607 2125
rect 573 2057 607 2069
rect 573 2035 607 2057
rect 573 1989 607 1997
rect 573 1963 607 1989
rect 573 1921 607 1925
rect 573 1891 607 1921
rect 573 1819 607 1853
rect 573 1751 607 1781
rect 573 1747 607 1751
rect 573 1683 607 1709
rect 573 1675 607 1683
rect 573 1615 607 1637
rect 573 1603 607 1615
rect 573 1547 607 1565
rect 573 1531 607 1547
rect 573 1479 607 1493
rect 573 1459 607 1479
rect 573 1411 607 1421
rect 573 1387 607 1411
rect 573 1343 607 1349
rect 573 1315 607 1343
rect 573 1275 607 1277
rect 573 1243 607 1275
rect 573 1173 607 1205
rect 573 1171 607 1173
rect 573 1105 607 1133
rect 573 1099 607 1105
rect 573 1037 607 1061
rect 573 1027 607 1037
rect 573 969 607 989
rect 573 955 607 969
rect 573 901 607 917
rect 573 883 607 901
rect 573 833 607 845
rect 573 811 607 833
rect 573 765 607 773
rect 573 739 607 765
rect 573 697 607 701
rect 573 667 607 697
rect 573 595 607 629
rect 573 527 607 557
rect 573 523 607 527
rect 573 459 607 485
rect 573 451 607 459
rect 573 391 607 413
rect 573 379 607 391
rect 573 323 607 341
rect 573 307 607 323
rect 573 255 607 269
rect 573 235 607 255
rect 573 187 607 197
rect 573 163 607 187
rect 573 119 607 125
rect 573 91 607 119
rect 573 51 607 53
rect 573 19 607 51
rect 573 -51 607 -19
rect 573 -53 607 -51
rect 573 -119 607 -91
rect 573 -125 607 -119
rect 573 -187 607 -163
rect 573 -197 607 -187
rect 573 -255 607 -235
rect 573 -269 607 -255
rect 573 -323 607 -307
rect 573 -341 607 -323
rect 573 -391 607 -379
rect 573 -413 607 -391
rect 573 -459 607 -451
rect 573 -485 607 -459
rect 573 -527 607 -523
rect 573 -557 607 -527
rect 573 -629 607 -595
rect 573 -697 607 -667
rect 573 -701 607 -697
rect 573 -765 607 -739
rect 573 -773 607 -765
rect 573 -833 607 -811
rect 573 -845 607 -833
rect 573 -901 607 -883
rect 573 -917 607 -901
rect 573 -969 607 -955
rect 573 -989 607 -969
rect 573 -1037 607 -1027
rect 573 -1061 607 -1037
rect 573 -1105 607 -1099
rect 573 -1133 607 -1105
rect 573 -1173 607 -1171
rect 573 -1205 607 -1173
rect 573 -1275 607 -1243
rect 573 -1277 607 -1275
rect 573 -1343 607 -1315
rect 573 -1349 607 -1343
rect 573 -1411 607 -1387
rect 573 -1421 607 -1411
rect 573 -1479 607 -1459
rect 573 -1493 607 -1479
rect 573 -1547 607 -1531
rect 573 -1565 607 -1547
rect 573 -1615 607 -1603
rect 573 -1637 607 -1615
rect 573 -1683 607 -1675
rect 573 -1709 607 -1683
rect 573 -1751 607 -1747
rect 573 -1781 607 -1751
rect 573 -1853 607 -1819
rect 573 -1921 607 -1891
rect 573 -1925 607 -1921
rect 573 -1989 607 -1963
rect 573 -1997 607 -1989
rect 573 -2057 607 -2035
rect 573 -2069 607 -2057
rect 573 -2125 607 -2107
rect 573 -2141 607 -2125
rect 573 -2193 607 -2179
rect 573 -2213 607 -2193
rect 573 -2261 607 -2251
rect 573 -2285 607 -2261
rect 573 -2329 607 -2323
rect 573 -2357 607 -2329
rect 573 -2397 607 -2395
rect 573 -2429 607 -2397
rect 573 -2499 607 -2467
rect 573 -2501 607 -2499
rect 573 -2567 607 -2539
rect 573 -2573 607 -2567
rect 573 -2635 607 -2611
rect 573 -2645 607 -2635
rect 573 -2703 607 -2683
rect 573 -2717 607 -2703
rect 573 -2771 607 -2755
rect 573 -2789 607 -2771
rect 573 -2839 607 -2827
rect 573 -2861 607 -2839
rect 573 -2907 607 -2899
rect 573 -2933 607 -2907
rect 573 -2975 607 -2971
rect 573 -3005 607 -2975
rect 573 -3077 607 -3043
rect 573 -3145 607 -3115
rect 573 -3149 607 -3145
rect 573 -3213 607 -3187
rect 573 -3221 607 -3213
rect 573 -3281 607 -3259
rect 573 -3293 607 -3281
rect 573 -3349 607 -3331
rect 573 -3365 607 -3349
rect 573 -3417 607 -3403
rect 573 -3437 607 -3417
rect 573 -3485 607 -3475
rect 573 -3509 607 -3485
rect 573 -3553 607 -3547
rect 573 -3581 607 -3553
rect 573 -3621 607 -3619
rect 573 -3653 607 -3621
rect 573 -3723 607 -3691
rect 573 -3725 607 -3723
rect 573 -3791 607 -3763
rect 573 -3797 607 -3791
rect 573 -3859 607 -3835
rect 573 -3869 607 -3859
rect 573 -3927 607 -3907
rect 573 -3941 607 -3927
rect 573 -3995 607 -3979
rect 573 -4013 607 -3995
rect 573 -4063 607 -4051
rect 573 -4085 607 -4063
rect 573 -4131 607 -4123
rect 573 -4157 607 -4131
rect 573 -4199 607 -4195
rect 573 -4229 607 -4199
rect 573 -4301 607 -4267
rect 573 -4369 607 -4339
rect 573 -4373 607 -4369
rect 573 -4437 607 -4411
rect 573 -4445 607 -4437
rect 573 -4505 607 -4483
rect 573 -4517 607 -4505
rect 573 -4573 607 -4555
rect 573 -4589 607 -4573
rect 573 -4641 607 -4627
rect 573 -4661 607 -4641
rect 573 -4709 607 -4699
rect 573 -4733 607 -4709
rect 573 -4777 607 -4771
rect 573 -4805 607 -4777
rect 573 -4845 607 -4843
rect 573 -4877 607 -4845
rect 573 -4947 607 -4915
rect 573 -4949 607 -4947
rect 573 -5015 607 -4987
rect 573 -5021 607 -5015
rect 573 -5083 607 -5059
rect 573 -5093 607 -5083
rect 573 -5151 607 -5131
rect 573 -5165 607 -5151
rect 573 -5219 607 -5203
rect 573 -5237 607 -5219
rect 573 -5287 607 -5275
rect 573 -5309 607 -5287
rect 573 -5355 607 -5347
rect 573 -5381 607 -5355
rect 573 -5423 607 -5419
rect 573 -5453 607 -5423
rect 573 -5525 607 -5491
rect 573 -5593 607 -5563
rect 573 -5597 607 -5593
rect 573 -5661 607 -5635
rect 573 -5669 607 -5661
rect 573 -5729 607 -5707
rect 573 -5741 607 -5729
rect 573 -5797 607 -5779
rect 573 -5813 607 -5797
rect 573 -5865 607 -5851
rect 573 -5885 607 -5865
rect 573 -5933 607 -5923
rect 573 -5957 607 -5933
<< metal1 >>
rect -560 6072 -502 6078
rect -560 6038 -548 6072
rect -514 6038 -502 6072
rect -560 6032 -502 6038
rect -613 5957 -567 6000
rect -613 5923 -607 5957
rect -573 5923 -567 5957
rect -613 5885 -567 5923
rect -613 5851 -607 5885
rect -573 5851 -567 5885
rect -613 5813 -567 5851
rect -613 5779 -607 5813
rect -573 5779 -567 5813
rect -613 5741 -567 5779
rect -613 5707 -607 5741
rect -573 5707 -567 5741
rect -613 5669 -567 5707
rect -613 5635 -607 5669
rect -573 5635 -567 5669
rect -613 5597 -567 5635
rect -613 5563 -607 5597
rect -573 5563 -567 5597
rect -613 5525 -567 5563
rect -613 5491 -607 5525
rect -573 5491 -567 5525
rect -613 5453 -567 5491
rect -613 5419 -607 5453
rect -573 5419 -567 5453
rect -613 5381 -567 5419
rect -613 5347 -607 5381
rect -573 5347 -567 5381
rect -613 5309 -567 5347
rect -613 5275 -607 5309
rect -573 5275 -567 5309
rect -613 5237 -567 5275
rect -613 5203 -607 5237
rect -573 5203 -567 5237
rect -613 5165 -567 5203
rect -613 5131 -607 5165
rect -573 5131 -567 5165
rect -613 5093 -567 5131
rect -613 5059 -607 5093
rect -573 5059 -567 5093
rect -613 5021 -567 5059
rect -613 4987 -607 5021
rect -573 4987 -567 5021
rect -613 4949 -567 4987
rect -613 4915 -607 4949
rect -573 4915 -567 4949
rect -613 4877 -567 4915
rect -613 4843 -607 4877
rect -573 4843 -567 4877
rect -613 4805 -567 4843
rect -613 4771 -607 4805
rect -573 4771 -567 4805
rect -613 4733 -567 4771
rect -613 4699 -607 4733
rect -573 4699 -567 4733
rect -613 4661 -567 4699
rect -613 4627 -607 4661
rect -573 4627 -567 4661
rect -613 4589 -567 4627
rect -613 4555 -607 4589
rect -573 4555 -567 4589
rect -613 4517 -567 4555
rect -613 4483 -607 4517
rect -573 4483 -567 4517
rect -613 4445 -567 4483
rect -613 4411 -607 4445
rect -573 4411 -567 4445
rect -613 4373 -567 4411
rect -613 4339 -607 4373
rect -573 4339 -567 4373
rect -613 4301 -567 4339
rect -613 4267 -607 4301
rect -573 4267 -567 4301
rect -613 4229 -567 4267
rect -613 4195 -607 4229
rect -573 4195 -567 4229
rect -613 4157 -567 4195
rect -613 4123 -607 4157
rect -573 4123 -567 4157
rect -613 4085 -567 4123
rect -613 4051 -607 4085
rect -573 4051 -567 4085
rect -613 4013 -567 4051
rect -613 3979 -607 4013
rect -573 3979 -567 4013
rect -613 3941 -567 3979
rect -613 3907 -607 3941
rect -573 3907 -567 3941
rect -613 3869 -567 3907
rect -613 3835 -607 3869
rect -573 3835 -567 3869
rect -613 3797 -567 3835
rect -613 3763 -607 3797
rect -573 3763 -567 3797
rect -613 3725 -567 3763
rect -613 3691 -607 3725
rect -573 3691 -567 3725
rect -613 3653 -567 3691
rect -613 3619 -607 3653
rect -573 3619 -567 3653
rect -613 3581 -567 3619
rect -613 3547 -607 3581
rect -573 3547 -567 3581
rect -613 3509 -567 3547
rect -613 3475 -607 3509
rect -573 3475 -567 3509
rect -613 3437 -567 3475
rect -613 3403 -607 3437
rect -573 3403 -567 3437
rect -613 3365 -567 3403
rect -613 3331 -607 3365
rect -573 3331 -567 3365
rect -613 3293 -567 3331
rect -613 3259 -607 3293
rect -573 3259 -567 3293
rect -613 3221 -567 3259
rect -613 3187 -607 3221
rect -573 3187 -567 3221
rect -613 3149 -567 3187
rect -613 3115 -607 3149
rect -573 3115 -567 3149
rect -613 3077 -567 3115
rect -613 3043 -607 3077
rect -573 3043 -567 3077
rect -613 3005 -567 3043
rect -613 2971 -607 3005
rect -573 2971 -567 3005
rect -613 2933 -567 2971
rect -613 2899 -607 2933
rect -573 2899 -567 2933
rect -613 2861 -567 2899
rect -613 2827 -607 2861
rect -573 2827 -567 2861
rect -613 2789 -567 2827
rect -613 2755 -607 2789
rect -573 2755 -567 2789
rect -613 2717 -567 2755
rect -613 2683 -607 2717
rect -573 2683 -567 2717
rect -613 2645 -567 2683
rect -613 2611 -607 2645
rect -573 2611 -567 2645
rect -613 2573 -567 2611
rect -613 2539 -607 2573
rect -573 2539 -567 2573
rect -613 2501 -567 2539
rect -613 2467 -607 2501
rect -573 2467 -567 2501
rect -613 2429 -567 2467
rect -613 2395 -607 2429
rect -573 2395 -567 2429
rect -613 2357 -567 2395
rect -613 2323 -607 2357
rect -573 2323 -567 2357
rect -613 2285 -567 2323
rect -613 2251 -607 2285
rect -573 2251 -567 2285
rect -613 2213 -567 2251
rect -613 2179 -607 2213
rect -573 2179 -567 2213
rect -613 2141 -567 2179
rect -613 2107 -607 2141
rect -573 2107 -567 2141
rect -613 2069 -567 2107
rect -613 2035 -607 2069
rect -573 2035 -567 2069
rect -613 1997 -567 2035
rect -613 1963 -607 1997
rect -573 1963 -567 1997
rect -613 1925 -567 1963
rect -613 1891 -607 1925
rect -573 1891 -567 1925
rect -613 1853 -567 1891
rect -613 1819 -607 1853
rect -573 1819 -567 1853
rect -613 1781 -567 1819
rect -613 1747 -607 1781
rect -573 1747 -567 1781
rect -613 1709 -567 1747
rect -613 1675 -607 1709
rect -573 1675 -567 1709
rect -613 1637 -567 1675
rect -613 1603 -607 1637
rect -573 1603 -567 1637
rect -613 1565 -567 1603
rect -613 1531 -607 1565
rect -573 1531 -567 1565
rect -613 1493 -567 1531
rect -613 1459 -607 1493
rect -573 1459 -567 1493
rect -613 1421 -567 1459
rect -613 1387 -607 1421
rect -573 1387 -567 1421
rect -613 1349 -567 1387
rect -613 1315 -607 1349
rect -573 1315 -567 1349
rect -613 1277 -567 1315
rect -613 1243 -607 1277
rect -573 1243 -567 1277
rect -613 1205 -567 1243
rect -613 1171 -607 1205
rect -573 1171 -567 1205
rect -613 1133 -567 1171
rect -613 1099 -607 1133
rect -573 1099 -567 1133
rect -613 1061 -567 1099
rect -613 1027 -607 1061
rect -573 1027 -567 1061
rect -613 989 -567 1027
rect -613 955 -607 989
rect -573 955 -567 989
rect -613 917 -567 955
rect -613 883 -607 917
rect -573 883 -567 917
rect -613 845 -567 883
rect -613 811 -607 845
rect -573 811 -567 845
rect -613 773 -567 811
rect -613 739 -607 773
rect -573 739 -567 773
rect -613 701 -567 739
rect -613 667 -607 701
rect -573 667 -567 701
rect -613 629 -567 667
rect -613 595 -607 629
rect -573 595 -567 629
rect -613 557 -567 595
rect -613 523 -607 557
rect -573 523 -567 557
rect -613 485 -567 523
rect -613 451 -607 485
rect -573 451 -567 485
rect -613 413 -567 451
rect -613 379 -607 413
rect -573 379 -567 413
rect -613 341 -567 379
rect -613 307 -607 341
rect -573 307 -567 341
rect -613 269 -567 307
rect -613 235 -607 269
rect -573 235 -567 269
rect -613 197 -567 235
rect -613 163 -607 197
rect -573 163 -567 197
rect -613 125 -567 163
rect -613 91 -607 125
rect -573 91 -567 125
rect -613 53 -567 91
rect -613 19 -607 53
rect -573 19 -567 53
rect -613 -19 -567 19
rect -613 -53 -607 -19
rect -573 -53 -567 -19
rect -613 -91 -567 -53
rect -613 -125 -607 -91
rect -573 -125 -567 -91
rect -613 -163 -567 -125
rect -613 -197 -607 -163
rect -573 -197 -567 -163
rect -613 -235 -567 -197
rect -613 -269 -607 -235
rect -573 -269 -567 -235
rect -613 -307 -567 -269
rect -613 -341 -607 -307
rect -573 -341 -567 -307
rect -613 -379 -567 -341
rect -613 -413 -607 -379
rect -573 -413 -567 -379
rect -613 -451 -567 -413
rect -613 -485 -607 -451
rect -573 -485 -567 -451
rect -613 -523 -567 -485
rect -613 -557 -607 -523
rect -573 -557 -567 -523
rect -613 -595 -567 -557
rect -613 -629 -607 -595
rect -573 -629 -567 -595
rect -613 -667 -567 -629
rect -613 -701 -607 -667
rect -573 -701 -567 -667
rect -613 -739 -567 -701
rect -613 -773 -607 -739
rect -573 -773 -567 -739
rect -613 -811 -567 -773
rect -613 -845 -607 -811
rect -573 -845 -567 -811
rect -613 -883 -567 -845
rect -613 -917 -607 -883
rect -573 -917 -567 -883
rect -613 -955 -567 -917
rect -613 -989 -607 -955
rect -573 -989 -567 -955
rect -613 -1027 -567 -989
rect -613 -1061 -607 -1027
rect -573 -1061 -567 -1027
rect -613 -1099 -567 -1061
rect -613 -1133 -607 -1099
rect -573 -1133 -567 -1099
rect -613 -1171 -567 -1133
rect -613 -1205 -607 -1171
rect -573 -1205 -567 -1171
rect -613 -1243 -567 -1205
rect -613 -1277 -607 -1243
rect -573 -1277 -567 -1243
rect -613 -1315 -567 -1277
rect -613 -1349 -607 -1315
rect -573 -1349 -567 -1315
rect -613 -1387 -567 -1349
rect -613 -1421 -607 -1387
rect -573 -1421 -567 -1387
rect -613 -1459 -567 -1421
rect -613 -1493 -607 -1459
rect -573 -1493 -567 -1459
rect -613 -1531 -567 -1493
rect -613 -1565 -607 -1531
rect -573 -1565 -567 -1531
rect -613 -1603 -567 -1565
rect -613 -1637 -607 -1603
rect -573 -1637 -567 -1603
rect -613 -1675 -567 -1637
rect -613 -1709 -607 -1675
rect -573 -1709 -567 -1675
rect -613 -1747 -567 -1709
rect -613 -1781 -607 -1747
rect -573 -1781 -567 -1747
rect -613 -1819 -567 -1781
rect -613 -1853 -607 -1819
rect -573 -1853 -567 -1819
rect -613 -1891 -567 -1853
rect -613 -1925 -607 -1891
rect -573 -1925 -567 -1891
rect -613 -1963 -567 -1925
rect -613 -1997 -607 -1963
rect -573 -1997 -567 -1963
rect -613 -2035 -567 -1997
rect -613 -2069 -607 -2035
rect -573 -2069 -567 -2035
rect -613 -2107 -567 -2069
rect -613 -2141 -607 -2107
rect -573 -2141 -567 -2107
rect -613 -2179 -567 -2141
rect -613 -2213 -607 -2179
rect -573 -2213 -567 -2179
rect -613 -2251 -567 -2213
rect -613 -2285 -607 -2251
rect -573 -2285 -567 -2251
rect -613 -2323 -567 -2285
rect -613 -2357 -607 -2323
rect -573 -2357 -567 -2323
rect -613 -2395 -567 -2357
rect -613 -2429 -607 -2395
rect -573 -2429 -567 -2395
rect -613 -2467 -567 -2429
rect -613 -2501 -607 -2467
rect -573 -2501 -567 -2467
rect -613 -2539 -567 -2501
rect -613 -2573 -607 -2539
rect -573 -2573 -567 -2539
rect -613 -2611 -567 -2573
rect -613 -2645 -607 -2611
rect -573 -2645 -567 -2611
rect -613 -2683 -567 -2645
rect -613 -2717 -607 -2683
rect -573 -2717 -567 -2683
rect -613 -2755 -567 -2717
rect -613 -2789 -607 -2755
rect -573 -2789 -567 -2755
rect -613 -2827 -567 -2789
rect -613 -2861 -607 -2827
rect -573 -2861 -567 -2827
rect -613 -2899 -567 -2861
rect -613 -2933 -607 -2899
rect -573 -2933 -567 -2899
rect -613 -2971 -567 -2933
rect -613 -3005 -607 -2971
rect -573 -3005 -567 -2971
rect -613 -3043 -567 -3005
rect -613 -3077 -607 -3043
rect -573 -3077 -567 -3043
rect -613 -3115 -567 -3077
rect -613 -3149 -607 -3115
rect -573 -3149 -567 -3115
rect -613 -3187 -567 -3149
rect -613 -3221 -607 -3187
rect -573 -3221 -567 -3187
rect -613 -3259 -567 -3221
rect -613 -3293 -607 -3259
rect -573 -3293 -567 -3259
rect -613 -3331 -567 -3293
rect -613 -3365 -607 -3331
rect -573 -3365 -567 -3331
rect -613 -3403 -567 -3365
rect -613 -3437 -607 -3403
rect -573 -3437 -567 -3403
rect -613 -3475 -567 -3437
rect -613 -3509 -607 -3475
rect -573 -3509 -567 -3475
rect -613 -3547 -567 -3509
rect -613 -3581 -607 -3547
rect -573 -3581 -567 -3547
rect -613 -3619 -567 -3581
rect -613 -3653 -607 -3619
rect -573 -3653 -567 -3619
rect -613 -3691 -567 -3653
rect -613 -3725 -607 -3691
rect -573 -3725 -567 -3691
rect -613 -3763 -567 -3725
rect -613 -3797 -607 -3763
rect -573 -3797 -567 -3763
rect -613 -3835 -567 -3797
rect -613 -3869 -607 -3835
rect -573 -3869 -567 -3835
rect -613 -3907 -567 -3869
rect -613 -3941 -607 -3907
rect -573 -3941 -567 -3907
rect -613 -3979 -567 -3941
rect -613 -4013 -607 -3979
rect -573 -4013 -567 -3979
rect -613 -4051 -567 -4013
rect -613 -4085 -607 -4051
rect -573 -4085 -567 -4051
rect -613 -4123 -567 -4085
rect -613 -4157 -607 -4123
rect -573 -4157 -567 -4123
rect -613 -4195 -567 -4157
rect -613 -4229 -607 -4195
rect -573 -4229 -567 -4195
rect -613 -4267 -567 -4229
rect -613 -4301 -607 -4267
rect -573 -4301 -567 -4267
rect -613 -4339 -567 -4301
rect -613 -4373 -607 -4339
rect -573 -4373 -567 -4339
rect -613 -4411 -567 -4373
rect -613 -4445 -607 -4411
rect -573 -4445 -567 -4411
rect -613 -4483 -567 -4445
rect -613 -4517 -607 -4483
rect -573 -4517 -567 -4483
rect -613 -4555 -567 -4517
rect -613 -4589 -607 -4555
rect -573 -4589 -567 -4555
rect -613 -4627 -567 -4589
rect -613 -4661 -607 -4627
rect -573 -4661 -567 -4627
rect -613 -4699 -567 -4661
rect -613 -4733 -607 -4699
rect -573 -4733 -567 -4699
rect -613 -4771 -567 -4733
rect -613 -4805 -607 -4771
rect -573 -4805 -567 -4771
rect -613 -4843 -567 -4805
rect -613 -4877 -607 -4843
rect -573 -4877 -567 -4843
rect -613 -4915 -567 -4877
rect -613 -4949 -607 -4915
rect -573 -4949 -567 -4915
rect -613 -4987 -567 -4949
rect -613 -5021 -607 -4987
rect -573 -5021 -567 -4987
rect -613 -5059 -567 -5021
rect -613 -5093 -607 -5059
rect -573 -5093 -567 -5059
rect -613 -5131 -567 -5093
rect -613 -5165 -607 -5131
rect -573 -5165 -567 -5131
rect -613 -5203 -567 -5165
rect -613 -5237 -607 -5203
rect -573 -5237 -567 -5203
rect -613 -5275 -567 -5237
rect -613 -5309 -607 -5275
rect -573 -5309 -567 -5275
rect -613 -5347 -567 -5309
rect -613 -5381 -607 -5347
rect -573 -5381 -567 -5347
rect -613 -5419 -567 -5381
rect -613 -5453 -607 -5419
rect -573 -5453 -567 -5419
rect -613 -5491 -567 -5453
rect -613 -5525 -607 -5491
rect -573 -5525 -567 -5491
rect -613 -5563 -567 -5525
rect -613 -5597 -607 -5563
rect -573 -5597 -567 -5563
rect -613 -5635 -567 -5597
rect -613 -5669 -607 -5635
rect -573 -5669 -567 -5635
rect -613 -5707 -567 -5669
rect -613 -5741 -607 -5707
rect -573 -5741 -567 -5707
rect -613 -5779 -567 -5741
rect -613 -5813 -607 -5779
rect -573 -5813 -567 -5779
rect -613 -5851 -567 -5813
rect -613 -5885 -607 -5851
rect -573 -5885 -567 -5851
rect -613 -5923 -567 -5885
rect -613 -5957 -607 -5923
rect -573 -5957 -567 -5923
rect -613 -6000 -567 -5957
rect -495 5957 -449 6000
rect -495 5923 -489 5957
rect -455 5923 -449 5957
rect -495 5885 -449 5923
rect -495 5851 -489 5885
rect -455 5851 -449 5885
rect -495 5813 -449 5851
rect -495 5779 -489 5813
rect -455 5779 -449 5813
rect -495 5741 -449 5779
rect -495 5707 -489 5741
rect -455 5707 -449 5741
rect -495 5669 -449 5707
rect -495 5635 -489 5669
rect -455 5635 -449 5669
rect -495 5597 -449 5635
rect -495 5563 -489 5597
rect -455 5563 -449 5597
rect -495 5525 -449 5563
rect -495 5491 -489 5525
rect -455 5491 -449 5525
rect -495 5453 -449 5491
rect -495 5419 -489 5453
rect -455 5419 -449 5453
rect -495 5381 -449 5419
rect -495 5347 -489 5381
rect -455 5347 -449 5381
rect -495 5309 -449 5347
rect -495 5275 -489 5309
rect -455 5275 -449 5309
rect -495 5237 -449 5275
rect -495 5203 -489 5237
rect -455 5203 -449 5237
rect -495 5165 -449 5203
rect -495 5131 -489 5165
rect -455 5131 -449 5165
rect -495 5093 -449 5131
rect -495 5059 -489 5093
rect -455 5059 -449 5093
rect -495 5021 -449 5059
rect -495 4987 -489 5021
rect -455 4987 -449 5021
rect -495 4949 -449 4987
rect -495 4915 -489 4949
rect -455 4915 -449 4949
rect -495 4877 -449 4915
rect -495 4843 -489 4877
rect -455 4843 -449 4877
rect -495 4805 -449 4843
rect -495 4771 -489 4805
rect -455 4771 -449 4805
rect -495 4733 -449 4771
rect -495 4699 -489 4733
rect -455 4699 -449 4733
rect -495 4661 -449 4699
rect -495 4627 -489 4661
rect -455 4627 -449 4661
rect -495 4589 -449 4627
rect -495 4555 -489 4589
rect -455 4555 -449 4589
rect -495 4517 -449 4555
rect -495 4483 -489 4517
rect -455 4483 -449 4517
rect -495 4445 -449 4483
rect -495 4411 -489 4445
rect -455 4411 -449 4445
rect -495 4373 -449 4411
rect -495 4339 -489 4373
rect -455 4339 -449 4373
rect -495 4301 -449 4339
rect -495 4267 -489 4301
rect -455 4267 -449 4301
rect -495 4229 -449 4267
rect -495 4195 -489 4229
rect -455 4195 -449 4229
rect -495 4157 -449 4195
rect -495 4123 -489 4157
rect -455 4123 -449 4157
rect -495 4085 -449 4123
rect -495 4051 -489 4085
rect -455 4051 -449 4085
rect -495 4013 -449 4051
rect -495 3979 -489 4013
rect -455 3979 -449 4013
rect -495 3941 -449 3979
rect -495 3907 -489 3941
rect -455 3907 -449 3941
rect -495 3869 -449 3907
rect -495 3835 -489 3869
rect -455 3835 -449 3869
rect -495 3797 -449 3835
rect -495 3763 -489 3797
rect -455 3763 -449 3797
rect -495 3725 -449 3763
rect -495 3691 -489 3725
rect -455 3691 -449 3725
rect -495 3653 -449 3691
rect -495 3619 -489 3653
rect -455 3619 -449 3653
rect -495 3581 -449 3619
rect -495 3547 -489 3581
rect -455 3547 -449 3581
rect -495 3509 -449 3547
rect -495 3475 -489 3509
rect -455 3475 -449 3509
rect -495 3437 -449 3475
rect -495 3403 -489 3437
rect -455 3403 -449 3437
rect -495 3365 -449 3403
rect -495 3331 -489 3365
rect -455 3331 -449 3365
rect -495 3293 -449 3331
rect -495 3259 -489 3293
rect -455 3259 -449 3293
rect -495 3221 -449 3259
rect -495 3187 -489 3221
rect -455 3187 -449 3221
rect -495 3149 -449 3187
rect -495 3115 -489 3149
rect -455 3115 -449 3149
rect -495 3077 -449 3115
rect -495 3043 -489 3077
rect -455 3043 -449 3077
rect -495 3005 -449 3043
rect -495 2971 -489 3005
rect -455 2971 -449 3005
rect -495 2933 -449 2971
rect -495 2899 -489 2933
rect -455 2899 -449 2933
rect -495 2861 -449 2899
rect -495 2827 -489 2861
rect -455 2827 -449 2861
rect -495 2789 -449 2827
rect -495 2755 -489 2789
rect -455 2755 -449 2789
rect -495 2717 -449 2755
rect -495 2683 -489 2717
rect -455 2683 -449 2717
rect -495 2645 -449 2683
rect -495 2611 -489 2645
rect -455 2611 -449 2645
rect -495 2573 -449 2611
rect -495 2539 -489 2573
rect -455 2539 -449 2573
rect -495 2501 -449 2539
rect -495 2467 -489 2501
rect -455 2467 -449 2501
rect -495 2429 -449 2467
rect -495 2395 -489 2429
rect -455 2395 -449 2429
rect -495 2357 -449 2395
rect -495 2323 -489 2357
rect -455 2323 -449 2357
rect -495 2285 -449 2323
rect -495 2251 -489 2285
rect -455 2251 -449 2285
rect -495 2213 -449 2251
rect -495 2179 -489 2213
rect -455 2179 -449 2213
rect -495 2141 -449 2179
rect -495 2107 -489 2141
rect -455 2107 -449 2141
rect -495 2069 -449 2107
rect -495 2035 -489 2069
rect -455 2035 -449 2069
rect -495 1997 -449 2035
rect -495 1963 -489 1997
rect -455 1963 -449 1997
rect -495 1925 -449 1963
rect -495 1891 -489 1925
rect -455 1891 -449 1925
rect -495 1853 -449 1891
rect -495 1819 -489 1853
rect -455 1819 -449 1853
rect -495 1781 -449 1819
rect -495 1747 -489 1781
rect -455 1747 -449 1781
rect -495 1709 -449 1747
rect -495 1675 -489 1709
rect -455 1675 -449 1709
rect -495 1637 -449 1675
rect -495 1603 -489 1637
rect -455 1603 -449 1637
rect -495 1565 -449 1603
rect -495 1531 -489 1565
rect -455 1531 -449 1565
rect -495 1493 -449 1531
rect -495 1459 -489 1493
rect -455 1459 -449 1493
rect -495 1421 -449 1459
rect -495 1387 -489 1421
rect -455 1387 -449 1421
rect -495 1349 -449 1387
rect -495 1315 -489 1349
rect -455 1315 -449 1349
rect -495 1277 -449 1315
rect -495 1243 -489 1277
rect -455 1243 -449 1277
rect -495 1205 -449 1243
rect -495 1171 -489 1205
rect -455 1171 -449 1205
rect -495 1133 -449 1171
rect -495 1099 -489 1133
rect -455 1099 -449 1133
rect -495 1061 -449 1099
rect -495 1027 -489 1061
rect -455 1027 -449 1061
rect -495 989 -449 1027
rect -495 955 -489 989
rect -455 955 -449 989
rect -495 917 -449 955
rect -495 883 -489 917
rect -455 883 -449 917
rect -495 845 -449 883
rect -495 811 -489 845
rect -455 811 -449 845
rect -495 773 -449 811
rect -495 739 -489 773
rect -455 739 -449 773
rect -495 701 -449 739
rect -495 667 -489 701
rect -455 667 -449 701
rect -495 629 -449 667
rect -495 595 -489 629
rect -455 595 -449 629
rect -495 557 -449 595
rect -495 523 -489 557
rect -455 523 -449 557
rect -495 485 -449 523
rect -495 451 -489 485
rect -455 451 -449 485
rect -495 413 -449 451
rect -495 379 -489 413
rect -455 379 -449 413
rect -495 341 -449 379
rect -495 307 -489 341
rect -455 307 -449 341
rect -495 269 -449 307
rect -495 235 -489 269
rect -455 235 -449 269
rect -495 197 -449 235
rect -495 163 -489 197
rect -455 163 -449 197
rect -495 125 -449 163
rect -495 91 -489 125
rect -455 91 -449 125
rect -495 53 -449 91
rect -495 19 -489 53
rect -455 19 -449 53
rect -495 -19 -449 19
rect -495 -53 -489 -19
rect -455 -53 -449 -19
rect -495 -91 -449 -53
rect -495 -125 -489 -91
rect -455 -125 -449 -91
rect -495 -163 -449 -125
rect -495 -197 -489 -163
rect -455 -197 -449 -163
rect -495 -235 -449 -197
rect -495 -269 -489 -235
rect -455 -269 -449 -235
rect -495 -307 -449 -269
rect -495 -341 -489 -307
rect -455 -341 -449 -307
rect -495 -379 -449 -341
rect -495 -413 -489 -379
rect -455 -413 -449 -379
rect -495 -451 -449 -413
rect -495 -485 -489 -451
rect -455 -485 -449 -451
rect -495 -523 -449 -485
rect -495 -557 -489 -523
rect -455 -557 -449 -523
rect -495 -595 -449 -557
rect -495 -629 -489 -595
rect -455 -629 -449 -595
rect -495 -667 -449 -629
rect -495 -701 -489 -667
rect -455 -701 -449 -667
rect -495 -739 -449 -701
rect -495 -773 -489 -739
rect -455 -773 -449 -739
rect -495 -811 -449 -773
rect -495 -845 -489 -811
rect -455 -845 -449 -811
rect -495 -883 -449 -845
rect -495 -917 -489 -883
rect -455 -917 -449 -883
rect -495 -955 -449 -917
rect -495 -989 -489 -955
rect -455 -989 -449 -955
rect -495 -1027 -449 -989
rect -495 -1061 -489 -1027
rect -455 -1061 -449 -1027
rect -495 -1099 -449 -1061
rect -495 -1133 -489 -1099
rect -455 -1133 -449 -1099
rect -495 -1171 -449 -1133
rect -495 -1205 -489 -1171
rect -455 -1205 -449 -1171
rect -495 -1243 -449 -1205
rect -495 -1277 -489 -1243
rect -455 -1277 -449 -1243
rect -495 -1315 -449 -1277
rect -495 -1349 -489 -1315
rect -455 -1349 -449 -1315
rect -495 -1387 -449 -1349
rect -495 -1421 -489 -1387
rect -455 -1421 -449 -1387
rect -495 -1459 -449 -1421
rect -495 -1493 -489 -1459
rect -455 -1493 -449 -1459
rect -495 -1531 -449 -1493
rect -495 -1565 -489 -1531
rect -455 -1565 -449 -1531
rect -495 -1603 -449 -1565
rect -495 -1637 -489 -1603
rect -455 -1637 -449 -1603
rect -495 -1675 -449 -1637
rect -495 -1709 -489 -1675
rect -455 -1709 -449 -1675
rect -495 -1747 -449 -1709
rect -495 -1781 -489 -1747
rect -455 -1781 -449 -1747
rect -495 -1819 -449 -1781
rect -495 -1853 -489 -1819
rect -455 -1853 -449 -1819
rect -495 -1891 -449 -1853
rect -495 -1925 -489 -1891
rect -455 -1925 -449 -1891
rect -495 -1963 -449 -1925
rect -495 -1997 -489 -1963
rect -455 -1997 -449 -1963
rect -495 -2035 -449 -1997
rect -495 -2069 -489 -2035
rect -455 -2069 -449 -2035
rect -495 -2107 -449 -2069
rect -495 -2141 -489 -2107
rect -455 -2141 -449 -2107
rect -495 -2179 -449 -2141
rect -495 -2213 -489 -2179
rect -455 -2213 -449 -2179
rect -495 -2251 -449 -2213
rect -495 -2285 -489 -2251
rect -455 -2285 -449 -2251
rect -495 -2323 -449 -2285
rect -495 -2357 -489 -2323
rect -455 -2357 -449 -2323
rect -495 -2395 -449 -2357
rect -495 -2429 -489 -2395
rect -455 -2429 -449 -2395
rect -495 -2467 -449 -2429
rect -495 -2501 -489 -2467
rect -455 -2501 -449 -2467
rect -495 -2539 -449 -2501
rect -495 -2573 -489 -2539
rect -455 -2573 -449 -2539
rect -495 -2611 -449 -2573
rect -495 -2645 -489 -2611
rect -455 -2645 -449 -2611
rect -495 -2683 -449 -2645
rect -495 -2717 -489 -2683
rect -455 -2717 -449 -2683
rect -495 -2755 -449 -2717
rect -495 -2789 -489 -2755
rect -455 -2789 -449 -2755
rect -495 -2827 -449 -2789
rect -495 -2861 -489 -2827
rect -455 -2861 -449 -2827
rect -495 -2899 -449 -2861
rect -495 -2933 -489 -2899
rect -455 -2933 -449 -2899
rect -495 -2971 -449 -2933
rect -495 -3005 -489 -2971
rect -455 -3005 -449 -2971
rect -495 -3043 -449 -3005
rect -495 -3077 -489 -3043
rect -455 -3077 -449 -3043
rect -495 -3115 -449 -3077
rect -495 -3149 -489 -3115
rect -455 -3149 -449 -3115
rect -495 -3187 -449 -3149
rect -495 -3221 -489 -3187
rect -455 -3221 -449 -3187
rect -495 -3259 -449 -3221
rect -495 -3293 -489 -3259
rect -455 -3293 -449 -3259
rect -495 -3331 -449 -3293
rect -495 -3365 -489 -3331
rect -455 -3365 -449 -3331
rect -495 -3403 -449 -3365
rect -495 -3437 -489 -3403
rect -455 -3437 -449 -3403
rect -495 -3475 -449 -3437
rect -495 -3509 -489 -3475
rect -455 -3509 -449 -3475
rect -495 -3547 -449 -3509
rect -495 -3581 -489 -3547
rect -455 -3581 -449 -3547
rect -495 -3619 -449 -3581
rect -495 -3653 -489 -3619
rect -455 -3653 -449 -3619
rect -495 -3691 -449 -3653
rect -495 -3725 -489 -3691
rect -455 -3725 -449 -3691
rect -495 -3763 -449 -3725
rect -495 -3797 -489 -3763
rect -455 -3797 -449 -3763
rect -495 -3835 -449 -3797
rect -495 -3869 -489 -3835
rect -455 -3869 -449 -3835
rect -495 -3907 -449 -3869
rect -495 -3941 -489 -3907
rect -455 -3941 -449 -3907
rect -495 -3979 -449 -3941
rect -495 -4013 -489 -3979
rect -455 -4013 -449 -3979
rect -495 -4051 -449 -4013
rect -495 -4085 -489 -4051
rect -455 -4085 -449 -4051
rect -495 -4123 -449 -4085
rect -495 -4157 -489 -4123
rect -455 -4157 -449 -4123
rect -495 -4195 -449 -4157
rect -495 -4229 -489 -4195
rect -455 -4229 -449 -4195
rect -495 -4267 -449 -4229
rect -495 -4301 -489 -4267
rect -455 -4301 -449 -4267
rect -495 -4339 -449 -4301
rect -495 -4373 -489 -4339
rect -455 -4373 -449 -4339
rect -495 -4411 -449 -4373
rect -495 -4445 -489 -4411
rect -455 -4445 -449 -4411
rect -495 -4483 -449 -4445
rect -495 -4517 -489 -4483
rect -455 -4517 -449 -4483
rect -495 -4555 -449 -4517
rect -495 -4589 -489 -4555
rect -455 -4589 -449 -4555
rect -495 -4627 -449 -4589
rect -495 -4661 -489 -4627
rect -455 -4661 -449 -4627
rect -495 -4699 -449 -4661
rect -495 -4733 -489 -4699
rect -455 -4733 -449 -4699
rect -495 -4771 -449 -4733
rect -495 -4805 -489 -4771
rect -455 -4805 -449 -4771
rect -495 -4843 -449 -4805
rect -495 -4877 -489 -4843
rect -455 -4877 -449 -4843
rect -495 -4915 -449 -4877
rect -495 -4949 -489 -4915
rect -455 -4949 -449 -4915
rect -495 -4987 -449 -4949
rect -495 -5021 -489 -4987
rect -455 -5021 -449 -4987
rect -495 -5059 -449 -5021
rect -495 -5093 -489 -5059
rect -455 -5093 -449 -5059
rect -495 -5131 -449 -5093
rect -495 -5165 -489 -5131
rect -455 -5165 -449 -5131
rect -495 -5203 -449 -5165
rect -495 -5237 -489 -5203
rect -455 -5237 -449 -5203
rect -495 -5275 -449 -5237
rect -495 -5309 -489 -5275
rect -455 -5309 -449 -5275
rect -495 -5347 -449 -5309
rect -495 -5381 -489 -5347
rect -455 -5381 -449 -5347
rect -495 -5419 -449 -5381
rect -495 -5453 -489 -5419
rect -455 -5453 -449 -5419
rect -495 -5491 -449 -5453
rect -495 -5525 -489 -5491
rect -455 -5525 -449 -5491
rect -495 -5563 -449 -5525
rect -495 -5597 -489 -5563
rect -455 -5597 -449 -5563
rect -495 -5635 -449 -5597
rect -495 -5669 -489 -5635
rect -455 -5669 -449 -5635
rect -495 -5707 -449 -5669
rect -495 -5741 -489 -5707
rect -455 -5741 -449 -5707
rect -495 -5779 -449 -5741
rect -495 -5813 -489 -5779
rect -455 -5813 -449 -5779
rect -495 -5851 -449 -5813
rect -495 -5885 -489 -5851
rect -455 -5885 -449 -5851
rect -495 -5923 -449 -5885
rect -495 -5957 -489 -5923
rect -455 -5957 -449 -5923
rect -495 -6000 -449 -5957
rect -377 5957 -331 6000
rect -377 5923 -371 5957
rect -337 5923 -331 5957
rect -377 5885 -331 5923
rect -377 5851 -371 5885
rect -337 5851 -331 5885
rect -377 5813 -331 5851
rect -377 5779 -371 5813
rect -337 5779 -331 5813
rect -377 5741 -331 5779
rect -377 5707 -371 5741
rect -337 5707 -331 5741
rect -377 5669 -331 5707
rect -377 5635 -371 5669
rect -337 5635 -331 5669
rect -377 5597 -331 5635
rect -377 5563 -371 5597
rect -337 5563 -331 5597
rect -377 5525 -331 5563
rect -377 5491 -371 5525
rect -337 5491 -331 5525
rect -377 5453 -331 5491
rect -377 5419 -371 5453
rect -337 5419 -331 5453
rect -377 5381 -331 5419
rect -377 5347 -371 5381
rect -337 5347 -331 5381
rect -377 5309 -331 5347
rect -377 5275 -371 5309
rect -337 5275 -331 5309
rect -377 5237 -331 5275
rect -377 5203 -371 5237
rect -337 5203 -331 5237
rect -377 5165 -331 5203
rect -377 5131 -371 5165
rect -337 5131 -331 5165
rect -377 5093 -331 5131
rect -377 5059 -371 5093
rect -337 5059 -331 5093
rect -377 5021 -331 5059
rect -377 4987 -371 5021
rect -337 4987 -331 5021
rect -377 4949 -331 4987
rect -377 4915 -371 4949
rect -337 4915 -331 4949
rect -377 4877 -331 4915
rect -377 4843 -371 4877
rect -337 4843 -331 4877
rect -377 4805 -331 4843
rect -377 4771 -371 4805
rect -337 4771 -331 4805
rect -377 4733 -331 4771
rect -377 4699 -371 4733
rect -337 4699 -331 4733
rect -377 4661 -331 4699
rect -377 4627 -371 4661
rect -337 4627 -331 4661
rect -377 4589 -331 4627
rect -377 4555 -371 4589
rect -337 4555 -331 4589
rect -377 4517 -331 4555
rect -377 4483 -371 4517
rect -337 4483 -331 4517
rect -377 4445 -331 4483
rect -377 4411 -371 4445
rect -337 4411 -331 4445
rect -377 4373 -331 4411
rect -377 4339 -371 4373
rect -337 4339 -331 4373
rect -377 4301 -331 4339
rect -377 4267 -371 4301
rect -337 4267 -331 4301
rect -377 4229 -331 4267
rect -377 4195 -371 4229
rect -337 4195 -331 4229
rect -377 4157 -331 4195
rect -377 4123 -371 4157
rect -337 4123 -331 4157
rect -377 4085 -331 4123
rect -377 4051 -371 4085
rect -337 4051 -331 4085
rect -377 4013 -331 4051
rect -377 3979 -371 4013
rect -337 3979 -331 4013
rect -377 3941 -331 3979
rect -377 3907 -371 3941
rect -337 3907 -331 3941
rect -377 3869 -331 3907
rect -377 3835 -371 3869
rect -337 3835 -331 3869
rect -377 3797 -331 3835
rect -377 3763 -371 3797
rect -337 3763 -331 3797
rect -377 3725 -331 3763
rect -377 3691 -371 3725
rect -337 3691 -331 3725
rect -377 3653 -331 3691
rect -377 3619 -371 3653
rect -337 3619 -331 3653
rect -377 3581 -331 3619
rect -377 3547 -371 3581
rect -337 3547 -331 3581
rect -377 3509 -331 3547
rect -377 3475 -371 3509
rect -337 3475 -331 3509
rect -377 3437 -331 3475
rect -377 3403 -371 3437
rect -337 3403 -331 3437
rect -377 3365 -331 3403
rect -377 3331 -371 3365
rect -337 3331 -331 3365
rect -377 3293 -331 3331
rect -377 3259 -371 3293
rect -337 3259 -331 3293
rect -377 3221 -331 3259
rect -377 3187 -371 3221
rect -337 3187 -331 3221
rect -377 3149 -331 3187
rect -377 3115 -371 3149
rect -337 3115 -331 3149
rect -377 3077 -331 3115
rect -377 3043 -371 3077
rect -337 3043 -331 3077
rect -377 3005 -331 3043
rect -377 2971 -371 3005
rect -337 2971 -331 3005
rect -377 2933 -331 2971
rect -377 2899 -371 2933
rect -337 2899 -331 2933
rect -377 2861 -331 2899
rect -377 2827 -371 2861
rect -337 2827 -331 2861
rect -377 2789 -331 2827
rect -377 2755 -371 2789
rect -337 2755 -331 2789
rect -377 2717 -331 2755
rect -377 2683 -371 2717
rect -337 2683 -331 2717
rect -377 2645 -331 2683
rect -377 2611 -371 2645
rect -337 2611 -331 2645
rect -377 2573 -331 2611
rect -377 2539 -371 2573
rect -337 2539 -331 2573
rect -377 2501 -331 2539
rect -377 2467 -371 2501
rect -337 2467 -331 2501
rect -377 2429 -331 2467
rect -377 2395 -371 2429
rect -337 2395 -331 2429
rect -377 2357 -331 2395
rect -377 2323 -371 2357
rect -337 2323 -331 2357
rect -377 2285 -331 2323
rect -377 2251 -371 2285
rect -337 2251 -331 2285
rect -377 2213 -331 2251
rect -377 2179 -371 2213
rect -337 2179 -331 2213
rect -377 2141 -331 2179
rect -377 2107 -371 2141
rect -337 2107 -331 2141
rect -377 2069 -331 2107
rect -377 2035 -371 2069
rect -337 2035 -331 2069
rect -377 1997 -331 2035
rect -377 1963 -371 1997
rect -337 1963 -331 1997
rect -377 1925 -331 1963
rect -377 1891 -371 1925
rect -337 1891 -331 1925
rect -377 1853 -331 1891
rect -377 1819 -371 1853
rect -337 1819 -331 1853
rect -377 1781 -331 1819
rect -377 1747 -371 1781
rect -337 1747 -331 1781
rect -377 1709 -331 1747
rect -377 1675 -371 1709
rect -337 1675 -331 1709
rect -377 1637 -331 1675
rect -377 1603 -371 1637
rect -337 1603 -331 1637
rect -377 1565 -331 1603
rect -377 1531 -371 1565
rect -337 1531 -331 1565
rect -377 1493 -331 1531
rect -377 1459 -371 1493
rect -337 1459 -331 1493
rect -377 1421 -331 1459
rect -377 1387 -371 1421
rect -337 1387 -331 1421
rect -377 1349 -331 1387
rect -377 1315 -371 1349
rect -337 1315 -331 1349
rect -377 1277 -331 1315
rect -377 1243 -371 1277
rect -337 1243 -331 1277
rect -377 1205 -331 1243
rect -377 1171 -371 1205
rect -337 1171 -331 1205
rect -377 1133 -331 1171
rect -377 1099 -371 1133
rect -337 1099 -331 1133
rect -377 1061 -331 1099
rect -377 1027 -371 1061
rect -337 1027 -331 1061
rect -377 989 -331 1027
rect -377 955 -371 989
rect -337 955 -331 989
rect -377 917 -331 955
rect -377 883 -371 917
rect -337 883 -331 917
rect -377 845 -331 883
rect -377 811 -371 845
rect -337 811 -331 845
rect -377 773 -331 811
rect -377 739 -371 773
rect -337 739 -331 773
rect -377 701 -331 739
rect -377 667 -371 701
rect -337 667 -331 701
rect -377 629 -331 667
rect -377 595 -371 629
rect -337 595 -331 629
rect -377 557 -331 595
rect -377 523 -371 557
rect -337 523 -331 557
rect -377 485 -331 523
rect -377 451 -371 485
rect -337 451 -331 485
rect -377 413 -331 451
rect -377 379 -371 413
rect -337 379 -331 413
rect -377 341 -331 379
rect -377 307 -371 341
rect -337 307 -331 341
rect -377 269 -331 307
rect -377 235 -371 269
rect -337 235 -331 269
rect -377 197 -331 235
rect -377 163 -371 197
rect -337 163 -331 197
rect -377 125 -331 163
rect -377 91 -371 125
rect -337 91 -331 125
rect -377 53 -331 91
rect -377 19 -371 53
rect -337 19 -331 53
rect -377 -19 -331 19
rect -377 -53 -371 -19
rect -337 -53 -331 -19
rect -377 -91 -331 -53
rect -377 -125 -371 -91
rect -337 -125 -331 -91
rect -377 -163 -331 -125
rect -377 -197 -371 -163
rect -337 -197 -331 -163
rect -377 -235 -331 -197
rect -377 -269 -371 -235
rect -337 -269 -331 -235
rect -377 -307 -331 -269
rect -377 -341 -371 -307
rect -337 -341 -331 -307
rect -377 -379 -331 -341
rect -377 -413 -371 -379
rect -337 -413 -331 -379
rect -377 -451 -331 -413
rect -377 -485 -371 -451
rect -337 -485 -331 -451
rect -377 -523 -331 -485
rect -377 -557 -371 -523
rect -337 -557 -331 -523
rect -377 -595 -331 -557
rect -377 -629 -371 -595
rect -337 -629 -331 -595
rect -377 -667 -331 -629
rect -377 -701 -371 -667
rect -337 -701 -331 -667
rect -377 -739 -331 -701
rect -377 -773 -371 -739
rect -337 -773 -331 -739
rect -377 -811 -331 -773
rect -377 -845 -371 -811
rect -337 -845 -331 -811
rect -377 -883 -331 -845
rect -377 -917 -371 -883
rect -337 -917 -331 -883
rect -377 -955 -331 -917
rect -377 -989 -371 -955
rect -337 -989 -331 -955
rect -377 -1027 -331 -989
rect -377 -1061 -371 -1027
rect -337 -1061 -331 -1027
rect -377 -1099 -331 -1061
rect -377 -1133 -371 -1099
rect -337 -1133 -331 -1099
rect -377 -1171 -331 -1133
rect -377 -1205 -371 -1171
rect -337 -1205 -331 -1171
rect -377 -1243 -331 -1205
rect -377 -1277 -371 -1243
rect -337 -1277 -331 -1243
rect -377 -1315 -331 -1277
rect -377 -1349 -371 -1315
rect -337 -1349 -331 -1315
rect -377 -1387 -331 -1349
rect -377 -1421 -371 -1387
rect -337 -1421 -331 -1387
rect -377 -1459 -331 -1421
rect -377 -1493 -371 -1459
rect -337 -1493 -331 -1459
rect -377 -1531 -331 -1493
rect -377 -1565 -371 -1531
rect -337 -1565 -331 -1531
rect -377 -1603 -331 -1565
rect -377 -1637 -371 -1603
rect -337 -1637 -331 -1603
rect -377 -1675 -331 -1637
rect -377 -1709 -371 -1675
rect -337 -1709 -331 -1675
rect -377 -1747 -331 -1709
rect -377 -1781 -371 -1747
rect -337 -1781 -331 -1747
rect -377 -1819 -331 -1781
rect -377 -1853 -371 -1819
rect -337 -1853 -331 -1819
rect -377 -1891 -331 -1853
rect -377 -1925 -371 -1891
rect -337 -1925 -331 -1891
rect -377 -1963 -331 -1925
rect -377 -1997 -371 -1963
rect -337 -1997 -331 -1963
rect -377 -2035 -331 -1997
rect -377 -2069 -371 -2035
rect -337 -2069 -331 -2035
rect -377 -2107 -331 -2069
rect -377 -2141 -371 -2107
rect -337 -2141 -331 -2107
rect -377 -2179 -331 -2141
rect -377 -2213 -371 -2179
rect -337 -2213 -331 -2179
rect -377 -2251 -331 -2213
rect -377 -2285 -371 -2251
rect -337 -2285 -331 -2251
rect -377 -2323 -331 -2285
rect -377 -2357 -371 -2323
rect -337 -2357 -331 -2323
rect -377 -2395 -331 -2357
rect -377 -2429 -371 -2395
rect -337 -2429 -331 -2395
rect -377 -2467 -331 -2429
rect -377 -2501 -371 -2467
rect -337 -2501 -331 -2467
rect -377 -2539 -331 -2501
rect -377 -2573 -371 -2539
rect -337 -2573 -331 -2539
rect -377 -2611 -331 -2573
rect -377 -2645 -371 -2611
rect -337 -2645 -331 -2611
rect -377 -2683 -331 -2645
rect -377 -2717 -371 -2683
rect -337 -2717 -331 -2683
rect -377 -2755 -331 -2717
rect -377 -2789 -371 -2755
rect -337 -2789 -331 -2755
rect -377 -2827 -331 -2789
rect -377 -2861 -371 -2827
rect -337 -2861 -331 -2827
rect -377 -2899 -331 -2861
rect -377 -2933 -371 -2899
rect -337 -2933 -331 -2899
rect -377 -2971 -331 -2933
rect -377 -3005 -371 -2971
rect -337 -3005 -331 -2971
rect -377 -3043 -331 -3005
rect -377 -3077 -371 -3043
rect -337 -3077 -331 -3043
rect -377 -3115 -331 -3077
rect -377 -3149 -371 -3115
rect -337 -3149 -331 -3115
rect -377 -3187 -331 -3149
rect -377 -3221 -371 -3187
rect -337 -3221 -331 -3187
rect -377 -3259 -331 -3221
rect -377 -3293 -371 -3259
rect -337 -3293 -331 -3259
rect -377 -3331 -331 -3293
rect -377 -3365 -371 -3331
rect -337 -3365 -331 -3331
rect -377 -3403 -331 -3365
rect -377 -3437 -371 -3403
rect -337 -3437 -331 -3403
rect -377 -3475 -331 -3437
rect -377 -3509 -371 -3475
rect -337 -3509 -331 -3475
rect -377 -3547 -331 -3509
rect -377 -3581 -371 -3547
rect -337 -3581 -331 -3547
rect -377 -3619 -331 -3581
rect -377 -3653 -371 -3619
rect -337 -3653 -331 -3619
rect -377 -3691 -331 -3653
rect -377 -3725 -371 -3691
rect -337 -3725 -331 -3691
rect -377 -3763 -331 -3725
rect -377 -3797 -371 -3763
rect -337 -3797 -331 -3763
rect -377 -3835 -331 -3797
rect -377 -3869 -371 -3835
rect -337 -3869 -331 -3835
rect -377 -3907 -331 -3869
rect -377 -3941 -371 -3907
rect -337 -3941 -331 -3907
rect -377 -3979 -331 -3941
rect -377 -4013 -371 -3979
rect -337 -4013 -331 -3979
rect -377 -4051 -331 -4013
rect -377 -4085 -371 -4051
rect -337 -4085 -331 -4051
rect -377 -4123 -331 -4085
rect -377 -4157 -371 -4123
rect -337 -4157 -331 -4123
rect -377 -4195 -331 -4157
rect -377 -4229 -371 -4195
rect -337 -4229 -331 -4195
rect -377 -4267 -331 -4229
rect -377 -4301 -371 -4267
rect -337 -4301 -331 -4267
rect -377 -4339 -331 -4301
rect -377 -4373 -371 -4339
rect -337 -4373 -331 -4339
rect -377 -4411 -331 -4373
rect -377 -4445 -371 -4411
rect -337 -4445 -331 -4411
rect -377 -4483 -331 -4445
rect -377 -4517 -371 -4483
rect -337 -4517 -331 -4483
rect -377 -4555 -331 -4517
rect -377 -4589 -371 -4555
rect -337 -4589 -331 -4555
rect -377 -4627 -331 -4589
rect -377 -4661 -371 -4627
rect -337 -4661 -331 -4627
rect -377 -4699 -331 -4661
rect -377 -4733 -371 -4699
rect -337 -4733 -331 -4699
rect -377 -4771 -331 -4733
rect -377 -4805 -371 -4771
rect -337 -4805 -331 -4771
rect -377 -4843 -331 -4805
rect -377 -4877 -371 -4843
rect -337 -4877 -331 -4843
rect -377 -4915 -331 -4877
rect -377 -4949 -371 -4915
rect -337 -4949 -331 -4915
rect -377 -4987 -331 -4949
rect -377 -5021 -371 -4987
rect -337 -5021 -331 -4987
rect -377 -5059 -331 -5021
rect -377 -5093 -371 -5059
rect -337 -5093 -331 -5059
rect -377 -5131 -331 -5093
rect -377 -5165 -371 -5131
rect -337 -5165 -331 -5131
rect -377 -5203 -331 -5165
rect -377 -5237 -371 -5203
rect -337 -5237 -331 -5203
rect -377 -5275 -331 -5237
rect -377 -5309 -371 -5275
rect -337 -5309 -331 -5275
rect -377 -5347 -331 -5309
rect -377 -5381 -371 -5347
rect -337 -5381 -331 -5347
rect -377 -5419 -331 -5381
rect -377 -5453 -371 -5419
rect -337 -5453 -331 -5419
rect -377 -5491 -331 -5453
rect -377 -5525 -371 -5491
rect -337 -5525 -331 -5491
rect -377 -5563 -331 -5525
rect -377 -5597 -371 -5563
rect -337 -5597 -331 -5563
rect -377 -5635 -331 -5597
rect -377 -5669 -371 -5635
rect -337 -5669 -331 -5635
rect -377 -5707 -331 -5669
rect -377 -5741 -371 -5707
rect -337 -5741 -331 -5707
rect -377 -5779 -331 -5741
rect -377 -5813 -371 -5779
rect -337 -5813 -331 -5779
rect -377 -5851 -331 -5813
rect -377 -5885 -371 -5851
rect -337 -5885 -331 -5851
rect -377 -5923 -331 -5885
rect -377 -5957 -371 -5923
rect -337 -5957 -331 -5923
rect -377 -6000 -331 -5957
rect -259 5957 -213 6000
rect -259 5923 -253 5957
rect -219 5923 -213 5957
rect -259 5885 -213 5923
rect -259 5851 -253 5885
rect -219 5851 -213 5885
rect -259 5813 -213 5851
rect -259 5779 -253 5813
rect -219 5779 -213 5813
rect -259 5741 -213 5779
rect -259 5707 -253 5741
rect -219 5707 -213 5741
rect -259 5669 -213 5707
rect -259 5635 -253 5669
rect -219 5635 -213 5669
rect -259 5597 -213 5635
rect -259 5563 -253 5597
rect -219 5563 -213 5597
rect -259 5525 -213 5563
rect -259 5491 -253 5525
rect -219 5491 -213 5525
rect -259 5453 -213 5491
rect -259 5419 -253 5453
rect -219 5419 -213 5453
rect -259 5381 -213 5419
rect -259 5347 -253 5381
rect -219 5347 -213 5381
rect -259 5309 -213 5347
rect -259 5275 -253 5309
rect -219 5275 -213 5309
rect -259 5237 -213 5275
rect -259 5203 -253 5237
rect -219 5203 -213 5237
rect -259 5165 -213 5203
rect -259 5131 -253 5165
rect -219 5131 -213 5165
rect -259 5093 -213 5131
rect -259 5059 -253 5093
rect -219 5059 -213 5093
rect -259 5021 -213 5059
rect -259 4987 -253 5021
rect -219 4987 -213 5021
rect -259 4949 -213 4987
rect -259 4915 -253 4949
rect -219 4915 -213 4949
rect -259 4877 -213 4915
rect -259 4843 -253 4877
rect -219 4843 -213 4877
rect -259 4805 -213 4843
rect -259 4771 -253 4805
rect -219 4771 -213 4805
rect -259 4733 -213 4771
rect -259 4699 -253 4733
rect -219 4699 -213 4733
rect -259 4661 -213 4699
rect -259 4627 -253 4661
rect -219 4627 -213 4661
rect -259 4589 -213 4627
rect -259 4555 -253 4589
rect -219 4555 -213 4589
rect -259 4517 -213 4555
rect -259 4483 -253 4517
rect -219 4483 -213 4517
rect -259 4445 -213 4483
rect -259 4411 -253 4445
rect -219 4411 -213 4445
rect -259 4373 -213 4411
rect -259 4339 -253 4373
rect -219 4339 -213 4373
rect -259 4301 -213 4339
rect -259 4267 -253 4301
rect -219 4267 -213 4301
rect -259 4229 -213 4267
rect -259 4195 -253 4229
rect -219 4195 -213 4229
rect -259 4157 -213 4195
rect -259 4123 -253 4157
rect -219 4123 -213 4157
rect -259 4085 -213 4123
rect -259 4051 -253 4085
rect -219 4051 -213 4085
rect -259 4013 -213 4051
rect -259 3979 -253 4013
rect -219 3979 -213 4013
rect -259 3941 -213 3979
rect -259 3907 -253 3941
rect -219 3907 -213 3941
rect -259 3869 -213 3907
rect -259 3835 -253 3869
rect -219 3835 -213 3869
rect -259 3797 -213 3835
rect -259 3763 -253 3797
rect -219 3763 -213 3797
rect -259 3725 -213 3763
rect -259 3691 -253 3725
rect -219 3691 -213 3725
rect -259 3653 -213 3691
rect -259 3619 -253 3653
rect -219 3619 -213 3653
rect -259 3581 -213 3619
rect -259 3547 -253 3581
rect -219 3547 -213 3581
rect -259 3509 -213 3547
rect -259 3475 -253 3509
rect -219 3475 -213 3509
rect -259 3437 -213 3475
rect -259 3403 -253 3437
rect -219 3403 -213 3437
rect -259 3365 -213 3403
rect -259 3331 -253 3365
rect -219 3331 -213 3365
rect -259 3293 -213 3331
rect -259 3259 -253 3293
rect -219 3259 -213 3293
rect -259 3221 -213 3259
rect -259 3187 -253 3221
rect -219 3187 -213 3221
rect -259 3149 -213 3187
rect -259 3115 -253 3149
rect -219 3115 -213 3149
rect -259 3077 -213 3115
rect -259 3043 -253 3077
rect -219 3043 -213 3077
rect -259 3005 -213 3043
rect -259 2971 -253 3005
rect -219 2971 -213 3005
rect -259 2933 -213 2971
rect -259 2899 -253 2933
rect -219 2899 -213 2933
rect -259 2861 -213 2899
rect -259 2827 -253 2861
rect -219 2827 -213 2861
rect -259 2789 -213 2827
rect -259 2755 -253 2789
rect -219 2755 -213 2789
rect -259 2717 -213 2755
rect -259 2683 -253 2717
rect -219 2683 -213 2717
rect -259 2645 -213 2683
rect -259 2611 -253 2645
rect -219 2611 -213 2645
rect -259 2573 -213 2611
rect -259 2539 -253 2573
rect -219 2539 -213 2573
rect -259 2501 -213 2539
rect -259 2467 -253 2501
rect -219 2467 -213 2501
rect -259 2429 -213 2467
rect -259 2395 -253 2429
rect -219 2395 -213 2429
rect -259 2357 -213 2395
rect -259 2323 -253 2357
rect -219 2323 -213 2357
rect -259 2285 -213 2323
rect -259 2251 -253 2285
rect -219 2251 -213 2285
rect -259 2213 -213 2251
rect -259 2179 -253 2213
rect -219 2179 -213 2213
rect -259 2141 -213 2179
rect -259 2107 -253 2141
rect -219 2107 -213 2141
rect -259 2069 -213 2107
rect -259 2035 -253 2069
rect -219 2035 -213 2069
rect -259 1997 -213 2035
rect -259 1963 -253 1997
rect -219 1963 -213 1997
rect -259 1925 -213 1963
rect -259 1891 -253 1925
rect -219 1891 -213 1925
rect -259 1853 -213 1891
rect -259 1819 -253 1853
rect -219 1819 -213 1853
rect -259 1781 -213 1819
rect -259 1747 -253 1781
rect -219 1747 -213 1781
rect -259 1709 -213 1747
rect -259 1675 -253 1709
rect -219 1675 -213 1709
rect -259 1637 -213 1675
rect -259 1603 -253 1637
rect -219 1603 -213 1637
rect -259 1565 -213 1603
rect -259 1531 -253 1565
rect -219 1531 -213 1565
rect -259 1493 -213 1531
rect -259 1459 -253 1493
rect -219 1459 -213 1493
rect -259 1421 -213 1459
rect -259 1387 -253 1421
rect -219 1387 -213 1421
rect -259 1349 -213 1387
rect -259 1315 -253 1349
rect -219 1315 -213 1349
rect -259 1277 -213 1315
rect -259 1243 -253 1277
rect -219 1243 -213 1277
rect -259 1205 -213 1243
rect -259 1171 -253 1205
rect -219 1171 -213 1205
rect -259 1133 -213 1171
rect -259 1099 -253 1133
rect -219 1099 -213 1133
rect -259 1061 -213 1099
rect -259 1027 -253 1061
rect -219 1027 -213 1061
rect -259 989 -213 1027
rect -259 955 -253 989
rect -219 955 -213 989
rect -259 917 -213 955
rect -259 883 -253 917
rect -219 883 -213 917
rect -259 845 -213 883
rect -259 811 -253 845
rect -219 811 -213 845
rect -259 773 -213 811
rect -259 739 -253 773
rect -219 739 -213 773
rect -259 701 -213 739
rect -259 667 -253 701
rect -219 667 -213 701
rect -259 629 -213 667
rect -259 595 -253 629
rect -219 595 -213 629
rect -259 557 -213 595
rect -259 523 -253 557
rect -219 523 -213 557
rect -259 485 -213 523
rect -259 451 -253 485
rect -219 451 -213 485
rect -259 413 -213 451
rect -259 379 -253 413
rect -219 379 -213 413
rect -259 341 -213 379
rect -259 307 -253 341
rect -219 307 -213 341
rect -259 269 -213 307
rect -259 235 -253 269
rect -219 235 -213 269
rect -259 197 -213 235
rect -259 163 -253 197
rect -219 163 -213 197
rect -259 125 -213 163
rect -259 91 -253 125
rect -219 91 -213 125
rect -259 53 -213 91
rect -259 19 -253 53
rect -219 19 -213 53
rect -259 -19 -213 19
rect -259 -53 -253 -19
rect -219 -53 -213 -19
rect -259 -91 -213 -53
rect -259 -125 -253 -91
rect -219 -125 -213 -91
rect -259 -163 -213 -125
rect -259 -197 -253 -163
rect -219 -197 -213 -163
rect -259 -235 -213 -197
rect -259 -269 -253 -235
rect -219 -269 -213 -235
rect -259 -307 -213 -269
rect -259 -341 -253 -307
rect -219 -341 -213 -307
rect -259 -379 -213 -341
rect -259 -413 -253 -379
rect -219 -413 -213 -379
rect -259 -451 -213 -413
rect -259 -485 -253 -451
rect -219 -485 -213 -451
rect -259 -523 -213 -485
rect -259 -557 -253 -523
rect -219 -557 -213 -523
rect -259 -595 -213 -557
rect -259 -629 -253 -595
rect -219 -629 -213 -595
rect -259 -667 -213 -629
rect -259 -701 -253 -667
rect -219 -701 -213 -667
rect -259 -739 -213 -701
rect -259 -773 -253 -739
rect -219 -773 -213 -739
rect -259 -811 -213 -773
rect -259 -845 -253 -811
rect -219 -845 -213 -811
rect -259 -883 -213 -845
rect -259 -917 -253 -883
rect -219 -917 -213 -883
rect -259 -955 -213 -917
rect -259 -989 -253 -955
rect -219 -989 -213 -955
rect -259 -1027 -213 -989
rect -259 -1061 -253 -1027
rect -219 -1061 -213 -1027
rect -259 -1099 -213 -1061
rect -259 -1133 -253 -1099
rect -219 -1133 -213 -1099
rect -259 -1171 -213 -1133
rect -259 -1205 -253 -1171
rect -219 -1205 -213 -1171
rect -259 -1243 -213 -1205
rect -259 -1277 -253 -1243
rect -219 -1277 -213 -1243
rect -259 -1315 -213 -1277
rect -259 -1349 -253 -1315
rect -219 -1349 -213 -1315
rect -259 -1387 -213 -1349
rect -259 -1421 -253 -1387
rect -219 -1421 -213 -1387
rect -259 -1459 -213 -1421
rect -259 -1493 -253 -1459
rect -219 -1493 -213 -1459
rect -259 -1531 -213 -1493
rect -259 -1565 -253 -1531
rect -219 -1565 -213 -1531
rect -259 -1603 -213 -1565
rect -259 -1637 -253 -1603
rect -219 -1637 -213 -1603
rect -259 -1675 -213 -1637
rect -259 -1709 -253 -1675
rect -219 -1709 -213 -1675
rect -259 -1747 -213 -1709
rect -259 -1781 -253 -1747
rect -219 -1781 -213 -1747
rect -259 -1819 -213 -1781
rect -259 -1853 -253 -1819
rect -219 -1853 -213 -1819
rect -259 -1891 -213 -1853
rect -259 -1925 -253 -1891
rect -219 -1925 -213 -1891
rect -259 -1963 -213 -1925
rect -259 -1997 -253 -1963
rect -219 -1997 -213 -1963
rect -259 -2035 -213 -1997
rect -259 -2069 -253 -2035
rect -219 -2069 -213 -2035
rect -259 -2107 -213 -2069
rect -259 -2141 -253 -2107
rect -219 -2141 -213 -2107
rect -259 -2179 -213 -2141
rect -259 -2213 -253 -2179
rect -219 -2213 -213 -2179
rect -259 -2251 -213 -2213
rect -259 -2285 -253 -2251
rect -219 -2285 -213 -2251
rect -259 -2323 -213 -2285
rect -259 -2357 -253 -2323
rect -219 -2357 -213 -2323
rect -259 -2395 -213 -2357
rect -259 -2429 -253 -2395
rect -219 -2429 -213 -2395
rect -259 -2467 -213 -2429
rect -259 -2501 -253 -2467
rect -219 -2501 -213 -2467
rect -259 -2539 -213 -2501
rect -259 -2573 -253 -2539
rect -219 -2573 -213 -2539
rect -259 -2611 -213 -2573
rect -259 -2645 -253 -2611
rect -219 -2645 -213 -2611
rect -259 -2683 -213 -2645
rect -259 -2717 -253 -2683
rect -219 -2717 -213 -2683
rect -259 -2755 -213 -2717
rect -259 -2789 -253 -2755
rect -219 -2789 -213 -2755
rect -259 -2827 -213 -2789
rect -259 -2861 -253 -2827
rect -219 -2861 -213 -2827
rect -259 -2899 -213 -2861
rect -259 -2933 -253 -2899
rect -219 -2933 -213 -2899
rect -259 -2971 -213 -2933
rect -259 -3005 -253 -2971
rect -219 -3005 -213 -2971
rect -259 -3043 -213 -3005
rect -259 -3077 -253 -3043
rect -219 -3077 -213 -3043
rect -259 -3115 -213 -3077
rect -259 -3149 -253 -3115
rect -219 -3149 -213 -3115
rect -259 -3187 -213 -3149
rect -259 -3221 -253 -3187
rect -219 -3221 -213 -3187
rect -259 -3259 -213 -3221
rect -259 -3293 -253 -3259
rect -219 -3293 -213 -3259
rect -259 -3331 -213 -3293
rect -259 -3365 -253 -3331
rect -219 -3365 -213 -3331
rect -259 -3403 -213 -3365
rect -259 -3437 -253 -3403
rect -219 -3437 -213 -3403
rect -259 -3475 -213 -3437
rect -259 -3509 -253 -3475
rect -219 -3509 -213 -3475
rect -259 -3547 -213 -3509
rect -259 -3581 -253 -3547
rect -219 -3581 -213 -3547
rect -259 -3619 -213 -3581
rect -259 -3653 -253 -3619
rect -219 -3653 -213 -3619
rect -259 -3691 -213 -3653
rect -259 -3725 -253 -3691
rect -219 -3725 -213 -3691
rect -259 -3763 -213 -3725
rect -259 -3797 -253 -3763
rect -219 -3797 -213 -3763
rect -259 -3835 -213 -3797
rect -259 -3869 -253 -3835
rect -219 -3869 -213 -3835
rect -259 -3907 -213 -3869
rect -259 -3941 -253 -3907
rect -219 -3941 -213 -3907
rect -259 -3979 -213 -3941
rect -259 -4013 -253 -3979
rect -219 -4013 -213 -3979
rect -259 -4051 -213 -4013
rect -259 -4085 -253 -4051
rect -219 -4085 -213 -4051
rect -259 -4123 -213 -4085
rect -259 -4157 -253 -4123
rect -219 -4157 -213 -4123
rect -259 -4195 -213 -4157
rect -259 -4229 -253 -4195
rect -219 -4229 -213 -4195
rect -259 -4267 -213 -4229
rect -259 -4301 -253 -4267
rect -219 -4301 -213 -4267
rect -259 -4339 -213 -4301
rect -259 -4373 -253 -4339
rect -219 -4373 -213 -4339
rect -259 -4411 -213 -4373
rect -259 -4445 -253 -4411
rect -219 -4445 -213 -4411
rect -259 -4483 -213 -4445
rect -259 -4517 -253 -4483
rect -219 -4517 -213 -4483
rect -259 -4555 -213 -4517
rect -259 -4589 -253 -4555
rect -219 -4589 -213 -4555
rect -259 -4627 -213 -4589
rect -259 -4661 -253 -4627
rect -219 -4661 -213 -4627
rect -259 -4699 -213 -4661
rect -259 -4733 -253 -4699
rect -219 -4733 -213 -4699
rect -259 -4771 -213 -4733
rect -259 -4805 -253 -4771
rect -219 -4805 -213 -4771
rect -259 -4843 -213 -4805
rect -259 -4877 -253 -4843
rect -219 -4877 -213 -4843
rect -259 -4915 -213 -4877
rect -259 -4949 -253 -4915
rect -219 -4949 -213 -4915
rect -259 -4987 -213 -4949
rect -259 -5021 -253 -4987
rect -219 -5021 -213 -4987
rect -259 -5059 -213 -5021
rect -259 -5093 -253 -5059
rect -219 -5093 -213 -5059
rect -259 -5131 -213 -5093
rect -259 -5165 -253 -5131
rect -219 -5165 -213 -5131
rect -259 -5203 -213 -5165
rect -259 -5237 -253 -5203
rect -219 -5237 -213 -5203
rect -259 -5275 -213 -5237
rect -259 -5309 -253 -5275
rect -219 -5309 -213 -5275
rect -259 -5347 -213 -5309
rect -259 -5381 -253 -5347
rect -219 -5381 -213 -5347
rect -259 -5419 -213 -5381
rect -259 -5453 -253 -5419
rect -219 -5453 -213 -5419
rect -259 -5491 -213 -5453
rect -259 -5525 -253 -5491
rect -219 -5525 -213 -5491
rect -259 -5563 -213 -5525
rect -259 -5597 -253 -5563
rect -219 -5597 -213 -5563
rect -259 -5635 -213 -5597
rect -259 -5669 -253 -5635
rect -219 -5669 -213 -5635
rect -259 -5707 -213 -5669
rect -259 -5741 -253 -5707
rect -219 -5741 -213 -5707
rect -259 -5779 -213 -5741
rect -259 -5813 -253 -5779
rect -219 -5813 -213 -5779
rect -259 -5851 -213 -5813
rect -259 -5885 -253 -5851
rect -219 -5885 -213 -5851
rect -259 -5923 -213 -5885
rect -259 -5957 -253 -5923
rect -219 -5957 -213 -5923
rect -259 -6000 -213 -5957
rect -141 5957 -95 6000
rect -141 5923 -135 5957
rect -101 5923 -95 5957
rect -141 5885 -95 5923
rect -141 5851 -135 5885
rect -101 5851 -95 5885
rect -141 5813 -95 5851
rect -141 5779 -135 5813
rect -101 5779 -95 5813
rect -141 5741 -95 5779
rect -141 5707 -135 5741
rect -101 5707 -95 5741
rect -141 5669 -95 5707
rect -141 5635 -135 5669
rect -101 5635 -95 5669
rect -141 5597 -95 5635
rect -141 5563 -135 5597
rect -101 5563 -95 5597
rect -141 5525 -95 5563
rect -141 5491 -135 5525
rect -101 5491 -95 5525
rect -141 5453 -95 5491
rect -141 5419 -135 5453
rect -101 5419 -95 5453
rect -141 5381 -95 5419
rect -141 5347 -135 5381
rect -101 5347 -95 5381
rect -141 5309 -95 5347
rect -141 5275 -135 5309
rect -101 5275 -95 5309
rect -141 5237 -95 5275
rect -141 5203 -135 5237
rect -101 5203 -95 5237
rect -141 5165 -95 5203
rect -141 5131 -135 5165
rect -101 5131 -95 5165
rect -141 5093 -95 5131
rect -141 5059 -135 5093
rect -101 5059 -95 5093
rect -141 5021 -95 5059
rect -141 4987 -135 5021
rect -101 4987 -95 5021
rect -141 4949 -95 4987
rect -141 4915 -135 4949
rect -101 4915 -95 4949
rect -141 4877 -95 4915
rect -141 4843 -135 4877
rect -101 4843 -95 4877
rect -141 4805 -95 4843
rect -141 4771 -135 4805
rect -101 4771 -95 4805
rect -141 4733 -95 4771
rect -141 4699 -135 4733
rect -101 4699 -95 4733
rect -141 4661 -95 4699
rect -141 4627 -135 4661
rect -101 4627 -95 4661
rect -141 4589 -95 4627
rect -141 4555 -135 4589
rect -101 4555 -95 4589
rect -141 4517 -95 4555
rect -141 4483 -135 4517
rect -101 4483 -95 4517
rect -141 4445 -95 4483
rect -141 4411 -135 4445
rect -101 4411 -95 4445
rect -141 4373 -95 4411
rect -141 4339 -135 4373
rect -101 4339 -95 4373
rect -141 4301 -95 4339
rect -141 4267 -135 4301
rect -101 4267 -95 4301
rect -141 4229 -95 4267
rect -141 4195 -135 4229
rect -101 4195 -95 4229
rect -141 4157 -95 4195
rect -141 4123 -135 4157
rect -101 4123 -95 4157
rect -141 4085 -95 4123
rect -141 4051 -135 4085
rect -101 4051 -95 4085
rect -141 4013 -95 4051
rect -141 3979 -135 4013
rect -101 3979 -95 4013
rect -141 3941 -95 3979
rect -141 3907 -135 3941
rect -101 3907 -95 3941
rect -141 3869 -95 3907
rect -141 3835 -135 3869
rect -101 3835 -95 3869
rect -141 3797 -95 3835
rect -141 3763 -135 3797
rect -101 3763 -95 3797
rect -141 3725 -95 3763
rect -141 3691 -135 3725
rect -101 3691 -95 3725
rect -141 3653 -95 3691
rect -141 3619 -135 3653
rect -101 3619 -95 3653
rect -141 3581 -95 3619
rect -141 3547 -135 3581
rect -101 3547 -95 3581
rect -141 3509 -95 3547
rect -141 3475 -135 3509
rect -101 3475 -95 3509
rect -141 3437 -95 3475
rect -141 3403 -135 3437
rect -101 3403 -95 3437
rect -141 3365 -95 3403
rect -141 3331 -135 3365
rect -101 3331 -95 3365
rect -141 3293 -95 3331
rect -141 3259 -135 3293
rect -101 3259 -95 3293
rect -141 3221 -95 3259
rect -141 3187 -135 3221
rect -101 3187 -95 3221
rect -141 3149 -95 3187
rect -141 3115 -135 3149
rect -101 3115 -95 3149
rect -141 3077 -95 3115
rect -141 3043 -135 3077
rect -101 3043 -95 3077
rect -141 3005 -95 3043
rect -141 2971 -135 3005
rect -101 2971 -95 3005
rect -141 2933 -95 2971
rect -141 2899 -135 2933
rect -101 2899 -95 2933
rect -141 2861 -95 2899
rect -141 2827 -135 2861
rect -101 2827 -95 2861
rect -141 2789 -95 2827
rect -141 2755 -135 2789
rect -101 2755 -95 2789
rect -141 2717 -95 2755
rect -141 2683 -135 2717
rect -101 2683 -95 2717
rect -141 2645 -95 2683
rect -141 2611 -135 2645
rect -101 2611 -95 2645
rect -141 2573 -95 2611
rect -141 2539 -135 2573
rect -101 2539 -95 2573
rect -141 2501 -95 2539
rect -141 2467 -135 2501
rect -101 2467 -95 2501
rect -141 2429 -95 2467
rect -141 2395 -135 2429
rect -101 2395 -95 2429
rect -141 2357 -95 2395
rect -141 2323 -135 2357
rect -101 2323 -95 2357
rect -141 2285 -95 2323
rect -141 2251 -135 2285
rect -101 2251 -95 2285
rect -141 2213 -95 2251
rect -141 2179 -135 2213
rect -101 2179 -95 2213
rect -141 2141 -95 2179
rect -141 2107 -135 2141
rect -101 2107 -95 2141
rect -141 2069 -95 2107
rect -141 2035 -135 2069
rect -101 2035 -95 2069
rect -141 1997 -95 2035
rect -141 1963 -135 1997
rect -101 1963 -95 1997
rect -141 1925 -95 1963
rect -141 1891 -135 1925
rect -101 1891 -95 1925
rect -141 1853 -95 1891
rect -141 1819 -135 1853
rect -101 1819 -95 1853
rect -141 1781 -95 1819
rect -141 1747 -135 1781
rect -101 1747 -95 1781
rect -141 1709 -95 1747
rect -141 1675 -135 1709
rect -101 1675 -95 1709
rect -141 1637 -95 1675
rect -141 1603 -135 1637
rect -101 1603 -95 1637
rect -141 1565 -95 1603
rect -141 1531 -135 1565
rect -101 1531 -95 1565
rect -141 1493 -95 1531
rect -141 1459 -135 1493
rect -101 1459 -95 1493
rect -141 1421 -95 1459
rect -141 1387 -135 1421
rect -101 1387 -95 1421
rect -141 1349 -95 1387
rect -141 1315 -135 1349
rect -101 1315 -95 1349
rect -141 1277 -95 1315
rect -141 1243 -135 1277
rect -101 1243 -95 1277
rect -141 1205 -95 1243
rect -141 1171 -135 1205
rect -101 1171 -95 1205
rect -141 1133 -95 1171
rect -141 1099 -135 1133
rect -101 1099 -95 1133
rect -141 1061 -95 1099
rect -141 1027 -135 1061
rect -101 1027 -95 1061
rect -141 989 -95 1027
rect -141 955 -135 989
rect -101 955 -95 989
rect -141 917 -95 955
rect -141 883 -135 917
rect -101 883 -95 917
rect -141 845 -95 883
rect -141 811 -135 845
rect -101 811 -95 845
rect -141 773 -95 811
rect -141 739 -135 773
rect -101 739 -95 773
rect -141 701 -95 739
rect -141 667 -135 701
rect -101 667 -95 701
rect -141 629 -95 667
rect -141 595 -135 629
rect -101 595 -95 629
rect -141 557 -95 595
rect -141 523 -135 557
rect -101 523 -95 557
rect -141 485 -95 523
rect -141 451 -135 485
rect -101 451 -95 485
rect -141 413 -95 451
rect -141 379 -135 413
rect -101 379 -95 413
rect -141 341 -95 379
rect -141 307 -135 341
rect -101 307 -95 341
rect -141 269 -95 307
rect -141 235 -135 269
rect -101 235 -95 269
rect -141 197 -95 235
rect -141 163 -135 197
rect -101 163 -95 197
rect -141 125 -95 163
rect -141 91 -135 125
rect -101 91 -95 125
rect -141 53 -95 91
rect -141 19 -135 53
rect -101 19 -95 53
rect -141 -19 -95 19
rect -141 -53 -135 -19
rect -101 -53 -95 -19
rect -141 -91 -95 -53
rect -141 -125 -135 -91
rect -101 -125 -95 -91
rect -141 -163 -95 -125
rect -141 -197 -135 -163
rect -101 -197 -95 -163
rect -141 -235 -95 -197
rect -141 -269 -135 -235
rect -101 -269 -95 -235
rect -141 -307 -95 -269
rect -141 -341 -135 -307
rect -101 -341 -95 -307
rect -141 -379 -95 -341
rect -141 -413 -135 -379
rect -101 -413 -95 -379
rect -141 -451 -95 -413
rect -141 -485 -135 -451
rect -101 -485 -95 -451
rect -141 -523 -95 -485
rect -141 -557 -135 -523
rect -101 -557 -95 -523
rect -141 -595 -95 -557
rect -141 -629 -135 -595
rect -101 -629 -95 -595
rect -141 -667 -95 -629
rect -141 -701 -135 -667
rect -101 -701 -95 -667
rect -141 -739 -95 -701
rect -141 -773 -135 -739
rect -101 -773 -95 -739
rect -141 -811 -95 -773
rect -141 -845 -135 -811
rect -101 -845 -95 -811
rect -141 -883 -95 -845
rect -141 -917 -135 -883
rect -101 -917 -95 -883
rect -141 -955 -95 -917
rect -141 -989 -135 -955
rect -101 -989 -95 -955
rect -141 -1027 -95 -989
rect -141 -1061 -135 -1027
rect -101 -1061 -95 -1027
rect -141 -1099 -95 -1061
rect -141 -1133 -135 -1099
rect -101 -1133 -95 -1099
rect -141 -1171 -95 -1133
rect -141 -1205 -135 -1171
rect -101 -1205 -95 -1171
rect -141 -1243 -95 -1205
rect -141 -1277 -135 -1243
rect -101 -1277 -95 -1243
rect -141 -1315 -95 -1277
rect -141 -1349 -135 -1315
rect -101 -1349 -95 -1315
rect -141 -1387 -95 -1349
rect -141 -1421 -135 -1387
rect -101 -1421 -95 -1387
rect -141 -1459 -95 -1421
rect -141 -1493 -135 -1459
rect -101 -1493 -95 -1459
rect -141 -1531 -95 -1493
rect -141 -1565 -135 -1531
rect -101 -1565 -95 -1531
rect -141 -1603 -95 -1565
rect -141 -1637 -135 -1603
rect -101 -1637 -95 -1603
rect -141 -1675 -95 -1637
rect -141 -1709 -135 -1675
rect -101 -1709 -95 -1675
rect -141 -1747 -95 -1709
rect -141 -1781 -135 -1747
rect -101 -1781 -95 -1747
rect -141 -1819 -95 -1781
rect -141 -1853 -135 -1819
rect -101 -1853 -95 -1819
rect -141 -1891 -95 -1853
rect -141 -1925 -135 -1891
rect -101 -1925 -95 -1891
rect -141 -1963 -95 -1925
rect -141 -1997 -135 -1963
rect -101 -1997 -95 -1963
rect -141 -2035 -95 -1997
rect -141 -2069 -135 -2035
rect -101 -2069 -95 -2035
rect -141 -2107 -95 -2069
rect -141 -2141 -135 -2107
rect -101 -2141 -95 -2107
rect -141 -2179 -95 -2141
rect -141 -2213 -135 -2179
rect -101 -2213 -95 -2179
rect -141 -2251 -95 -2213
rect -141 -2285 -135 -2251
rect -101 -2285 -95 -2251
rect -141 -2323 -95 -2285
rect -141 -2357 -135 -2323
rect -101 -2357 -95 -2323
rect -141 -2395 -95 -2357
rect -141 -2429 -135 -2395
rect -101 -2429 -95 -2395
rect -141 -2467 -95 -2429
rect -141 -2501 -135 -2467
rect -101 -2501 -95 -2467
rect -141 -2539 -95 -2501
rect -141 -2573 -135 -2539
rect -101 -2573 -95 -2539
rect -141 -2611 -95 -2573
rect -141 -2645 -135 -2611
rect -101 -2645 -95 -2611
rect -141 -2683 -95 -2645
rect -141 -2717 -135 -2683
rect -101 -2717 -95 -2683
rect -141 -2755 -95 -2717
rect -141 -2789 -135 -2755
rect -101 -2789 -95 -2755
rect -141 -2827 -95 -2789
rect -141 -2861 -135 -2827
rect -101 -2861 -95 -2827
rect -141 -2899 -95 -2861
rect -141 -2933 -135 -2899
rect -101 -2933 -95 -2899
rect -141 -2971 -95 -2933
rect -141 -3005 -135 -2971
rect -101 -3005 -95 -2971
rect -141 -3043 -95 -3005
rect -141 -3077 -135 -3043
rect -101 -3077 -95 -3043
rect -141 -3115 -95 -3077
rect -141 -3149 -135 -3115
rect -101 -3149 -95 -3115
rect -141 -3187 -95 -3149
rect -141 -3221 -135 -3187
rect -101 -3221 -95 -3187
rect -141 -3259 -95 -3221
rect -141 -3293 -135 -3259
rect -101 -3293 -95 -3259
rect -141 -3331 -95 -3293
rect -141 -3365 -135 -3331
rect -101 -3365 -95 -3331
rect -141 -3403 -95 -3365
rect -141 -3437 -135 -3403
rect -101 -3437 -95 -3403
rect -141 -3475 -95 -3437
rect -141 -3509 -135 -3475
rect -101 -3509 -95 -3475
rect -141 -3547 -95 -3509
rect -141 -3581 -135 -3547
rect -101 -3581 -95 -3547
rect -141 -3619 -95 -3581
rect -141 -3653 -135 -3619
rect -101 -3653 -95 -3619
rect -141 -3691 -95 -3653
rect -141 -3725 -135 -3691
rect -101 -3725 -95 -3691
rect -141 -3763 -95 -3725
rect -141 -3797 -135 -3763
rect -101 -3797 -95 -3763
rect -141 -3835 -95 -3797
rect -141 -3869 -135 -3835
rect -101 -3869 -95 -3835
rect -141 -3907 -95 -3869
rect -141 -3941 -135 -3907
rect -101 -3941 -95 -3907
rect -141 -3979 -95 -3941
rect -141 -4013 -135 -3979
rect -101 -4013 -95 -3979
rect -141 -4051 -95 -4013
rect -141 -4085 -135 -4051
rect -101 -4085 -95 -4051
rect -141 -4123 -95 -4085
rect -141 -4157 -135 -4123
rect -101 -4157 -95 -4123
rect -141 -4195 -95 -4157
rect -141 -4229 -135 -4195
rect -101 -4229 -95 -4195
rect -141 -4267 -95 -4229
rect -141 -4301 -135 -4267
rect -101 -4301 -95 -4267
rect -141 -4339 -95 -4301
rect -141 -4373 -135 -4339
rect -101 -4373 -95 -4339
rect -141 -4411 -95 -4373
rect -141 -4445 -135 -4411
rect -101 -4445 -95 -4411
rect -141 -4483 -95 -4445
rect -141 -4517 -135 -4483
rect -101 -4517 -95 -4483
rect -141 -4555 -95 -4517
rect -141 -4589 -135 -4555
rect -101 -4589 -95 -4555
rect -141 -4627 -95 -4589
rect -141 -4661 -135 -4627
rect -101 -4661 -95 -4627
rect -141 -4699 -95 -4661
rect -141 -4733 -135 -4699
rect -101 -4733 -95 -4699
rect -141 -4771 -95 -4733
rect -141 -4805 -135 -4771
rect -101 -4805 -95 -4771
rect -141 -4843 -95 -4805
rect -141 -4877 -135 -4843
rect -101 -4877 -95 -4843
rect -141 -4915 -95 -4877
rect -141 -4949 -135 -4915
rect -101 -4949 -95 -4915
rect -141 -4987 -95 -4949
rect -141 -5021 -135 -4987
rect -101 -5021 -95 -4987
rect -141 -5059 -95 -5021
rect -141 -5093 -135 -5059
rect -101 -5093 -95 -5059
rect -141 -5131 -95 -5093
rect -141 -5165 -135 -5131
rect -101 -5165 -95 -5131
rect -141 -5203 -95 -5165
rect -141 -5237 -135 -5203
rect -101 -5237 -95 -5203
rect -141 -5275 -95 -5237
rect -141 -5309 -135 -5275
rect -101 -5309 -95 -5275
rect -141 -5347 -95 -5309
rect -141 -5381 -135 -5347
rect -101 -5381 -95 -5347
rect -141 -5419 -95 -5381
rect -141 -5453 -135 -5419
rect -101 -5453 -95 -5419
rect -141 -5491 -95 -5453
rect -141 -5525 -135 -5491
rect -101 -5525 -95 -5491
rect -141 -5563 -95 -5525
rect -141 -5597 -135 -5563
rect -101 -5597 -95 -5563
rect -141 -5635 -95 -5597
rect -141 -5669 -135 -5635
rect -101 -5669 -95 -5635
rect -141 -5707 -95 -5669
rect -141 -5741 -135 -5707
rect -101 -5741 -95 -5707
rect -141 -5779 -95 -5741
rect -141 -5813 -135 -5779
rect -101 -5813 -95 -5779
rect -141 -5851 -95 -5813
rect -141 -5885 -135 -5851
rect -101 -5885 -95 -5851
rect -141 -5923 -95 -5885
rect -141 -5957 -135 -5923
rect -101 -5957 -95 -5923
rect -141 -6000 -95 -5957
rect -23 5957 23 6000
rect -23 5923 -17 5957
rect 17 5923 23 5957
rect -23 5885 23 5923
rect -23 5851 -17 5885
rect 17 5851 23 5885
rect -23 5813 23 5851
rect -23 5779 -17 5813
rect 17 5779 23 5813
rect -23 5741 23 5779
rect -23 5707 -17 5741
rect 17 5707 23 5741
rect -23 5669 23 5707
rect -23 5635 -17 5669
rect 17 5635 23 5669
rect -23 5597 23 5635
rect -23 5563 -17 5597
rect 17 5563 23 5597
rect -23 5525 23 5563
rect -23 5491 -17 5525
rect 17 5491 23 5525
rect -23 5453 23 5491
rect -23 5419 -17 5453
rect 17 5419 23 5453
rect -23 5381 23 5419
rect -23 5347 -17 5381
rect 17 5347 23 5381
rect -23 5309 23 5347
rect -23 5275 -17 5309
rect 17 5275 23 5309
rect -23 5237 23 5275
rect -23 5203 -17 5237
rect 17 5203 23 5237
rect -23 5165 23 5203
rect -23 5131 -17 5165
rect 17 5131 23 5165
rect -23 5093 23 5131
rect -23 5059 -17 5093
rect 17 5059 23 5093
rect -23 5021 23 5059
rect -23 4987 -17 5021
rect 17 4987 23 5021
rect -23 4949 23 4987
rect -23 4915 -17 4949
rect 17 4915 23 4949
rect -23 4877 23 4915
rect -23 4843 -17 4877
rect 17 4843 23 4877
rect -23 4805 23 4843
rect -23 4771 -17 4805
rect 17 4771 23 4805
rect -23 4733 23 4771
rect -23 4699 -17 4733
rect 17 4699 23 4733
rect -23 4661 23 4699
rect -23 4627 -17 4661
rect 17 4627 23 4661
rect -23 4589 23 4627
rect -23 4555 -17 4589
rect 17 4555 23 4589
rect -23 4517 23 4555
rect -23 4483 -17 4517
rect 17 4483 23 4517
rect -23 4445 23 4483
rect -23 4411 -17 4445
rect 17 4411 23 4445
rect -23 4373 23 4411
rect -23 4339 -17 4373
rect 17 4339 23 4373
rect -23 4301 23 4339
rect -23 4267 -17 4301
rect 17 4267 23 4301
rect -23 4229 23 4267
rect -23 4195 -17 4229
rect 17 4195 23 4229
rect -23 4157 23 4195
rect -23 4123 -17 4157
rect 17 4123 23 4157
rect -23 4085 23 4123
rect -23 4051 -17 4085
rect 17 4051 23 4085
rect -23 4013 23 4051
rect -23 3979 -17 4013
rect 17 3979 23 4013
rect -23 3941 23 3979
rect -23 3907 -17 3941
rect 17 3907 23 3941
rect -23 3869 23 3907
rect -23 3835 -17 3869
rect 17 3835 23 3869
rect -23 3797 23 3835
rect -23 3763 -17 3797
rect 17 3763 23 3797
rect -23 3725 23 3763
rect -23 3691 -17 3725
rect 17 3691 23 3725
rect -23 3653 23 3691
rect -23 3619 -17 3653
rect 17 3619 23 3653
rect -23 3581 23 3619
rect -23 3547 -17 3581
rect 17 3547 23 3581
rect -23 3509 23 3547
rect -23 3475 -17 3509
rect 17 3475 23 3509
rect -23 3437 23 3475
rect -23 3403 -17 3437
rect 17 3403 23 3437
rect -23 3365 23 3403
rect -23 3331 -17 3365
rect 17 3331 23 3365
rect -23 3293 23 3331
rect -23 3259 -17 3293
rect 17 3259 23 3293
rect -23 3221 23 3259
rect -23 3187 -17 3221
rect 17 3187 23 3221
rect -23 3149 23 3187
rect -23 3115 -17 3149
rect 17 3115 23 3149
rect -23 3077 23 3115
rect -23 3043 -17 3077
rect 17 3043 23 3077
rect -23 3005 23 3043
rect -23 2971 -17 3005
rect 17 2971 23 3005
rect -23 2933 23 2971
rect -23 2899 -17 2933
rect 17 2899 23 2933
rect -23 2861 23 2899
rect -23 2827 -17 2861
rect 17 2827 23 2861
rect -23 2789 23 2827
rect -23 2755 -17 2789
rect 17 2755 23 2789
rect -23 2717 23 2755
rect -23 2683 -17 2717
rect 17 2683 23 2717
rect -23 2645 23 2683
rect -23 2611 -17 2645
rect 17 2611 23 2645
rect -23 2573 23 2611
rect -23 2539 -17 2573
rect 17 2539 23 2573
rect -23 2501 23 2539
rect -23 2467 -17 2501
rect 17 2467 23 2501
rect -23 2429 23 2467
rect -23 2395 -17 2429
rect 17 2395 23 2429
rect -23 2357 23 2395
rect -23 2323 -17 2357
rect 17 2323 23 2357
rect -23 2285 23 2323
rect -23 2251 -17 2285
rect 17 2251 23 2285
rect -23 2213 23 2251
rect -23 2179 -17 2213
rect 17 2179 23 2213
rect -23 2141 23 2179
rect -23 2107 -17 2141
rect 17 2107 23 2141
rect -23 2069 23 2107
rect -23 2035 -17 2069
rect 17 2035 23 2069
rect -23 1997 23 2035
rect -23 1963 -17 1997
rect 17 1963 23 1997
rect -23 1925 23 1963
rect -23 1891 -17 1925
rect 17 1891 23 1925
rect -23 1853 23 1891
rect -23 1819 -17 1853
rect 17 1819 23 1853
rect -23 1781 23 1819
rect -23 1747 -17 1781
rect 17 1747 23 1781
rect -23 1709 23 1747
rect -23 1675 -17 1709
rect 17 1675 23 1709
rect -23 1637 23 1675
rect -23 1603 -17 1637
rect 17 1603 23 1637
rect -23 1565 23 1603
rect -23 1531 -17 1565
rect 17 1531 23 1565
rect -23 1493 23 1531
rect -23 1459 -17 1493
rect 17 1459 23 1493
rect -23 1421 23 1459
rect -23 1387 -17 1421
rect 17 1387 23 1421
rect -23 1349 23 1387
rect -23 1315 -17 1349
rect 17 1315 23 1349
rect -23 1277 23 1315
rect -23 1243 -17 1277
rect 17 1243 23 1277
rect -23 1205 23 1243
rect -23 1171 -17 1205
rect 17 1171 23 1205
rect -23 1133 23 1171
rect -23 1099 -17 1133
rect 17 1099 23 1133
rect -23 1061 23 1099
rect -23 1027 -17 1061
rect 17 1027 23 1061
rect -23 989 23 1027
rect -23 955 -17 989
rect 17 955 23 989
rect -23 917 23 955
rect -23 883 -17 917
rect 17 883 23 917
rect -23 845 23 883
rect -23 811 -17 845
rect 17 811 23 845
rect -23 773 23 811
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -811 23 -773
rect -23 -845 -17 -811
rect 17 -845 23 -811
rect -23 -883 23 -845
rect -23 -917 -17 -883
rect 17 -917 23 -883
rect -23 -955 23 -917
rect -23 -989 -17 -955
rect 17 -989 23 -955
rect -23 -1027 23 -989
rect -23 -1061 -17 -1027
rect 17 -1061 23 -1027
rect -23 -1099 23 -1061
rect -23 -1133 -17 -1099
rect 17 -1133 23 -1099
rect -23 -1171 23 -1133
rect -23 -1205 -17 -1171
rect 17 -1205 23 -1171
rect -23 -1243 23 -1205
rect -23 -1277 -17 -1243
rect 17 -1277 23 -1243
rect -23 -1315 23 -1277
rect -23 -1349 -17 -1315
rect 17 -1349 23 -1315
rect -23 -1387 23 -1349
rect -23 -1421 -17 -1387
rect 17 -1421 23 -1387
rect -23 -1459 23 -1421
rect -23 -1493 -17 -1459
rect 17 -1493 23 -1459
rect -23 -1531 23 -1493
rect -23 -1565 -17 -1531
rect 17 -1565 23 -1531
rect -23 -1603 23 -1565
rect -23 -1637 -17 -1603
rect 17 -1637 23 -1603
rect -23 -1675 23 -1637
rect -23 -1709 -17 -1675
rect 17 -1709 23 -1675
rect -23 -1747 23 -1709
rect -23 -1781 -17 -1747
rect 17 -1781 23 -1747
rect -23 -1819 23 -1781
rect -23 -1853 -17 -1819
rect 17 -1853 23 -1819
rect -23 -1891 23 -1853
rect -23 -1925 -17 -1891
rect 17 -1925 23 -1891
rect -23 -1963 23 -1925
rect -23 -1997 -17 -1963
rect 17 -1997 23 -1963
rect -23 -2035 23 -1997
rect -23 -2069 -17 -2035
rect 17 -2069 23 -2035
rect -23 -2107 23 -2069
rect -23 -2141 -17 -2107
rect 17 -2141 23 -2107
rect -23 -2179 23 -2141
rect -23 -2213 -17 -2179
rect 17 -2213 23 -2179
rect -23 -2251 23 -2213
rect -23 -2285 -17 -2251
rect 17 -2285 23 -2251
rect -23 -2323 23 -2285
rect -23 -2357 -17 -2323
rect 17 -2357 23 -2323
rect -23 -2395 23 -2357
rect -23 -2429 -17 -2395
rect 17 -2429 23 -2395
rect -23 -2467 23 -2429
rect -23 -2501 -17 -2467
rect 17 -2501 23 -2467
rect -23 -2539 23 -2501
rect -23 -2573 -17 -2539
rect 17 -2573 23 -2539
rect -23 -2611 23 -2573
rect -23 -2645 -17 -2611
rect 17 -2645 23 -2611
rect -23 -2683 23 -2645
rect -23 -2717 -17 -2683
rect 17 -2717 23 -2683
rect -23 -2755 23 -2717
rect -23 -2789 -17 -2755
rect 17 -2789 23 -2755
rect -23 -2827 23 -2789
rect -23 -2861 -17 -2827
rect 17 -2861 23 -2827
rect -23 -2899 23 -2861
rect -23 -2933 -17 -2899
rect 17 -2933 23 -2899
rect -23 -2971 23 -2933
rect -23 -3005 -17 -2971
rect 17 -3005 23 -2971
rect -23 -3043 23 -3005
rect -23 -3077 -17 -3043
rect 17 -3077 23 -3043
rect -23 -3115 23 -3077
rect -23 -3149 -17 -3115
rect 17 -3149 23 -3115
rect -23 -3187 23 -3149
rect -23 -3221 -17 -3187
rect 17 -3221 23 -3187
rect -23 -3259 23 -3221
rect -23 -3293 -17 -3259
rect 17 -3293 23 -3259
rect -23 -3331 23 -3293
rect -23 -3365 -17 -3331
rect 17 -3365 23 -3331
rect -23 -3403 23 -3365
rect -23 -3437 -17 -3403
rect 17 -3437 23 -3403
rect -23 -3475 23 -3437
rect -23 -3509 -17 -3475
rect 17 -3509 23 -3475
rect -23 -3547 23 -3509
rect -23 -3581 -17 -3547
rect 17 -3581 23 -3547
rect -23 -3619 23 -3581
rect -23 -3653 -17 -3619
rect 17 -3653 23 -3619
rect -23 -3691 23 -3653
rect -23 -3725 -17 -3691
rect 17 -3725 23 -3691
rect -23 -3763 23 -3725
rect -23 -3797 -17 -3763
rect 17 -3797 23 -3763
rect -23 -3835 23 -3797
rect -23 -3869 -17 -3835
rect 17 -3869 23 -3835
rect -23 -3907 23 -3869
rect -23 -3941 -17 -3907
rect 17 -3941 23 -3907
rect -23 -3979 23 -3941
rect -23 -4013 -17 -3979
rect 17 -4013 23 -3979
rect -23 -4051 23 -4013
rect -23 -4085 -17 -4051
rect 17 -4085 23 -4051
rect -23 -4123 23 -4085
rect -23 -4157 -17 -4123
rect 17 -4157 23 -4123
rect -23 -4195 23 -4157
rect -23 -4229 -17 -4195
rect 17 -4229 23 -4195
rect -23 -4267 23 -4229
rect -23 -4301 -17 -4267
rect 17 -4301 23 -4267
rect -23 -4339 23 -4301
rect -23 -4373 -17 -4339
rect 17 -4373 23 -4339
rect -23 -4411 23 -4373
rect -23 -4445 -17 -4411
rect 17 -4445 23 -4411
rect -23 -4483 23 -4445
rect -23 -4517 -17 -4483
rect 17 -4517 23 -4483
rect -23 -4555 23 -4517
rect -23 -4589 -17 -4555
rect 17 -4589 23 -4555
rect -23 -4627 23 -4589
rect -23 -4661 -17 -4627
rect 17 -4661 23 -4627
rect -23 -4699 23 -4661
rect -23 -4733 -17 -4699
rect 17 -4733 23 -4699
rect -23 -4771 23 -4733
rect -23 -4805 -17 -4771
rect 17 -4805 23 -4771
rect -23 -4843 23 -4805
rect -23 -4877 -17 -4843
rect 17 -4877 23 -4843
rect -23 -4915 23 -4877
rect -23 -4949 -17 -4915
rect 17 -4949 23 -4915
rect -23 -4987 23 -4949
rect -23 -5021 -17 -4987
rect 17 -5021 23 -4987
rect -23 -5059 23 -5021
rect -23 -5093 -17 -5059
rect 17 -5093 23 -5059
rect -23 -5131 23 -5093
rect -23 -5165 -17 -5131
rect 17 -5165 23 -5131
rect -23 -5203 23 -5165
rect -23 -5237 -17 -5203
rect 17 -5237 23 -5203
rect -23 -5275 23 -5237
rect -23 -5309 -17 -5275
rect 17 -5309 23 -5275
rect -23 -5347 23 -5309
rect -23 -5381 -17 -5347
rect 17 -5381 23 -5347
rect -23 -5419 23 -5381
rect -23 -5453 -17 -5419
rect 17 -5453 23 -5419
rect -23 -5491 23 -5453
rect -23 -5525 -17 -5491
rect 17 -5525 23 -5491
rect -23 -5563 23 -5525
rect -23 -5597 -17 -5563
rect 17 -5597 23 -5563
rect -23 -5635 23 -5597
rect -23 -5669 -17 -5635
rect 17 -5669 23 -5635
rect -23 -5707 23 -5669
rect -23 -5741 -17 -5707
rect 17 -5741 23 -5707
rect -23 -5779 23 -5741
rect -23 -5813 -17 -5779
rect 17 -5813 23 -5779
rect -23 -5851 23 -5813
rect -23 -5885 -17 -5851
rect 17 -5885 23 -5851
rect -23 -5923 23 -5885
rect -23 -5957 -17 -5923
rect 17 -5957 23 -5923
rect -23 -6000 23 -5957
rect 95 5957 141 6000
rect 95 5923 101 5957
rect 135 5923 141 5957
rect 95 5885 141 5923
rect 95 5851 101 5885
rect 135 5851 141 5885
rect 95 5813 141 5851
rect 95 5779 101 5813
rect 135 5779 141 5813
rect 95 5741 141 5779
rect 95 5707 101 5741
rect 135 5707 141 5741
rect 95 5669 141 5707
rect 95 5635 101 5669
rect 135 5635 141 5669
rect 95 5597 141 5635
rect 95 5563 101 5597
rect 135 5563 141 5597
rect 95 5525 141 5563
rect 95 5491 101 5525
rect 135 5491 141 5525
rect 95 5453 141 5491
rect 95 5419 101 5453
rect 135 5419 141 5453
rect 95 5381 141 5419
rect 95 5347 101 5381
rect 135 5347 141 5381
rect 95 5309 141 5347
rect 95 5275 101 5309
rect 135 5275 141 5309
rect 95 5237 141 5275
rect 95 5203 101 5237
rect 135 5203 141 5237
rect 95 5165 141 5203
rect 95 5131 101 5165
rect 135 5131 141 5165
rect 95 5093 141 5131
rect 95 5059 101 5093
rect 135 5059 141 5093
rect 95 5021 141 5059
rect 95 4987 101 5021
rect 135 4987 141 5021
rect 95 4949 141 4987
rect 95 4915 101 4949
rect 135 4915 141 4949
rect 95 4877 141 4915
rect 95 4843 101 4877
rect 135 4843 141 4877
rect 95 4805 141 4843
rect 95 4771 101 4805
rect 135 4771 141 4805
rect 95 4733 141 4771
rect 95 4699 101 4733
rect 135 4699 141 4733
rect 95 4661 141 4699
rect 95 4627 101 4661
rect 135 4627 141 4661
rect 95 4589 141 4627
rect 95 4555 101 4589
rect 135 4555 141 4589
rect 95 4517 141 4555
rect 95 4483 101 4517
rect 135 4483 141 4517
rect 95 4445 141 4483
rect 95 4411 101 4445
rect 135 4411 141 4445
rect 95 4373 141 4411
rect 95 4339 101 4373
rect 135 4339 141 4373
rect 95 4301 141 4339
rect 95 4267 101 4301
rect 135 4267 141 4301
rect 95 4229 141 4267
rect 95 4195 101 4229
rect 135 4195 141 4229
rect 95 4157 141 4195
rect 95 4123 101 4157
rect 135 4123 141 4157
rect 95 4085 141 4123
rect 95 4051 101 4085
rect 135 4051 141 4085
rect 95 4013 141 4051
rect 95 3979 101 4013
rect 135 3979 141 4013
rect 95 3941 141 3979
rect 95 3907 101 3941
rect 135 3907 141 3941
rect 95 3869 141 3907
rect 95 3835 101 3869
rect 135 3835 141 3869
rect 95 3797 141 3835
rect 95 3763 101 3797
rect 135 3763 141 3797
rect 95 3725 141 3763
rect 95 3691 101 3725
rect 135 3691 141 3725
rect 95 3653 141 3691
rect 95 3619 101 3653
rect 135 3619 141 3653
rect 95 3581 141 3619
rect 95 3547 101 3581
rect 135 3547 141 3581
rect 95 3509 141 3547
rect 95 3475 101 3509
rect 135 3475 141 3509
rect 95 3437 141 3475
rect 95 3403 101 3437
rect 135 3403 141 3437
rect 95 3365 141 3403
rect 95 3331 101 3365
rect 135 3331 141 3365
rect 95 3293 141 3331
rect 95 3259 101 3293
rect 135 3259 141 3293
rect 95 3221 141 3259
rect 95 3187 101 3221
rect 135 3187 141 3221
rect 95 3149 141 3187
rect 95 3115 101 3149
rect 135 3115 141 3149
rect 95 3077 141 3115
rect 95 3043 101 3077
rect 135 3043 141 3077
rect 95 3005 141 3043
rect 95 2971 101 3005
rect 135 2971 141 3005
rect 95 2933 141 2971
rect 95 2899 101 2933
rect 135 2899 141 2933
rect 95 2861 141 2899
rect 95 2827 101 2861
rect 135 2827 141 2861
rect 95 2789 141 2827
rect 95 2755 101 2789
rect 135 2755 141 2789
rect 95 2717 141 2755
rect 95 2683 101 2717
rect 135 2683 141 2717
rect 95 2645 141 2683
rect 95 2611 101 2645
rect 135 2611 141 2645
rect 95 2573 141 2611
rect 95 2539 101 2573
rect 135 2539 141 2573
rect 95 2501 141 2539
rect 95 2467 101 2501
rect 135 2467 141 2501
rect 95 2429 141 2467
rect 95 2395 101 2429
rect 135 2395 141 2429
rect 95 2357 141 2395
rect 95 2323 101 2357
rect 135 2323 141 2357
rect 95 2285 141 2323
rect 95 2251 101 2285
rect 135 2251 141 2285
rect 95 2213 141 2251
rect 95 2179 101 2213
rect 135 2179 141 2213
rect 95 2141 141 2179
rect 95 2107 101 2141
rect 135 2107 141 2141
rect 95 2069 141 2107
rect 95 2035 101 2069
rect 135 2035 141 2069
rect 95 1997 141 2035
rect 95 1963 101 1997
rect 135 1963 141 1997
rect 95 1925 141 1963
rect 95 1891 101 1925
rect 135 1891 141 1925
rect 95 1853 141 1891
rect 95 1819 101 1853
rect 135 1819 141 1853
rect 95 1781 141 1819
rect 95 1747 101 1781
rect 135 1747 141 1781
rect 95 1709 141 1747
rect 95 1675 101 1709
rect 135 1675 141 1709
rect 95 1637 141 1675
rect 95 1603 101 1637
rect 135 1603 141 1637
rect 95 1565 141 1603
rect 95 1531 101 1565
rect 135 1531 141 1565
rect 95 1493 141 1531
rect 95 1459 101 1493
rect 135 1459 141 1493
rect 95 1421 141 1459
rect 95 1387 101 1421
rect 135 1387 141 1421
rect 95 1349 141 1387
rect 95 1315 101 1349
rect 135 1315 141 1349
rect 95 1277 141 1315
rect 95 1243 101 1277
rect 135 1243 141 1277
rect 95 1205 141 1243
rect 95 1171 101 1205
rect 135 1171 141 1205
rect 95 1133 141 1171
rect 95 1099 101 1133
rect 135 1099 141 1133
rect 95 1061 141 1099
rect 95 1027 101 1061
rect 135 1027 141 1061
rect 95 989 141 1027
rect 95 955 101 989
rect 135 955 141 989
rect 95 917 141 955
rect 95 883 101 917
rect 135 883 141 917
rect 95 845 141 883
rect 95 811 101 845
rect 135 811 141 845
rect 95 773 141 811
rect 95 739 101 773
rect 135 739 141 773
rect 95 701 141 739
rect 95 667 101 701
rect 135 667 141 701
rect 95 629 141 667
rect 95 595 101 629
rect 135 595 141 629
rect 95 557 141 595
rect 95 523 101 557
rect 135 523 141 557
rect 95 485 141 523
rect 95 451 101 485
rect 135 451 141 485
rect 95 413 141 451
rect 95 379 101 413
rect 135 379 141 413
rect 95 341 141 379
rect 95 307 101 341
rect 135 307 141 341
rect 95 269 141 307
rect 95 235 101 269
rect 135 235 141 269
rect 95 197 141 235
rect 95 163 101 197
rect 135 163 141 197
rect 95 125 141 163
rect 95 91 101 125
rect 135 91 141 125
rect 95 53 141 91
rect 95 19 101 53
rect 135 19 141 53
rect 95 -19 141 19
rect 95 -53 101 -19
rect 135 -53 141 -19
rect 95 -91 141 -53
rect 95 -125 101 -91
rect 135 -125 141 -91
rect 95 -163 141 -125
rect 95 -197 101 -163
rect 135 -197 141 -163
rect 95 -235 141 -197
rect 95 -269 101 -235
rect 135 -269 141 -235
rect 95 -307 141 -269
rect 95 -341 101 -307
rect 135 -341 141 -307
rect 95 -379 141 -341
rect 95 -413 101 -379
rect 135 -413 141 -379
rect 95 -451 141 -413
rect 95 -485 101 -451
rect 135 -485 141 -451
rect 95 -523 141 -485
rect 95 -557 101 -523
rect 135 -557 141 -523
rect 95 -595 141 -557
rect 95 -629 101 -595
rect 135 -629 141 -595
rect 95 -667 141 -629
rect 95 -701 101 -667
rect 135 -701 141 -667
rect 95 -739 141 -701
rect 95 -773 101 -739
rect 135 -773 141 -739
rect 95 -811 141 -773
rect 95 -845 101 -811
rect 135 -845 141 -811
rect 95 -883 141 -845
rect 95 -917 101 -883
rect 135 -917 141 -883
rect 95 -955 141 -917
rect 95 -989 101 -955
rect 135 -989 141 -955
rect 95 -1027 141 -989
rect 95 -1061 101 -1027
rect 135 -1061 141 -1027
rect 95 -1099 141 -1061
rect 95 -1133 101 -1099
rect 135 -1133 141 -1099
rect 95 -1171 141 -1133
rect 95 -1205 101 -1171
rect 135 -1205 141 -1171
rect 95 -1243 141 -1205
rect 95 -1277 101 -1243
rect 135 -1277 141 -1243
rect 95 -1315 141 -1277
rect 95 -1349 101 -1315
rect 135 -1349 141 -1315
rect 95 -1387 141 -1349
rect 95 -1421 101 -1387
rect 135 -1421 141 -1387
rect 95 -1459 141 -1421
rect 95 -1493 101 -1459
rect 135 -1493 141 -1459
rect 95 -1531 141 -1493
rect 95 -1565 101 -1531
rect 135 -1565 141 -1531
rect 95 -1603 141 -1565
rect 95 -1637 101 -1603
rect 135 -1637 141 -1603
rect 95 -1675 141 -1637
rect 95 -1709 101 -1675
rect 135 -1709 141 -1675
rect 95 -1747 141 -1709
rect 95 -1781 101 -1747
rect 135 -1781 141 -1747
rect 95 -1819 141 -1781
rect 95 -1853 101 -1819
rect 135 -1853 141 -1819
rect 95 -1891 141 -1853
rect 95 -1925 101 -1891
rect 135 -1925 141 -1891
rect 95 -1963 141 -1925
rect 95 -1997 101 -1963
rect 135 -1997 141 -1963
rect 95 -2035 141 -1997
rect 95 -2069 101 -2035
rect 135 -2069 141 -2035
rect 95 -2107 141 -2069
rect 95 -2141 101 -2107
rect 135 -2141 141 -2107
rect 95 -2179 141 -2141
rect 95 -2213 101 -2179
rect 135 -2213 141 -2179
rect 95 -2251 141 -2213
rect 95 -2285 101 -2251
rect 135 -2285 141 -2251
rect 95 -2323 141 -2285
rect 95 -2357 101 -2323
rect 135 -2357 141 -2323
rect 95 -2395 141 -2357
rect 95 -2429 101 -2395
rect 135 -2429 141 -2395
rect 95 -2467 141 -2429
rect 95 -2501 101 -2467
rect 135 -2501 141 -2467
rect 95 -2539 141 -2501
rect 95 -2573 101 -2539
rect 135 -2573 141 -2539
rect 95 -2611 141 -2573
rect 95 -2645 101 -2611
rect 135 -2645 141 -2611
rect 95 -2683 141 -2645
rect 95 -2717 101 -2683
rect 135 -2717 141 -2683
rect 95 -2755 141 -2717
rect 95 -2789 101 -2755
rect 135 -2789 141 -2755
rect 95 -2827 141 -2789
rect 95 -2861 101 -2827
rect 135 -2861 141 -2827
rect 95 -2899 141 -2861
rect 95 -2933 101 -2899
rect 135 -2933 141 -2899
rect 95 -2971 141 -2933
rect 95 -3005 101 -2971
rect 135 -3005 141 -2971
rect 95 -3043 141 -3005
rect 95 -3077 101 -3043
rect 135 -3077 141 -3043
rect 95 -3115 141 -3077
rect 95 -3149 101 -3115
rect 135 -3149 141 -3115
rect 95 -3187 141 -3149
rect 95 -3221 101 -3187
rect 135 -3221 141 -3187
rect 95 -3259 141 -3221
rect 95 -3293 101 -3259
rect 135 -3293 141 -3259
rect 95 -3331 141 -3293
rect 95 -3365 101 -3331
rect 135 -3365 141 -3331
rect 95 -3403 141 -3365
rect 95 -3437 101 -3403
rect 135 -3437 141 -3403
rect 95 -3475 141 -3437
rect 95 -3509 101 -3475
rect 135 -3509 141 -3475
rect 95 -3547 141 -3509
rect 95 -3581 101 -3547
rect 135 -3581 141 -3547
rect 95 -3619 141 -3581
rect 95 -3653 101 -3619
rect 135 -3653 141 -3619
rect 95 -3691 141 -3653
rect 95 -3725 101 -3691
rect 135 -3725 141 -3691
rect 95 -3763 141 -3725
rect 95 -3797 101 -3763
rect 135 -3797 141 -3763
rect 95 -3835 141 -3797
rect 95 -3869 101 -3835
rect 135 -3869 141 -3835
rect 95 -3907 141 -3869
rect 95 -3941 101 -3907
rect 135 -3941 141 -3907
rect 95 -3979 141 -3941
rect 95 -4013 101 -3979
rect 135 -4013 141 -3979
rect 95 -4051 141 -4013
rect 95 -4085 101 -4051
rect 135 -4085 141 -4051
rect 95 -4123 141 -4085
rect 95 -4157 101 -4123
rect 135 -4157 141 -4123
rect 95 -4195 141 -4157
rect 95 -4229 101 -4195
rect 135 -4229 141 -4195
rect 95 -4267 141 -4229
rect 95 -4301 101 -4267
rect 135 -4301 141 -4267
rect 95 -4339 141 -4301
rect 95 -4373 101 -4339
rect 135 -4373 141 -4339
rect 95 -4411 141 -4373
rect 95 -4445 101 -4411
rect 135 -4445 141 -4411
rect 95 -4483 141 -4445
rect 95 -4517 101 -4483
rect 135 -4517 141 -4483
rect 95 -4555 141 -4517
rect 95 -4589 101 -4555
rect 135 -4589 141 -4555
rect 95 -4627 141 -4589
rect 95 -4661 101 -4627
rect 135 -4661 141 -4627
rect 95 -4699 141 -4661
rect 95 -4733 101 -4699
rect 135 -4733 141 -4699
rect 95 -4771 141 -4733
rect 95 -4805 101 -4771
rect 135 -4805 141 -4771
rect 95 -4843 141 -4805
rect 95 -4877 101 -4843
rect 135 -4877 141 -4843
rect 95 -4915 141 -4877
rect 95 -4949 101 -4915
rect 135 -4949 141 -4915
rect 95 -4987 141 -4949
rect 95 -5021 101 -4987
rect 135 -5021 141 -4987
rect 95 -5059 141 -5021
rect 95 -5093 101 -5059
rect 135 -5093 141 -5059
rect 95 -5131 141 -5093
rect 95 -5165 101 -5131
rect 135 -5165 141 -5131
rect 95 -5203 141 -5165
rect 95 -5237 101 -5203
rect 135 -5237 141 -5203
rect 95 -5275 141 -5237
rect 95 -5309 101 -5275
rect 135 -5309 141 -5275
rect 95 -5347 141 -5309
rect 95 -5381 101 -5347
rect 135 -5381 141 -5347
rect 95 -5419 141 -5381
rect 95 -5453 101 -5419
rect 135 -5453 141 -5419
rect 95 -5491 141 -5453
rect 95 -5525 101 -5491
rect 135 -5525 141 -5491
rect 95 -5563 141 -5525
rect 95 -5597 101 -5563
rect 135 -5597 141 -5563
rect 95 -5635 141 -5597
rect 95 -5669 101 -5635
rect 135 -5669 141 -5635
rect 95 -5707 141 -5669
rect 95 -5741 101 -5707
rect 135 -5741 141 -5707
rect 95 -5779 141 -5741
rect 95 -5813 101 -5779
rect 135 -5813 141 -5779
rect 95 -5851 141 -5813
rect 95 -5885 101 -5851
rect 135 -5885 141 -5851
rect 95 -5923 141 -5885
rect 95 -5957 101 -5923
rect 135 -5957 141 -5923
rect 95 -6000 141 -5957
rect 213 5957 259 6000
rect 213 5923 219 5957
rect 253 5923 259 5957
rect 213 5885 259 5923
rect 213 5851 219 5885
rect 253 5851 259 5885
rect 213 5813 259 5851
rect 213 5779 219 5813
rect 253 5779 259 5813
rect 213 5741 259 5779
rect 213 5707 219 5741
rect 253 5707 259 5741
rect 213 5669 259 5707
rect 213 5635 219 5669
rect 253 5635 259 5669
rect 213 5597 259 5635
rect 213 5563 219 5597
rect 253 5563 259 5597
rect 213 5525 259 5563
rect 213 5491 219 5525
rect 253 5491 259 5525
rect 213 5453 259 5491
rect 213 5419 219 5453
rect 253 5419 259 5453
rect 213 5381 259 5419
rect 213 5347 219 5381
rect 253 5347 259 5381
rect 213 5309 259 5347
rect 213 5275 219 5309
rect 253 5275 259 5309
rect 213 5237 259 5275
rect 213 5203 219 5237
rect 253 5203 259 5237
rect 213 5165 259 5203
rect 213 5131 219 5165
rect 253 5131 259 5165
rect 213 5093 259 5131
rect 213 5059 219 5093
rect 253 5059 259 5093
rect 213 5021 259 5059
rect 213 4987 219 5021
rect 253 4987 259 5021
rect 213 4949 259 4987
rect 213 4915 219 4949
rect 253 4915 259 4949
rect 213 4877 259 4915
rect 213 4843 219 4877
rect 253 4843 259 4877
rect 213 4805 259 4843
rect 213 4771 219 4805
rect 253 4771 259 4805
rect 213 4733 259 4771
rect 213 4699 219 4733
rect 253 4699 259 4733
rect 213 4661 259 4699
rect 213 4627 219 4661
rect 253 4627 259 4661
rect 213 4589 259 4627
rect 213 4555 219 4589
rect 253 4555 259 4589
rect 213 4517 259 4555
rect 213 4483 219 4517
rect 253 4483 259 4517
rect 213 4445 259 4483
rect 213 4411 219 4445
rect 253 4411 259 4445
rect 213 4373 259 4411
rect 213 4339 219 4373
rect 253 4339 259 4373
rect 213 4301 259 4339
rect 213 4267 219 4301
rect 253 4267 259 4301
rect 213 4229 259 4267
rect 213 4195 219 4229
rect 253 4195 259 4229
rect 213 4157 259 4195
rect 213 4123 219 4157
rect 253 4123 259 4157
rect 213 4085 259 4123
rect 213 4051 219 4085
rect 253 4051 259 4085
rect 213 4013 259 4051
rect 213 3979 219 4013
rect 253 3979 259 4013
rect 213 3941 259 3979
rect 213 3907 219 3941
rect 253 3907 259 3941
rect 213 3869 259 3907
rect 213 3835 219 3869
rect 253 3835 259 3869
rect 213 3797 259 3835
rect 213 3763 219 3797
rect 253 3763 259 3797
rect 213 3725 259 3763
rect 213 3691 219 3725
rect 253 3691 259 3725
rect 213 3653 259 3691
rect 213 3619 219 3653
rect 253 3619 259 3653
rect 213 3581 259 3619
rect 213 3547 219 3581
rect 253 3547 259 3581
rect 213 3509 259 3547
rect 213 3475 219 3509
rect 253 3475 259 3509
rect 213 3437 259 3475
rect 213 3403 219 3437
rect 253 3403 259 3437
rect 213 3365 259 3403
rect 213 3331 219 3365
rect 253 3331 259 3365
rect 213 3293 259 3331
rect 213 3259 219 3293
rect 253 3259 259 3293
rect 213 3221 259 3259
rect 213 3187 219 3221
rect 253 3187 259 3221
rect 213 3149 259 3187
rect 213 3115 219 3149
rect 253 3115 259 3149
rect 213 3077 259 3115
rect 213 3043 219 3077
rect 253 3043 259 3077
rect 213 3005 259 3043
rect 213 2971 219 3005
rect 253 2971 259 3005
rect 213 2933 259 2971
rect 213 2899 219 2933
rect 253 2899 259 2933
rect 213 2861 259 2899
rect 213 2827 219 2861
rect 253 2827 259 2861
rect 213 2789 259 2827
rect 213 2755 219 2789
rect 253 2755 259 2789
rect 213 2717 259 2755
rect 213 2683 219 2717
rect 253 2683 259 2717
rect 213 2645 259 2683
rect 213 2611 219 2645
rect 253 2611 259 2645
rect 213 2573 259 2611
rect 213 2539 219 2573
rect 253 2539 259 2573
rect 213 2501 259 2539
rect 213 2467 219 2501
rect 253 2467 259 2501
rect 213 2429 259 2467
rect 213 2395 219 2429
rect 253 2395 259 2429
rect 213 2357 259 2395
rect 213 2323 219 2357
rect 253 2323 259 2357
rect 213 2285 259 2323
rect 213 2251 219 2285
rect 253 2251 259 2285
rect 213 2213 259 2251
rect 213 2179 219 2213
rect 253 2179 259 2213
rect 213 2141 259 2179
rect 213 2107 219 2141
rect 253 2107 259 2141
rect 213 2069 259 2107
rect 213 2035 219 2069
rect 253 2035 259 2069
rect 213 1997 259 2035
rect 213 1963 219 1997
rect 253 1963 259 1997
rect 213 1925 259 1963
rect 213 1891 219 1925
rect 253 1891 259 1925
rect 213 1853 259 1891
rect 213 1819 219 1853
rect 253 1819 259 1853
rect 213 1781 259 1819
rect 213 1747 219 1781
rect 253 1747 259 1781
rect 213 1709 259 1747
rect 213 1675 219 1709
rect 253 1675 259 1709
rect 213 1637 259 1675
rect 213 1603 219 1637
rect 253 1603 259 1637
rect 213 1565 259 1603
rect 213 1531 219 1565
rect 253 1531 259 1565
rect 213 1493 259 1531
rect 213 1459 219 1493
rect 253 1459 259 1493
rect 213 1421 259 1459
rect 213 1387 219 1421
rect 253 1387 259 1421
rect 213 1349 259 1387
rect 213 1315 219 1349
rect 253 1315 259 1349
rect 213 1277 259 1315
rect 213 1243 219 1277
rect 253 1243 259 1277
rect 213 1205 259 1243
rect 213 1171 219 1205
rect 253 1171 259 1205
rect 213 1133 259 1171
rect 213 1099 219 1133
rect 253 1099 259 1133
rect 213 1061 259 1099
rect 213 1027 219 1061
rect 253 1027 259 1061
rect 213 989 259 1027
rect 213 955 219 989
rect 253 955 259 989
rect 213 917 259 955
rect 213 883 219 917
rect 253 883 259 917
rect 213 845 259 883
rect 213 811 219 845
rect 253 811 259 845
rect 213 773 259 811
rect 213 739 219 773
rect 253 739 259 773
rect 213 701 259 739
rect 213 667 219 701
rect 253 667 259 701
rect 213 629 259 667
rect 213 595 219 629
rect 253 595 259 629
rect 213 557 259 595
rect 213 523 219 557
rect 253 523 259 557
rect 213 485 259 523
rect 213 451 219 485
rect 253 451 259 485
rect 213 413 259 451
rect 213 379 219 413
rect 253 379 259 413
rect 213 341 259 379
rect 213 307 219 341
rect 253 307 259 341
rect 213 269 259 307
rect 213 235 219 269
rect 253 235 259 269
rect 213 197 259 235
rect 213 163 219 197
rect 253 163 259 197
rect 213 125 259 163
rect 213 91 219 125
rect 253 91 259 125
rect 213 53 259 91
rect 213 19 219 53
rect 253 19 259 53
rect 213 -19 259 19
rect 213 -53 219 -19
rect 253 -53 259 -19
rect 213 -91 259 -53
rect 213 -125 219 -91
rect 253 -125 259 -91
rect 213 -163 259 -125
rect 213 -197 219 -163
rect 253 -197 259 -163
rect 213 -235 259 -197
rect 213 -269 219 -235
rect 253 -269 259 -235
rect 213 -307 259 -269
rect 213 -341 219 -307
rect 253 -341 259 -307
rect 213 -379 259 -341
rect 213 -413 219 -379
rect 253 -413 259 -379
rect 213 -451 259 -413
rect 213 -485 219 -451
rect 253 -485 259 -451
rect 213 -523 259 -485
rect 213 -557 219 -523
rect 253 -557 259 -523
rect 213 -595 259 -557
rect 213 -629 219 -595
rect 253 -629 259 -595
rect 213 -667 259 -629
rect 213 -701 219 -667
rect 253 -701 259 -667
rect 213 -739 259 -701
rect 213 -773 219 -739
rect 253 -773 259 -739
rect 213 -811 259 -773
rect 213 -845 219 -811
rect 253 -845 259 -811
rect 213 -883 259 -845
rect 213 -917 219 -883
rect 253 -917 259 -883
rect 213 -955 259 -917
rect 213 -989 219 -955
rect 253 -989 259 -955
rect 213 -1027 259 -989
rect 213 -1061 219 -1027
rect 253 -1061 259 -1027
rect 213 -1099 259 -1061
rect 213 -1133 219 -1099
rect 253 -1133 259 -1099
rect 213 -1171 259 -1133
rect 213 -1205 219 -1171
rect 253 -1205 259 -1171
rect 213 -1243 259 -1205
rect 213 -1277 219 -1243
rect 253 -1277 259 -1243
rect 213 -1315 259 -1277
rect 213 -1349 219 -1315
rect 253 -1349 259 -1315
rect 213 -1387 259 -1349
rect 213 -1421 219 -1387
rect 253 -1421 259 -1387
rect 213 -1459 259 -1421
rect 213 -1493 219 -1459
rect 253 -1493 259 -1459
rect 213 -1531 259 -1493
rect 213 -1565 219 -1531
rect 253 -1565 259 -1531
rect 213 -1603 259 -1565
rect 213 -1637 219 -1603
rect 253 -1637 259 -1603
rect 213 -1675 259 -1637
rect 213 -1709 219 -1675
rect 253 -1709 259 -1675
rect 213 -1747 259 -1709
rect 213 -1781 219 -1747
rect 253 -1781 259 -1747
rect 213 -1819 259 -1781
rect 213 -1853 219 -1819
rect 253 -1853 259 -1819
rect 213 -1891 259 -1853
rect 213 -1925 219 -1891
rect 253 -1925 259 -1891
rect 213 -1963 259 -1925
rect 213 -1997 219 -1963
rect 253 -1997 259 -1963
rect 213 -2035 259 -1997
rect 213 -2069 219 -2035
rect 253 -2069 259 -2035
rect 213 -2107 259 -2069
rect 213 -2141 219 -2107
rect 253 -2141 259 -2107
rect 213 -2179 259 -2141
rect 213 -2213 219 -2179
rect 253 -2213 259 -2179
rect 213 -2251 259 -2213
rect 213 -2285 219 -2251
rect 253 -2285 259 -2251
rect 213 -2323 259 -2285
rect 213 -2357 219 -2323
rect 253 -2357 259 -2323
rect 213 -2395 259 -2357
rect 213 -2429 219 -2395
rect 253 -2429 259 -2395
rect 213 -2467 259 -2429
rect 213 -2501 219 -2467
rect 253 -2501 259 -2467
rect 213 -2539 259 -2501
rect 213 -2573 219 -2539
rect 253 -2573 259 -2539
rect 213 -2611 259 -2573
rect 213 -2645 219 -2611
rect 253 -2645 259 -2611
rect 213 -2683 259 -2645
rect 213 -2717 219 -2683
rect 253 -2717 259 -2683
rect 213 -2755 259 -2717
rect 213 -2789 219 -2755
rect 253 -2789 259 -2755
rect 213 -2827 259 -2789
rect 213 -2861 219 -2827
rect 253 -2861 259 -2827
rect 213 -2899 259 -2861
rect 213 -2933 219 -2899
rect 253 -2933 259 -2899
rect 213 -2971 259 -2933
rect 213 -3005 219 -2971
rect 253 -3005 259 -2971
rect 213 -3043 259 -3005
rect 213 -3077 219 -3043
rect 253 -3077 259 -3043
rect 213 -3115 259 -3077
rect 213 -3149 219 -3115
rect 253 -3149 259 -3115
rect 213 -3187 259 -3149
rect 213 -3221 219 -3187
rect 253 -3221 259 -3187
rect 213 -3259 259 -3221
rect 213 -3293 219 -3259
rect 253 -3293 259 -3259
rect 213 -3331 259 -3293
rect 213 -3365 219 -3331
rect 253 -3365 259 -3331
rect 213 -3403 259 -3365
rect 213 -3437 219 -3403
rect 253 -3437 259 -3403
rect 213 -3475 259 -3437
rect 213 -3509 219 -3475
rect 253 -3509 259 -3475
rect 213 -3547 259 -3509
rect 213 -3581 219 -3547
rect 253 -3581 259 -3547
rect 213 -3619 259 -3581
rect 213 -3653 219 -3619
rect 253 -3653 259 -3619
rect 213 -3691 259 -3653
rect 213 -3725 219 -3691
rect 253 -3725 259 -3691
rect 213 -3763 259 -3725
rect 213 -3797 219 -3763
rect 253 -3797 259 -3763
rect 213 -3835 259 -3797
rect 213 -3869 219 -3835
rect 253 -3869 259 -3835
rect 213 -3907 259 -3869
rect 213 -3941 219 -3907
rect 253 -3941 259 -3907
rect 213 -3979 259 -3941
rect 213 -4013 219 -3979
rect 253 -4013 259 -3979
rect 213 -4051 259 -4013
rect 213 -4085 219 -4051
rect 253 -4085 259 -4051
rect 213 -4123 259 -4085
rect 213 -4157 219 -4123
rect 253 -4157 259 -4123
rect 213 -4195 259 -4157
rect 213 -4229 219 -4195
rect 253 -4229 259 -4195
rect 213 -4267 259 -4229
rect 213 -4301 219 -4267
rect 253 -4301 259 -4267
rect 213 -4339 259 -4301
rect 213 -4373 219 -4339
rect 253 -4373 259 -4339
rect 213 -4411 259 -4373
rect 213 -4445 219 -4411
rect 253 -4445 259 -4411
rect 213 -4483 259 -4445
rect 213 -4517 219 -4483
rect 253 -4517 259 -4483
rect 213 -4555 259 -4517
rect 213 -4589 219 -4555
rect 253 -4589 259 -4555
rect 213 -4627 259 -4589
rect 213 -4661 219 -4627
rect 253 -4661 259 -4627
rect 213 -4699 259 -4661
rect 213 -4733 219 -4699
rect 253 -4733 259 -4699
rect 213 -4771 259 -4733
rect 213 -4805 219 -4771
rect 253 -4805 259 -4771
rect 213 -4843 259 -4805
rect 213 -4877 219 -4843
rect 253 -4877 259 -4843
rect 213 -4915 259 -4877
rect 213 -4949 219 -4915
rect 253 -4949 259 -4915
rect 213 -4987 259 -4949
rect 213 -5021 219 -4987
rect 253 -5021 259 -4987
rect 213 -5059 259 -5021
rect 213 -5093 219 -5059
rect 253 -5093 259 -5059
rect 213 -5131 259 -5093
rect 213 -5165 219 -5131
rect 253 -5165 259 -5131
rect 213 -5203 259 -5165
rect 213 -5237 219 -5203
rect 253 -5237 259 -5203
rect 213 -5275 259 -5237
rect 213 -5309 219 -5275
rect 253 -5309 259 -5275
rect 213 -5347 259 -5309
rect 213 -5381 219 -5347
rect 253 -5381 259 -5347
rect 213 -5419 259 -5381
rect 213 -5453 219 -5419
rect 253 -5453 259 -5419
rect 213 -5491 259 -5453
rect 213 -5525 219 -5491
rect 253 -5525 259 -5491
rect 213 -5563 259 -5525
rect 213 -5597 219 -5563
rect 253 -5597 259 -5563
rect 213 -5635 259 -5597
rect 213 -5669 219 -5635
rect 253 -5669 259 -5635
rect 213 -5707 259 -5669
rect 213 -5741 219 -5707
rect 253 -5741 259 -5707
rect 213 -5779 259 -5741
rect 213 -5813 219 -5779
rect 253 -5813 259 -5779
rect 213 -5851 259 -5813
rect 213 -5885 219 -5851
rect 253 -5885 259 -5851
rect 213 -5923 259 -5885
rect 213 -5957 219 -5923
rect 253 -5957 259 -5923
rect 213 -6000 259 -5957
rect 331 5957 377 6000
rect 331 5923 337 5957
rect 371 5923 377 5957
rect 331 5885 377 5923
rect 331 5851 337 5885
rect 371 5851 377 5885
rect 331 5813 377 5851
rect 331 5779 337 5813
rect 371 5779 377 5813
rect 331 5741 377 5779
rect 331 5707 337 5741
rect 371 5707 377 5741
rect 331 5669 377 5707
rect 331 5635 337 5669
rect 371 5635 377 5669
rect 331 5597 377 5635
rect 331 5563 337 5597
rect 371 5563 377 5597
rect 331 5525 377 5563
rect 331 5491 337 5525
rect 371 5491 377 5525
rect 331 5453 377 5491
rect 331 5419 337 5453
rect 371 5419 377 5453
rect 331 5381 377 5419
rect 331 5347 337 5381
rect 371 5347 377 5381
rect 331 5309 377 5347
rect 331 5275 337 5309
rect 371 5275 377 5309
rect 331 5237 377 5275
rect 331 5203 337 5237
rect 371 5203 377 5237
rect 331 5165 377 5203
rect 331 5131 337 5165
rect 371 5131 377 5165
rect 331 5093 377 5131
rect 331 5059 337 5093
rect 371 5059 377 5093
rect 331 5021 377 5059
rect 331 4987 337 5021
rect 371 4987 377 5021
rect 331 4949 377 4987
rect 331 4915 337 4949
rect 371 4915 377 4949
rect 331 4877 377 4915
rect 331 4843 337 4877
rect 371 4843 377 4877
rect 331 4805 377 4843
rect 331 4771 337 4805
rect 371 4771 377 4805
rect 331 4733 377 4771
rect 331 4699 337 4733
rect 371 4699 377 4733
rect 331 4661 377 4699
rect 331 4627 337 4661
rect 371 4627 377 4661
rect 331 4589 377 4627
rect 331 4555 337 4589
rect 371 4555 377 4589
rect 331 4517 377 4555
rect 331 4483 337 4517
rect 371 4483 377 4517
rect 331 4445 377 4483
rect 331 4411 337 4445
rect 371 4411 377 4445
rect 331 4373 377 4411
rect 331 4339 337 4373
rect 371 4339 377 4373
rect 331 4301 377 4339
rect 331 4267 337 4301
rect 371 4267 377 4301
rect 331 4229 377 4267
rect 331 4195 337 4229
rect 371 4195 377 4229
rect 331 4157 377 4195
rect 331 4123 337 4157
rect 371 4123 377 4157
rect 331 4085 377 4123
rect 331 4051 337 4085
rect 371 4051 377 4085
rect 331 4013 377 4051
rect 331 3979 337 4013
rect 371 3979 377 4013
rect 331 3941 377 3979
rect 331 3907 337 3941
rect 371 3907 377 3941
rect 331 3869 377 3907
rect 331 3835 337 3869
rect 371 3835 377 3869
rect 331 3797 377 3835
rect 331 3763 337 3797
rect 371 3763 377 3797
rect 331 3725 377 3763
rect 331 3691 337 3725
rect 371 3691 377 3725
rect 331 3653 377 3691
rect 331 3619 337 3653
rect 371 3619 377 3653
rect 331 3581 377 3619
rect 331 3547 337 3581
rect 371 3547 377 3581
rect 331 3509 377 3547
rect 331 3475 337 3509
rect 371 3475 377 3509
rect 331 3437 377 3475
rect 331 3403 337 3437
rect 371 3403 377 3437
rect 331 3365 377 3403
rect 331 3331 337 3365
rect 371 3331 377 3365
rect 331 3293 377 3331
rect 331 3259 337 3293
rect 371 3259 377 3293
rect 331 3221 377 3259
rect 331 3187 337 3221
rect 371 3187 377 3221
rect 331 3149 377 3187
rect 331 3115 337 3149
rect 371 3115 377 3149
rect 331 3077 377 3115
rect 331 3043 337 3077
rect 371 3043 377 3077
rect 331 3005 377 3043
rect 331 2971 337 3005
rect 371 2971 377 3005
rect 331 2933 377 2971
rect 331 2899 337 2933
rect 371 2899 377 2933
rect 331 2861 377 2899
rect 331 2827 337 2861
rect 371 2827 377 2861
rect 331 2789 377 2827
rect 331 2755 337 2789
rect 371 2755 377 2789
rect 331 2717 377 2755
rect 331 2683 337 2717
rect 371 2683 377 2717
rect 331 2645 377 2683
rect 331 2611 337 2645
rect 371 2611 377 2645
rect 331 2573 377 2611
rect 331 2539 337 2573
rect 371 2539 377 2573
rect 331 2501 377 2539
rect 331 2467 337 2501
rect 371 2467 377 2501
rect 331 2429 377 2467
rect 331 2395 337 2429
rect 371 2395 377 2429
rect 331 2357 377 2395
rect 331 2323 337 2357
rect 371 2323 377 2357
rect 331 2285 377 2323
rect 331 2251 337 2285
rect 371 2251 377 2285
rect 331 2213 377 2251
rect 331 2179 337 2213
rect 371 2179 377 2213
rect 331 2141 377 2179
rect 331 2107 337 2141
rect 371 2107 377 2141
rect 331 2069 377 2107
rect 331 2035 337 2069
rect 371 2035 377 2069
rect 331 1997 377 2035
rect 331 1963 337 1997
rect 371 1963 377 1997
rect 331 1925 377 1963
rect 331 1891 337 1925
rect 371 1891 377 1925
rect 331 1853 377 1891
rect 331 1819 337 1853
rect 371 1819 377 1853
rect 331 1781 377 1819
rect 331 1747 337 1781
rect 371 1747 377 1781
rect 331 1709 377 1747
rect 331 1675 337 1709
rect 371 1675 377 1709
rect 331 1637 377 1675
rect 331 1603 337 1637
rect 371 1603 377 1637
rect 331 1565 377 1603
rect 331 1531 337 1565
rect 371 1531 377 1565
rect 331 1493 377 1531
rect 331 1459 337 1493
rect 371 1459 377 1493
rect 331 1421 377 1459
rect 331 1387 337 1421
rect 371 1387 377 1421
rect 331 1349 377 1387
rect 331 1315 337 1349
rect 371 1315 377 1349
rect 331 1277 377 1315
rect 331 1243 337 1277
rect 371 1243 377 1277
rect 331 1205 377 1243
rect 331 1171 337 1205
rect 371 1171 377 1205
rect 331 1133 377 1171
rect 331 1099 337 1133
rect 371 1099 377 1133
rect 331 1061 377 1099
rect 331 1027 337 1061
rect 371 1027 377 1061
rect 331 989 377 1027
rect 331 955 337 989
rect 371 955 377 989
rect 331 917 377 955
rect 331 883 337 917
rect 371 883 377 917
rect 331 845 377 883
rect 331 811 337 845
rect 371 811 377 845
rect 331 773 377 811
rect 331 739 337 773
rect 371 739 377 773
rect 331 701 377 739
rect 331 667 337 701
rect 371 667 377 701
rect 331 629 377 667
rect 331 595 337 629
rect 371 595 377 629
rect 331 557 377 595
rect 331 523 337 557
rect 371 523 377 557
rect 331 485 377 523
rect 331 451 337 485
rect 371 451 377 485
rect 331 413 377 451
rect 331 379 337 413
rect 371 379 377 413
rect 331 341 377 379
rect 331 307 337 341
rect 371 307 377 341
rect 331 269 377 307
rect 331 235 337 269
rect 371 235 377 269
rect 331 197 377 235
rect 331 163 337 197
rect 371 163 377 197
rect 331 125 377 163
rect 331 91 337 125
rect 371 91 377 125
rect 331 53 377 91
rect 331 19 337 53
rect 371 19 377 53
rect 331 -19 377 19
rect 331 -53 337 -19
rect 371 -53 377 -19
rect 331 -91 377 -53
rect 331 -125 337 -91
rect 371 -125 377 -91
rect 331 -163 377 -125
rect 331 -197 337 -163
rect 371 -197 377 -163
rect 331 -235 377 -197
rect 331 -269 337 -235
rect 371 -269 377 -235
rect 331 -307 377 -269
rect 331 -341 337 -307
rect 371 -341 377 -307
rect 331 -379 377 -341
rect 331 -413 337 -379
rect 371 -413 377 -379
rect 331 -451 377 -413
rect 331 -485 337 -451
rect 371 -485 377 -451
rect 331 -523 377 -485
rect 331 -557 337 -523
rect 371 -557 377 -523
rect 331 -595 377 -557
rect 331 -629 337 -595
rect 371 -629 377 -595
rect 331 -667 377 -629
rect 331 -701 337 -667
rect 371 -701 377 -667
rect 331 -739 377 -701
rect 331 -773 337 -739
rect 371 -773 377 -739
rect 331 -811 377 -773
rect 331 -845 337 -811
rect 371 -845 377 -811
rect 331 -883 377 -845
rect 331 -917 337 -883
rect 371 -917 377 -883
rect 331 -955 377 -917
rect 331 -989 337 -955
rect 371 -989 377 -955
rect 331 -1027 377 -989
rect 331 -1061 337 -1027
rect 371 -1061 377 -1027
rect 331 -1099 377 -1061
rect 331 -1133 337 -1099
rect 371 -1133 377 -1099
rect 331 -1171 377 -1133
rect 331 -1205 337 -1171
rect 371 -1205 377 -1171
rect 331 -1243 377 -1205
rect 331 -1277 337 -1243
rect 371 -1277 377 -1243
rect 331 -1315 377 -1277
rect 331 -1349 337 -1315
rect 371 -1349 377 -1315
rect 331 -1387 377 -1349
rect 331 -1421 337 -1387
rect 371 -1421 377 -1387
rect 331 -1459 377 -1421
rect 331 -1493 337 -1459
rect 371 -1493 377 -1459
rect 331 -1531 377 -1493
rect 331 -1565 337 -1531
rect 371 -1565 377 -1531
rect 331 -1603 377 -1565
rect 331 -1637 337 -1603
rect 371 -1637 377 -1603
rect 331 -1675 377 -1637
rect 331 -1709 337 -1675
rect 371 -1709 377 -1675
rect 331 -1747 377 -1709
rect 331 -1781 337 -1747
rect 371 -1781 377 -1747
rect 331 -1819 377 -1781
rect 331 -1853 337 -1819
rect 371 -1853 377 -1819
rect 331 -1891 377 -1853
rect 331 -1925 337 -1891
rect 371 -1925 377 -1891
rect 331 -1963 377 -1925
rect 331 -1997 337 -1963
rect 371 -1997 377 -1963
rect 331 -2035 377 -1997
rect 331 -2069 337 -2035
rect 371 -2069 377 -2035
rect 331 -2107 377 -2069
rect 331 -2141 337 -2107
rect 371 -2141 377 -2107
rect 331 -2179 377 -2141
rect 331 -2213 337 -2179
rect 371 -2213 377 -2179
rect 331 -2251 377 -2213
rect 331 -2285 337 -2251
rect 371 -2285 377 -2251
rect 331 -2323 377 -2285
rect 331 -2357 337 -2323
rect 371 -2357 377 -2323
rect 331 -2395 377 -2357
rect 331 -2429 337 -2395
rect 371 -2429 377 -2395
rect 331 -2467 377 -2429
rect 331 -2501 337 -2467
rect 371 -2501 377 -2467
rect 331 -2539 377 -2501
rect 331 -2573 337 -2539
rect 371 -2573 377 -2539
rect 331 -2611 377 -2573
rect 331 -2645 337 -2611
rect 371 -2645 377 -2611
rect 331 -2683 377 -2645
rect 331 -2717 337 -2683
rect 371 -2717 377 -2683
rect 331 -2755 377 -2717
rect 331 -2789 337 -2755
rect 371 -2789 377 -2755
rect 331 -2827 377 -2789
rect 331 -2861 337 -2827
rect 371 -2861 377 -2827
rect 331 -2899 377 -2861
rect 331 -2933 337 -2899
rect 371 -2933 377 -2899
rect 331 -2971 377 -2933
rect 331 -3005 337 -2971
rect 371 -3005 377 -2971
rect 331 -3043 377 -3005
rect 331 -3077 337 -3043
rect 371 -3077 377 -3043
rect 331 -3115 377 -3077
rect 331 -3149 337 -3115
rect 371 -3149 377 -3115
rect 331 -3187 377 -3149
rect 331 -3221 337 -3187
rect 371 -3221 377 -3187
rect 331 -3259 377 -3221
rect 331 -3293 337 -3259
rect 371 -3293 377 -3259
rect 331 -3331 377 -3293
rect 331 -3365 337 -3331
rect 371 -3365 377 -3331
rect 331 -3403 377 -3365
rect 331 -3437 337 -3403
rect 371 -3437 377 -3403
rect 331 -3475 377 -3437
rect 331 -3509 337 -3475
rect 371 -3509 377 -3475
rect 331 -3547 377 -3509
rect 331 -3581 337 -3547
rect 371 -3581 377 -3547
rect 331 -3619 377 -3581
rect 331 -3653 337 -3619
rect 371 -3653 377 -3619
rect 331 -3691 377 -3653
rect 331 -3725 337 -3691
rect 371 -3725 377 -3691
rect 331 -3763 377 -3725
rect 331 -3797 337 -3763
rect 371 -3797 377 -3763
rect 331 -3835 377 -3797
rect 331 -3869 337 -3835
rect 371 -3869 377 -3835
rect 331 -3907 377 -3869
rect 331 -3941 337 -3907
rect 371 -3941 377 -3907
rect 331 -3979 377 -3941
rect 331 -4013 337 -3979
rect 371 -4013 377 -3979
rect 331 -4051 377 -4013
rect 331 -4085 337 -4051
rect 371 -4085 377 -4051
rect 331 -4123 377 -4085
rect 331 -4157 337 -4123
rect 371 -4157 377 -4123
rect 331 -4195 377 -4157
rect 331 -4229 337 -4195
rect 371 -4229 377 -4195
rect 331 -4267 377 -4229
rect 331 -4301 337 -4267
rect 371 -4301 377 -4267
rect 331 -4339 377 -4301
rect 331 -4373 337 -4339
rect 371 -4373 377 -4339
rect 331 -4411 377 -4373
rect 331 -4445 337 -4411
rect 371 -4445 377 -4411
rect 331 -4483 377 -4445
rect 331 -4517 337 -4483
rect 371 -4517 377 -4483
rect 331 -4555 377 -4517
rect 331 -4589 337 -4555
rect 371 -4589 377 -4555
rect 331 -4627 377 -4589
rect 331 -4661 337 -4627
rect 371 -4661 377 -4627
rect 331 -4699 377 -4661
rect 331 -4733 337 -4699
rect 371 -4733 377 -4699
rect 331 -4771 377 -4733
rect 331 -4805 337 -4771
rect 371 -4805 377 -4771
rect 331 -4843 377 -4805
rect 331 -4877 337 -4843
rect 371 -4877 377 -4843
rect 331 -4915 377 -4877
rect 331 -4949 337 -4915
rect 371 -4949 377 -4915
rect 331 -4987 377 -4949
rect 331 -5021 337 -4987
rect 371 -5021 377 -4987
rect 331 -5059 377 -5021
rect 331 -5093 337 -5059
rect 371 -5093 377 -5059
rect 331 -5131 377 -5093
rect 331 -5165 337 -5131
rect 371 -5165 377 -5131
rect 331 -5203 377 -5165
rect 331 -5237 337 -5203
rect 371 -5237 377 -5203
rect 331 -5275 377 -5237
rect 331 -5309 337 -5275
rect 371 -5309 377 -5275
rect 331 -5347 377 -5309
rect 331 -5381 337 -5347
rect 371 -5381 377 -5347
rect 331 -5419 377 -5381
rect 331 -5453 337 -5419
rect 371 -5453 377 -5419
rect 331 -5491 377 -5453
rect 331 -5525 337 -5491
rect 371 -5525 377 -5491
rect 331 -5563 377 -5525
rect 331 -5597 337 -5563
rect 371 -5597 377 -5563
rect 331 -5635 377 -5597
rect 331 -5669 337 -5635
rect 371 -5669 377 -5635
rect 331 -5707 377 -5669
rect 331 -5741 337 -5707
rect 371 -5741 377 -5707
rect 331 -5779 377 -5741
rect 331 -5813 337 -5779
rect 371 -5813 377 -5779
rect 331 -5851 377 -5813
rect 331 -5885 337 -5851
rect 371 -5885 377 -5851
rect 331 -5923 377 -5885
rect 331 -5957 337 -5923
rect 371 -5957 377 -5923
rect 331 -6000 377 -5957
rect 449 5957 495 6000
rect 449 5923 455 5957
rect 489 5923 495 5957
rect 449 5885 495 5923
rect 449 5851 455 5885
rect 489 5851 495 5885
rect 449 5813 495 5851
rect 449 5779 455 5813
rect 489 5779 495 5813
rect 449 5741 495 5779
rect 449 5707 455 5741
rect 489 5707 495 5741
rect 449 5669 495 5707
rect 449 5635 455 5669
rect 489 5635 495 5669
rect 449 5597 495 5635
rect 449 5563 455 5597
rect 489 5563 495 5597
rect 449 5525 495 5563
rect 449 5491 455 5525
rect 489 5491 495 5525
rect 449 5453 495 5491
rect 449 5419 455 5453
rect 489 5419 495 5453
rect 449 5381 495 5419
rect 449 5347 455 5381
rect 489 5347 495 5381
rect 449 5309 495 5347
rect 449 5275 455 5309
rect 489 5275 495 5309
rect 449 5237 495 5275
rect 449 5203 455 5237
rect 489 5203 495 5237
rect 449 5165 495 5203
rect 449 5131 455 5165
rect 489 5131 495 5165
rect 449 5093 495 5131
rect 449 5059 455 5093
rect 489 5059 495 5093
rect 449 5021 495 5059
rect 449 4987 455 5021
rect 489 4987 495 5021
rect 449 4949 495 4987
rect 449 4915 455 4949
rect 489 4915 495 4949
rect 449 4877 495 4915
rect 449 4843 455 4877
rect 489 4843 495 4877
rect 449 4805 495 4843
rect 449 4771 455 4805
rect 489 4771 495 4805
rect 449 4733 495 4771
rect 449 4699 455 4733
rect 489 4699 495 4733
rect 449 4661 495 4699
rect 449 4627 455 4661
rect 489 4627 495 4661
rect 449 4589 495 4627
rect 449 4555 455 4589
rect 489 4555 495 4589
rect 449 4517 495 4555
rect 449 4483 455 4517
rect 489 4483 495 4517
rect 449 4445 495 4483
rect 449 4411 455 4445
rect 489 4411 495 4445
rect 449 4373 495 4411
rect 449 4339 455 4373
rect 489 4339 495 4373
rect 449 4301 495 4339
rect 449 4267 455 4301
rect 489 4267 495 4301
rect 449 4229 495 4267
rect 449 4195 455 4229
rect 489 4195 495 4229
rect 449 4157 495 4195
rect 449 4123 455 4157
rect 489 4123 495 4157
rect 449 4085 495 4123
rect 449 4051 455 4085
rect 489 4051 495 4085
rect 449 4013 495 4051
rect 449 3979 455 4013
rect 489 3979 495 4013
rect 449 3941 495 3979
rect 449 3907 455 3941
rect 489 3907 495 3941
rect 449 3869 495 3907
rect 449 3835 455 3869
rect 489 3835 495 3869
rect 449 3797 495 3835
rect 449 3763 455 3797
rect 489 3763 495 3797
rect 449 3725 495 3763
rect 449 3691 455 3725
rect 489 3691 495 3725
rect 449 3653 495 3691
rect 449 3619 455 3653
rect 489 3619 495 3653
rect 449 3581 495 3619
rect 449 3547 455 3581
rect 489 3547 495 3581
rect 449 3509 495 3547
rect 449 3475 455 3509
rect 489 3475 495 3509
rect 449 3437 495 3475
rect 449 3403 455 3437
rect 489 3403 495 3437
rect 449 3365 495 3403
rect 449 3331 455 3365
rect 489 3331 495 3365
rect 449 3293 495 3331
rect 449 3259 455 3293
rect 489 3259 495 3293
rect 449 3221 495 3259
rect 449 3187 455 3221
rect 489 3187 495 3221
rect 449 3149 495 3187
rect 449 3115 455 3149
rect 489 3115 495 3149
rect 449 3077 495 3115
rect 449 3043 455 3077
rect 489 3043 495 3077
rect 449 3005 495 3043
rect 449 2971 455 3005
rect 489 2971 495 3005
rect 449 2933 495 2971
rect 449 2899 455 2933
rect 489 2899 495 2933
rect 449 2861 495 2899
rect 449 2827 455 2861
rect 489 2827 495 2861
rect 449 2789 495 2827
rect 449 2755 455 2789
rect 489 2755 495 2789
rect 449 2717 495 2755
rect 449 2683 455 2717
rect 489 2683 495 2717
rect 449 2645 495 2683
rect 449 2611 455 2645
rect 489 2611 495 2645
rect 449 2573 495 2611
rect 449 2539 455 2573
rect 489 2539 495 2573
rect 449 2501 495 2539
rect 449 2467 455 2501
rect 489 2467 495 2501
rect 449 2429 495 2467
rect 449 2395 455 2429
rect 489 2395 495 2429
rect 449 2357 495 2395
rect 449 2323 455 2357
rect 489 2323 495 2357
rect 449 2285 495 2323
rect 449 2251 455 2285
rect 489 2251 495 2285
rect 449 2213 495 2251
rect 449 2179 455 2213
rect 489 2179 495 2213
rect 449 2141 495 2179
rect 449 2107 455 2141
rect 489 2107 495 2141
rect 449 2069 495 2107
rect 449 2035 455 2069
rect 489 2035 495 2069
rect 449 1997 495 2035
rect 449 1963 455 1997
rect 489 1963 495 1997
rect 449 1925 495 1963
rect 449 1891 455 1925
rect 489 1891 495 1925
rect 449 1853 495 1891
rect 449 1819 455 1853
rect 489 1819 495 1853
rect 449 1781 495 1819
rect 449 1747 455 1781
rect 489 1747 495 1781
rect 449 1709 495 1747
rect 449 1675 455 1709
rect 489 1675 495 1709
rect 449 1637 495 1675
rect 449 1603 455 1637
rect 489 1603 495 1637
rect 449 1565 495 1603
rect 449 1531 455 1565
rect 489 1531 495 1565
rect 449 1493 495 1531
rect 449 1459 455 1493
rect 489 1459 495 1493
rect 449 1421 495 1459
rect 449 1387 455 1421
rect 489 1387 495 1421
rect 449 1349 495 1387
rect 449 1315 455 1349
rect 489 1315 495 1349
rect 449 1277 495 1315
rect 449 1243 455 1277
rect 489 1243 495 1277
rect 449 1205 495 1243
rect 449 1171 455 1205
rect 489 1171 495 1205
rect 449 1133 495 1171
rect 449 1099 455 1133
rect 489 1099 495 1133
rect 449 1061 495 1099
rect 449 1027 455 1061
rect 489 1027 495 1061
rect 449 989 495 1027
rect 449 955 455 989
rect 489 955 495 989
rect 449 917 495 955
rect 449 883 455 917
rect 489 883 495 917
rect 449 845 495 883
rect 449 811 455 845
rect 489 811 495 845
rect 449 773 495 811
rect 449 739 455 773
rect 489 739 495 773
rect 449 701 495 739
rect 449 667 455 701
rect 489 667 495 701
rect 449 629 495 667
rect 449 595 455 629
rect 489 595 495 629
rect 449 557 495 595
rect 449 523 455 557
rect 489 523 495 557
rect 449 485 495 523
rect 449 451 455 485
rect 489 451 495 485
rect 449 413 495 451
rect 449 379 455 413
rect 489 379 495 413
rect 449 341 495 379
rect 449 307 455 341
rect 489 307 495 341
rect 449 269 495 307
rect 449 235 455 269
rect 489 235 495 269
rect 449 197 495 235
rect 449 163 455 197
rect 489 163 495 197
rect 449 125 495 163
rect 449 91 455 125
rect 489 91 495 125
rect 449 53 495 91
rect 449 19 455 53
rect 489 19 495 53
rect 449 -19 495 19
rect 449 -53 455 -19
rect 489 -53 495 -19
rect 449 -91 495 -53
rect 449 -125 455 -91
rect 489 -125 495 -91
rect 449 -163 495 -125
rect 449 -197 455 -163
rect 489 -197 495 -163
rect 449 -235 495 -197
rect 449 -269 455 -235
rect 489 -269 495 -235
rect 449 -307 495 -269
rect 449 -341 455 -307
rect 489 -341 495 -307
rect 449 -379 495 -341
rect 449 -413 455 -379
rect 489 -413 495 -379
rect 449 -451 495 -413
rect 449 -485 455 -451
rect 489 -485 495 -451
rect 449 -523 495 -485
rect 449 -557 455 -523
rect 489 -557 495 -523
rect 449 -595 495 -557
rect 449 -629 455 -595
rect 489 -629 495 -595
rect 449 -667 495 -629
rect 449 -701 455 -667
rect 489 -701 495 -667
rect 449 -739 495 -701
rect 449 -773 455 -739
rect 489 -773 495 -739
rect 449 -811 495 -773
rect 449 -845 455 -811
rect 489 -845 495 -811
rect 449 -883 495 -845
rect 449 -917 455 -883
rect 489 -917 495 -883
rect 449 -955 495 -917
rect 449 -989 455 -955
rect 489 -989 495 -955
rect 449 -1027 495 -989
rect 449 -1061 455 -1027
rect 489 -1061 495 -1027
rect 449 -1099 495 -1061
rect 449 -1133 455 -1099
rect 489 -1133 495 -1099
rect 449 -1171 495 -1133
rect 449 -1205 455 -1171
rect 489 -1205 495 -1171
rect 449 -1243 495 -1205
rect 449 -1277 455 -1243
rect 489 -1277 495 -1243
rect 449 -1315 495 -1277
rect 449 -1349 455 -1315
rect 489 -1349 495 -1315
rect 449 -1387 495 -1349
rect 449 -1421 455 -1387
rect 489 -1421 495 -1387
rect 449 -1459 495 -1421
rect 449 -1493 455 -1459
rect 489 -1493 495 -1459
rect 449 -1531 495 -1493
rect 449 -1565 455 -1531
rect 489 -1565 495 -1531
rect 449 -1603 495 -1565
rect 449 -1637 455 -1603
rect 489 -1637 495 -1603
rect 449 -1675 495 -1637
rect 449 -1709 455 -1675
rect 489 -1709 495 -1675
rect 449 -1747 495 -1709
rect 449 -1781 455 -1747
rect 489 -1781 495 -1747
rect 449 -1819 495 -1781
rect 449 -1853 455 -1819
rect 489 -1853 495 -1819
rect 449 -1891 495 -1853
rect 449 -1925 455 -1891
rect 489 -1925 495 -1891
rect 449 -1963 495 -1925
rect 449 -1997 455 -1963
rect 489 -1997 495 -1963
rect 449 -2035 495 -1997
rect 449 -2069 455 -2035
rect 489 -2069 495 -2035
rect 449 -2107 495 -2069
rect 449 -2141 455 -2107
rect 489 -2141 495 -2107
rect 449 -2179 495 -2141
rect 449 -2213 455 -2179
rect 489 -2213 495 -2179
rect 449 -2251 495 -2213
rect 449 -2285 455 -2251
rect 489 -2285 495 -2251
rect 449 -2323 495 -2285
rect 449 -2357 455 -2323
rect 489 -2357 495 -2323
rect 449 -2395 495 -2357
rect 449 -2429 455 -2395
rect 489 -2429 495 -2395
rect 449 -2467 495 -2429
rect 449 -2501 455 -2467
rect 489 -2501 495 -2467
rect 449 -2539 495 -2501
rect 449 -2573 455 -2539
rect 489 -2573 495 -2539
rect 449 -2611 495 -2573
rect 449 -2645 455 -2611
rect 489 -2645 495 -2611
rect 449 -2683 495 -2645
rect 449 -2717 455 -2683
rect 489 -2717 495 -2683
rect 449 -2755 495 -2717
rect 449 -2789 455 -2755
rect 489 -2789 495 -2755
rect 449 -2827 495 -2789
rect 449 -2861 455 -2827
rect 489 -2861 495 -2827
rect 449 -2899 495 -2861
rect 449 -2933 455 -2899
rect 489 -2933 495 -2899
rect 449 -2971 495 -2933
rect 449 -3005 455 -2971
rect 489 -3005 495 -2971
rect 449 -3043 495 -3005
rect 449 -3077 455 -3043
rect 489 -3077 495 -3043
rect 449 -3115 495 -3077
rect 449 -3149 455 -3115
rect 489 -3149 495 -3115
rect 449 -3187 495 -3149
rect 449 -3221 455 -3187
rect 489 -3221 495 -3187
rect 449 -3259 495 -3221
rect 449 -3293 455 -3259
rect 489 -3293 495 -3259
rect 449 -3331 495 -3293
rect 449 -3365 455 -3331
rect 489 -3365 495 -3331
rect 449 -3403 495 -3365
rect 449 -3437 455 -3403
rect 489 -3437 495 -3403
rect 449 -3475 495 -3437
rect 449 -3509 455 -3475
rect 489 -3509 495 -3475
rect 449 -3547 495 -3509
rect 449 -3581 455 -3547
rect 489 -3581 495 -3547
rect 449 -3619 495 -3581
rect 449 -3653 455 -3619
rect 489 -3653 495 -3619
rect 449 -3691 495 -3653
rect 449 -3725 455 -3691
rect 489 -3725 495 -3691
rect 449 -3763 495 -3725
rect 449 -3797 455 -3763
rect 489 -3797 495 -3763
rect 449 -3835 495 -3797
rect 449 -3869 455 -3835
rect 489 -3869 495 -3835
rect 449 -3907 495 -3869
rect 449 -3941 455 -3907
rect 489 -3941 495 -3907
rect 449 -3979 495 -3941
rect 449 -4013 455 -3979
rect 489 -4013 495 -3979
rect 449 -4051 495 -4013
rect 449 -4085 455 -4051
rect 489 -4085 495 -4051
rect 449 -4123 495 -4085
rect 449 -4157 455 -4123
rect 489 -4157 495 -4123
rect 449 -4195 495 -4157
rect 449 -4229 455 -4195
rect 489 -4229 495 -4195
rect 449 -4267 495 -4229
rect 449 -4301 455 -4267
rect 489 -4301 495 -4267
rect 449 -4339 495 -4301
rect 449 -4373 455 -4339
rect 489 -4373 495 -4339
rect 449 -4411 495 -4373
rect 449 -4445 455 -4411
rect 489 -4445 495 -4411
rect 449 -4483 495 -4445
rect 449 -4517 455 -4483
rect 489 -4517 495 -4483
rect 449 -4555 495 -4517
rect 449 -4589 455 -4555
rect 489 -4589 495 -4555
rect 449 -4627 495 -4589
rect 449 -4661 455 -4627
rect 489 -4661 495 -4627
rect 449 -4699 495 -4661
rect 449 -4733 455 -4699
rect 489 -4733 495 -4699
rect 449 -4771 495 -4733
rect 449 -4805 455 -4771
rect 489 -4805 495 -4771
rect 449 -4843 495 -4805
rect 449 -4877 455 -4843
rect 489 -4877 495 -4843
rect 449 -4915 495 -4877
rect 449 -4949 455 -4915
rect 489 -4949 495 -4915
rect 449 -4987 495 -4949
rect 449 -5021 455 -4987
rect 489 -5021 495 -4987
rect 449 -5059 495 -5021
rect 449 -5093 455 -5059
rect 489 -5093 495 -5059
rect 449 -5131 495 -5093
rect 449 -5165 455 -5131
rect 489 -5165 495 -5131
rect 449 -5203 495 -5165
rect 449 -5237 455 -5203
rect 489 -5237 495 -5203
rect 449 -5275 495 -5237
rect 449 -5309 455 -5275
rect 489 -5309 495 -5275
rect 449 -5347 495 -5309
rect 449 -5381 455 -5347
rect 489 -5381 495 -5347
rect 449 -5419 495 -5381
rect 449 -5453 455 -5419
rect 489 -5453 495 -5419
rect 449 -5491 495 -5453
rect 449 -5525 455 -5491
rect 489 -5525 495 -5491
rect 449 -5563 495 -5525
rect 449 -5597 455 -5563
rect 489 -5597 495 -5563
rect 449 -5635 495 -5597
rect 449 -5669 455 -5635
rect 489 -5669 495 -5635
rect 449 -5707 495 -5669
rect 449 -5741 455 -5707
rect 489 -5741 495 -5707
rect 449 -5779 495 -5741
rect 449 -5813 455 -5779
rect 489 -5813 495 -5779
rect 449 -5851 495 -5813
rect 449 -5885 455 -5851
rect 489 -5885 495 -5851
rect 449 -5923 495 -5885
rect 449 -5957 455 -5923
rect 489 -5957 495 -5923
rect 449 -6000 495 -5957
rect 567 5957 613 6000
rect 567 5923 573 5957
rect 607 5923 613 5957
rect 567 5885 613 5923
rect 567 5851 573 5885
rect 607 5851 613 5885
rect 567 5813 613 5851
rect 567 5779 573 5813
rect 607 5779 613 5813
rect 567 5741 613 5779
rect 567 5707 573 5741
rect 607 5707 613 5741
rect 567 5669 613 5707
rect 567 5635 573 5669
rect 607 5635 613 5669
rect 567 5597 613 5635
rect 567 5563 573 5597
rect 607 5563 613 5597
rect 567 5525 613 5563
rect 567 5491 573 5525
rect 607 5491 613 5525
rect 567 5453 613 5491
rect 567 5419 573 5453
rect 607 5419 613 5453
rect 567 5381 613 5419
rect 567 5347 573 5381
rect 607 5347 613 5381
rect 567 5309 613 5347
rect 567 5275 573 5309
rect 607 5275 613 5309
rect 567 5237 613 5275
rect 567 5203 573 5237
rect 607 5203 613 5237
rect 567 5165 613 5203
rect 567 5131 573 5165
rect 607 5131 613 5165
rect 567 5093 613 5131
rect 567 5059 573 5093
rect 607 5059 613 5093
rect 567 5021 613 5059
rect 567 4987 573 5021
rect 607 4987 613 5021
rect 567 4949 613 4987
rect 567 4915 573 4949
rect 607 4915 613 4949
rect 567 4877 613 4915
rect 567 4843 573 4877
rect 607 4843 613 4877
rect 567 4805 613 4843
rect 567 4771 573 4805
rect 607 4771 613 4805
rect 567 4733 613 4771
rect 567 4699 573 4733
rect 607 4699 613 4733
rect 567 4661 613 4699
rect 567 4627 573 4661
rect 607 4627 613 4661
rect 567 4589 613 4627
rect 567 4555 573 4589
rect 607 4555 613 4589
rect 567 4517 613 4555
rect 567 4483 573 4517
rect 607 4483 613 4517
rect 567 4445 613 4483
rect 567 4411 573 4445
rect 607 4411 613 4445
rect 567 4373 613 4411
rect 567 4339 573 4373
rect 607 4339 613 4373
rect 567 4301 613 4339
rect 567 4267 573 4301
rect 607 4267 613 4301
rect 567 4229 613 4267
rect 567 4195 573 4229
rect 607 4195 613 4229
rect 567 4157 613 4195
rect 567 4123 573 4157
rect 607 4123 613 4157
rect 567 4085 613 4123
rect 567 4051 573 4085
rect 607 4051 613 4085
rect 567 4013 613 4051
rect 567 3979 573 4013
rect 607 3979 613 4013
rect 567 3941 613 3979
rect 567 3907 573 3941
rect 607 3907 613 3941
rect 567 3869 613 3907
rect 567 3835 573 3869
rect 607 3835 613 3869
rect 567 3797 613 3835
rect 567 3763 573 3797
rect 607 3763 613 3797
rect 567 3725 613 3763
rect 567 3691 573 3725
rect 607 3691 613 3725
rect 567 3653 613 3691
rect 567 3619 573 3653
rect 607 3619 613 3653
rect 567 3581 613 3619
rect 567 3547 573 3581
rect 607 3547 613 3581
rect 567 3509 613 3547
rect 567 3475 573 3509
rect 607 3475 613 3509
rect 567 3437 613 3475
rect 567 3403 573 3437
rect 607 3403 613 3437
rect 567 3365 613 3403
rect 567 3331 573 3365
rect 607 3331 613 3365
rect 567 3293 613 3331
rect 567 3259 573 3293
rect 607 3259 613 3293
rect 567 3221 613 3259
rect 567 3187 573 3221
rect 607 3187 613 3221
rect 567 3149 613 3187
rect 567 3115 573 3149
rect 607 3115 613 3149
rect 567 3077 613 3115
rect 567 3043 573 3077
rect 607 3043 613 3077
rect 567 3005 613 3043
rect 567 2971 573 3005
rect 607 2971 613 3005
rect 567 2933 613 2971
rect 567 2899 573 2933
rect 607 2899 613 2933
rect 567 2861 613 2899
rect 567 2827 573 2861
rect 607 2827 613 2861
rect 567 2789 613 2827
rect 567 2755 573 2789
rect 607 2755 613 2789
rect 567 2717 613 2755
rect 567 2683 573 2717
rect 607 2683 613 2717
rect 567 2645 613 2683
rect 567 2611 573 2645
rect 607 2611 613 2645
rect 567 2573 613 2611
rect 567 2539 573 2573
rect 607 2539 613 2573
rect 567 2501 613 2539
rect 567 2467 573 2501
rect 607 2467 613 2501
rect 567 2429 613 2467
rect 567 2395 573 2429
rect 607 2395 613 2429
rect 567 2357 613 2395
rect 567 2323 573 2357
rect 607 2323 613 2357
rect 567 2285 613 2323
rect 567 2251 573 2285
rect 607 2251 613 2285
rect 567 2213 613 2251
rect 567 2179 573 2213
rect 607 2179 613 2213
rect 567 2141 613 2179
rect 567 2107 573 2141
rect 607 2107 613 2141
rect 567 2069 613 2107
rect 567 2035 573 2069
rect 607 2035 613 2069
rect 567 1997 613 2035
rect 567 1963 573 1997
rect 607 1963 613 1997
rect 567 1925 613 1963
rect 567 1891 573 1925
rect 607 1891 613 1925
rect 567 1853 613 1891
rect 567 1819 573 1853
rect 607 1819 613 1853
rect 567 1781 613 1819
rect 567 1747 573 1781
rect 607 1747 613 1781
rect 567 1709 613 1747
rect 567 1675 573 1709
rect 607 1675 613 1709
rect 567 1637 613 1675
rect 567 1603 573 1637
rect 607 1603 613 1637
rect 567 1565 613 1603
rect 567 1531 573 1565
rect 607 1531 613 1565
rect 567 1493 613 1531
rect 567 1459 573 1493
rect 607 1459 613 1493
rect 567 1421 613 1459
rect 567 1387 573 1421
rect 607 1387 613 1421
rect 567 1349 613 1387
rect 567 1315 573 1349
rect 607 1315 613 1349
rect 567 1277 613 1315
rect 567 1243 573 1277
rect 607 1243 613 1277
rect 567 1205 613 1243
rect 567 1171 573 1205
rect 607 1171 613 1205
rect 567 1133 613 1171
rect 567 1099 573 1133
rect 607 1099 613 1133
rect 567 1061 613 1099
rect 567 1027 573 1061
rect 607 1027 613 1061
rect 567 989 613 1027
rect 567 955 573 989
rect 607 955 613 989
rect 567 917 613 955
rect 567 883 573 917
rect 607 883 613 917
rect 567 845 613 883
rect 567 811 573 845
rect 607 811 613 845
rect 567 773 613 811
rect 567 739 573 773
rect 607 739 613 773
rect 567 701 613 739
rect 567 667 573 701
rect 607 667 613 701
rect 567 629 613 667
rect 567 595 573 629
rect 607 595 613 629
rect 567 557 613 595
rect 567 523 573 557
rect 607 523 613 557
rect 567 485 613 523
rect 567 451 573 485
rect 607 451 613 485
rect 567 413 613 451
rect 567 379 573 413
rect 607 379 613 413
rect 567 341 613 379
rect 567 307 573 341
rect 607 307 613 341
rect 567 269 613 307
rect 567 235 573 269
rect 607 235 613 269
rect 567 197 613 235
rect 567 163 573 197
rect 607 163 613 197
rect 567 125 613 163
rect 567 91 573 125
rect 607 91 613 125
rect 567 53 613 91
rect 567 19 573 53
rect 607 19 613 53
rect 567 -19 613 19
rect 567 -53 573 -19
rect 607 -53 613 -19
rect 567 -91 613 -53
rect 567 -125 573 -91
rect 607 -125 613 -91
rect 567 -163 613 -125
rect 567 -197 573 -163
rect 607 -197 613 -163
rect 567 -235 613 -197
rect 567 -269 573 -235
rect 607 -269 613 -235
rect 567 -307 613 -269
rect 567 -341 573 -307
rect 607 -341 613 -307
rect 567 -379 613 -341
rect 567 -413 573 -379
rect 607 -413 613 -379
rect 567 -451 613 -413
rect 567 -485 573 -451
rect 607 -485 613 -451
rect 567 -523 613 -485
rect 567 -557 573 -523
rect 607 -557 613 -523
rect 567 -595 613 -557
rect 567 -629 573 -595
rect 607 -629 613 -595
rect 567 -667 613 -629
rect 567 -701 573 -667
rect 607 -701 613 -667
rect 567 -739 613 -701
rect 567 -773 573 -739
rect 607 -773 613 -739
rect 567 -811 613 -773
rect 567 -845 573 -811
rect 607 -845 613 -811
rect 567 -883 613 -845
rect 567 -917 573 -883
rect 607 -917 613 -883
rect 567 -955 613 -917
rect 567 -989 573 -955
rect 607 -989 613 -955
rect 567 -1027 613 -989
rect 567 -1061 573 -1027
rect 607 -1061 613 -1027
rect 567 -1099 613 -1061
rect 567 -1133 573 -1099
rect 607 -1133 613 -1099
rect 567 -1171 613 -1133
rect 567 -1205 573 -1171
rect 607 -1205 613 -1171
rect 567 -1243 613 -1205
rect 567 -1277 573 -1243
rect 607 -1277 613 -1243
rect 567 -1315 613 -1277
rect 567 -1349 573 -1315
rect 607 -1349 613 -1315
rect 567 -1387 613 -1349
rect 567 -1421 573 -1387
rect 607 -1421 613 -1387
rect 567 -1459 613 -1421
rect 567 -1493 573 -1459
rect 607 -1493 613 -1459
rect 567 -1531 613 -1493
rect 567 -1565 573 -1531
rect 607 -1565 613 -1531
rect 567 -1603 613 -1565
rect 567 -1637 573 -1603
rect 607 -1637 613 -1603
rect 567 -1675 613 -1637
rect 567 -1709 573 -1675
rect 607 -1709 613 -1675
rect 567 -1747 613 -1709
rect 567 -1781 573 -1747
rect 607 -1781 613 -1747
rect 567 -1819 613 -1781
rect 567 -1853 573 -1819
rect 607 -1853 613 -1819
rect 567 -1891 613 -1853
rect 567 -1925 573 -1891
rect 607 -1925 613 -1891
rect 567 -1963 613 -1925
rect 567 -1997 573 -1963
rect 607 -1997 613 -1963
rect 567 -2035 613 -1997
rect 567 -2069 573 -2035
rect 607 -2069 613 -2035
rect 567 -2107 613 -2069
rect 567 -2141 573 -2107
rect 607 -2141 613 -2107
rect 567 -2179 613 -2141
rect 567 -2213 573 -2179
rect 607 -2213 613 -2179
rect 567 -2251 613 -2213
rect 567 -2285 573 -2251
rect 607 -2285 613 -2251
rect 567 -2323 613 -2285
rect 567 -2357 573 -2323
rect 607 -2357 613 -2323
rect 567 -2395 613 -2357
rect 567 -2429 573 -2395
rect 607 -2429 613 -2395
rect 567 -2467 613 -2429
rect 567 -2501 573 -2467
rect 607 -2501 613 -2467
rect 567 -2539 613 -2501
rect 567 -2573 573 -2539
rect 607 -2573 613 -2539
rect 567 -2611 613 -2573
rect 567 -2645 573 -2611
rect 607 -2645 613 -2611
rect 567 -2683 613 -2645
rect 567 -2717 573 -2683
rect 607 -2717 613 -2683
rect 567 -2755 613 -2717
rect 567 -2789 573 -2755
rect 607 -2789 613 -2755
rect 567 -2827 613 -2789
rect 567 -2861 573 -2827
rect 607 -2861 613 -2827
rect 567 -2899 613 -2861
rect 567 -2933 573 -2899
rect 607 -2933 613 -2899
rect 567 -2971 613 -2933
rect 567 -3005 573 -2971
rect 607 -3005 613 -2971
rect 567 -3043 613 -3005
rect 567 -3077 573 -3043
rect 607 -3077 613 -3043
rect 567 -3115 613 -3077
rect 567 -3149 573 -3115
rect 607 -3149 613 -3115
rect 567 -3187 613 -3149
rect 567 -3221 573 -3187
rect 607 -3221 613 -3187
rect 567 -3259 613 -3221
rect 567 -3293 573 -3259
rect 607 -3293 613 -3259
rect 567 -3331 613 -3293
rect 567 -3365 573 -3331
rect 607 -3365 613 -3331
rect 567 -3403 613 -3365
rect 567 -3437 573 -3403
rect 607 -3437 613 -3403
rect 567 -3475 613 -3437
rect 567 -3509 573 -3475
rect 607 -3509 613 -3475
rect 567 -3547 613 -3509
rect 567 -3581 573 -3547
rect 607 -3581 613 -3547
rect 567 -3619 613 -3581
rect 567 -3653 573 -3619
rect 607 -3653 613 -3619
rect 567 -3691 613 -3653
rect 567 -3725 573 -3691
rect 607 -3725 613 -3691
rect 567 -3763 613 -3725
rect 567 -3797 573 -3763
rect 607 -3797 613 -3763
rect 567 -3835 613 -3797
rect 567 -3869 573 -3835
rect 607 -3869 613 -3835
rect 567 -3907 613 -3869
rect 567 -3941 573 -3907
rect 607 -3941 613 -3907
rect 567 -3979 613 -3941
rect 567 -4013 573 -3979
rect 607 -4013 613 -3979
rect 567 -4051 613 -4013
rect 567 -4085 573 -4051
rect 607 -4085 613 -4051
rect 567 -4123 613 -4085
rect 567 -4157 573 -4123
rect 607 -4157 613 -4123
rect 567 -4195 613 -4157
rect 567 -4229 573 -4195
rect 607 -4229 613 -4195
rect 567 -4267 613 -4229
rect 567 -4301 573 -4267
rect 607 -4301 613 -4267
rect 567 -4339 613 -4301
rect 567 -4373 573 -4339
rect 607 -4373 613 -4339
rect 567 -4411 613 -4373
rect 567 -4445 573 -4411
rect 607 -4445 613 -4411
rect 567 -4483 613 -4445
rect 567 -4517 573 -4483
rect 607 -4517 613 -4483
rect 567 -4555 613 -4517
rect 567 -4589 573 -4555
rect 607 -4589 613 -4555
rect 567 -4627 613 -4589
rect 567 -4661 573 -4627
rect 607 -4661 613 -4627
rect 567 -4699 613 -4661
rect 567 -4733 573 -4699
rect 607 -4733 613 -4699
rect 567 -4771 613 -4733
rect 567 -4805 573 -4771
rect 607 -4805 613 -4771
rect 567 -4843 613 -4805
rect 567 -4877 573 -4843
rect 607 -4877 613 -4843
rect 567 -4915 613 -4877
rect 567 -4949 573 -4915
rect 607 -4949 613 -4915
rect 567 -4987 613 -4949
rect 567 -5021 573 -4987
rect 607 -5021 613 -4987
rect 567 -5059 613 -5021
rect 567 -5093 573 -5059
rect 607 -5093 613 -5059
rect 567 -5131 613 -5093
rect 567 -5165 573 -5131
rect 607 -5165 613 -5131
rect 567 -5203 613 -5165
rect 567 -5237 573 -5203
rect 607 -5237 613 -5203
rect 567 -5275 613 -5237
rect 567 -5309 573 -5275
rect 607 -5309 613 -5275
rect 567 -5347 613 -5309
rect 567 -5381 573 -5347
rect 607 -5381 613 -5347
rect 567 -5419 613 -5381
rect 567 -5453 573 -5419
rect 607 -5453 613 -5419
rect 567 -5491 613 -5453
rect 567 -5525 573 -5491
rect 607 -5525 613 -5491
rect 567 -5563 613 -5525
rect 567 -5597 573 -5563
rect 607 -5597 613 -5563
rect 567 -5635 613 -5597
rect 567 -5669 573 -5635
rect 607 -5669 613 -5635
rect 567 -5707 613 -5669
rect 567 -5741 573 -5707
rect 607 -5741 613 -5707
rect 567 -5779 613 -5741
rect 567 -5813 573 -5779
rect 607 -5813 613 -5779
rect 567 -5851 613 -5813
rect 567 -5885 573 -5851
rect 607 -5885 613 -5851
rect 567 -5923 613 -5885
rect 567 -5957 573 -5923
rect 607 -5957 613 -5923
rect 567 -6000 613 -5957
<< end >>
