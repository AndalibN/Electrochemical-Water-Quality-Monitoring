magic
tech sky130A
magscale 1 2
timestamp 1665001199
<< nmos >>
rect -200 109 200 2109
rect -200 -2109 200 -109
<< ndiff >>
rect -258 2097 -200 2109
rect -258 121 -246 2097
rect -212 121 -200 2097
rect -258 109 -200 121
rect 200 2097 258 2109
rect 200 121 212 2097
rect 246 121 258 2097
rect 200 109 258 121
rect -258 -121 -200 -109
rect -258 -2097 -246 -121
rect -212 -2097 -200 -121
rect -258 -2109 -200 -2097
rect 200 -121 258 -109
rect 200 -2097 212 -121
rect 246 -2097 258 -121
rect 200 -2109 258 -2097
<< ndiffc >>
rect -246 121 -212 2097
rect 212 121 246 2097
rect -246 -2097 -212 -121
rect 212 -2097 246 -121
<< poly >>
rect -200 2181 200 2197
rect -200 2147 -184 2181
rect 184 2147 200 2181
rect -200 2109 200 2147
rect -200 71 200 109
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -109 200 -71
rect -200 -2147 200 -2109
rect -200 -2181 -184 -2147
rect 184 -2181 200 -2147
rect -200 -2197 200 -2181
<< polycont >>
rect -184 2147 184 2181
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -2181 184 -2147
<< locali >>
rect -200 2147 -184 2181
rect 184 2147 200 2181
rect -246 2097 -212 2113
rect -246 105 -212 121
rect 212 2097 246 2113
rect 212 105 246 121
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -121 -212 -105
rect -246 -2113 -212 -2097
rect 212 -121 246 -105
rect 212 -2113 246 -2097
rect -200 -2181 -184 -2147
rect 184 -2181 200 -2147
<< viali >>
rect -184 2147 184 2181
rect -246 121 -212 2097
rect 212 121 246 2097
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -2097 -212 -121
rect 212 -2097 246 -121
rect -184 -2181 184 -2147
<< metal1 >>
rect -196 2181 196 2187
rect -196 2147 -184 2181
rect 184 2147 196 2181
rect -196 2141 196 2147
rect -252 2097 -206 2109
rect -252 121 -246 2097
rect -212 121 -206 2097
rect -252 109 -206 121
rect 206 2097 252 2109
rect 206 121 212 2097
rect 246 121 252 2097
rect 206 109 252 121
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -121 -206 -109
rect -252 -2097 -246 -121
rect -212 -2097 -206 -121
rect -252 -2109 -206 -2097
rect 206 -121 252 -109
rect 206 -2097 212 -121
rect 246 -2097 252 -121
rect 206 -2109 252 -2097
rect -196 -2147 196 -2141
rect -196 -2181 -184 -2147
rect 184 -2181 196 -2147
rect -196 -2187 196 -2181
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 2 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
