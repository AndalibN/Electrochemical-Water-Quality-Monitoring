magic
tech sky130A
magscale 1 2
timestamp 1668702877
<< pwell >>
rect -256 -84191 256 84191
<< nmos >>
rect -60 67381 60 83981
rect -60 50563 60 67163
rect -60 33745 60 50345
rect -60 16927 60 33527
rect -60 109 60 16709
rect -60 -16709 60 -109
rect -60 -33527 60 -16927
rect -60 -50345 60 -33745
rect -60 -67163 60 -50563
rect -60 -83981 60 -67381
<< ndiff >>
rect -118 83969 -60 83981
rect -118 67393 -106 83969
rect -72 67393 -60 83969
rect -118 67381 -60 67393
rect 60 83969 118 83981
rect 60 67393 72 83969
rect 106 67393 118 83969
rect 60 67381 118 67393
rect -118 67151 -60 67163
rect -118 50575 -106 67151
rect -72 50575 -60 67151
rect -118 50563 -60 50575
rect 60 67151 118 67163
rect 60 50575 72 67151
rect 106 50575 118 67151
rect 60 50563 118 50575
rect -118 50333 -60 50345
rect -118 33757 -106 50333
rect -72 33757 -60 50333
rect -118 33745 -60 33757
rect 60 50333 118 50345
rect 60 33757 72 50333
rect 106 33757 118 50333
rect 60 33745 118 33757
rect -118 33515 -60 33527
rect -118 16939 -106 33515
rect -72 16939 -60 33515
rect -118 16927 -60 16939
rect 60 33515 118 33527
rect 60 16939 72 33515
rect 106 16939 118 33515
rect 60 16927 118 16939
rect -118 16697 -60 16709
rect -118 121 -106 16697
rect -72 121 -60 16697
rect -118 109 -60 121
rect 60 16697 118 16709
rect 60 121 72 16697
rect 106 121 118 16697
rect 60 109 118 121
rect -118 -121 -60 -109
rect -118 -16697 -106 -121
rect -72 -16697 -60 -121
rect -118 -16709 -60 -16697
rect 60 -121 118 -109
rect 60 -16697 72 -121
rect 106 -16697 118 -121
rect 60 -16709 118 -16697
rect -118 -16939 -60 -16927
rect -118 -33515 -106 -16939
rect -72 -33515 -60 -16939
rect -118 -33527 -60 -33515
rect 60 -16939 118 -16927
rect 60 -33515 72 -16939
rect 106 -33515 118 -16939
rect 60 -33527 118 -33515
rect -118 -33757 -60 -33745
rect -118 -50333 -106 -33757
rect -72 -50333 -60 -33757
rect -118 -50345 -60 -50333
rect 60 -33757 118 -33745
rect 60 -50333 72 -33757
rect 106 -50333 118 -33757
rect 60 -50345 118 -50333
rect -118 -50575 -60 -50563
rect -118 -67151 -106 -50575
rect -72 -67151 -60 -50575
rect -118 -67163 -60 -67151
rect 60 -50575 118 -50563
rect 60 -67151 72 -50575
rect 106 -67151 118 -50575
rect 60 -67163 118 -67151
rect -118 -67393 -60 -67381
rect -118 -83969 -106 -67393
rect -72 -83969 -60 -67393
rect -118 -83981 -60 -83969
rect 60 -67393 118 -67381
rect 60 -83969 72 -67393
rect 106 -83969 118 -67393
rect 60 -83981 118 -83969
<< ndiffc >>
rect -106 67393 -72 83969
rect 72 67393 106 83969
rect -106 50575 -72 67151
rect 72 50575 106 67151
rect -106 33757 -72 50333
rect 72 33757 106 50333
rect -106 16939 -72 33515
rect 72 16939 106 33515
rect -106 121 -72 16697
rect 72 121 106 16697
rect -106 -16697 -72 -121
rect 72 -16697 106 -121
rect -106 -33515 -72 -16939
rect 72 -33515 106 -16939
rect -106 -50333 -72 -33757
rect 72 -50333 106 -33757
rect -106 -67151 -72 -50575
rect 72 -67151 106 -50575
rect -106 -83969 -72 -67393
rect 72 -83969 106 -67393
<< psubdiff >>
rect -220 84121 -124 84155
rect 124 84121 220 84155
rect -220 84059 -186 84121
rect 186 84059 220 84121
rect -220 -84121 -186 -84059
rect 186 -84121 220 -84059
rect -220 -84155 -124 -84121
rect 124 -84155 220 -84121
<< psubdiffcont >>
rect -124 84121 124 84155
rect -220 -84059 -186 84059
rect 186 -84059 220 84059
rect -124 -84155 124 -84121
<< poly >>
rect -60 84053 60 84069
rect -60 84019 -44 84053
rect 44 84019 60 84053
rect -60 83981 60 84019
rect -60 67343 60 67381
rect -60 67309 -44 67343
rect 44 67309 60 67343
rect -60 67293 60 67309
rect -60 67235 60 67251
rect -60 67201 -44 67235
rect 44 67201 60 67235
rect -60 67163 60 67201
rect -60 50525 60 50563
rect -60 50491 -44 50525
rect 44 50491 60 50525
rect -60 50475 60 50491
rect -60 50417 60 50433
rect -60 50383 -44 50417
rect 44 50383 60 50417
rect -60 50345 60 50383
rect -60 33707 60 33745
rect -60 33673 -44 33707
rect 44 33673 60 33707
rect -60 33657 60 33673
rect -60 33599 60 33615
rect -60 33565 -44 33599
rect 44 33565 60 33599
rect -60 33527 60 33565
rect -60 16889 60 16927
rect -60 16855 -44 16889
rect 44 16855 60 16889
rect -60 16839 60 16855
rect -60 16781 60 16797
rect -60 16747 -44 16781
rect 44 16747 60 16781
rect -60 16709 60 16747
rect -60 71 60 109
rect -60 37 -44 71
rect 44 37 60 71
rect -60 21 60 37
rect -60 -37 60 -21
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect -60 -109 60 -71
rect -60 -16747 60 -16709
rect -60 -16781 -44 -16747
rect 44 -16781 60 -16747
rect -60 -16797 60 -16781
rect -60 -16855 60 -16839
rect -60 -16889 -44 -16855
rect 44 -16889 60 -16855
rect -60 -16927 60 -16889
rect -60 -33565 60 -33527
rect -60 -33599 -44 -33565
rect 44 -33599 60 -33565
rect -60 -33615 60 -33599
rect -60 -33673 60 -33657
rect -60 -33707 -44 -33673
rect 44 -33707 60 -33673
rect -60 -33745 60 -33707
rect -60 -50383 60 -50345
rect -60 -50417 -44 -50383
rect 44 -50417 60 -50383
rect -60 -50433 60 -50417
rect -60 -50491 60 -50475
rect -60 -50525 -44 -50491
rect 44 -50525 60 -50491
rect -60 -50563 60 -50525
rect -60 -67201 60 -67163
rect -60 -67235 -44 -67201
rect 44 -67235 60 -67201
rect -60 -67251 60 -67235
rect -60 -67309 60 -67293
rect -60 -67343 -44 -67309
rect 44 -67343 60 -67309
rect -60 -67381 60 -67343
rect -60 -84019 60 -83981
rect -60 -84053 -44 -84019
rect 44 -84053 60 -84019
rect -60 -84069 60 -84053
<< polycont >>
rect -44 84019 44 84053
rect -44 67309 44 67343
rect -44 67201 44 67235
rect -44 50491 44 50525
rect -44 50383 44 50417
rect -44 33673 44 33707
rect -44 33565 44 33599
rect -44 16855 44 16889
rect -44 16747 44 16781
rect -44 37 44 71
rect -44 -71 44 -37
rect -44 -16781 44 -16747
rect -44 -16889 44 -16855
rect -44 -33599 44 -33565
rect -44 -33707 44 -33673
rect -44 -50417 44 -50383
rect -44 -50525 44 -50491
rect -44 -67235 44 -67201
rect -44 -67343 44 -67309
rect -44 -84053 44 -84019
<< locali >>
rect -220 84121 -124 84155
rect 124 84121 220 84155
rect -220 84059 -186 84121
rect 186 84059 220 84121
rect -60 84019 -44 84053
rect 44 84019 60 84053
rect -106 83969 -72 83985
rect -106 67377 -72 67393
rect 72 83969 106 83985
rect 72 67377 106 67393
rect -60 67309 -44 67343
rect 44 67309 60 67343
rect -60 67201 -44 67235
rect 44 67201 60 67235
rect -106 67151 -72 67167
rect -106 50559 -72 50575
rect 72 67151 106 67167
rect 72 50559 106 50575
rect -60 50491 -44 50525
rect 44 50491 60 50525
rect -60 50383 -44 50417
rect 44 50383 60 50417
rect -106 50333 -72 50349
rect -106 33741 -72 33757
rect 72 50333 106 50349
rect 72 33741 106 33757
rect -60 33673 -44 33707
rect 44 33673 60 33707
rect -60 33565 -44 33599
rect 44 33565 60 33599
rect -106 33515 -72 33531
rect -106 16923 -72 16939
rect 72 33515 106 33531
rect 72 16923 106 16939
rect -60 16855 -44 16889
rect 44 16855 60 16889
rect -60 16747 -44 16781
rect 44 16747 60 16781
rect -106 16697 -72 16713
rect -106 105 -72 121
rect 72 16697 106 16713
rect 72 105 106 121
rect -60 37 -44 71
rect 44 37 60 71
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect -106 -121 -72 -105
rect -106 -16713 -72 -16697
rect 72 -121 106 -105
rect 72 -16713 106 -16697
rect -60 -16781 -44 -16747
rect 44 -16781 60 -16747
rect -60 -16889 -44 -16855
rect 44 -16889 60 -16855
rect -106 -16939 -72 -16923
rect -106 -33531 -72 -33515
rect 72 -16939 106 -16923
rect 72 -33531 106 -33515
rect -60 -33599 -44 -33565
rect 44 -33599 60 -33565
rect -60 -33707 -44 -33673
rect 44 -33707 60 -33673
rect -106 -33757 -72 -33741
rect -106 -50349 -72 -50333
rect 72 -33757 106 -33741
rect 72 -50349 106 -50333
rect -60 -50417 -44 -50383
rect 44 -50417 60 -50383
rect -60 -50525 -44 -50491
rect 44 -50525 60 -50491
rect -106 -50575 -72 -50559
rect -106 -67167 -72 -67151
rect 72 -50575 106 -50559
rect 72 -67167 106 -67151
rect -60 -67235 -44 -67201
rect 44 -67235 60 -67201
rect -60 -67343 -44 -67309
rect 44 -67343 60 -67309
rect -106 -67393 -72 -67377
rect -106 -83985 -72 -83969
rect 72 -67393 106 -67377
rect 72 -83985 106 -83969
rect -60 -84053 -44 -84019
rect 44 -84053 60 -84019
rect -220 -84121 -186 -84059
rect 186 -84121 220 -84059
rect -220 -84155 -124 -84121
rect 124 -84155 220 -84121
<< viali >>
rect -44 84019 44 84053
rect -106 67393 -72 83969
rect 72 67393 106 83969
rect -44 67309 44 67343
rect -44 67201 44 67235
rect -106 50575 -72 67151
rect 72 50575 106 67151
rect -44 50491 44 50525
rect -44 50383 44 50417
rect -106 33757 -72 50333
rect 72 33757 106 50333
rect -44 33673 44 33707
rect -44 33565 44 33599
rect -106 16939 -72 33515
rect 72 16939 106 33515
rect -44 16855 44 16889
rect -44 16747 44 16781
rect -106 121 -72 16697
rect 72 121 106 16697
rect -44 37 44 71
rect -44 -71 44 -37
rect -106 -16697 -72 -121
rect 72 -16697 106 -121
rect -44 -16781 44 -16747
rect -44 -16889 44 -16855
rect -106 -33515 -72 -16939
rect 72 -33515 106 -16939
rect -44 -33599 44 -33565
rect -44 -33707 44 -33673
rect -106 -50333 -72 -33757
rect 72 -50333 106 -33757
rect -44 -50417 44 -50383
rect -44 -50525 44 -50491
rect -106 -67151 -72 -50575
rect 72 -67151 106 -50575
rect -44 -67235 44 -67201
rect -44 -67343 44 -67309
rect -106 -83969 -72 -67393
rect 72 -83969 106 -67393
rect -44 -84053 44 -84019
<< metal1 >>
rect -56 84053 56 84059
rect -56 84019 -44 84053
rect 44 84019 56 84053
rect -56 84013 56 84019
rect -112 83969 -66 83981
rect -112 67393 -106 83969
rect -72 67393 -66 83969
rect -112 67381 -66 67393
rect 66 83969 112 83981
rect 66 67393 72 83969
rect 106 67393 112 83969
rect 66 67381 112 67393
rect -56 67343 56 67349
rect -56 67309 -44 67343
rect 44 67309 56 67343
rect -56 67303 56 67309
rect -56 67235 56 67241
rect -56 67201 -44 67235
rect 44 67201 56 67235
rect -56 67195 56 67201
rect -112 67151 -66 67163
rect -112 50575 -106 67151
rect -72 50575 -66 67151
rect -112 50563 -66 50575
rect 66 67151 112 67163
rect 66 50575 72 67151
rect 106 50575 112 67151
rect 66 50563 112 50575
rect -56 50525 56 50531
rect -56 50491 -44 50525
rect 44 50491 56 50525
rect -56 50485 56 50491
rect -56 50417 56 50423
rect -56 50383 -44 50417
rect 44 50383 56 50417
rect -56 50377 56 50383
rect -112 50333 -66 50345
rect -112 33757 -106 50333
rect -72 33757 -66 50333
rect -112 33745 -66 33757
rect 66 50333 112 50345
rect 66 33757 72 50333
rect 106 33757 112 50333
rect 66 33745 112 33757
rect -56 33707 56 33713
rect -56 33673 -44 33707
rect 44 33673 56 33707
rect -56 33667 56 33673
rect -56 33599 56 33605
rect -56 33565 -44 33599
rect 44 33565 56 33599
rect -56 33559 56 33565
rect -112 33515 -66 33527
rect -112 16939 -106 33515
rect -72 16939 -66 33515
rect -112 16927 -66 16939
rect 66 33515 112 33527
rect 66 16939 72 33515
rect 106 16939 112 33515
rect 66 16927 112 16939
rect -56 16889 56 16895
rect -56 16855 -44 16889
rect 44 16855 56 16889
rect -56 16849 56 16855
rect -56 16781 56 16787
rect -56 16747 -44 16781
rect 44 16747 56 16781
rect -56 16741 56 16747
rect -112 16697 -66 16709
rect -112 121 -106 16697
rect -72 121 -66 16697
rect -112 109 -66 121
rect 66 16697 112 16709
rect 66 121 72 16697
rect 106 121 112 16697
rect 66 109 112 121
rect -56 71 56 77
rect -56 37 -44 71
rect 44 37 56 71
rect -56 31 56 37
rect -56 -37 56 -31
rect -56 -71 -44 -37
rect 44 -71 56 -37
rect -56 -77 56 -71
rect -112 -121 -66 -109
rect -112 -16697 -106 -121
rect -72 -16697 -66 -121
rect -112 -16709 -66 -16697
rect 66 -121 112 -109
rect 66 -16697 72 -121
rect 106 -16697 112 -121
rect 66 -16709 112 -16697
rect -56 -16747 56 -16741
rect -56 -16781 -44 -16747
rect 44 -16781 56 -16747
rect -56 -16787 56 -16781
rect -56 -16855 56 -16849
rect -56 -16889 -44 -16855
rect 44 -16889 56 -16855
rect -56 -16895 56 -16889
rect -112 -16939 -66 -16927
rect -112 -33515 -106 -16939
rect -72 -33515 -66 -16939
rect -112 -33527 -66 -33515
rect 66 -16939 112 -16927
rect 66 -33515 72 -16939
rect 106 -33515 112 -16939
rect 66 -33527 112 -33515
rect -56 -33565 56 -33559
rect -56 -33599 -44 -33565
rect 44 -33599 56 -33565
rect -56 -33605 56 -33599
rect -56 -33673 56 -33667
rect -56 -33707 -44 -33673
rect 44 -33707 56 -33673
rect -56 -33713 56 -33707
rect -112 -33757 -66 -33745
rect -112 -50333 -106 -33757
rect -72 -50333 -66 -33757
rect -112 -50345 -66 -50333
rect 66 -33757 112 -33745
rect 66 -50333 72 -33757
rect 106 -50333 112 -33757
rect 66 -50345 112 -50333
rect -56 -50383 56 -50377
rect -56 -50417 -44 -50383
rect 44 -50417 56 -50383
rect -56 -50423 56 -50417
rect -56 -50491 56 -50485
rect -56 -50525 -44 -50491
rect 44 -50525 56 -50491
rect -56 -50531 56 -50525
rect -112 -50575 -66 -50563
rect -112 -67151 -106 -50575
rect -72 -67151 -66 -50575
rect -112 -67163 -66 -67151
rect 66 -50575 112 -50563
rect 66 -67151 72 -50575
rect 106 -67151 112 -50575
rect 66 -67163 112 -67151
rect -56 -67201 56 -67195
rect -56 -67235 -44 -67201
rect 44 -67235 56 -67201
rect -56 -67241 56 -67235
rect -56 -67309 56 -67303
rect -56 -67343 -44 -67309
rect 44 -67343 56 -67309
rect -56 -67349 56 -67343
rect -112 -67393 -66 -67381
rect -112 -83969 -106 -67393
rect -72 -83969 -66 -67393
rect -112 -83981 -66 -83969
rect 66 -67393 112 -67381
rect 66 -83969 72 -67393
rect 106 -83969 112 -67393
rect 66 -83981 112 -83969
rect -56 -84019 56 -84013
rect -56 -84053 -44 -84019
rect 44 -84053 56 -84019
rect -56 -84059 56 -84053
<< properties >>
string FIXED_BBOX -203 -84138 203 84138
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 83.0 l 0.6 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
