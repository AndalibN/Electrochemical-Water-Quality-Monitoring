magic
tech sky130A
magscale 1 2
timestamp 1666102132
<< nwell >>
rect -246 -1337 246 1337
<< pmos >>
rect -50 118 50 1118
rect -50 -1118 50 -118
<< pdiff >>
rect -108 1106 -50 1118
rect -108 130 -96 1106
rect -62 130 -50 1106
rect -108 118 -50 130
rect 50 1106 108 1118
rect 50 130 62 1106
rect 96 130 108 1106
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -1106 -96 -130
rect -62 -1106 -50 -130
rect -108 -1118 -50 -1106
rect 50 -130 108 -118
rect 50 -1106 62 -130
rect 96 -1106 108 -130
rect 50 -1118 108 -1106
<< pdiffc >>
rect -96 130 -62 1106
rect 62 130 96 1106
rect -96 -1106 -62 -130
rect 62 -1106 96 -130
<< nsubdiff >>
rect -210 1267 -114 1301
rect 114 1267 210 1301
rect -210 1205 -176 1267
rect 176 1205 210 1267
rect -210 -1267 -176 -1205
rect 176 -1267 210 -1205
rect -210 -1301 -114 -1267
rect 114 -1301 210 -1267
<< nsubdiffcont >>
rect -114 1267 114 1301
rect -210 -1205 -176 1205
rect 176 -1205 210 1205
rect -114 -1301 114 -1267
<< poly >>
rect -50 1199 50 1215
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -50 1118 50 1165
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -1165 50 -1118
rect -50 -1199 -34 -1165
rect 34 -1199 50 -1165
rect -50 -1215 50 -1199
<< polycont >>
rect -34 1165 34 1199
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1199 34 -1165
<< locali >>
rect -210 1267 -114 1301
rect 114 1267 210 1301
rect -210 1205 -176 1267
rect 176 1205 210 1267
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -96 1106 -62 1122
rect -96 114 -62 130
rect 62 1106 96 1122
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -1122 -62 -1106
rect 62 -130 96 -114
rect 62 -1122 96 -1106
rect -50 -1199 -34 -1165
rect 34 -1199 50 -1165
rect -210 -1267 -176 -1205
rect 176 -1267 210 -1205
rect -210 -1301 -114 -1267
rect 114 -1301 210 -1267
<< viali >>
rect -34 1165 34 1199
rect -96 130 -62 1106
rect 62 130 96 1106
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1106 -62 -130
rect 62 -1106 96 -130
rect -34 -1199 34 -1165
<< metal1 >>
rect -46 1199 46 1205
rect -46 1165 -34 1199
rect 34 1165 46 1199
rect -46 1159 46 1165
rect -102 1106 -56 1118
rect -102 130 -96 1106
rect -62 130 -56 1106
rect -102 118 -56 130
rect 56 1106 102 1118
rect 56 130 62 1106
rect 96 130 102 1106
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -1106 -96 -130
rect -62 -1106 -56 -130
rect -102 -1118 -56 -1106
rect 56 -130 102 -118
rect 56 -1106 62 -130
rect 96 -1106 102 -130
rect 56 -1118 102 -1106
rect -46 -1165 46 -1159
rect -46 -1199 -34 -1165
rect 34 -1199 46 -1165
rect -46 -1205 46 -1199
<< properties >>
string FIXED_BBOX -193 -1284 193 1284
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
