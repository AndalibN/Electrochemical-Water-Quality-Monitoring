magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 3000 35 3432
rect -35 -3432 35 -3000
<< xpolyres >>
rect -35 -3000 35 3000
<< viali >>
rect -17 3378 17 3412
rect -17 3306 17 3340
rect -17 3234 17 3268
rect -17 3162 17 3196
rect -17 3090 17 3124
rect -17 3018 17 3052
rect -17 -3053 17 -3019
rect -17 -3125 17 -3091
rect -17 -3197 17 -3163
rect -17 -3269 17 -3235
rect -17 -3341 17 -3307
rect -17 -3413 17 -3379
<< metal1 >>
rect -25 3412 25 3426
rect -25 3378 -17 3412
rect 17 3378 25 3412
rect -25 3340 25 3378
rect -25 3306 -17 3340
rect 17 3306 25 3340
rect -25 3268 25 3306
rect -25 3234 -17 3268
rect 17 3234 25 3268
rect -25 3196 25 3234
rect -25 3162 -17 3196
rect 17 3162 25 3196
rect -25 3124 25 3162
rect -25 3090 -17 3124
rect 17 3090 25 3124
rect -25 3052 25 3090
rect -25 3018 -17 3052
rect 17 3018 25 3052
rect -25 3005 25 3018
rect -25 -3019 25 -3005
rect -25 -3053 -17 -3019
rect 17 -3053 25 -3019
rect -25 -3091 25 -3053
rect -25 -3125 -17 -3091
rect 17 -3125 25 -3091
rect -25 -3163 25 -3125
rect -25 -3197 -17 -3163
rect 17 -3197 25 -3163
rect -25 -3235 25 -3197
rect -25 -3269 -17 -3235
rect 17 -3269 25 -3235
rect -25 -3307 25 -3269
rect -25 -3341 -17 -3307
rect 17 -3341 25 -3307
rect -25 -3379 25 -3341
rect -25 -3413 -17 -3379
rect 17 -3413 25 -3379
rect -25 -3426 25 -3413
<< end >>
