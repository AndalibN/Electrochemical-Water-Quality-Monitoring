magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -184 -757 184 695
<< nmos >>
rect -100 -731 100 669
<< ndiff >>
rect -158 632 -100 669
rect -158 598 -146 632
rect -112 598 -100 632
rect -158 564 -100 598
rect -158 530 -146 564
rect -112 530 -100 564
rect -158 496 -100 530
rect -158 462 -146 496
rect -112 462 -100 496
rect -158 428 -100 462
rect -158 394 -146 428
rect -112 394 -100 428
rect -158 360 -100 394
rect -158 326 -146 360
rect -112 326 -100 360
rect -158 292 -100 326
rect -158 258 -146 292
rect -112 258 -100 292
rect -158 224 -100 258
rect -158 190 -146 224
rect -112 190 -100 224
rect -158 156 -100 190
rect -158 122 -146 156
rect -112 122 -100 156
rect -158 88 -100 122
rect -158 54 -146 88
rect -112 54 -100 88
rect -158 20 -100 54
rect -158 -14 -146 20
rect -112 -14 -100 20
rect -158 -48 -100 -14
rect -158 -82 -146 -48
rect -112 -82 -100 -48
rect -158 -116 -100 -82
rect -158 -150 -146 -116
rect -112 -150 -100 -116
rect -158 -184 -100 -150
rect -158 -218 -146 -184
rect -112 -218 -100 -184
rect -158 -252 -100 -218
rect -158 -286 -146 -252
rect -112 -286 -100 -252
rect -158 -320 -100 -286
rect -158 -354 -146 -320
rect -112 -354 -100 -320
rect -158 -388 -100 -354
rect -158 -422 -146 -388
rect -112 -422 -100 -388
rect -158 -456 -100 -422
rect -158 -490 -146 -456
rect -112 -490 -100 -456
rect -158 -524 -100 -490
rect -158 -558 -146 -524
rect -112 -558 -100 -524
rect -158 -592 -100 -558
rect -158 -626 -146 -592
rect -112 -626 -100 -592
rect -158 -660 -100 -626
rect -158 -694 -146 -660
rect -112 -694 -100 -660
rect -158 -731 -100 -694
rect 100 632 158 669
rect 100 598 112 632
rect 146 598 158 632
rect 100 564 158 598
rect 100 530 112 564
rect 146 530 158 564
rect 100 496 158 530
rect 100 462 112 496
rect 146 462 158 496
rect 100 428 158 462
rect 100 394 112 428
rect 146 394 158 428
rect 100 360 158 394
rect 100 326 112 360
rect 146 326 158 360
rect 100 292 158 326
rect 100 258 112 292
rect 146 258 158 292
rect 100 224 158 258
rect 100 190 112 224
rect 146 190 158 224
rect 100 156 158 190
rect 100 122 112 156
rect 146 122 158 156
rect 100 88 158 122
rect 100 54 112 88
rect 146 54 158 88
rect 100 20 158 54
rect 100 -14 112 20
rect 146 -14 158 20
rect 100 -48 158 -14
rect 100 -82 112 -48
rect 146 -82 158 -48
rect 100 -116 158 -82
rect 100 -150 112 -116
rect 146 -150 158 -116
rect 100 -184 158 -150
rect 100 -218 112 -184
rect 146 -218 158 -184
rect 100 -252 158 -218
rect 100 -286 112 -252
rect 146 -286 158 -252
rect 100 -320 158 -286
rect 100 -354 112 -320
rect 146 -354 158 -320
rect 100 -388 158 -354
rect 100 -422 112 -388
rect 146 -422 158 -388
rect 100 -456 158 -422
rect 100 -490 112 -456
rect 146 -490 158 -456
rect 100 -524 158 -490
rect 100 -558 112 -524
rect 146 -558 158 -524
rect 100 -592 158 -558
rect 100 -626 112 -592
rect 146 -626 158 -592
rect 100 -660 158 -626
rect 100 -694 112 -660
rect 146 -694 158 -660
rect 100 -731 158 -694
<< ndiffc >>
rect -146 598 -112 632
rect -146 530 -112 564
rect -146 462 -112 496
rect -146 394 -112 428
rect -146 326 -112 360
rect -146 258 -112 292
rect -146 190 -112 224
rect -146 122 -112 156
rect -146 54 -112 88
rect -146 -14 -112 20
rect -146 -82 -112 -48
rect -146 -150 -112 -116
rect -146 -218 -112 -184
rect -146 -286 -112 -252
rect -146 -354 -112 -320
rect -146 -422 -112 -388
rect -146 -490 -112 -456
rect -146 -558 -112 -524
rect -146 -626 -112 -592
rect -146 -694 -112 -660
rect 112 598 146 632
rect 112 530 146 564
rect 112 462 146 496
rect 112 394 146 428
rect 112 326 146 360
rect 112 258 146 292
rect 112 190 146 224
rect 112 122 146 156
rect 112 54 146 88
rect 112 -14 146 20
rect 112 -82 146 -48
rect 112 -150 146 -116
rect 112 -218 146 -184
rect 112 -286 146 -252
rect 112 -354 146 -320
rect 112 -422 146 -388
rect 112 -490 146 -456
rect 112 -558 146 -524
rect 112 -626 146 -592
rect 112 -694 146 -660
<< poly >>
rect -100 741 100 757
rect -100 707 -51 741
rect -17 707 17 741
rect 51 707 100 741
rect -100 669 100 707
rect -100 -757 100 -731
<< polycont >>
rect -51 707 -17 741
rect 17 707 51 741
<< locali >>
rect -100 707 -53 741
rect -17 707 17 741
rect 53 707 100 741
rect -146 634 -112 673
rect -146 564 -112 598
rect -146 496 -112 528
rect -146 428 -112 456
rect -146 360 -112 384
rect -146 292 -112 312
rect -146 224 -112 240
rect -146 156 -112 168
rect -146 88 -112 96
rect -146 20 -112 24
rect -146 -86 -112 -82
rect -146 -158 -112 -150
rect -146 -230 -112 -218
rect -146 -302 -112 -286
rect -146 -374 -112 -354
rect -146 -446 -112 -422
rect -146 -518 -112 -490
rect -146 -590 -112 -558
rect -146 -660 -112 -626
rect -146 -735 -112 -696
rect 112 634 146 673
rect 112 564 146 598
rect 112 496 146 528
rect 112 428 146 456
rect 112 360 146 384
rect 112 292 146 312
rect 112 224 146 240
rect 112 156 146 168
rect 112 88 146 96
rect 112 20 146 24
rect 112 -86 146 -82
rect 112 -158 146 -150
rect 112 -230 146 -218
rect 112 -302 146 -286
rect 112 -374 146 -354
rect 112 -446 146 -422
rect 112 -518 146 -490
rect 112 -590 146 -558
rect 112 -660 146 -626
rect 112 -735 146 -696
<< viali >>
rect -53 707 -51 741
rect -51 707 -19 741
rect 19 707 51 741
rect 51 707 53 741
rect -146 632 -112 634
rect -146 600 -112 632
rect -146 530 -112 562
rect -146 528 -112 530
rect -146 462 -112 490
rect -146 456 -112 462
rect -146 394 -112 418
rect -146 384 -112 394
rect -146 326 -112 346
rect -146 312 -112 326
rect -146 258 -112 274
rect -146 240 -112 258
rect -146 190 -112 202
rect -146 168 -112 190
rect -146 122 -112 130
rect -146 96 -112 122
rect -146 54 -112 58
rect -146 24 -112 54
rect -146 -48 -112 -14
rect -146 -116 -112 -86
rect -146 -120 -112 -116
rect -146 -184 -112 -158
rect -146 -192 -112 -184
rect -146 -252 -112 -230
rect -146 -264 -112 -252
rect -146 -320 -112 -302
rect -146 -336 -112 -320
rect -146 -388 -112 -374
rect -146 -408 -112 -388
rect -146 -456 -112 -446
rect -146 -480 -112 -456
rect -146 -524 -112 -518
rect -146 -552 -112 -524
rect -146 -592 -112 -590
rect -146 -624 -112 -592
rect -146 -694 -112 -662
rect -146 -696 -112 -694
rect 112 632 146 634
rect 112 600 146 632
rect 112 530 146 562
rect 112 528 146 530
rect 112 462 146 490
rect 112 456 146 462
rect 112 394 146 418
rect 112 384 146 394
rect 112 326 146 346
rect 112 312 146 326
rect 112 258 146 274
rect 112 240 146 258
rect 112 190 146 202
rect 112 168 146 190
rect 112 122 146 130
rect 112 96 146 122
rect 112 54 146 58
rect 112 24 146 54
rect 112 -48 146 -14
rect 112 -116 146 -86
rect 112 -120 146 -116
rect 112 -184 146 -158
rect 112 -192 146 -184
rect 112 -252 146 -230
rect 112 -264 146 -252
rect 112 -320 146 -302
rect 112 -336 146 -320
rect 112 -388 146 -374
rect 112 -408 146 -388
rect 112 -456 146 -446
rect 112 -480 146 -456
rect 112 -524 146 -518
rect 112 -552 146 -524
rect 112 -592 146 -590
rect 112 -624 146 -592
rect 112 -694 146 -662
rect 112 -696 146 -694
<< metal1 >>
rect -96 741 96 747
rect -96 707 -53 741
rect -19 707 19 741
rect 53 707 96 741
rect -96 701 96 707
rect -152 634 -106 669
rect -152 600 -146 634
rect -112 600 -106 634
rect -152 562 -106 600
rect -152 528 -146 562
rect -112 528 -106 562
rect -152 490 -106 528
rect -152 456 -146 490
rect -112 456 -106 490
rect -152 418 -106 456
rect -152 384 -146 418
rect -112 384 -106 418
rect -152 346 -106 384
rect -152 312 -146 346
rect -112 312 -106 346
rect -152 274 -106 312
rect -152 240 -146 274
rect -112 240 -106 274
rect -152 202 -106 240
rect -152 168 -146 202
rect -112 168 -106 202
rect -152 130 -106 168
rect -152 96 -146 130
rect -112 96 -106 130
rect -152 58 -106 96
rect -152 24 -146 58
rect -112 24 -106 58
rect -152 -14 -106 24
rect -152 -48 -146 -14
rect -112 -48 -106 -14
rect -152 -86 -106 -48
rect -152 -120 -146 -86
rect -112 -120 -106 -86
rect -152 -158 -106 -120
rect -152 -192 -146 -158
rect -112 -192 -106 -158
rect -152 -230 -106 -192
rect -152 -264 -146 -230
rect -112 -264 -106 -230
rect -152 -302 -106 -264
rect -152 -336 -146 -302
rect -112 -336 -106 -302
rect -152 -374 -106 -336
rect -152 -408 -146 -374
rect -112 -408 -106 -374
rect -152 -446 -106 -408
rect -152 -480 -146 -446
rect -112 -480 -106 -446
rect -152 -518 -106 -480
rect -152 -552 -146 -518
rect -112 -552 -106 -518
rect -152 -590 -106 -552
rect -152 -624 -146 -590
rect -112 -624 -106 -590
rect -152 -662 -106 -624
rect -152 -696 -146 -662
rect -112 -696 -106 -662
rect -152 -731 -106 -696
rect 106 634 152 669
rect 106 600 112 634
rect 146 600 152 634
rect 106 562 152 600
rect 106 528 112 562
rect 146 528 152 562
rect 106 490 152 528
rect 106 456 112 490
rect 146 456 152 490
rect 106 418 152 456
rect 106 384 112 418
rect 146 384 152 418
rect 106 346 152 384
rect 106 312 112 346
rect 146 312 152 346
rect 106 274 152 312
rect 106 240 112 274
rect 146 240 152 274
rect 106 202 152 240
rect 106 168 112 202
rect 146 168 152 202
rect 106 130 152 168
rect 106 96 112 130
rect 146 96 152 130
rect 106 58 152 96
rect 106 24 112 58
rect 146 24 152 58
rect 106 -14 152 24
rect 106 -48 112 -14
rect 146 -48 152 -14
rect 106 -86 152 -48
rect 106 -120 112 -86
rect 146 -120 152 -86
rect 106 -158 152 -120
rect 106 -192 112 -158
rect 146 -192 152 -158
rect 106 -230 152 -192
rect 106 -264 112 -230
rect 146 -264 152 -230
rect 106 -302 152 -264
rect 106 -336 112 -302
rect 146 -336 152 -302
rect 106 -374 152 -336
rect 106 -408 112 -374
rect 146 -408 152 -374
rect 106 -446 152 -408
rect 106 -480 112 -446
rect 146 -480 152 -446
rect 106 -518 152 -480
rect 106 -552 112 -518
rect 146 -552 152 -518
rect 106 -590 152 -552
rect 106 -624 112 -590
rect 146 -624 152 -590
rect 106 -662 152 -624
rect 106 -696 112 -662
rect 146 -696 152 -662
rect 106 -731 152 -696
<< end >>
