magic
tech sky130A
timestamp 1668374365
<< nmos >>
rect -537 -3000 -507 3000
rect -421 -3000 -391 3000
rect -305 -3000 -275 3000
rect -189 -3000 -159 3000
rect -73 -3000 -43 3000
rect 43 -3000 73 3000
rect 159 -3000 189 3000
rect 275 -3000 305 3000
rect 391 -3000 421 3000
rect 507 -3000 537 3000
<< ndiff >>
rect -566 2994 -537 3000
rect -566 -2994 -560 2994
rect -543 -2994 -537 2994
rect -566 -3000 -537 -2994
rect -507 2994 -478 3000
rect -507 -2994 -501 2994
rect -484 -2994 -478 2994
rect -507 -3000 -478 -2994
rect -450 2994 -421 3000
rect -450 -2994 -444 2994
rect -427 -2994 -421 2994
rect -450 -3000 -421 -2994
rect -391 2994 -362 3000
rect -391 -2994 -385 2994
rect -368 -2994 -362 2994
rect -391 -3000 -362 -2994
rect -334 2994 -305 3000
rect -334 -2994 -328 2994
rect -311 -2994 -305 2994
rect -334 -3000 -305 -2994
rect -275 2994 -246 3000
rect -275 -2994 -269 2994
rect -252 -2994 -246 2994
rect -275 -3000 -246 -2994
rect -218 2994 -189 3000
rect -218 -2994 -212 2994
rect -195 -2994 -189 2994
rect -218 -3000 -189 -2994
rect -159 2994 -130 3000
rect -159 -2994 -153 2994
rect -136 -2994 -130 2994
rect -159 -3000 -130 -2994
rect -102 2994 -73 3000
rect -102 -2994 -96 2994
rect -79 -2994 -73 2994
rect -102 -3000 -73 -2994
rect -43 2994 -14 3000
rect -43 -2994 -37 2994
rect -20 -2994 -14 2994
rect -43 -3000 -14 -2994
rect 14 2994 43 3000
rect 14 -2994 20 2994
rect 37 -2994 43 2994
rect 14 -3000 43 -2994
rect 73 2994 102 3000
rect 73 -2994 79 2994
rect 96 -2994 102 2994
rect 73 -3000 102 -2994
rect 130 2994 159 3000
rect 130 -2994 136 2994
rect 153 -2994 159 2994
rect 130 -3000 159 -2994
rect 189 2994 218 3000
rect 189 -2994 195 2994
rect 212 -2994 218 2994
rect 189 -3000 218 -2994
rect 246 2994 275 3000
rect 246 -2994 252 2994
rect 269 -2994 275 2994
rect 246 -3000 275 -2994
rect 305 2994 334 3000
rect 305 -2994 311 2994
rect 328 -2994 334 2994
rect 305 -3000 334 -2994
rect 362 2994 391 3000
rect 362 -2994 368 2994
rect 385 -2994 391 2994
rect 362 -3000 391 -2994
rect 421 2994 450 3000
rect 421 -2994 427 2994
rect 444 -2994 450 2994
rect 421 -3000 450 -2994
rect 478 2994 507 3000
rect 478 -2994 484 2994
rect 501 -2994 507 2994
rect 478 -3000 507 -2994
rect 537 2994 566 3000
rect 537 -2994 543 2994
rect 560 -2994 566 2994
rect 537 -3000 566 -2994
<< ndiffc >>
rect -560 -2994 -543 2994
rect -501 -2994 -484 2994
rect -444 -2994 -427 2994
rect -385 -2994 -368 2994
rect -328 -2994 -311 2994
rect -269 -2994 -252 2994
rect -212 -2994 -195 2994
rect -153 -2994 -136 2994
rect -96 -2994 -79 2994
rect -37 -2994 -20 2994
rect 20 -2994 37 2994
rect 79 -2994 96 2994
rect 136 -2994 153 2994
rect 195 -2994 212 2994
rect 252 -2994 269 2994
rect 311 -2994 328 2994
rect 368 -2994 385 2994
rect 427 -2994 444 2994
rect 484 -2994 501 2994
rect 543 -2994 560 2994
<< poly >>
rect -537 3000 -507 3013
rect -421 3000 -391 3013
rect -305 3000 -275 3013
rect -189 3000 -159 3013
rect -73 3000 -43 3013
rect 43 3000 73 3013
rect 159 3000 189 3013
rect 275 3000 305 3013
rect 391 3000 421 3013
rect 507 3000 537 3013
rect -537 -3013 -507 -3000
rect -421 -3013 -391 -3000
rect -305 -3013 -275 -3000
rect -189 -3013 -159 -3000
rect -73 -3013 -43 -3000
rect 43 -3013 73 -3000
rect 159 -3013 189 -3000
rect 275 -3013 305 -3000
rect 391 -3013 421 -3000
rect 507 -3013 537 -3000
<< locali >>
rect -560 2994 -543 3002
rect -560 -3002 -543 -2994
rect -501 2994 -484 3002
rect -501 -3002 -484 -2994
rect -444 2994 -427 3002
rect -444 -3002 -427 -2994
rect -385 2994 -368 3002
rect -385 -3002 -368 -2994
rect -328 2994 -311 3002
rect -328 -3002 -311 -2994
rect -269 2994 -252 3002
rect -269 -3002 -252 -2994
rect -212 2994 -195 3002
rect -212 -3002 -195 -2994
rect -153 2994 -136 3002
rect -153 -3002 -136 -2994
rect -96 2994 -79 3002
rect -96 -3002 -79 -2994
rect -37 2994 -20 3002
rect -37 -3002 -20 -2994
rect 20 2994 37 3002
rect 20 -3002 37 -2994
rect 79 2994 96 3002
rect 79 -3002 96 -2994
rect 136 2994 153 3002
rect 136 -3002 153 -2994
rect 195 2994 212 3002
rect 195 -3002 212 -2994
rect 252 2994 269 3002
rect 252 -3002 269 -2994
rect 311 2994 328 3002
rect 311 -3002 328 -2994
rect 368 2994 385 3002
rect 368 -3002 385 -2994
rect 427 2994 444 3002
rect 427 -3002 444 -2994
rect 484 2994 501 3002
rect 484 -3002 501 -2994
rect 543 2994 560 3002
rect 543 -3002 560 -2994
<< viali >>
rect -560 -2994 -543 2994
rect -501 -2994 -484 2994
rect -444 -2994 -427 2994
rect -385 -2994 -368 2994
rect -328 -2994 -311 2994
rect -269 -2994 -252 2994
rect -212 -2994 -195 2994
rect -153 -2994 -136 2994
rect -96 -2994 -79 2994
rect -37 -2994 -20 2994
rect 20 -2994 37 2994
rect 79 -2994 96 2994
rect 136 -2994 153 2994
rect 195 -2994 212 2994
rect 252 -2994 269 2994
rect 311 -2994 328 2994
rect 368 -2994 385 2994
rect 427 -2994 444 2994
rect 484 -2994 501 2994
rect 543 -2994 560 2994
<< metal1 >>
rect -563 2994 -540 3000
rect -563 -2994 -560 2994
rect -543 -2994 -540 2994
rect -563 -3000 -540 -2994
rect -504 2994 -481 3000
rect -504 -2994 -501 2994
rect -484 -2994 -481 2994
rect -504 -3000 -481 -2994
rect -447 2994 -424 3000
rect -447 -2994 -444 2994
rect -427 -2994 -424 2994
rect -447 -3000 -424 -2994
rect -388 2994 -365 3000
rect -388 -2994 -385 2994
rect -368 -2994 -365 2994
rect -388 -3000 -365 -2994
rect -331 2994 -308 3000
rect -331 -2994 -328 2994
rect -311 -2994 -308 2994
rect -331 -3000 -308 -2994
rect -272 2994 -249 3000
rect -272 -2994 -269 2994
rect -252 -2994 -249 2994
rect -272 -3000 -249 -2994
rect -215 2994 -192 3000
rect -215 -2994 -212 2994
rect -195 -2994 -192 2994
rect -215 -3000 -192 -2994
rect -156 2994 -133 3000
rect -156 -2994 -153 2994
rect -136 -2994 -133 2994
rect -156 -3000 -133 -2994
rect -99 2994 -76 3000
rect -99 -2994 -96 2994
rect -79 -2994 -76 2994
rect -99 -3000 -76 -2994
rect -40 2994 -17 3000
rect -40 -2994 -37 2994
rect -20 -2994 -17 2994
rect -40 -3000 -17 -2994
rect 17 2994 40 3000
rect 17 -2994 20 2994
rect 37 -2994 40 2994
rect 17 -3000 40 -2994
rect 76 2994 99 3000
rect 76 -2994 79 2994
rect 96 -2994 99 2994
rect 76 -3000 99 -2994
rect 133 2994 156 3000
rect 133 -2994 136 2994
rect 153 -2994 156 2994
rect 133 -3000 156 -2994
rect 192 2994 215 3000
rect 192 -2994 195 2994
rect 212 -2994 215 2994
rect 192 -3000 215 -2994
rect 249 2994 272 3000
rect 249 -2994 252 2994
rect 269 -2994 272 2994
rect 249 -3000 272 -2994
rect 308 2994 331 3000
rect 308 -2994 311 2994
rect 328 -2994 331 2994
rect 308 -3000 331 -2994
rect 365 2994 388 3000
rect 365 -2994 368 2994
rect 385 -2994 388 2994
rect 365 -3000 388 -2994
rect 424 2994 447 3000
rect 424 -2994 427 2994
rect 444 -2994 447 2994
rect 424 -3000 447 -2994
rect 481 2994 504 3000
rect 481 -2994 484 2994
rect 501 -2994 504 2994
rect 481 -3000 504 -2994
rect 540 2994 563 3000
rect 540 -2994 543 2994
rect 560 -2994 563 2994
rect 540 -3000 563 -2994
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 60 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
