magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 510 35 942
rect -35 -942 35 -510
<< xpolyres >>
rect -35 -510 35 510
<< viali >>
rect -17 888 17 922
rect -17 816 17 850
rect -17 744 17 778
rect -17 672 17 706
rect -17 600 17 634
rect -17 528 17 562
rect -17 -563 17 -529
rect -17 -635 17 -601
rect -17 -707 17 -673
rect -17 -779 17 -745
rect -17 -851 17 -817
rect -17 -923 17 -889
<< metal1 >>
rect -25 922 25 936
rect -25 888 -17 922
rect 17 888 25 922
rect -25 850 25 888
rect -25 816 -17 850
rect 17 816 25 850
rect -25 778 25 816
rect -25 744 -17 778
rect 17 744 25 778
rect -25 706 25 744
rect -25 672 -17 706
rect 17 672 25 706
rect -25 634 25 672
rect -25 600 -17 634
rect 17 600 25 634
rect -25 562 25 600
rect -25 528 -17 562
rect 17 528 25 562
rect -25 515 25 528
rect -25 -529 25 -515
rect -25 -563 -17 -529
rect 17 -563 25 -529
rect -25 -601 25 -563
rect -25 -635 -17 -601
rect 17 -635 25 -601
rect -25 -673 25 -635
rect -25 -707 -17 -673
rect 17 -707 25 -673
rect -25 -745 25 -707
rect -25 -779 -17 -745
rect 17 -779 25 -745
rect -25 -817 25 -779
rect -25 -851 -17 -817
rect 17 -851 25 -817
rect -25 -889 25 -851
rect -25 -923 -17 -889
rect 17 -923 25 -889
rect -25 -936 25 -923
<< end >>
