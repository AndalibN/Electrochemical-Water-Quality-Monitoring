magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nmos >>
rect -603 -1250 -503 1250
rect -445 -1250 -345 1250
rect -287 -1250 -187 1250
rect -129 -1250 -29 1250
rect 29 -1250 129 1250
rect 187 -1250 287 1250
rect 345 -1250 445 1250
rect 503 -1250 603 1250
<< ndiff >>
rect -661 1238 -603 1250
rect -661 -1238 -649 1238
rect -615 -1238 -603 1238
rect -661 -1250 -603 -1238
rect -503 1238 -445 1250
rect -503 -1238 -491 1238
rect -457 -1238 -445 1238
rect -503 -1250 -445 -1238
rect -345 1238 -287 1250
rect -345 -1238 -333 1238
rect -299 -1238 -287 1238
rect -345 -1250 -287 -1238
rect -187 1238 -129 1250
rect -187 -1238 -175 1238
rect -141 -1238 -129 1238
rect -187 -1250 -129 -1238
rect -29 1238 29 1250
rect -29 -1238 -17 1238
rect 17 -1238 29 1238
rect -29 -1250 29 -1238
rect 129 1238 187 1250
rect 129 -1238 141 1238
rect 175 -1238 187 1238
rect 129 -1250 187 -1238
rect 287 1238 345 1250
rect 287 -1238 299 1238
rect 333 -1238 345 1238
rect 287 -1250 345 -1238
rect 445 1238 503 1250
rect 445 -1238 457 1238
rect 491 -1238 503 1238
rect 445 -1250 503 -1238
rect 603 1238 661 1250
rect 603 -1238 615 1238
rect 649 -1238 661 1238
rect 603 -1250 661 -1238
<< ndiffc >>
rect -649 -1238 -615 1238
rect -491 -1238 -457 1238
rect -333 -1238 -299 1238
rect -175 -1238 -141 1238
rect -17 -1238 17 1238
rect 141 -1238 175 1238
rect 299 -1238 333 1238
rect 457 -1238 491 1238
rect 615 -1238 649 1238
<< poly >>
rect -603 1322 -503 1338
rect -603 1288 -587 1322
rect -519 1288 -503 1322
rect -603 1250 -503 1288
rect -445 1322 -345 1338
rect -445 1288 -429 1322
rect -361 1288 -345 1322
rect -445 1250 -345 1288
rect -287 1322 -187 1338
rect -287 1288 -271 1322
rect -203 1288 -187 1322
rect -287 1250 -187 1288
rect -129 1322 -29 1338
rect -129 1288 -113 1322
rect -45 1288 -29 1322
rect -129 1250 -29 1288
rect 29 1322 129 1338
rect 29 1288 45 1322
rect 113 1288 129 1322
rect 29 1250 129 1288
rect 187 1322 287 1338
rect 187 1288 203 1322
rect 271 1288 287 1322
rect 187 1250 287 1288
rect 345 1322 445 1338
rect 345 1288 361 1322
rect 429 1288 445 1322
rect 345 1250 445 1288
rect 503 1322 603 1338
rect 503 1288 519 1322
rect 587 1288 603 1322
rect 503 1250 603 1288
rect -603 -1288 -503 -1250
rect -603 -1322 -587 -1288
rect -519 -1322 -503 -1288
rect -603 -1338 -503 -1322
rect -445 -1288 -345 -1250
rect -445 -1322 -429 -1288
rect -361 -1322 -345 -1288
rect -445 -1338 -345 -1322
rect -287 -1288 -187 -1250
rect -287 -1322 -271 -1288
rect -203 -1322 -187 -1288
rect -287 -1338 -187 -1322
rect -129 -1288 -29 -1250
rect -129 -1322 -113 -1288
rect -45 -1322 -29 -1288
rect -129 -1338 -29 -1322
rect 29 -1288 129 -1250
rect 29 -1322 45 -1288
rect 113 -1322 129 -1288
rect 29 -1338 129 -1322
rect 187 -1288 287 -1250
rect 187 -1322 203 -1288
rect 271 -1322 287 -1288
rect 187 -1338 287 -1322
rect 345 -1288 445 -1250
rect 345 -1322 361 -1288
rect 429 -1322 445 -1288
rect 345 -1338 445 -1322
rect 503 -1288 603 -1250
rect 503 -1322 519 -1288
rect 587 -1322 603 -1288
rect 503 -1338 603 -1322
<< polycont >>
rect -587 1288 -519 1322
rect -429 1288 -361 1322
rect -271 1288 -203 1322
rect -113 1288 -45 1322
rect 45 1288 113 1322
rect 203 1288 271 1322
rect 361 1288 429 1322
rect 519 1288 587 1322
rect -587 -1322 -519 -1288
rect -429 -1322 -361 -1288
rect -271 -1322 -203 -1288
rect -113 -1322 -45 -1288
rect 45 -1322 113 -1288
rect 203 -1322 271 -1288
rect 361 -1322 429 -1288
rect 519 -1322 587 -1288
<< locali >>
rect -603 1288 -587 1322
rect -519 1288 -503 1322
rect -445 1288 -429 1322
rect -361 1288 -345 1322
rect -287 1288 -271 1322
rect -203 1288 -187 1322
rect -129 1288 -113 1322
rect -45 1288 -29 1322
rect 29 1288 45 1322
rect 113 1288 129 1322
rect 187 1288 203 1322
rect 271 1288 287 1322
rect 345 1288 361 1322
rect 429 1288 445 1322
rect 503 1288 519 1322
rect 587 1288 603 1322
rect -649 1238 -615 1254
rect -649 -1254 -615 -1238
rect -491 1238 -457 1254
rect -491 -1254 -457 -1238
rect -333 1238 -299 1254
rect -333 -1254 -299 -1238
rect -175 1238 -141 1254
rect -175 -1254 -141 -1238
rect -17 1238 17 1254
rect -17 -1254 17 -1238
rect 141 1238 175 1254
rect 141 -1254 175 -1238
rect 299 1238 333 1254
rect 299 -1254 333 -1238
rect 457 1238 491 1254
rect 457 -1254 491 -1238
rect 615 1238 649 1254
rect 615 -1254 649 -1238
rect -603 -1322 -587 -1288
rect -519 -1322 -503 -1288
rect -445 -1322 -429 -1288
rect -361 -1322 -345 -1288
rect -287 -1322 -271 -1288
rect -203 -1322 -187 -1288
rect -129 -1322 -113 -1288
rect -45 -1322 -29 -1288
rect 29 -1322 45 -1288
rect 113 -1322 129 -1288
rect 187 -1322 203 -1288
rect 271 -1322 287 -1288
rect 345 -1322 361 -1288
rect 429 -1322 445 -1288
rect 503 -1322 519 -1288
rect 587 -1322 603 -1288
<< viali >>
rect -587 1288 -519 1322
rect -429 1288 -361 1322
rect -271 1288 -203 1322
rect -113 1288 -45 1322
rect 45 1288 113 1322
rect 203 1288 271 1322
rect 361 1288 429 1322
rect 519 1288 587 1322
rect -649 -1238 -615 1238
rect -491 -1238 -457 1238
rect -333 -1238 -299 1238
rect -175 -1238 -141 1238
rect -17 -1238 17 1238
rect 141 -1238 175 1238
rect 299 -1238 333 1238
rect 457 -1238 491 1238
rect 615 -1238 649 1238
rect -587 -1322 -519 -1288
rect -429 -1322 -361 -1288
rect -271 -1322 -203 -1288
rect -113 -1322 -45 -1288
rect 45 -1322 113 -1288
rect 203 -1322 271 -1288
rect 361 -1322 429 -1288
rect 519 -1322 587 -1288
<< metal1 >>
rect -599 1322 -507 1328
rect -599 1288 -587 1322
rect -519 1288 -507 1322
rect -599 1282 -507 1288
rect -441 1322 -349 1328
rect -441 1288 -429 1322
rect -361 1288 -349 1322
rect -441 1282 -349 1288
rect -283 1322 -191 1328
rect -283 1288 -271 1322
rect -203 1288 -191 1322
rect -283 1282 -191 1288
rect -125 1322 -33 1328
rect -125 1288 -113 1322
rect -45 1288 -33 1322
rect -125 1282 -33 1288
rect 33 1322 125 1328
rect 33 1288 45 1322
rect 113 1288 125 1322
rect 33 1282 125 1288
rect 191 1322 283 1328
rect 191 1288 203 1322
rect 271 1288 283 1322
rect 191 1282 283 1288
rect 349 1322 441 1328
rect 349 1288 361 1322
rect 429 1288 441 1322
rect 349 1282 441 1288
rect 507 1322 599 1328
rect 507 1288 519 1322
rect 587 1288 599 1322
rect 507 1282 599 1288
rect -655 1238 -609 1250
rect -655 -1238 -649 1238
rect -615 -1238 -609 1238
rect -655 -1250 -609 -1238
rect -497 1238 -451 1250
rect -497 -1238 -491 1238
rect -457 -1238 -451 1238
rect -497 -1250 -451 -1238
rect -339 1238 -293 1250
rect -339 -1238 -333 1238
rect -299 -1238 -293 1238
rect -339 -1250 -293 -1238
rect -181 1238 -135 1250
rect -181 -1238 -175 1238
rect -141 -1238 -135 1238
rect -181 -1250 -135 -1238
rect -23 1238 23 1250
rect -23 -1238 -17 1238
rect 17 -1238 23 1238
rect -23 -1250 23 -1238
rect 135 1238 181 1250
rect 135 -1238 141 1238
rect 175 -1238 181 1238
rect 135 -1250 181 -1238
rect 293 1238 339 1250
rect 293 -1238 299 1238
rect 333 -1238 339 1238
rect 293 -1250 339 -1238
rect 451 1238 497 1250
rect 451 -1238 457 1238
rect 491 -1238 497 1238
rect 451 -1250 497 -1238
rect 609 1238 655 1250
rect 609 -1238 615 1238
rect 649 -1238 655 1238
rect 609 -1250 655 -1238
rect -599 -1288 -507 -1282
rect -599 -1322 -587 -1288
rect -519 -1322 -507 -1288
rect -599 -1328 -507 -1322
rect -441 -1288 -349 -1282
rect -441 -1322 -429 -1288
rect -361 -1322 -349 -1288
rect -441 -1328 -349 -1322
rect -283 -1288 -191 -1282
rect -283 -1322 -271 -1288
rect -203 -1322 -191 -1288
rect -283 -1328 -191 -1322
rect -125 -1288 -33 -1282
rect -125 -1322 -113 -1288
rect -45 -1322 -33 -1288
rect -125 -1328 -33 -1322
rect 33 -1288 125 -1282
rect 33 -1322 45 -1288
rect 113 -1322 125 -1288
rect 33 -1328 125 -1322
rect 191 -1288 283 -1282
rect 191 -1322 203 -1288
rect 271 -1322 283 -1288
rect 191 -1328 283 -1322
rect 349 -1288 441 -1282
rect 349 -1322 361 -1288
rect 429 -1322 441 -1288
rect 349 -1328 441 -1322
rect 507 -1288 599 -1282
rect 507 -1322 519 -1288
rect 587 -1322 599 -1288
rect 507 -1328 599 -1322
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 12.5 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
