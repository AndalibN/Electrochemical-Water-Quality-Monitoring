magic
tech sky130A
magscale 1 2
timestamp 1666965119
<< nwell >>
rect -523 -800 523 800
<< pmos >>
rect -429 -700 -29 700
rect 29 -700 429 700
<< pdiff >>
rect -487 688 -429 700
rect -487 -688 -475 688
rect -441 -688 -429 688
rect -487 -700 -429 -688
rect -29 688 29 700
rect -29 -688 -17 688
rect 17 -688 29 688
rect -29 -700 29 -688
rect 429 688 487 700
rect 429 -688 441 688
rect 475 -688 487 688
rect 429 -700 487 -688
<< pdiffc >>
rect -475 -688 -441 688
rect -17 -688 17 688
rect 441 -688 475 688
<< poly >>
rect -429 781 -29 797
rect -429 747 -413 781
rect -45 747 -29 781
rect -429 700 -29 747
rect 29 781 429 797
rect 29 747 45 781
rect 413 747 429 781
rect 29 700 429 747
rect -429 -747 -29 -700
rect -429 -781 -413 -747
rect -45 -781 -29 -747
rect -429 -797 -29 -781
rect 29 -747 429 -700
rect 29 -781 45 -747
rect 413 -781 429 -747
rect 29 -797 429 -781
<< polycont >>
rect -413 747 -45 781
rect 45 747 413 781
rect -413 -781 -45 -747
rect 45 -781 413 -747
<< locali >>
rect -429 747 -413 781
rect -45 747 -29 781
rect 29 747 45 781
rect 413 747 429 781
rect -475 688 -441 704
rect -475 -704 -441 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 441 688 475 704
rect 441 -704 475 -688
rect -429 -781 -413 -747
rect -45 -781 -29 -747
rect 29 -781 45 -747
rect 413 -781 429 -747
<< viali >>
rect -413 747 -45 781
rect 45 747 413 781
rect -475 -688 -441 688
rect -17 -688 17 688
rect 441 -688 475 688
rect -413 -781 -45 -747
rect 45 -781 413 -747
<< metal1 >>
rect -425 781 -33 787
rect -425 747 -413 781
rect -45 747 -33 781
rect -425 741 -33 747
rect 33 781 425 787
rect 33 747 45 781
rect 413 747 425 781
rect 33 741 425 747
rect -481 688 -435 700
rect -481 -688 -475 688
rect -441 -688 -435 688
rect -481 -700 -435 -688
rect -23 688 23 700
rect -23 -688 -17 688
rect 17 -688 23 688
rect -23 -700 23 -688
rect 435 688 481 700
rect 435 -688 441 688
rect 475 -688 481 688
rect 435 -700 481 -688
rect -425 -747 -33 -741
rect -425 -781 -413 -747
rect -45 -781 -33 -747
rect -425 -787 -33 -781
rect 33 -747 425 -741
rect 33 -781 45 -747
rect 413 -781 425 -747
rect 33 -787 425 -781
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 2.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
