magic
tech sky130A
magscale 1 2
timestamp 1667856991
<< error_p >>
rect -2588 2530 -2528 3670
rect -2508 2530 -2448 3670
rect -1329 2530 -1269 3670
rect -1249 2530 -1189 3670
rect -70 2530 -10 3670
rect 10 2530 70 3670
rect 1189 2530 1249 3670
rect 1269 2530 1329 3670
rect 2448 2530 2508 3670
rect 2528 2530 2588 3670
rect -2588 1290 -2528 2430
rect -2508 1290 -2448 2430
rect -1329 1290 -1269 2430
rect -1249 1290 -1189 2430
rect -70 1290 -10 2430
rect 10 1290 70 2430
rect 1189 1290 1249 2430
rect 1269 1290 1329 2430
rect 2448 1290 2508 2430
rect 2528 1290 2588 2430
rect -2588 50 -2528 1190
rect -2508 50 -2448 1190
rect -1329 50 -1269 1190
rect -1249 50 -1189 1190
rect -70 50 -10 1190
rect 10 50 70 1190
rect 1189 50 1249 1190
rect 1269 50 1329 1190
rect 2448 50 2508 1190
rect 2528 50 2588 1190
rect -2588 -1190 -2528 -50
rect -2508 -1190 -2448 -50
rect -1329 -1190 -1269 -50
rect -1249 -1190 -1189 -50
rect -70 -1190 -10 -50
rect 10 -1190 70 -50
rect 1189 -1190 1249 -50
rect 1269 -1190 1329 -50
rect 2448 -1190 2508 -50
rect 2528 -1190 2588 -50
rect -2588 -2430 -2528 -1290
rect -2508 -2430 -2448 -1290
rect -1329 -2430 -1269 -1290
rect -1249 -2430 -1189 -1290
rect -70 -2430 -10 -1290
rect 10 -2430 70 -1290
rect 1189 -2430 1249 -1290
rect 1269 -2430 1329 -1290
rect 2448 -2430 2508 -1290
rect 2528 -2430 2588 -1290
rect -2588 -3670 -2528 -2530
rect -2508 -3670 -2448 -2530
rect -1329 -3670 -1269 -2530
rect -1249 -3670 -1189 -2530
rect -70 -3670 -10 -2530
rect 10 -3670 70 -2530
rect 1189 -3670 1249 -2530
rect 1269 -3670 1329 -2530
rect 2448 -3670 2508 -2530
rect 2528 -3670 2588 -2530
<< metal3 >>
rect -3767 3642 -2528 3670
rect -3767 2558 -2612 3642
rect -2548 2558 -2528 3642
rect -3767 2530 -2528 2558
rect -2508 3642 -1269 3670
rect -2508 2558 -1353 3642
rect -1289 2558 -1269 3642
rect -2508 2530 -1269 2558
rect -1249 3642 -10 3670
rect -1249 2558 -94 3642
rect -30 2558 -10 3642
rect -1249 2530 -10 2558
rect 10 3642 1249 3670
rect 10 2558 1165 3642
rect 1229 2558 1249 3642
rect 10 2530 1249 2558
rect 1269 3642 2508 3670
rect 1269 2558 2424 3642
rect 2488 2558 2508 3642
rect 1269 2530 2508 2558
rect 2528 3642 3767 3670
rect 2528 2558 3683 3642
rect 3747 2558 3767 3642
rect 2528 2530 3767 2558
rect -3767 2402 -2528 2430
rect -3767 1318 -2612 2402
rect -2548 1318 -2528 2402
rect -3767 1290 -2528 1318
rect -2508 2402 -1269 2430
rect -2508 1318 -1353 2402
rect -1289 1318 -1269 2402
rect -2508 1290 -1269 1318
rect -1249 2402 -10 2430
rect -1249 1318 -94 2402
rect -30 1318 -10 2402
rect -1249 1290 -10 1318
rect 10 2402 1249 2430
rect 10 1318 1165 2402
rect 1229 1318 1249 2402
rect 10 1290 1249 1318
rect 1269 2402 2508 2430
rect 1269 1318 2424 2402
rect 2488 1318 2508 2402
rect 1269 1290 2508 1318
rect 2528 2402 3767 2430
rect 2528 1318 3683 2402
rect 3747 1318 3767 2402
rect 2528 1290 3767 1318
rect -3767 1162 -2528 1190
rect -3767 78 -2612 1162
rect -2548 78 -2528 1162
rect -3767 50 -2528 78
rect -2508 1162 -1269 1190
rect -2508 78 -1353 1162
rect -1289 78 -1269 1162
rect -2508 50 -1269 78
rect -1249 1162 -10 1190
rect -1249 78 -94 1162
rect -30 78 -10 1162
rect -1249 50 -10 78
rect 10 1162 1249 1190
rect 10 78 1165 1162
rect 1229 78 1249 1162
rect 10 50 1249 78
rect 1269 1162 2508 1190
rect 1269 78 2424 1162
rect 2488 78 2508 1162
rect 1269 50 2508 78
rect 2528 1162 3767 1190
rect 2528 78 3683 1162
rect 3747 78 3767 1162
rect 2528 50 3767 78
rect -3767 -78 -2528 -50
rect -3767 -1162 -2612 -78
rect -2548 -1162 -2528 -78
rect -3767 -1190 -2528 -1162
rect -2508 -78 -1269 -50
rect -2508 -1162 -1353 -78
rect -1289 -1162 -1269 -78
rect -2508 -1190 -1269 -1162
rect -1249 -78 -10 -50
rect -1249 -1162 -94 -78
rect -30 -1162 -10 -78
rect -1249 -1190 -10 -1162
rect 10 -78 1249 -50
rect 10 -1162 1165 -78
rect 1229 -1162 1249 -78
rect 10 -1190 1249 -1162
rect 1269 -78 2508 -50
rect 1269 -1162 2424 -78
rect 2488 -1162 2508 -78
rect 1269 -1190 2508 -1162
rect 2528 -78 3767 -50
rect 2528 -1162 3683 -78
rect 3747 -1162 3767 -78
rect 2528 -1190 3767 -1162
rect -3767 -1318 -2528 -1290
rect -3767 -2402 -2612 -1318
rect -2548 -2402 -2528 -1318
rect -3767 -2430 -2528 -2402
rect -2508 -1318 -1269 -1290
rect -2508 -2402 -1353 -1318
rect -1289 -2402 -1269 -1318
rect -2508 -2430 -1269 -2402
rect -1249 -1318 -10 -1290
rect -1249 -2402 -94 -1318
rect -30 -2402 -10 -1318
rect -1249 -2430 -10 -2402
rect 10 -1318 1249 -1290
rect 10 -2402 1165 -1318
rect 1229 -2402 1249 -1318
rect 10 -2430 1249 -2402
rect 1269 -1318 2508 -1290
rect 1269 -2402 2424 -1318
rect 2488 -2402 2508 -1318
rect 1269 -2430 2508 -2402
rect 2528 -1318 3767 -1290
rect 2528 -2402 3683 -1318
rect 3747 -2402 3767 -1318
rect 2528 -2430 3767 -2402
rect -3767 -2558 -2528 -2530
rect -3767 -3642 -2612 -2558
rect -2548 -3642 -2528 -2558
rect -3767 -3670 -2528 -3642
rect -2508 -2558 -1269 -2530
rect -2508 -3642 -1353 -2558
rect -1289 -3642 -1269 -2558
rect -2508 -3670 -1269 -3642
rect -1249 -2558 -10 -2530
rect -1249 -3642 -94 -2558
rect -30 -3642 -10 -2558
rect -1249 -3670 -10 -3642
rect 10 -2558 1249 -2530
rect 10 -3642 1165 -2558
rect 1229 -3642 1249 -2558
rect 10 -3670 1249 -3642
rect 1269 -2558 2508 -2530
rect 1269 -3642 2424 -2558
rect 2488 -3642 2508 -2558
rect 1269 -3670 2508 -3642
rect 2528 -2558 3767 -2530
rect 2528 -3642 3683 -2558
rect 3747 -3642 3767 -2558
rect 2528 -3670 3767 -3642
<< via3 >>
rect -2612 2558 -2548 3642
rect -1353 2558 -1289 3642
rect -94 2558 -30 3642
rect 1165 2558 1229 3642
rect 2424 2558 2488 3642
rect 3683 2558 3747 3642
rect -2612 1318 -2548 2402
rect -1353 1318 -1289 2402
rect -94 1318 -30 2402
rect 1165 1318 1229 2402
rect 2424 1318 2488 2402
rect 3683 1318 3747 2402
rect -2612 78 -2548 1162
rect -1353 78 -1289 1162
rect -94 78 -30 1162
rect 1165 78 1229 1162
rect 2424 78 2488 1162
rect 3683 78 3747 1162
rect -2612 -1162 -2548 -78
rect -1353 -1162 -1289 -78
rect -94 -1162 -30 -78
rect 1165 -1162 1229 -78
rect 2424 -1162 2488 -78
rect 3683 -1162 3747 -78
rect -2612 -2402 -2548 -1318
rect -1353 -2402 -1289 -1318
rect -94 -2402 -30 -1318
rect 1165 -2402 1229 -1318
rect 2424 -2402 2488 -1318
rect 3683 -2402 3747 -1318
rect -2612 -3642 -2548 -2558
rect -1353 -3642 -1289 -2558
rect -94 -3642 -30 -2558
rect 1165 -3642 1229 -2558
rect 2424 -3642 2488 -2558
rect 3683 -3642 3747 -2558
<< mimcap >>
rect -3667 3530 -2727 3570
rect -3667 2670 -3627 3530
rect -2767 2670 -2727 3530
rect -3667 2630 -2727 2670
rect -2408 3530 -1468 3570
rect -2408 2670 -2368 3530
rect -1508 2670 -1468 3530
rect -2408 2630 -1468 2670
rect -1149 3530 -209 3570
rect -1149 2670 -1109 3530
rect -249 2670 -209 3530
rect -1149 2630 -209 2670
rect 110 3530 1050 3570
rect 110 2670 150 3530
rect 1010 2670 1050 3530
rect 110 2630 1050 2670
rect 1369 3530 2309 3570
rect 1369 2670 1409 3530
rect 2269 2670 2309 3530
rect 1369 2630 2309 2670
rect 2628 3530 3568 3570
rect 2628 2670 2668 3530
rect 3528 2670 3568 3530
rect 2628 2630 3568 2670
rect -3667 2290 -2727 2330
rect -3667 1430 -3627 2290
rect -2767 1430 -2727 2290
rect -3667 1390 -2727 1430
rect -2408 2290 -1468 2330
rect -2408 1430 -2368 2290
rect -1508 1430 -1468 2290
rect -2408 1390 -1468 1430
rect -1149 2290 -209 2330
rect -1149 1430 -1109 2290
rect -249 1430 -209 2290
rect -1149 1390 -209 1430
rect 110 2290 1050 2330
rect 110 1430 150 2290
rect 1010 1430 1050 2290
rect 110 1390 1050 1430
rect 1369 2290 2309 2330
rect 1369 1430 1409 2290
rect 2269 1430 2309 2290
rect 1369 1390 2309 1430
rect 2628 2290 3568 2330
rect 2628 1430 2668 2290
rect 3528 1430 3568 2290
rect 2628 1390 3568 1430
rect -3667 1050 -2727 1090
rect -3667 190 -3627 1050
rect -2767 190 -2727 1050
rect -3667 150 -2727 190
rect -2408 1050 -1468 1090
rect -2408 190 -2368 1050
rect -1508 190 -1468 1050
rect -2408 150 -1468 190
rect -1149 1050 -209 1090
rect -1149 190 -1109 1050
rect -249 190 -209 1050
rect -1149 150 -209 190
rect 110 1050 1050 1090
rect 110 190 150 1050
rect 1010 190 1050 1050
rect 110 150 1050 190
rect 1369 1050 2309 1090
rect 1369 190 1409 1050
rect 2269 190 2309 1050
rect 1369 150 2309 190
rect 2628 1050 3568 1090
rect 2628 190 2668 1050
rect 3528 190 3568 1050
rect 2628 150 3568 190
rect -3667 -190 -2727 -150
rect -3667 -1050 -3627 -190
rect -2767 -1050 -2727 -190
rect -3667 -1090 -2727 -1050
rect -2408 -190 -1468 -150
rect -2408 -1050 -2368 -190
rect -1508 -1050 -1468 -190
rect -2408 -1090 -1468 -1050
rect -1149 -190 -209 -150
rect -1149 -1050 -1109 -190
rect -249 -1050 -209 -190
rect -1149 -1090 -209 -1050
rect 110 -190 1050 -150
rect 110 -1050 150 -190
rect 1010 -1050 1050 -190
rect 110 -1090 1050 -1050
rect 1369 -190 2309 -150
rect 1369 -1050 1409 -190
rect 2269 -1050 2309 -190
rect 1369 -1090 2309 -1050
rect 2628 -190 3568 -150
rect 2628 -1050 2668 -190
rect 3528 -1050 3568 -190
rect 2628 -1090 3568 -1050
rect -3667 -1430 -2727 -1390
rect -3667 -2290 -3627 -1430
rect -2767 -2290 -2727 -1430
rect -3667 -2330 -2727 -2290
rect -2408 -1430 -1468 -1390
rect -2408 -2290 -2368 -1430
rect -1508 -2290 -1468 -1430
rect -2408 -2330 -1468 -2290
rect -1149 -1430 -209 -1390
rect -1149 -2290 -1109 -1430
rect -249 -2290 -209 -1430
rect -1149 -2330 -209 -2290
rect 110 -1430 1050 -1390
rect 110 -2290 150 -1430
rect 1010 -2290 1050 -1430
rect 110 -2330 1050 -2290
rect 1369 -1430 2309 -1390
rect 1369 -2290 1409 -1430
rect 2269 -2290 2309 -1430
rect 1369 -2330 2309 -2290
rect 2628 -1430 3568 -1390
rect 2628 -2290 2668 -1430
rect 3528 -2290 3568 -1430
rect 2628 -2330 3568 -2290
rect -3667 -2670 -2727 -2630
rect -3667 -3530 -3627 -2670
rect -2767 -3530 -2727 -2670
rect -3667 -3570 -2727 -3530
rect -2408 -2670 -1468 -2630
rect -2408 -3530 -2368 -2670
rect -1508 -3530 -1468 -2670
rect -2408 -3570 -1468 -3530
rect -1149 -2670 -209 -2630
rect -1149 -3530 -1109 -2670
rect -249 -3530 -209 -2670
rect -1149 -3570 -209 -3530
rect 110 -2670 1050 -2630
rect 110 -3530 150 -2670
rect 1010 -3530 1050 -2670
rect 110 -3570 1050 -3530
rect 1369 -2670 2309 -2630
rect 1369 -3530 1409 -2670
rect 2269 -3530 2309 -2670
rect 1369 -3570 2309 -3530
rect 2628 -2670 3568 -2630
rect 2628 -3530 2668 -2670
rect 3528 -3530 3568 -2670
rect 2628 -3570 3568 -3530
<< mimcapcontact >>
rect -3627 2670 -2767 3530
rect -2368 2670 -1508 3530
rect -1109 2670 -249 3530
rect 150 2670 1010 3530
rect 1409 2670 2269 3530
rect 2668 2670 3528 3530
rect -3627 1430 -2767 2290
rect -2368 1430 -1508 2290
rect -1109 1430 -249 2290
rect 150 1430 1010 2290
rect 1409 1430 2269 2290
rect 2668 1430 3528 2290
rect -3627 190 -2767 1050
rect -2368 190 -1508 1050
rect -1109 190 -249 1050
rect 150 190 1010 1050
rect 1409 190 2269 1050
rect 2668 190 3528 1050
rect -3627 -1050 -2767 -190
rect -2368 -1050 -1508 -190
rect -1109 -1050 -249 -190
rect 150 -1050 1010 -190
rect 1409 -1050 2269 -190
rect 2668 -1050 3528 -190
rect -3627 -2290 -2767 -1430
rect -2368 -2290 -1508 -1430
rect -1109 -2290 -249 -1430
rect 150 -2290 1010 -1430
rect 1409 -2290 2269 -1430
rect 2668 -2290 3528 -1430
rect -3627 -3530 -2767 -2670
rect -2368 -3530 -1508 -2670
rect -1109 -3530 -249 -2670
rect 150 -3530 1010 -2670
rect 1409 -3530 2269 -2670
rect 2668 -3530 3528 -2670
<< metal4 >>
rect -3249 3531 -3145 3720
rect -2659 3658 -2555 3720
rect -2659 3642 -2532 3658
rect -3628 3530 -2766 3531
rect -3628 2670 -3627 3530
rect -2767 2670 -2766 3530
rect -3628 2669 -2766 2670
rect -3249 2291 -3145 2669
rect -2659 2558 -2612 3642
rect -2548 2558 -2532 3642
rect -1990 3531 -1886 3720
rect -1400 3658 -1296 3720
rect -1400 3642 -1273 3658
rect -2369 3530 -1507 3531
rect -2369 2670 -2368 3530
rect -1508 2670 -1507 3530
rect -2369 2669 -1507 2670
rect -2659 2542 -2532 2558
rect -2659 2418 -2555 2542
rect -2659 2402 -2532 2418
rect -3628 2290 -2766 2291
rect -3628 1430 -3627 2290
rect -2767 1430 -2766 2290
rect -3628 1429 -2766 1430
rect -3249 1051 -3145 1429
rect -2659 1318 -2612 2402
rect -2548 1318 -2532 2402
rect -1990 2291 -1886 2669
rect -1400 2558 -1353 3642
rect -1289 2558 -1273 3642
rect -731 3531 -627 3720
rect -141 3658 -37 3720
rect -141 3642 -14 3658
rect -1110 3530 -248 3531
rect -1110 2670 -1109 3530
rect -249 2670 -248 3530
rect -1110 2669 -248 2670
rect -1400 2542 -1273 2558
rect -1400 2418 -1296 2542
rect -1400 2402 -1273 2418
rect -2369 2290 -1507 2291
rect -2369 1430 -2368 2290
rect -1508 1430 -1507 2290
rect -2369 1429 -1507 1430
rect -2659 1302 -2532 1318
rect -2659 1178 -2555 1302
rect -2659 1162 -2532 1178
rect -3628 1050 -2766 1051
rect -3628 190 -3627 1050
rect -2767 190 -2766 1050
rect -3628 189 -2766 190
rect -3249 -189 -3145 189
rect -2659 78 -2612 1162
rect -2548 78 -2532 1162
rect -1990 1051 -1886 1429
rect -1400 1318 -1353 2402
rect -1289 1318 -1273 2402
rect -731 2291 -627 2669
rect -141 2558 -94 3642
rect -30 2558 -14 3642
rect 528 3531 632 3720
rect 1118 3658 1222 3720
rect 1118 3642 1245 3658
rect 149 3530 1011 3531
rect 149 2670 150 3530
rect 1010 2670 1011 3530
rect 149 2669 1011 2670
rect -141 2542 -14 2558
rect -141 2418 -37 2542
rect -141 2402 -14 2418
rect -1110 2290 -248 2291
rect -1110 1430 -1109 2290
rect -249 1430 -248 2290
rect -1110 1429 -248 1430
rect -1400 1302 -1273 1318
rect -1400 1178 -1296 1302
rect -1400 1162 -1273 1178
rect -2369 1050 -1507 1051
rect -2369 190 -2368 1050
rect -1508 190 -1507 1050
rect -2369 189 -1507 190
rect -2659 62 -2532 78
rect -2659 -62 -2555 62
rect -2659 -78 -2532 -62
rect -3628 -190 -2766 -189
rect -3628 -1050 -3627 -190
rect -2767 -1050 -2766 -190
rect -3628 -1051 -2766 -1050
rect -3249 -1429 -3145 -1051
rect -2659 -1162 -2612 -78
rect -2548 -1162 -2532 -78
rect -1990 -189 -1886 189
rect -1400 78 -1353 1162
rect -1289 78 -1273 1162
rect -731 1051 -627 1429
rect -141 1318 -94 2402
rect -30 1318 -14 2402
rect 528 2291 632 2669
rect 1118 2558 1165 3642
rect 1229 2558 1245 3642
rect 1787 3531 1891 3720
rect 2377 3658 2481 3720
rect 2377 3642 2504 3658
rect 1408 3530 2270 3531
rect 1408 2670 1409 3530
rect 2269 2670 2270 3530
rect 1408 2669 2270 2670
rect 1118 2542 1245 2558
rect 1118 2418 1222 2542
rect 1118 2402 1245 2418
rect 149 2290 1011 2291
rect 149 1430 150 2290
rect 1010 1430 1011 2290
rect 149 1429 1011 1430
rect -141 1302 -14 1318
rect -141 1178 -37 1302
rect -141 1162 -14 1178
rect -1110 1050 -248 1051
rect -1110 190 -1109 1050
rect -249 190 -248 1050
rect -1110 189 -248 190
rect -1400 62 -1273 78
rect -1400 -62 -1296 62
rect -1400 -78 -1273 -62
rect -2369 -190 -1507 -189
rect -2369 -1050 -2368 -190
rect -1508 -1050 -1507 -190
rect -2369 -1051 -1507 -1050
rect -2659 -1178 -2532 -1162
rect -2659 -1302 -2555 -1178
rect -2659 -1318 -2532 -1302
rect -3628 -1430 -2766 -1429
rect -3628 -2290 -3627 -1430
rect -2767 -2290 -2766 -1430
rect -3628 -2291 -2766 -2290
rect -3249 -2669 -3145 -2291
rect -2659 -2402 -2612 -1318
rect -2548 -2402 -2532 -1318
rect -1990 -1429 -1886 -1051
rect -1400 -1162 -1353 -78
rect -1289 -1162 -1273 -78
rect -731 -189 -627 189
rect -141 78 -94 1162
rect -30 78 -14 1162
rect 528 1051 632 1429
rect 1118 1318 1165 2402
rect 1229 1318 1245 2402
rect 1787 2291 1891 2669
rect 2377 2558 2424 3642
rect 2488 2558 2504 3642
rect 3046 3531 3150 3720
rect 3636 3658 3740 3720
rect 3636 3642 3763 3658
rect 2667 3530 3529 3531
rect 2667 2670 2668 3530
rect 3528 2670 3529 3530
rect 2667 2669 3529 2670
rect 2377 2542 2504 2558
rect 2377 2418 2481 2542
rect 2377 2402 2504 2418
rect 1408 2290 2270 2291
rect 1408 1430 1409 2290
rect 2269 1430 2270 2290
rect 1408 1429 2270 1430
rect 1118 1302 1245 1318
rect 1118 1178 1222 1302
rect 1118 1162 1245 1178
rect 149 1050 1011 1051
rect 149 190 150 1050
rect 1010 190 1011 1050
rect 149 189 1011 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -1110 -190 -248 -189
rect -1110 -1050 -1109 -190
rect -249 -1050 -248 -190
rect -1110 -1051 -248 -1050
rect -1400 -1178 -1273 -1162
rect -1400 -1302 -1296 -1178
rect -1400 -1318 -1273 -1302
rect -2369 -1430 -1507 -1429
rect -2369 -2290 -2368 -1430
rect -1508 -2290 -1507 -1430
rect -2369 -2291 -1507 -2290
rect -2659 -2418 -2532 -2402
rect -2659 -2542 -2555 -2418
rect -2659 -2558 -2532 -2542
rect -3628 -2670 -2766 -2669
rect -3628 -3530 -3627 -2670
rect -2767 -3530 -2766 -2670
rect -3628 -3531 -2766 -3530
rect -3249 -3720 -3145 -3531
rect -2659 -3642 -2612 -2558
rect -2548 -3642 -2532 -2558
rect -1990 -2669 -1886 -2291
rect -1400 -2402 -1353 -1318
rect -1289 -2402 -1273 -1318
rect -731 -1429 -627 -1051
rect -141 -1162 -94 -78
rect -30 -1162 -14 -78
rect 528 -189 632 189
rect 1118 78 1165 1162
rect 1229 78 1245 1162
rect 1787 1051 1891 1429
rect 2377 1318 2424 2402
rect 2488 1318 2504 2402
rect 3046 2291 3150 2669
rect 3636 2558 3683 3642
rect 3747 2558 3763 3642
rect 3636 2542 3763 2558
rect 3636 2418 3740 2542
rect 3636 2402 3763 2418
rect 2667 2290 3529 2291
rect 2667 1430 2668 2290
rect 3528 1430 3529 2290
rect 2667 1429 3529 1430
rect 2377 1302 2504 1318
rect 2377 1178 2481 1302
rect 2377 1162 2504 1178
rect 1408 1050 2270 1051
rect 1408 190 1409 1050
rect 2269 190 2270 1050
rect 1408 189 2270 190
rect 1118 62 1245 78
rect 1118 -62 1222 62
rect 1118 -78 1245 -62
rect 149 -190 1011 -189
rect 149 -1050 150 -190
rect 1010 -1050 1011 -190
rect 149 -1051 1011 -1050
rect -141 -1178 -14 -1162
rect -141 -1302 -37 -1178
rect -141 -1318 -14 -1302
rect -1110 -1430 -248 -1429
rect -1110 -2290 -1109 -1430
rect -249 -2290 -248 -1430
rect -1110 -2291 -248 -2290
rect -1400 -2418 -1273 -2402
rect -1400 -2542 -1296 -2418
rect -1400 -2558 -1273 -2542
rect -2369 -2670 -1507 -2669
rect -2369 -3530 -2368 -2670
rect -1508 -3530 -1507 -2670
rect -2369 -3531 -1507 -3530
rect -2659 -3658 -2532 -3642
rect -2659 -3720 -2555 -3658
rect -1990 -3720 -1886 -3531
rect -1400 -3642 -1353 -2558
rect -1289 -3642 -1273 -2558
rect -731 -2669 -627 -2291
rect -141 -2402 -94 -1318
rect -30 -2402 -14 -1318
rect 528 -1429 632 -1051
rect 1118 -1162 1165 -78
rect 1229 -1162 1245 -78
rect 1787 -189 1891 189
rect 2377 78 2424 1162
rect 2488 78 2504 1162
rect 3046 1051 3150 1429
rect 3636 1318 3683 2402
rect 3747 1318 3763 2402
rect 3636 1302 3763 1318
rect 3636 1178 3740 1302
rect 3636 1162 3763 1178
rect 2667 1050 3529 1051
rect 2667 190 2668 1050
rect 3528 190 3529 1050
rect 2667 189 3529 190
rect 2377 62 2504 78
rect 2377 -62 2481 62
rect 2377 -78 2504 -62
rect 1408 -190 2270 -189
rect 1408 -1050 1409 -190
rect 2269 -1050 2270 -190
rect 1408 -1051 2270 -1050
rect 1118 -1178 1245 -1162
rect 1118 -1302 1222 -1178
rect 1118 -1318 1245 -1302
rect 149 -1430 1011 -1429
rect 149 -2290 150 -1430
rect 1010 -2290 1011 -1430
rect 149 -2291 1011 -2290
rect -141 -2418 -14 -2402
rect -141 -2542 -37 -2418
rect -141 -2558 -14 -2542
rect -1110 -2670 -248 -2669
rect -1110 -3530 -1109 -2670
rect -249 -3530 -248 -2670
rect -1110 -3531 -248 -3530
rect -1400 -3658 -1273 -3642
rect -1400 -3720 -1296 -3658
rect -731 -3720 -627 -3531
rect -141 -3642 -94 -2558
rect -30 -3642 -14 -2558
rect 528 -2669 632 -2291
rect 1118 -2402 1165 -1318
rect 1229 -2402 1245 -1318
rect 1787 -1429 1891 -1051
rect 2377 -1162 2424 -78
rect 2488 -1162 2504 -78
rect 3046 -189 3150 189
rect 3636 78 3683 1162
rect 3747 78 3763 1162
rect 3636 62 3763 78
rect 3636 -62 3740 62
rect 3636 -78 3763 -62
rect 2667 -190 3529 -189
rect 2667 -1050 2668 -190
rect 3528 -1050 3529 -190
rect 2667 -1051 3529 -1050
rect 2377 -1178 2504 -1162
rect 2377 -1302 2481 -1178
rect 2377 -1318 2504 -1302
rect 1408 -1430 2270 -1429
rect 1408 -2290 1409 -1430
rect 2269 -2290 2270 -1430
rect 1408 -2291 2270 -2290
rect 1118 -2418 1245 -2402
rect 1118 -2542 1222 -2418
rect 1118 -2558 1245 -2542
rect 149 -2670 1011 -2669
rect 149 -3530 150 -2670
rect 1010 -3530 1011 -2670
rect 149 -3531 1011 -3530
rect -141 -3658 -14 -3642
rect -141 -3720 -37 -3658
rect 528 -3720 632 -3531
rect 1118 -3642 1165 -2558
rect 1229 -3642 1245 -2558
rect 1787 -2669 1891 -2291
rect 2377 -2402 2424 -1318
rect 2488 -2402 2504 -1318
rect 3046 -1429 3150 -1051
rect 3636 -1162 3683 -78
rect 3747 -1162 3763 -78
rect 3636 -1178 3763 -1162
rect 3636 -1302 3740 -1178
rect 3636 -1318 3763 -1302
rect 2667 -1430 3529 -1429
rect 2667 -2290 2668 -1430
rect 3528 -2290 3529 -1430
rect 2667 -2291 3529 -2290
rect 2377 -2418 2504 -2402
rect 2377 -2542 2481 -2418
rect 2377 -2558 2504 -2542
rect 1408 -2670 2270 -2669
rect 1408 -3530 1409 -2670
rect 2269 -3530 2270 -2670
rect 1408 -3531 2270 -3530
rect 1118 -3658 1245 -3642
rect 1118 -3720 1222 -3658
rect 1787 -3720 1891 -3531
rect 2377 -3642 2424 -2558
rect 2488 -3642 2504 -2558
rect 3046 -2669 3150 -2291
rect 3636 -2402 3683 -1318
rect 3747 -2402 3763 -1318
rect 3636 -2418 3763 -2402
rect 3636 -2542 3740 -2418
rect 3636 -2558 3763 -2542
rect 2667 -2670 3529 -2669
rect 2667 -3530 2668 -2670
rect 3528 -3530 3529 -2670
rect 2667 -3531 3529 -3530
rect 2377 -3658 2504 -3642
rect 2377 -3720 2481 -3658
rect 3046 -3720 3150 -3531
rect 3636 -3642 3683 -2558
rect 3747 -3642 3763 -2558
rect 3636 -3658 3763 -3642
rect 3636 -3720 3740 -3658
<< properties >>
string FIXED_BBOX 2528 2530 3668 3670
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.7 l 4.7 val 47.752 carea 2.00 cperi 0.19 nx 6 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
