magic
tech sky130A
magscale 1 2
timestamp 1668368552
<< error_p >>
rect -29 242579 29 242585
rect -29 242545 -17 242579
rect -29 242539 29 242545
rect -29 222469 29 222475
rect -29 222435 -17 222469
rect -29 222429 29 222435
rect -29 222361 29 222367
rect -29 222327 -17 222361
rect -29 222321 29 222327
rect -29 202251 29 202257
rect -29 202217 -17 202251
rect -29 202211 29 202217
rect -29 202143 29 202149
rect -29 202109 -17 202143
rect -29 202103 29 202109
rect -29 182033 29 182039
rect -29 181999 -17 182033
rect -29 181993 29 181999
rect -29 181925 29 181931
rect -29 181891 -17 181925
rect -29 181885 29 181891
rect -29 161815 29 161821
rect -29 161781 -17 161815
rect -29 161775 29 161781
rect -29 161707 29 161713
rect -29 161673 -17 161707
rect -29 161667 29 161673
rect -29 141597 29 141603
rect -29 141563 -17 141597
rect -29 141557 29 141563
rect -29 141489 29 141495
rect -29 141455 -17 141489
rect -29 141449 29 141455
rect -29 121379 29 121385
rect -29 121345 -17 121379
rect -29 121339 29 121345
rect -29 121271 29 121277
rect -29 121237 -17 121271
rect -29 121231 29 121237
rect -29 101161 29 101167
rect -29 101127 -17 101161
rect -29 101121 29 101127
rect -29 101053 29 101059
rect -29 101019 -17 101053
rect -29 101013 29 101019
rect -29 80943 29 80949
rect -29 80909 -17 80943
rect -29 80903 29 80909
rect -29 80835 29 80841
rect -29 80801 -17 80835
rect -29 80795 29 80801
rect -29 60725 29 60731
rect -29 60691 -17 60725
rect -29 60685 29 60691
rect -29 60617 29 60623
rect -29 60583 -17 60617
rect -29 60577 29 60583
rect -29 40507 29 40513
rect -29 40473 -17 40507
rect -29 40467 29 40473
rect -29 40399 29 40405
rect -29 40365 -17 40399
rect -29 40359 29 40365
rect -29 20289 29 20295
rect -29 20255 -17 20289
rect -29 20249 29 20255
rect -29 20181 29 20187
rect -29 20147 -17 20181
rect -29 20141 29 20147
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -20147 29 -20141
rect -29 -20181 -17 -20147
rect -29 -20187 29 -20181
rect -29 -20255 29 -20249
rect -29 -20289 -17 -20255
rect -29 -20295 29 -20289
rect -29 -40365 29 -40359
rect -29 -40399 -17 -40365
rect -29 -40405 29 -40399
rect -29 -40473 29 -40467
rect -29 -40507 -17 -40473
rect -29 -40513 29 -40507
rect -29 -60583 29 -60577
rect -29 -60617 -17 -60583
rect -29 -60623 29 -60617
rect -29 -60691 29 -60685
rect -29 -60725 -17 -60691
rect -29 -60731 29 -60725
rect -29 -80801 29 -80795
rect -29 -80835 -17 -80801
rect -29 -80841 29 -80835
rect -29 -80909 29 -80903
rect -29 -80943 -17 -80909
rect -29 -80949 29 -80943
rect -29 -101019 29 -101013
rect -29 -101053 -17 -101019
rect -29 -101059 29 -101053
rect -29 -101127 29 -101121
rect -29 -101161 -17 -101127
rect -29 -101167 29 -101161
rect -29 -121237 29 -121231
rect -29 -121271 -17 -121237
rect -29 -121277 29 -121271
rect -29 -121345 29 -121339
rect -29 -121379 -17 -121345
rect -29 -121385 29 -121379
rect -29 -141455 29 -141449
rect -29 -141489 -17 -141455
rect -29 -141495 29 -141489
rect -29 -141563 29 -141557
rect -29 -141597 -17 -141563
rect -29 -141603 29 -141597
rect -29 -161673 29 -161667
rect -29 -161707 -17 -161673
rect -29 -161713 29 -161707
rect -29 -161781 29 -161775
rect -29 -161815 -17 -161781
rect -29 -161821 29 -161815
rect -29 -181891 29 -181885
rect -29 -181925 -17 -181891
rect -29 -181931 29 -181925
rect -29 -181999 29 -181993
rect -29 -182033 -17 -181999
rect -29 -182039 29 -182033
rect -29 -202109 29 -202103
rect -29 -202143 -17 -202109
rect -29 -202149 29 -202143
rect -29 -202217 29 -202211
rect -29 -202251 -17 -202217
rect -29 -202257 29 -202251
rect -29 -222327 29 -222321
rect -29 -222361 -17 -222327
rect -29 -222367 29 -222361
rect -29 -222435 29 -222429
rect -29 -222469 -17 -222435
rect -29 -222475 29 -222469
rect -29 -242545 29 -242539
rect -29 -242579 -17 -242545
rect -29 -242585 29 -242579
<< pwell >>
rect -226 -242717 226 242717
<< nmos >>
rect -30 222507 30 242507
rect -30 202289 30 222289
rect -30 182071 30 202071
rect -30 161853 30 181853
rect -30 141635 30 161635
rect -30 121417 30 141417
rect -30 101199 30 121199
rect -30 80981 30 100981
rect -30 60763 30 80763
rect -30 40545 30 60545
rect -30 20327 30 40327
rect -30 109 30 20109
rect -30 -20109 30 -109
rect -30 -40327 30 -20327
rect -30 -60545 30 -40545
rect -30 -80763 30 -60763
rect -30 -100981 30 -80981
rect -30 -121199 30 -101199
rect -30 -141417 30 -121417
rect -30 -161635 30 -141635
rect -30 -181853 30 -161853
rect -30 -202071 30 -182071
rect -30 -222289 30 -202289
rect -30 -242507 30 -222507
<< ndiff >>
rect -88 242495 -30 242507
rect -88 222519 -76 242495
rect -42 222519 -30 242495
rect -88 222507 -30 222519
rect 30 242495 88 242507
rect 30 222519 42 242495
rect 76 222519 88 242495
rect 30 222507 88 222519
rect -88 222277 -30 222289
rect -88 202301 -76 222277
rect -42 202301 -30 222277
rect -88 202289 -30 202301
rect 30 222277 88 222289
rect 30 202301 42 222277
rect 76 202301 88 222277
rect 30 202289 88 202301
rect -88 202059 -30 202071
rect -88 182083 -76 202059
rect -42 182083 -30 202059
rect -88 182071 -30 182083
rect 30 202059 88 202071
rect 30 182083 42 202059
rect 76 182083 88 202059
rect 30 182071 88 182083
rect -88 181841 -30 181853
rect -88 161865 -76 181841
rect -42 161865 -30 181841
rect -88 161853 -30 161865
rect 30 181841 88 181853
rect 30 161865 42 181841
rect 76 161865 88 181841
rect 30 161853 88 161865
rect -88 161623 -30 161635
rect -88 141647 -76 161623
rect -42 141647 -30 161623
rect -88 141635 -30 141647
rect 30 161623 88 161635
rect 30 141647 42 161623
rect 76 141647 88 161623
rect 30 141635 88 141647
rect -88 141405 -30 141417
rect -88 121429 -76 141405
rect -42 121429 -30 141405
rect -88 121417 -30 121429
rect 30 141405 88 141417
rect 30 121429 42 141405
rect 76 121429 88 141405
rect 30 121417 88 121429
rect -88 121187 -30 121199
rect -88 101211 -76 121187
rect -42 101211 -30 121187
rect -88 101199 -30 101211
rect 30 121187 88 121199
rect 30 101211 42 121187
rect 76 101211 88 121187
rect 30 101199 88 101211
rect -88 100969 -30 100981
rect -88 80993 -76 100969
rect -42 80993 -30 100969
rect -88 80981 -30 80993
rect 30 100969 88 100981
rect 30 80993 42 100969
rect 76 80993 88 100969
rect 30 80981 88 80993
rect -88 80751 -30 80763
rect -88 60775 -76 80751
rect -42 60775 -30 80751
rect -88 60763 -30 60775
rect 30 80751 88 80763
rect 30 60775 42 80751
rect 76 60775 88 80751
rect 30 60763 88 60775
rect -88 60533 -30 60545
rect -88 40557 -76 60533
rect -42 40557 -30 60533
rect -88 40545 -30 40557
rect 30 60533 88 60545
rect 30 40557 42 60533
rect 76 40557 88 60533
rect 30 40545 88 40557
rect -88 40315 -30 40327
rect -88 20339 -76 40315
rect -42 20339 -30 40315
rect -88 20327 -30 20339
rect 30 40315 88 40327
rect 30 20339 42 40315
rect 76 20339 88 40315
rect 30 20327 88 20339
rect -88 20097 -30 20109
rect -88 121 -76 20097
rect -42 121 -30 20097
rect -88 109 -30 121
rect 30 20097 88 20109
rect 30 121 42 20097
rect 76 121 88 20097
rect 30 109 88 121
rect -88 -121 -30 -109
rect -88 -20097 -76 -121
rect -42 -20097 -30 -121
rect -88 -20109 -30 -20097
rect 30 -121 88 -109
rect 30 -20097 42 -121
rect 76 -20097 88 -121
rect 30 -20109 88 -20097
rect -88 -20339 -30 -20327
rect -88 -40315 -76 -20339
rect -42 -40315 -30 -20339
rect -88 -40327 -30 -40315
rect 30 -20339 88 -20327
rect 30 -40315 42 -20339
rect 76 -40315 88 -20339
rect 30 -40327 88 -40315
rect -88 -40557 -30 -40545
rect -88 -60533 -76 -40557
rect -42 -60533 -30 -40557
rect -88 -60545 -30 -60533
rect 30 -40557 88 -40545
rect 30 -60533 42 -40557
rect 76 -60533 88 -40557
rect 30 -60545 88 -60533
rect -88 -60775 -30 -60763
rect -88 -80751 -76 -60775
rect -42 -80751 -30 -60775
rect -88 -80763 -30 -80751
rect 30 -60775 88 -60763
rect 30 -80751 42 -60775
rect 76 -80751 88 -60775
rect 30 -80763 88 -80751
rect -88 -80993 -30 -80981
rect -88 -100969 -76 -80993
rect -42 -100969 -30 -80993
rect -88 -100981 -30 -100969
rect 30 -80993 88 -80981
rect 30 -100969 42 -80993
rect 76 -100969 88 -80993
rect 30 -100981 88 -100969
rect -88 -101211 -30 -101199
rect -88 -121187 -76 -101211
rect -42 -121187 -30 -101211
rect -88 -121199 -30 -121187
rect 30 -101211 88 -101199
rect 30 -121187 42 -101211
rect 76 -121187 88 -101211
rect 30 -121199 88 -121187
rect -88 -121429 -30 -121417
rect -88 -141405 -76 -121429
rect -42 -141405 -30 -121429
rect -88 -141417 -30 -141405
rect 30 -121429 88 -121417
rect 30 -141405 42 -121429
rect 76 -141405 88 -121429
rect 30 -141417 88 -141405
rect -88 -141647 -30 -141635
rect -88 -161623 -76 -141647
rect -42 -161623 -30 -141647
rect -88 -161635 -30 -161623
rect 30 -141647 88 -141635
rect 30 -161623 42 -141647
rect 76 -161623 88 -141647
rect 30 -161635 88 -161623
rect -88 -161865 -30 -161853
rect -88 -181841 -76 -161865
rect -42 -181841 -30 -161865
rect -88 -181853 -30 -181841
rect 30 -161865 88 -161853
rect 30 -181841 42 -161865
rect 76 -181841 88 -161865
rect 30 -181853 88 -181841
rect -88 -182083 -30 -182071
rect -88 -202059 -76 -182083
rect -42 -202059 -30 -182083
rect -88 -202071 -30 -202059
rect 30 -182083 88 -182071
rect 30 -202059 42 -182083
rect 76 -202059 88 -182083
rect 30 -202071 88 -202059
rect -88 -202301 -30 -202289
rect -88 -222277 -76 -202301
rect -42 -222277 -30 -202301
rect -88 -222289 -30 -222277
rect 30 -202301 88 -202289
rect 30 -222277 42 -202301
rect 76 -222277 88 -202301
rect 30 -222289 88 -222277
rect -88 -222519 -30 -222507
rect -88 -242495 -76 -222519
rect -42 -242495 -30 -222519
rect -88 -242507 -30 -242495
rect 30 -222519 88 -222507
rect 30 -242495 42 -222519
rect 76 -242495 88 -222519
rect 30 -242507 88 -242495
<< ndiffc >>
rect -76 222519 -42 242495
rect 42 222519 76 242495
rect -76 202301 -42 222277
rect 42 202301 76 222277
rect -76 182083 -42 202059
rect 42 182083 76 202059
rect -76 161865 -42 181841
rect 42 161865 76 181841
rect -76 141647 -42 161623
rect 42 141647 76 161623
rect -76 121429 -42 141405
rect 42 121429 76 141405
rect -76 101211 -42 121187
rect 42 101211 76 121187
rect -76 80993 -42 100969
rect 42 80993 76 100969
rect -76 60775 -42 80751
rect 42 60775 76 80751
rect -76 40557 -42 60533
rect 42 40557 76 60533
rect -76 20339 -42 40315
rect 42 20339 76 40315
rect -76 121 -42 20097
rect 42 121 76 20097
rect -76 -20097 -42 -121
rect 42 -20097 76 -121
rect -76 -40315 -42 -20339
rect 42 -40315 76 -20339
rect -76 -60533 -42 -40557
rect 42 -60533 76 -40557
rect -76 -80751 -42 -60775
rect 42 -80751 76 -60775
rect -76 -100969 -42 -80993
rect 42 -100969 76 -80993
rect -76 -121187 -42 -101211
rect 42 -121187 76 -101211
rect -76 -141405 -42 -121429
rect 42 -141405 76 -121429
rect -76 -161623 -42 -141647
rect 42 -161623 76 -141647
rect -76 -181841 -42 -161865
rect 42 -181841 76 -161865
rect -76 -202059 -42 -182083
rect 42 -202059 76 -182083
rect -76 -222277 -42 -202301
rect 42 -222277 76 -202301
rect -76 -242495 -42 -222519
rect 42 -242495 76 -222519
<< psubdiff >>
rect -190 242647 -94 242681
rect 94 242647 190 242681
rect -190 242585 -156 242647
rect 156 242585 190 242647
rect -190 -242647 -156 -242585
rect 156 -242647 190 -242585
rect -190 -242681 -94 -242647
rect 94 -242681 190 -242647
<< psubdiffcont >>
rect -94 242647 94 242681
rect -190 -242585 -156 242585
rect 156 -242585 190 242585
rect -94 -242681 94 -242647
<< poly >>
rect -33 242579 33 242595
rect -33 242545 -17 242579
rect 17 242545 33 242579
rect -33 242529 33 242545
rect -30 242507 30 242529
rect -30 222485 30 222507
rect -33 222469 33 222485
rect -33 222435 -17 222469
rect 17 222435 33 222469
rect -33 222419 33 222435
rect -33 222361 33 222377
rect -33 222327 -17 222361
rect 17 222327 33 222361
rect -33 222311 33 222327
rect -30 222289 30 222311
rect -30 202267 30 202289
rect -33 202251 33 202267
rect -33 202217 -17 202251
rect 17 202217 33 202251
rect -33 202201 33 202217
rect -33 202143 33 202159
rect -33 202109 -17 202143
rect 17 202109 33 202143
rect -33 202093 33 202109
rect -30 202071 30 202093
rect -30 182049 30 182071
rect -33 182033 33 182049
rect -33 181999 -17 182033
rect 17 181999 33 182033
rect -33 181983 33 181999
rect -33 181925 33 181941
rect -33 181891 -17 181925
rect 17 181891 33 181925
rect -33 181875 33 181891
rect -30 181853 30 181875
rect -30 161831 30 161853
rect -33 161815 33 161831
rect -33 161781 -17 161815
rect 17 161781 33 161815
rect -33 161765 33 161781
rect -33 161707 33 161723
rect -33 161673 -17 161707
rect 17 161673 33 161707
rect -33 161657 33 161673
rect -30 161635 30 161657
rect -30 141613 30 141635
rect -33 141597 33 141613
rect -33 141563 -17 141597
rect 17 141563 33 141597
rect -33 141547 33 141563
rect -33 141489 33 141505
rect -33 141455 -17 141489
rect 17 141455 33 141489
rect -33 141439 33 141455
rect -30 141417 30 141439
rect -30 121395 30 121417
rect -33 121379 33 121395
rect -33 121345 -17 121379
rect 17 121345 33 121379
rect -33 121329 33 121345
rect -33 121271 33 121287
rect -33 121237 -17 121271
rect 17 121237 33 121271
rect -33 121221 33 121237
rect -30 121199 30 121221
rect -30 101177 30 101199
rect -33 101161 33 101177
rect -33 101127 -17 101161
rect 17 101127 33 101161
rect -33 101111 33 101127
rect -33 101053 33 101069
rect -33 101019 -17 101053
rect 17 101019 33 101053
rect -33 101003 33 101019
rect -30 100981 30 101003
rect -30 80959 30 80981
rect -33 80943 33 80959
rect -33 80909 -17 80943
rect 17 80909 33 80943
rect -33 80893 33 80909
rect -33 80835 33 80851
rect -33 80801 -17 80835
rect 17 80801 33 80835
rect -33 80785 33 80801
rect -30 80763 30 80785
rect -30 60741 30 60763
rect -33 60725 33 60741
rect -33 60691 -17 60725
rect 17 60691 33 60725
rect -33 60675 33 60691
rect -33 60617 33 60633
rect -33 60583 -17 60617
rect 17 60583 33 60617
rect -33 60567 33 60583
rect -30 60545 30 60567
rect -30 40523 30 40545
rect -33 40507 33 40523
rect -33 40473 -17 40507
rect 17 40473 33 40507
rect -33 40457 33 40473
rect -33 40399 33 40415
rect -33 40365 -17 40399
rect 17 40365 33 40399
rect -33 40349 33 40365
rect -30 40327 30 40349
rect -30 20305 30 20327
rect -33 20289 33 20305
rect -33 20255 -17 20289
rect 17 20255 33 20289
rect -33 20239 33 20255
rect -33 20181 33 20197
rect -33 20147 -17 20181
rect 17 20147 33 20181
rect -33 20131 33 20147
rect -30 20109 30 20131
rect -30 87 30 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -109 30 -87
rect -30 -20131 30 -20109
rect -33 -20147 33 -20131
rect -33 -20181 -17 -20147
rect 17 -20181 33 -20147
rect -33 -20197 33 -20181
rect -33 -20255 33 -20239
rect -33 -20289 -17 -20255
rect 17 -20289 33 -20255
rect -33 -20305 33 -20289
rect -30 -20327 30 -20305
rect -30 -40349 30 -40327
rect -33 -40365 33 -40349
rect -33 -40399 -17 -40365
rect 17 -40399 33 -40365
rect -33 -40415 33 -40399
rect -33 -40473 33 -40457
rect -33 -40507 -17 -40473
rect 17 -40507 33 -40473
rect -33 -40523 33 -40507
rect -30 -40545 30 -40523
rect -30 -60567 30 -60545
rect -33 -60583 33 -60567
rect -33 -60617 -17 -60583
rect 17 -60617 33 -60583
rect -33 -60633 33 -60617
rect -33 -60691 33 -60675
rect -33 -60725 -17 -60691
rect 17 -60725 33 -60691
rect -33 -60741 33 -60725
rect -30 -60763 30 -60741
rect -30 -80785 30 -80763
rect -33 -80801 33 -80785
rect -33 -80835 -17 -80801
rect 17 -80835 33 -80801
rect -33 -80851 33 -80835
rect -33 -80909 33 -80893
rect -33 -80943 -17 -80909
rect 17 -80943 33 -80909
rect -33 -80959 33 -80943
rect -30 -80981 30 -80959
rect -30 -101003 30 -100981
rect -33 -101019 33 -101003
rect -33 -101053 -17 -101019
rect 17 -101053 33 -101019
rect -33 -101069 33 -101053
rect -33 -101127 33 -101111
rect -33 -101161 -17 -101127
rect 17 -101161 33 -101127
rect -33 -101177 33 -101161
rect -30 -101199 30 -101177
rect -30 -121221 30 -121199
rect -33 -121237 33 -121221
rect -33 -121271 -17 -121237
rect 17 -121271 33 -121237
rect -33 -121287 33 -121271
rect -33 -121345 33 -121329
rect -33 -121379 -17 -121345
rect 17 -121379 33 -121345
rect -33 -121395 33 -121379
rect -30 -121417 30 -121395
rect -30 -141439 30 -141417
rect -33 -141455 33 -141439
rect -33 -141489 -17 -141455
rect 17 -141489 33 -141455
rect -33 -141505 33 -141489
rect -33 -141563 33 -141547
rect -33 -141597 -17 -141563
rect 17 -141597 33 -141563
rect -33 -141613 33 -141597
rect -30 -141635 30 -141613
rect -30 -161657 30 -161635
rect -33 -161673 33 -161657
rect -33 -161707 -17 -161673
rect 17 -161707 33 -161673
rect -33 -161723 33 -161707
rect -33 -161781 33 -161765
rect -33 -161815 -17 -161781
rect 17 -161815 33 -161781
rect -33 -161831 33 -161815
rect -30 -161853 30 -161831
rect -30 -181875 30 -181853
rect -33 -181891 33 -181875
rect -33 -181925 -17 -181891
rect 17 -181925 33 -181891
rect -33 -181941 33 -181925
rect -33 -181999 33 -181983
rect -33 -182033 -17 -181999
rect 17 -182033 33 -181999
rect -33 -182049 33 -182033
rect -30 -182071 30 -182049
rect -30 -202093 30 -202071
rect -33 -202109 33 -202093
rect -33 -202143 -17 -202109
rect 17 -202143 33 -202109
rect -33 -202159 33 -202143
rect -33 -202217 33 -202201
rect -33 -202251 -17 -202217
rect 17 -202251 33 -202217
rect -33 -202267 33 -202251
rect -30 -202289 30 -202267
rect -30 -222311 30 -222289
rect -33 -222327 33 -222311
rect -33 -222361 -17 -222327
rect 17 -222361 33 -222327
rect -33 -222377 33 -222361
rect -33 -222435 33 -222419
rect -33 -222469 -17 -222435
rect 17 -222469 33 -222435
rect -33 -222485 33 -222469
rect -30 -222507 30 -222485
rect -30 -242529 30 -242507
rect -33 -242545 33 -242529
rect -33 -242579 -17 -242545
rect 17 -242579 33 -242545
rect -33 -242595 33 -242579
<< polycont >>
rect -17 242545 17 242579
rect -17 222435 17 222469
rect -17 222327 17 222361
rect -17 202217 17 202251
rect -17 202109 17 202143
rect -17 181999 17 182033
rect -17 181891 17 181925
rect -17 161781 17 161815
rect -17 161673 17 161707
rect -17 141563 17 141597
rect -17 141455 17 141489
rect -17 121345 17 121379
rect -17 121237 17 121271
rect -17 101127 17 101161
rect -17 101019 17 101053
rect -17 80909 17 80943
rect -17 80801 17 80835
rect -17 60691 17 60725
rect -17 60583 17 60617
rect -17 40473 17 40507
rect -17 40365 17 40399
rect -17 20255 17 20289
rect -17 20147 17 20181
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -20181 17 -20147
rect -17 -20289 17 -20255
rect -17 -40399 17 -40365
rect -17 -40507 17 -40473
rect -17 -60617 17 -60583
rect -17 -60725 17 -60691
rect -17 -80835 17 -80801
rect -17 -80943 17 -80909
rect -17 -101053 17 -101019
rect -17 -101161 17 -101127
rect -17 -121271 17 -121237
rect -17 -121379 17 -121345
rect -17 -141489 17 -141455
rect -17 -141597 17 -141563
rect -17 -161707 17 -161673
rect -17 -161815 17 -161781
rect -17 -181925 17 -181891
rect -17 -182033 17 -181999
rect -17 -202143 17 -202109
rect -17 -202251 17 -202217
rect -17 -222361 17 -222327
rect -17 -222469 17 -222435
rect -17 -242579 17 -242545
<< locali >>
rect -190 242647 -94 242681
rect 94 242647 190 242681
rect -190 242585 -156 242647
rect 156 242585 190 242647
rect -33 242545 -17 242579
rect 17 242545 33 242579
rect -76 242495 -42 242511
rect -76 222503 -42 222519
rect 42 242495 76 242511
rect 42 222503 76 222519
rect -33 222435 -17 222469
rect 17 222435 33 222469
rect -33 222327 -17 222361
rect 17 222327 33 222361
rect -76 222277 -42 222293
rect -76 202285 -42 202301
rect 42 222277 76 222293
rect 42 202285 76 202301
rect -33 202217 -17 202251
rect 17 202217 33 202251
rect -33 202109 -17 202143
rect 17 202109 33 202143
rect -76 202059 -42 202075
rect -76 182067 -42 182083
rect 42 202059 76 202075
rect 42 182067 76 182083
rect -33 181999 -17 182033
rect 17 181999 33 182033
rect -33 181891 -17 181925
rect 17 181891 33 181925
rect -76 181841 -42 181857
rect -76 161849 -42 161865
rect 42 181841 76 181857
rect 42 161849 76 161865
rect -33 161781 -17 161815
rect 17 161781 33 161815
rect -33 161673 -17 161707
rect 17 161673 33 161707
rect -76 161623 -42 161639
rect -76 141631 -42 141647
rect 42 161623 76 161639
rect 42 141631 76 141647
rect -33 141563 -17 141597
rect 17 141563 33 141597
rect -33 141455 -17 141489
rect 17 141455 33 141489
rect -76 141405 -42 141421
rect -76 121413 -42 121429
rect 42 141405 76 141421
rect 42 121413 76 121429
rect -33 121345 -17 121379
rect 17 121345 33 121379
rect -33 121237 -17 121271
rect 17 121237 33 121271
rect -76 121187 -42 121203
rect -76 101195 -42 101211
rect 42 121187 76 121203
rect 42 101195 76 101211
rect -33 101127 -17 101161
rect 17 101127 33 101161
rect -33 101019 -17 101053
rect 17 101019 33 101053
rect -76 100969 -42 100985
rect -76 80977 -42 80993
rect 42 100969 76 100985
rect 42 80977 76 80993
rect -33 80909 -17 80943
rect 17 80909 33 80943
rect -33 80801 -17 80835
rect 17 80801 33 80835
rect -76 80751 -42 80767
rect -76 60759 -42 60775
rect 42 80751 76 80767
rect 42 60759 76 60775
rect -33 60691 -17 60725
rect 17 60691 33 60725
rect -33 60583 -17 60617
rect 17 60583 33 60617
rect -76 60533 -42 60549
rect -76 40541 -42 40557
rect 42 60533 76 60549
rect 42 40541 76 40557
rect -33 40473 -17 40507
rect 17 40473 33 40507
rect -33 40365 -17 40399
rect 17 40365 33 40399
rect -76 40315 -42 40331
rect -76 20323 -42 20339
rect 42 40315 76 40331
rect 42 20323 76 20339
rect -33 20255 -17 20289
rect 17 20255 33 20289
rect -33 20147 -17 20181
rect 17 20147 33 20181
rect -76 20097 -42 20113
rect -76 105 -42 121
rect 42 20097 76 20113
rect 42 105 76 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -121 -42 -105
rect -76 -20113 -42 -20097
rect 42 -121 76 -105
rect 42 -20113 76 -20097
rect -33 -20181 -17 -20147
rect 17 -20181 33 -20147
rect -33 -20289 -17 -20255
rect 17 -20289 33 -20255
rect -76 -20339 -42 -20323
rect -76 -40331 -42 -40315
rect 42 -20339 76 -20323
rect 42 -40331 76 -40315
rect -33 -40399 -17 -40365
rect 17 -40399 33 -40365
rect -33 -40507 -17 -40473
rect 17 -40507 33 -40473
rect -76 -40557 -42 -40541
rect -76 -60549 -42 -60533
rect 42 -40557 76 -40541
rect 42 -60549 76 -60533
rect -33 -60617 -17 -60583
rect 17 -60617 33 -60583
rect -33 -60725 -17 -60691
rect 17 -60725 33 -60691
rect -76 -60775 -42 -60759
rect -76 -80767 -42 -80751
rect 42 -60775 76 -60759
rect 42 -80767 76 -80751
rect -33 -80835 -17 -80801
rect 17 -80835 33 -80801
rect -33 -80943 -17 -80909
rect 17 -80943 33 -80909
rect -76 -80993 -42 -80977
rect -76 -100985 -42 -100969
rect 42 -80993 76 -80977
rect 42 -100985 76 -100969
rect -33 -101053 -17 -101019
rect 17 -101053 33 -101019
rect -33 -101161 -17 -101127
rect 17 -101161 33 -101127
rect -76 -101211 -42 -101195
rect -76 -121203 -42 -121187
rect 42 -101211 76 -101195
rect 42 -121203 76 -121187
rect -33 -121271 -17 -121237
rect 17 -121271 33 -121237
rect -33 -121379 -17 -121345
rect 17 -121379 33 -121345
rect -76 -121429 -42 -121413
rect -76 -141421 -42 -141405
rect 42 -121429 76 -121413
rect 42 -141421 76 -141405
rect -33 -141489 -17 -141455
rect 17 -141489 33 -141455
rect -33 -141597 -17 -141563
rect 17 -141597 33 -141563
rect -76 -141647 -42 -141631
rect -76 -161639 -42 -161623
rect 42 -141647 76 -141631
rect 42 -161639 76 -161623
rect -33 -161707 -17 -161673
rect 17 -161707 33 -161673
rect -33 -161815 -17 -161781
rect 17 -161815 33 -161781
rect -76 -161865 -42 -161849
rect -76 -181857 -42 -181841
rect 42 -161865 76 -161849
rect 42 -181857 76 -181841
rect -33 -181925 -17 -181891
rect 17 -181925 33 -181891
rect -33 -182033 -17 -181999
rect 17 -182033 33 -181999
rect -76 -182083 -42 -182067
rect -76 -202075 -42 -202059
rect 42 -182083 76 -182067
rect 42 -202075 76 -202059
rect -33 -202143 -17 -202109
rect 17 -202143 33 -202109
rect -33 -202251 -17 -202217
rect 17 -202251 33 -202217
rect -76 -202301 -42 -202285
rect -76 -222293 -42 -222277
rect 42 -202301 76 -202285
rect 42 -222293 76 -222277
rect -33 -222361 -17 -222327
rect 17 -222361 33 -222327
rect -33 -222469 -17 -222435
rect 17 -222469 33 -222435
rect -76 -222519 -42 -222503
rect -76 -242511 -42 -242495
rect 42 -222519 76 -222503
rect 42 -242511 76 -242495
rect -33 -242579 -17 -242545
rect 17 -242579 33 -242545
rect -190 -242647 -156 -242585
rect 156 -242647 190 -242585
rect -190 -242681 -94 -242647
rect 94 -242681 190 -242647
<< viali >>
rect -17 242545 17 242579
rect -76 222519 -42 242495
rect 42 222519 76 242495
rect -17 222435 17 222469
rect -17 222327 17 222361
rect -76 202301 -42 222277
rect 42 202301 76 222277
rect -17 202217 17 202251
rect -17 202109 17 202143
rect -76 182083 -42 202059
rect 42 182083 76 202059
rect -17 181999 17 182033
rect -17 181891 17 181925
rect -76 161865 -42 181841
rect 42 161865 76 181841
rect -17 161781 17 161815
rect -17 161673 17 161707
rect -76 141647 -42 161623
rect 42 141647 76 161623
rect -17 141563 17 141597
rect -17 141455 17 141489
rect -76 121429 -42 141405
rect 42 121429 76 141405
rect -17 121345 17 121379
rect -17 121237 17 121271
rect -76 101211 -42 121187
rect 42 101211 76 121187
rect -17 101127 17 101161
rect -17 101019 17 101053
rect -76 80993 -42 100969
rect 42 80993 76 100969
rect -17 80909 17 80943
rect -17 80801 17 80835
rect -76 60775 -42 80751
rect 42 60775 76 80751
rect -17 60691 17 60725
rect -17 60583 17 60617
rect -76 40557 -42 60533
rect 42 40557 76 60533
rect -17 40473 17 40507
rect -17 40365 17 40399
rect -76 20339 -42 40315
rect 42 20339 76 40315
rect -17 20255 17 20289
rect -17 20147 17 20181
rect -76 121 -42 20097
rect 42 121 76 20097
rect -17 37 17 71
rect -17 -71 17 -37
rect -76 -20097 -42 -121
rect 42 -20097 76 -121
rect -17 -20181 17 -20147
rect -17 -20289 17 -20255
rect -76 -40315 -42 -20339
rect 42 -40315 76 -20339
rect -17 -40399 17 -40365
rect -17 -40507 17 -40473
rect -76 -60533 -42 -40557
rect 42 -60533 76 -40557
rect -17 -60617 17 -60583
rect -17 -60725 17 -60691
rect -76 -80751 -42 -60775
rect 42 -80751 76 -60775
rect -17 -80835 17 -80801
rect -17 -80943 17 -80909
rect -76 -100969 -42 -80993
rect 42 -100969 76 -80993
rect -17 -101053 17 -101019
rect -17 -101161 17 -101127
rect -76 -121187 -42 -101211
rect 42 -121187 76 -101211
rect -17 -121271 17 -121237
rect -17 -121379 17 -121345
rect -76 -141405 -42 -121429
rect 42 -141405 76 -121429
rect -17 -141489 17 -141455
rect -17 -141597 17 -141563
rect -76 -161623 -42 -141647
rect 42 -161623 76 -141647
rect -17 -161707 17 -161673
rect -17 -161815 17 -161781
rect -76 -181841 -42 -161865
rect 42 -181841 76 -161865
rect -17 -181925 17 -181891
rect -17 -182033 17 -181999
rect -76 -202059 -42 -182083
rect 42 -202059 76 -182083
rect -17 -202143 17 -202109
rect -17 -202251 17 -202217
rect -76 -222277 -42 -202301
rect 42 -222277 76 -202301
rect -17 -222361 17 -222327
rect -17 -222469 17 -222435
rect -76 -242495 -42 -222519
rect 42 -242495 76 -222519
rect -17 -242579 17 -242545
<< metal1 >>
rect -29 242579 29 242585
rect -29 242545 -17 242579
rect 17 242545 29 242579
rect -29 242539 29 242545
rect -82 242495 -36 242507
rect -82 222519 -76 242495
rect -42 222519 -36 242495
rect -82 222507 -36 222519
rect 36 242495 82 242507
rect 36 222519 42 242495
rect 76 222519 82 242495
rect 36 222507 82 222519
rect -29 222469 29 222475
rect -29 222435 -17 222469
rect 17 222435 29 222469
rect -29 222429 29 222435
rect -29 222361 29 222367
rect -29 222327 -17 222361
rect 17 222327 29 222361
rect -29 222321 29 222327
rect -82 222277 -36 222289
rect -82 202301 -76 222277
rect -42 202301 -36 222277
rect -82 202289 -36 202301
rect 36 222277 82 222289
rect 36 202301 42 222277
rect 76 202301 82 222277
rect 36 202289 82 202301
rect -29 202251 29 202257
rect -29 202217 -17 202251
rect 17 202217 29 202251
rect -29 202211 29 202217
rect -29 202143 29 202149
rect -29 202109 -17 202143
rect 17 202109 29 202143
rect -29 202103 29 202109
rect -82 202059 -36 202071
rect -82 182083 -76 202059
rect -42 182083 -36 202059
rect -82 182071 -36 182083
rect 36 202059 82 202071
rect 36 182083 42 202059
rect 76 182083 82 202059
rect 36 182071 82 182083
rect -29 182033 29 182039
rect -29 181999 -17 182033
rect 17 181999 29 182033
rect -29 181993 29 181999
rect -29 181925 29 181931
rect -29 181891 -17 181925
rect 17 181891 29 181925
rect -29 181885 29 181891
rect -82 181841 -36 181853
rect -82 161865 -76 181841
rect -42 161865 -36 181841
rect -82 161853 -36 161865
rect 36 181841 82 181853
rect 36 161865 42 181841
rect 76 161865 82 181841
rect 36 161853 82 161865
rect -29 161815 29 161821
rect -29 161781 -17 161815
rect 17 161781 29 161815
rect -29 161775 29 161781
rect -29 161707 29 161713
rect -29 161673 -17 161707
rect 17 161673 29 161707
rect -29 161667 29 161673
rect -82 161623 -36 161635
rect -82 141647 -76 161623
rect -42 141647 -36 161623
rect -82 141635 -36 141647
rect 36 161623 82 161635
rect 36 141647 42 161623
rect 76 141647 82 161623
rect 36 141635 82 141647
rect -29 141597 29 141603
rect -29 141563 -17 141597
rect 17 141563 29 141597
rect -29 141557 29 141563
rect -29 141489 29 141495
rect -29 141455 -17 141489
rect 17 141455 29 141489
rect -29 141449 29 141455
rect -82 141405 -36 141417
rect -82 121429 -76 141405
rect -42 121429 -36 141405
rect -82 121417 -36 121429
rect 36 141405 82 141417
rect 36 121429 42 141405
rect 76 121429 82 141405
rect 36 121417 82 121429
rect -29 121379 29 121385
rect -29 121345 -17 121379
rect 17 121345 29 121379
rect -29 121339 29 121345
rect -29 121271 29 121277
rect -29 121237 -17 121271
rect 17 121237 29 121271
rect -29 121231 29 121237
rect -82 121187 -36 121199
rect -82 101211 -76 121187
rect -42 101211 -36 121187
rect -82 101199 -36 101211
rect 36 121187 82 121199
rect 36 101211 42 121187
rect 76 101211 82 121187
rect 36 101199 82 101211
rect -29 101161 29 101167
rect -29 101127 -17 101161
rect 17 101127 29 101161
rect -29 101121 29 101127
rect -29 101053 29 101059
rect -29 101019 -17 101053
rect 17 101019 29 101053
rect -29 101013 29 101019
rect -82 100969 -36 100981
rect -82 80993 -76 100969
rect -42 80993 -36 100969
rect -82 80981 -36 80993
rect 36 100969 82 100981
rect 36 80993 42 100969
rect 76 80993 82 100969
rect 36 80981 82 80993
rect -29 80943 29 80949
rect -29 80909 -17 80943
rect 17 80909 29 80943
rect -29 80903 29 80909
rect -29 80835 29 80841
rect -29 80801 -17 80835
rect 17 80801 29 80835
rect -29 80795 29 80801
rect -82 80751 -36 80763
rect -82 60775 -76 80751
rect -42 60775 -36 80751
rect -82 60763 -36 60775
rect 36 80751 82 80763
rect 36 60775 42 80751
rect 76 60775 82 80751
rect 36 60763 82 60775
rect -29 60725 29 60731
rect -29 60691 -17 60725
rect 17 60691 29 60725
rect -29 60685 29 60691
rect -29 60617 29 60623
rect -29 60583 -17 60617
rect 17 60583 29 60617
rect -29 60577 29 60583
rect -82 60533 -36 60545
rect -82 40557 -76 60533
rect -42 40557 -36 60533
rect -82 40545 -36 40557
rect 36 60533 82 60545
rect 36 40557 42 60533
rect 76 40557 82 60533
rect 36 40545 82 40557
rect -29 40507 29 40513
rect -29 40473 -17 40507
rect 17 40473 29 40507
rect -29 40467 29 40473
rect -29 40399 29 40405
rect -29 40365 -17 40399
rect 17 40365 29 40399
rect -29 40359 29 40365
rect -82 40315 -36 40327
rect -82 20339 -76 40315
rect -42 20339 -36 40315
rect -82 20327 -36 20339
rect 36 40315 82 40327
rect 36 20339 42 40315
rect 76 20339 82 40315
rect 36 20327 82 20339
rect -29 20289 29 20295
rect -29 20255 -17 20289
rect 17 20255 29 20289
rect -29 20249 29 20255
rect -29 20181 29 20187
rect -29 20147 -17 20181
rect 17 20147 29 20181
rect -29 20141 29 20147
rect -82 20097 -36 20109
rect -82 121 -76 20097
rect -42 121 -36 20097
rect -82 109 -36 121
rect 36 20097 82 20109
rect 36 121 42 20097
rect 76 121 82 20097
rect 36 109 82 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -121 -36 -109
rect -82 -20097 -76 -121
rect -42 -20097 -36 -121
rect -82 -20109 -36 -20097
rect 36 -121 82 -109
rect 36 -20097 42 -121
rect 76 -20097 82 -121
rect 36 -20109 82 -20097
rect -29 -20147 29 -20141
rect -29 -20181 -17 -20147
rect 17 -20181 29 -20147
rect -29 -20187 29 -20181
rect -29 -20255 29 -20249
rect -29 -20289 -17 -20255
rect 17 -20289 29 -20255
rect -29 -20295 29 -20289
rect -82 -20339 -36 -20327
rect -82 -40315 -76 -20339
rect -42 -40315 -36 -20339
rect -82 -40327 -36 -40315
rect 36 -20339 82 -20327
rect 36 -40315 42 -20339
rect 76 -40315 82 -20339
rect 36 -40327 82 -40315
rect -29 -40365 29 -40359
rect -29 -40399 -17 -40365
rect 17 -40399 29 -40365
rect -29 -40405 29 -40399
rect -29 -40473 29 -40467
rect -29 -40507 -17 -40473
rect 17 -40507 29 -40473
rect -29 -40513 29 -40507
rect -82 -40557 -36 -40545
rect -82 -60533 -76 -40557
rect -42 -60533 -36 -40557
rect -82 -60545 -36 -60533
rect 36 -40557 82 -40545
rect 36 -60533 42 -40557
rect 76 -60533 82 -40557
rect 36 -60545 82 -60533
rect -29 -60583 29 -60577
rect -29 -60617 -17 -60583
rect 17 -60617 29 -60583
rect -29 -60623 29 -60617
rect -29 -60691 29 -60685
rect -29 -60725 -17 -60691
rect 17 -60725 29 -60691
rect -29 -60731 29 -60725
rect -82 -60775 -36 -60763
rect -82 -80751 -76 -60775
rect -42 -80751 -36 -60775
rect -82 -80763 -36 -80751
rect 36 -60775 82 -60763
rect 36 -80751 42 -60775
rect 76 -80751 82 -60775
rect 36 -80763 82 -80751
rect -29 -80801 29 -80795
rect -29 -80835 -17 -80801
rect 17 -80835 29 -80801
rect -29 -80841 29 -80835
rect -29 -80909 29 -80903
rect -29 -80943 -17 -80909
rect 17 -80943 29 -80909
rect -29 -80949 29 -80943
rect -82 -80993 -36 -80981
rect -82 -100969 -76 -80993
rect -42 -100969 -36 -80993
rect -82 -100981 -36 -100969
rect 36 -80993 82 -80981
rect 36 -100969 42 -80993
rect 76 -100969 82 -80993
rect 36 -100981 82 -100969
rect -29 -101019 29 -101013
rect -29 -101053 -17 -101019
rect 17 -101053 29 -101019
rect -29 -101059 29 -101053
rect -29 -101127 29 -101121
rect -29 -101161 -17 -101127
rect 17 -101161 29 -101127
rect -29 -101167 29 -101161
rect -82 -101211 -36 -101199
rect -82 -121187 -76 -101211
rect -42 -121187 -36 -101211
rect -82 -121199 -36 -121187
rect 36 -101211 82 -101199
rect 36 -121187 42 -101211
rect 76 -121187 82 -101211
rect 36 -121199 82 -121187
rect -29 -121237 29 -121231
rect -29 -121271 -17 -121237
rect 17 -121271 29 -121237
rect -29 -121277 29 -121271
rect -29 -121345 29 -121339
rect -29 -121379 -17 -121345
rect 17 -121379 29 -121345
rect -29 -121385 29 -121379
rect -82 -121429 -36 -121417
rect -82 -141405 -76 -121429
rect -42 -141405 -36 -121429
rect -82 -141417 -36 -141405
rect 36 -121429 82 -121417
rect 36 -141405 42 -121429
rect 76 -141405 82 -121429
rect 36 -141417 82 -141405
rect -29 -141455 29 -141449
rect -29 -141489 -17 -141455
rect 17 -141489 29 -141455
rect -29 -141495 29 -141489
rect -29 -141563 29 -141557
rect -29 -141597 -17 -141563
rect 17 -141597 29 -141563
rect -29 -141603 29 -141597
rect -82 -141647 -36 -141635
rect -82 -161623 -76 -141647
rect -42 -161623 -36 -141647
rect -82 -161635 -36 -161623
rect 36 -141647 82 -141635
rect 36 -161623 42 -141647
rect 76 -161623 82 -141647
rect 36 -161635 82 -161623
rect -29 -161673 29 -161667
rect -29 -161707 -17 -161673
rect 17 -161707 29 -161673
rect -29 -161713 29 -161707
rect -29 -161781 29 -161775
rect -29 -161815 -17 -161781
rect 17 -161815 29 -161781
rect -29 -161821 29 -161815
rect -82 -161865 -36 -161853
rect -82 -181841 -76 -161865
rect -42 -181841 -36 -161865
rect -82 -181853 -36 -181841
rect 36 -161865 82 -161853
rect 36 -181841 42 -161865
rect 76 -181841 82 -161865
rect 36 -181853 82 -181841
rect -29 -181891 29 -181885
rect -29 -181925 -17 -181891
rect 17 -181925 29 -181891
rect -29 -181931 29 -181925
rect -29 -181999 29 -181993
rect -29 -182033 -17 -181999
rect 17 -182033 29 -181999
rect -29 -182039 29 -182033
rect -82 -182083 -36 -182071
rect -82 -202059 -76 -182083
rect -42 -202059 -36 -182083
rect -82 -202071 -36 -202059
rect 36 -182083 82 -182071
rect 36 -202059 42 -182083
rect 76 -202059 82 -182083
rect 36 -202071 82 -202059
rect -29 -202109 29 -202103
rect -29 -202143 -17 -202109
rect 17 -202143 29 -202109
rect -29 -202149 29 -202143
rect -29 -202217 29 -202211
rect -29 -202251 -17 -202217
rect 17 -202251 29 -202217
rect -29 -202257 29 -202251
rect -82 -202301 -36 -202289
rect -82 -222277 -76 -202301
rect -42 -222277 -36 -202301
rect -82 -222289 -36 -222277
rect 36 -202301 82 -202289
rect 36 -222277 42 -202301
rect 76 -222277 82 -202301
rect 36 -222289 82 -222277
rect -29 -222327 29 -222321
rect -29 -222361 -17 -222327
rect 17 -222361 29 -222327
rect -29 -222367 29 -222361
rect -29 -222435 29 -222429
rect -29 -222469 -17 -222435
rect 17 -222469 29 -222435
rect -29 -222475 29 -222469
rect -82 -222519 -36 -222507
rect -82 -242495 -76 -222519
rect -42 -242495 -36 -222519
rect -82 -242507 -36 -242495
rect 36 -222519 82 -222507
rect 36 -242495 42 -222519
rect 76 -242495 82 -222519
rect 36 -242507 82 -242495
rect -29 -242545 29 -242539
rect -29 -242579 -17 -242545
rect 17 -242579 29 -242545
rect -29 -242585 29 -242579
<< properties >>
string FIXED_BBOX -173 -242664 173 242664
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 100.0 l 0.3 m 24 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
