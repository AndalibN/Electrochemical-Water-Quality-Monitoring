magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -124 -302 124 302
<< pmos >>
rect -30 -240 30 240
<< pdiff >>
rect -88 221 -30 240
rect -88 187 -76 221
rect -42 187 -30 221
rect -88 153 -30 187
rect -88 119 -76 153
rect -42 119 -30 153
rect -88 85 -30 119
rect -88 51 -76 85
rect -42 51 -30 85
rect -88 17 -30 51
rect -88 -17 -76 17
rect -42 -17 -30 17
rect -88 -51 -30 -17
rect -88 -85 -76 -51
rect -42 -85 -30 -51
rect -88 -119 -30 -85
rect -88 -153 -76 -119
rect -42 -153 -30 -119
rect -88 -187 -30 -153
rect -88 -221 -76 -187
rect -42 -221 -30 -187
rect -88 -240 -30 -221
rect 30 221 88 240
rect 30 187 42 221
rect 76 187 88 221
rect 30 153 88 187
rect 30 119 42 153
rect 76 119 88 153
rect 30 85 88 119
rect 30 51 42 85
rect 76 51 88 85
rect 30 17 88 51
rect 30 -17 42 17
rect 76 -17 88 17
rect 30 -51 88 -17
rect 30 -85 42 -51
rect 76 -85 88 -51
rect 30 -119 88 -85
rect 30 -153 42 -119
rect 76 -153 88 -119
rect 30 -187 88 -153
rect 30 -221 42 -187
rect 76 -221 88 -187
rect 30 -240 88 -221
<< pdiffc >>
rect -76 187 -42 221
rect -76 119 -42 153
rect -76 51 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -51
rect -76 -153 -42 -119
rect -76 -221 -42 -187
rect 42 187 76 221
rect 42 119 76 153
rect 42 51 76 85
rect 42 -17 76 17
rect 42 -85 76 -51
rect 42 -153 76 -119
rect 42 -221 76 -187
<< poly >>
rect -30 240 30 266
rect -30 -266 30 -240
<< locali >>
rect -76 221 -42 244
rect -76 153 -42 163
rect -76 85 -42 91
rect -76 17 -42 19
rect -76 -19 -42 -17
rect -76 -91 -42 -85
rect -76 -163 -42 -153
rect -76 -244 -42 -221
rect 42 221 76 244
rect 42 153 76 163
rect 42 85 76 91
rect 42 17 76 19
rect 42 -19 76 -17
rect 42 -91 76 -85
rect 42 -163 76 -153
rect 42 -244 76 -221
<< viali >>
rect -76 187 -42 197
rect -76 163 -42 187
rect -76 119 -42 125
rect -76 91 -42 119
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect -76 -119 -42 -91
rect -76 -125 -42 -119
rect -76 -187 -42 -163
rect -76 -197 -42 -187
rect 42 187 76 197
rect 42 163 76 187
rect 42 119 76 125
rect 42 91 76 119
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect 42 -119 76 -91
rect 42 -125 76 -119
rect 42 -187 76 -163
rect 42 -197 76 -187
<< metal1 >>
rect -82 197 -36 240
rect -82 163 -76 197
rect -42 163 -36 197
rect -82 125 -36 163
rect -82 91 -76 125
rect -42 91 -36 125
rect -82 53 -36 91
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -91 -36 -53
rect -82 -125 -76 -91
rect -42 -125 -36 -91
rect -82 -163 -36 -125
rect -82 -197 -76 -163
rect -42 -197 -36 -163
rect -82 -240 -36 -197
rect 36 197 82 240
rect 36 163 42 197
rect 76 163 82 197
rect 36 125 82 163
rect 36 91 42 125
rect 76 91 82 125
rect 36 53 82 91
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -91 82 -53
rect 36 -125 42 -91
rect 76 -125 82 -91
rect 36 -163 82 -125
rect 36 -197 42 -163
rect 76 -197 82 -163
rect 36 -240 82 -197
<< end >>
