magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_s >>
rect 1512 -1016 1602 -1012
rect -250 -1053 -194 -1040
rect -48 -1053 220 -1040
rect 1540 -1044 1630 -1040
rect -302 -1149 -296 -1145
rect -244 -1149 -238 -1145
rect -296 -1155 -290 -1149
rect -250 -1155 -244 -1149
<< nwell >>
rect -2498 1724 1462 2367
rect -2498 -716 1465 1724
<< pwell >>
rect -2730 -3066 2164 -2588
<< psubdiff >>
rect -2704 -2640 2138 -2614
rect -2704 -3014 -2680 -2640
rect 2114 -3014 2138 -2640
rect -2704 -3040 2138 -3014
<< nsubdiff >>
rect -2383 2126 1387 2229
rect -2383 2024 -2232 2126
rect 1270 2024 1387 2126
rect -2383 1895 1387 2024
<< psubdiffcont >>
rect -2680 -3014 2114 -2640
<< nsubdiffcont >>
rect -2232 2024 1270 2126
<< poly >>
rect -2634 1869 -2562 1888
rect -2634 1835 -2616 1869
rect -2582 1846 -2562 1869
rect -2582 1835 -982 1846
rect -2634 1816 -982 1835
rect -2628 1772 -2556 1773
rect -2628 1754 -1304 1772
rect -2628 1720 -2610 1754
rect -2576 1742 -1304 1754
rect -2576 1720 -2556 1742
rect -2628 1701 -2556 1720
rect -1348 1640 -1304 1742
rect -1012 1549 -982 1816
rect -733 1742 -653 1746
rect -733 1728 712 1742
rect -733 1694 -709 1728
rect -675 1694 712 1728
rect -733 1685 712 1694
rect -733 1676 -653 1685
rect -250 1615 -170 1628
rect -250 1610 482 1615
rect -250 1608 -226 1610
rect -535 1576 -226 1608
rect -192 1576 482 1610
rect -535 1566 482 1576
rect -535 1506 -475 1566
rect -417 1506 -357 1566
rect -250 1558 -170 1566
rect 422 1436 482 1566
rect 652 1457 712 1685
rect -653 -508 -593 -460
rect -299 -508 -239 -460
rect 40 -508 364 -507
rect -653 -548 364 -508
rect 899 -597 1083 -550
rect -289 -1053 1169 -1023
rect -289 -1147 -250 -1053
rect 499 -1159 557 -1053
rect 1113 -1156 1169 -1053
rect -1358 -1863 -1065 -1807
rect -534 -1874 -472 -1813
rect 115 -1874 175 -1809
rect -534 -1922 175 -1874
rect 116 -1935 175 -1922
rect 883 -1935 926 -1820
rect 116 -1979 926 -1935
<< polycont >>
rect -2616 1835 -2582 1869
rect -2610 1720 -2576 1754
rect -709 1694 -675 1728
rect -226 1576 -192 1610
<< locali >>
rect -2310 2140 1335 2190
rect -2310 2139 -965 2140
rect -2310 2132 -1403 2139
rect -2310 2126 -1520 2132
rect -1486 2126 -1403 2132
rect -1369 2126 -965 2139
rect -931 2129 1335 2140
rect -931 2127 483 2129
rect -931 2126 128 2127
rect 162 2126 483 2127
rect 517 2127 1335 2129
rect 517 2126 603 2127
rect 637 2126 964 2127
rect 998 2126 1335 2127
rect -2310 2024 -2232 2126
rect 1270 2024 1335 2126
rect -2310 1948 1335 2024
rect -2634 1869 -2562 1888
rect -2634 1835 -2616 1869
rect -2582 1835 -2562 1869
rect -2634 1816 -2562 1835
rect -2628 1754 -2556 1773
rect -2628 1720 -2610 1754
rect -2576 1720 -2556 1754
rect -2628 1701 -2556 1720
rect -733 1728 -653 1746
rect -733 1694 -709 1728
rect -675 1694 -653 1728
rect -733 1676 -653 1694
rect -250 1610 -170 1628
rect -2186 1531 -1944 1585
rect -250 1576 -226 1610
rect -192 1576 -170 1610
rect -250 1558 -170 1576
rect -2002 -818 -1944 1531
rect -1342 -566 -1308 -483
rect 258 -566 292 1419
rect -1342 -600 292 -566
rect 258 -708 292 -600
rect 818 -514 888 44
rect 1092 -513 1163 29
rect 818 -610 864 -514
rect 812 -625 864 -610
rect 812 -626 872 -625
rect 812 -660 824 -626
rect 858 -660 872 -626
rect 812 -668 872 -660
rect 812 -673 864 -668
rect 915 -708 949 -557
rect 1117 -614 1163 -513
rect 1116 -628 1170 -614
rect 1116 -662 1124 -628
rect 1158 -662 1170 -628
rect 1116 -674 1170 -662
rect 258 -742 949 -708
rect -2003 -828 -1944 -818
rect -2003 -862 -1991 -828
rect -1957 -836 -1944 -828
rect -1957 -862 44 -836
rect -2003 -870 44 -862
rect -2003 -872 -1944 -870
rect 9 -988 44 -870
rect 9 -1022 427 -988
rect 9 -1146 44 -1022
rect 393 -1153 427 -1022
rect -1171 -1894 -1137 -1197
rect -935 -1755 -901 -1165
rect -960 -1789 -901 -1755
rect -699 -1750 -665 -1181
rect 794 -1184 836 -742
rect 934 -823 992 -809
rect 934 -857 946 -823
rect 980 -857 992 -823
rect 934 -870 992 -857
rect 1117 -813 1163 -674
rect 1323 -813 1394 -801
rect 1117 -824 1394 -813
rect 1117 -858 1337 -824
rect 1371 -858 1394 -824
rect 1117 -859 1394 -858
rect -699 -1789 -640 -1750
rect -227 -1771 -193 -1195
rect 794 -1467 863 -1184
rect 940 -1329 986 -870
rect 1323 -873 1394 -859
rect 1331 -914 1378 -873
rect 1332 -1130 1378 -914
rect 1332 -1264 1414 -1130
rect -960 -1894 -926 -1789
rect -674 -1894 -640 -1789
rect -1171 -1928 -640 -1894
rect -2696 -2640 2130 -2614
rect -2696 -3014 -2680 -2640
rect 2114 -3014 2130 -2640
rect -2696 -3040 2130 -3014
<< viali >>
rect -1520 2126 -1486 2132
rect -1403 2126 -1369 2139
rect -965 2126 -931 2140
rect 128 2126 162 2127
rect 483 2126 517 2129
rect 603 2126 637 2127
rect 964 2126 998 2127
rect -1707 2069 -1673 2103
rect -1520 2098 -1486 2126
rect -1403 2105 -1369 2126
rect -965 2106 -931 2126
rect -463 2092 -429 2126
rect 128 2093 162 2126
rect 483 2095 517 2126
rect 603 2093 637 2126
rect 964 2093 998 2126
rect 1229 2090 1263 2124
rect -2616 1835 -2582 1869
rect -2610 1720 -2576 1754
rect -709 1694 -675 1728
rect -226 1576 -192 1610
rect 824 -660 858 -626
rect 1124 -662 1158 -628
rect -1991 -862 -1957 -828
rect -287 -1140 -253 -1106
rect 946 -857 980 -823
rect 1337 -858 1371 -824
rect -2392 -2831 -2358 -2797
rect -1861 -2830 -1827 -2796
rect -1419 -2836 -1385 -2802
rect -1053 -2836 -1019 -2802
rect -234 -2831 -200 -2797
rect 582 -2834 616 -2800
rect 1205 -2827 1239 -2793
rect 1613 -2822 1647 -2788
rect 1882 -2818 1916 -2784
rect -2519 -2876 -2485 -2842
<< metal1 >>
rect -1539 2132 -1465 2145
rect -1726 2103 -1652 2116
rect -1726 2069 -1707 2103
rect -1673 2069 -1652 2103
rect -1539 2098 -1520 2132
rect -1486 2098 -1465 2132
rect -1539 2082 -1465 2098
rect -1422 2139 -1348 2152
rect -1422 2105 -1403 2139
rect -1369 2105 -1348 2139
rect -1422 2089 -1348 2105
rect -984 2140 -910 2153
rect -984 2106 -965 2140
rect -931 2106 -910 2140
rect -984 2090 -910 2106
rect -482 2126 -408 2139
rect -482 2092 -463 2126
rect -429 2092 -408 2126
rect -1726 2050 -1652 2069
rect -2634 1879 -2562 1888
rect -2634 1827 -2622 1879
rect -2570 1827 -2562 1879
rect -2634 1816 -2562 1827
rect -2628 1764 -2556 1773
rect -2628 1712 -2616 1764
rect -2564 1712 -2556 1764
rect -2628 1701 -2556 1712
rect -5586 1586 -5458 1618
rect -5586 1580 -5546 1586
rect -5638 1534 -5546 1580
rect -5494 1580 -5458 1586
rect -3928 1595 -3800 1618
rect -3928 1586 -3790 1595
rect -3928 1580 -3888 1586
rect -5494 1534 -3888 1580
rect -3836 1580 -3790 1586
rect -2190 1583 -2127 1584
rect -2309 1580 -2242 1581
rect -3836 1534 -2242 1580
rect -5638 1530 -2242 1534
rect -5586 1502 -5458 1530
rect -4711 1276 -4648 1530
rect -3928 1528 -2242 1530
rect -3928 1517 -3790 1528
rect -3928 1502 -3800 1517
rect -3059 1295 -2988 1528
rect -2190 1526 -2126 1583
rect -2189 1525 -2126 1526
rect -1702 1322 -1668 2050
rect -1517 1707 -1483 2082
rect -1530 1700 -1467 1707
rect -1530 1648 -1524 1700
rect -1472 1648 -1467 1700
rect -1530 1640 -1467 1648
rect -1401 1345 -1367 2089
rect -962 1493 -928 2090
rect -482 2076 -408 2092
rect 109 2127 183 2140
rect 109 2093 128 2127
rect 162 2093 183 2127
rect 109 2077 183 2093
rect 464 2129 538 2142
rect 464 2095 483 2129
rect 517 2095 538 2129
rect 464 2079 538 2095
rect 584 2127 658 2140
rect 584 2093 603 2127
rect 637 2093 658 2127
rect -733 1728 -653 1746
rect -733 1694 -709 1728
rect -675 1694 -653 1728
rect -733 1676 -653 1694
rect -699 1561 -665 1676
rect -888 1527 -665 1561
rect -962 1465 -913 1493
rect -947 1331 -913 1465
rect -4976 478 -4879 781
rect -3318 541 -3212 844
rect -4976 371 -4878 478
rect -5384 243 -5326 251
rect -4972 247 -4878 371
rect -5384 191 -5378 243
rect -5326 226 -5311 243
rect -5326 198 -5309 226
rect -5326 191 -5311 198
rect -5384 183 -5311 191
rect -4972 195 -4958 247
rect -4906 195 -4878 247
rect -5384 182 -5326 183
rect -5378 -2848 -5326 182
rect -4972 171 -4878 195
rect -5268 42 -5140 74
rect -5268 36 -5228 42
rect -5282 -10 -5228 36
rect -5176 36 -5140 42
rect -4714 40 -4645 456
rect -3314 261 -3220 541
rect -3314 209 -3292 261
rect -3240 209 -3220 261
rect -3314 182 -3220 209
rect -3610 42 -3482 74
rect -4716 36 -4644 40
rect -3610 36 -3570 42
rect -5176 -10 -4644 36
rect -5282 -14 -4644 -10
rect -3624 -10 -3570 36
rect -3518 36 -3482 42
rect -3059 68 -2988 430
rect -3059 36 -2986 68
rect -3518 -10 -2986 36
rect -3624 -14 -2986 -10
rect -5268 -42 -5140 -14
rect -4982 -876 -4925 -14
rect -4714 -21 -4645 -14
rect -3610 -42 -3482 -14
rect -3216 -724 -3145 -14
rect -2369 -41 -2323 -40
rect -2369 -198 -2320 -41
rect -3218 -730 -3145 -724
rect -3218 -782 -3212 -730
rect -3160 -782 -3145 -730
rect -3218 -788 -3145 -782
rect -3215 -791 -3145 -788
rect -2368 -390 -2320 -198
rect -4986 -883 -4915 -876
rect -4988 -889 -4915 -883
rect -4988 -941 -4982 -889
rect -4930 -941 -4915 -889
rect -4988 -947 -4915 -941
rect -4985 -950 -4915 -947
rect -4982 -957 -4925 -950
rect -2368 -1229 -2333 -390
rect -2236 -484 -2202 -264
rect -2237 -492 -2174 -484
rect -2237 -544 -2232 -492
rect -2180 -544 -2174 -492
rect -2237 -550 -2174 -544
rect -2118 -1187 -2083 -130
rect -1866 -395 -1787 0
rect -1866 -492 -1802 -395
rect -1290 -406 -1236 -94
rect -1774 -483 -1711 -427
rect -1866 -544 -1859 -492
rect -1807 -544 -1802 -492
rect -1866 -550 -1802 -544
rect -1772 -601 -1716 -483
rect -1358 -496 -1292 -434
rect -1264 -524 -1236 -406
rect -1065 -474 -1031 612
rect -829 -474 -795 -145
rect -1065 -507 -783 -474
rect -1283 -550 -1236 -524
rect -1775 -612 -1711 -601
rect -1775 -664 -1768 -612
rect -1716 -664 -1711 -612
rect -1775 -670 -1711 -664
rect -2010 -810 -1938 -809
rect -2012 -816 -1938 -810
rect -2012 -868 -2000 -816
rect -1948 -868 -1938 -816
rect -2012 -879 -1938 -868
rect -2519 -1302 -2285 -1229
rect -2257 -1233 -1694 -1187
rect -2519 -1303 -2400 -1302
rect -2519 -1631 -2473 -1303
rect -2257 -1328 -2225 -1233
rect -2272 -1512 -2225 -1328
rect -2389 -2774 -2361 -1519
rect -1401 -1526 -1367 -1203
rect -1861 -1864 -1822 -1526
rect -1679 -1678 -1643 -1677
rect -1679 -1856 -1632 -1678
rect -1861 -2773 -1833 -1864
rect -1668 -1868 -1632 -1856
rect -1664 -1961 -1632 -1868
rect -1414 -1789 -1367 -1526
rect -1665 -1970 -1596 -1961
rect -1665 -2022 -1654 -1970
rect -1602 -2022 -1596 -1970
rect -1665 -2029 -1596 -2022
rect -2413 -2797 -2334 -2774
rect -2540 -2842 -2462 -2819
rect -2540 -2848 -2519 -2842
rect -5378 -2876 -2519 -2848
rect -2485 -2876 -2462 -2842
rect -2413 -2831 -2392 -2797
rect -2358 -2831 -2334 -2797
rect -2413 -2855 -2334 -2831
rect -1882 -2796 -1803 -2773
rect -1414 -2779 -1386 -1789
rect -1283 -1817 -1249 -550
rect -817 -731 -783 -507
rect -699 -635 -665 1527
rect -463 -428 -429 2076
rect -242 1610 -176 1623
rect -242 1576 -226 1610
rect -192 1576 -176 1610
rect -242 1563 -176 1576
rect -227 955 -193 1563
rect -228 -428 -193 955
rect -699 -669 -547 -635
rect -834 -737 -770 -731
rect -834 -789 -828 -737
rect -776 -789 -770 -737
rect -834 -795 -770 -789
rect -1053 -1482 -1019 -1197
rect -1358 -1857 -1249 -1817
rect -1358 -1863 -1292 -1857
rect -1054 -2186 -1019 -1482
rect -817 -1773 -783 -795
rect -581 -1773 -547 -669
rect -228 -939 -194 -428
rect -109 -492 -75 497
rect 129 -439 163 2077
rect 494 -477 528 2079
rect 584 2077 658 2093
rect 945 2127 1019 2140
rect 1242 2137 1276 2141
rect 945 2093 964 2127
rect 998 2093 1019 2127
rect 945 2077 1019 2093
rect 1210 2124 1284 2137
rect 1210 2090 1229 2124
rect 1263 2090 1284 2124
rect 606 -477 637 2077
rect 974 1405 1008 2077
rect 1210 2074 1284 2090
rect 1242 1551 1276 2074
rect 1229 1544 1292 1551
rect 1229 1492 1235 1544
rect 1287 1492 1292 1544
rect 1229 1484 1292 1492
rect 4339 -27 4488 12
rect 4339 -79 4386 -27
rect 4438 -79 4488 -27
rect 4339 -120 4488 -79
rect 4318 -278 4470 -248
rect 4141 -279 4470 -278
rect 1914 -291 4470 -279
rect -109 -538 113 -492
rect 69 -868 104 -538
rect 69 -904 353 -868
rect -228 -972 234 -939
rect -423 -996 -359 -990
rect -423 -1048 -417 -996
rect -365 -1048 -359 -996
rect -423 -1054 -359 -1048
rect -404 -1100 -370 -1054
rect -308 -1097 -231 -1088
rect -421 -1155 -353 -1100
rect -308 -1145 -296 -1097
rect -244 -1111 -231 -1097
rect -244 -1145 -77 -1111
rect -6 -1154 59 -1082
rect 187 -1097 234 -972
rect 114 -1152 234 -1097
rect 187 -1223 234 -1152
rect 325 -1187 353 -904
rect 723 -974 769 -304
rect 1914 -343 4368 -291
rect 4420 -343 4470 -291
rect 1914 -347 4470 -343
rect 899 -597 965 -543
rect 1018 -597 1084 -543
rect 812 -625 872 -610
rect 1116 -625 1170 -614
rect 812 -626 1170 -625
rect 812 -660 824 -626
rect 858 -628 1170 -626
rect 858 -660 1124 -628
rect 812 -662 1124 -660
rect 1158 -662 1170 -628
rect 812 -668 1170 -662
rect 812 -673 872 -668
rect 1116 -674 1170 -668
rect 1179 -772 1811 -744
rect 934 -821 992 -809
rect 1179 -821 1209 -772
rect 934 -823 1209 -821
rect 934 -857 946 -823
rect 980 -857 1209 -823
rect 1323 -807 1394 -801
rect 934 -870 992 -857
rect 1323 -859 1336 -807
rect 1388 -859 1394 -807
rect 1323 -873 1394 -859
rect 1771 -938 1811 -772
rect 1914 -797 1968 -347
rect 4318 -391 4470 -347
rect 1911 -803 1975 -797
rect 1911 -855 1917 -803
rect 1969 -855 1975 -803
rect 1911 -861 1975 -855
rect 1771 -974 2555 -938
rect 723 -1016 1602 -974
rect 1421 -1050 1490 -1044
rect 381 -1161 443 -1104
rect 499 -1161 561 -1104
rect 1112 -1158 1174 -1101
rect 1421 -1102 1430 -1050
rect 1482 -1102 1490 -1050
rect 1421 -1106 1490 -1102
rect 1540 -1104 1860 -1040
rect 1738 -1134 1768 -1104
rect 325 -1215 368 -1187
rect -469 -1725 -422 -1489
rect -469 -1782 -402 -1725
rect -892 -1865 -709 -1815
rect -818 -2038 -784 -1865
rect -538 -1870 -472 -1813
rect -831 -2045 -768 -2038
rect -831 -2097 -825 -2045
rect -773 -2097 -768 -2045
rect -831 -2105 -768 -2097
rect -1054 -2779 -1020 -2186
rect -442 -2389 -402 -1782
rect -452 -2395 -388 -2389
rect -452 -2447 -446 -2395
rect -394 -2447 -388 -2395
rect -452 -2453 -388 -2447
rect -227 -2774 -193 -1527
rect -52 -1750 -15 -1489
rect -52 -1964 -14 -1750
rect 187 -1771 221 -1223
rect 334 -1309 368 -1215
rect 570 -1791 620 -1400
rect 1738 -1418 1786 -1134
rect 1182 -1788 1236 -1513
rect 377 -1822 439 -1821
rect 377 -1878 443 -1822
rect 496 -1876 558 -1819
rect -60 -1971 5 -1964
rect -60 -2023 -54 -1971
rect -2 -2023 5 -1971
rect -60 -2030 5 -2023
rect -1882 -2830 -1861 -2796
rect -1827 -2830 -1803 -2796
rect -1882 -2854 -1803 -2830
rect -1440 -2802 -1361 -2779
rect -1440 -2836 -1419 -2802
rect -1385 -2836 -1361 -2802
rect -1440 -2860 -1361 -2836
rect -1074 -2802 -995 -2779
rect -1074 -2836 -1053 -2802
rect -1019 -2836 -995 -2802
rect -1074 -2860 -995 -2836
rect -255 -2797 -176 -2774
rect 586 -2777 620 -1791
rect 874 -1872 936 -1818
rect 992 -1872 1054 -1818
rect 1110 -1870 1172 -1816
rect 994 -2010 1052 -1872
rect 990 -2016 1054 -2010
rect 990 -2068 996 -2016
rect 1048 -2068 1054 -2016
rect 990 -2074 1054 -2068
rect 1202 -2770 1236 -1788
rect 1622 -2765 1656 -1511
rect 1876 -2761 1910 -1511
rect 2381 -2215 2555 -974
rect 2381 -2585 3665 -2215
rect -255 -2831 -234 -2797
rect -200 -2831 -176 -2797
rect -255 -2855 -176 -2831
rect 561 -2800 640 -2777
rect 561 -2834 582 -2800
rect 616 -2834 640 -2800
rect 561 -2858 640 -2834
rect 1184 -2793 1263 -2770
rect 1184 -2827 1205 -2793
rect 1239 -2827 1263 -2793
rect 1184 -2851 1263 -2827
rect 1592 -2788 1671 -2765
rect 1592 -2822 1613 -2788
rect 1647 -2822 1671 -2788
rect 1592 -2846 1671 -2822
rect 1861 -2784 1940 -2761
rect 1861 -2818 1882 -2784
rect 1916 -2818 1940 -2784
rect 1861 -2842 1940 -2818
rect -2540 -2899 -2462 -2876
<< via1 >>
rect -2622 1869 -2570 1879
rect -2622 1835 -2616 1869
rect -2616 1835 -2582 1869
rect -2582 1835 -2570 1869
rect -2622 1827 -2570 1835
rect -2616 1754 -2564 1764
rect -2616 1720 -2610 1754
rect -2610 1720 -2576 1754
rect -2576 1720 -2564 1754
rect -2616 1712 -2564 1720
rect -5546 1534 -5494 1586
rect -3888 1534 -3836 1586
rect -1524 1648 -1472 1700
rect -5378 191 -5326 243
rect -4958 195 -4906 247
rect -5228 -10 -5176 42
rect -3292 209 -3240 261
rect -3570 -10 -3518 42
rect -3212 -782 -3160 -730
rect -4982 -941 -4930 -889
rect -2232 -544 -2180 -492
rect -1859 -544 -1807 -492
rect -1768 -664 -1716 -612
rect -2000 -828 -1948 -816
rect -2000 -862 -1991 -828
rect -1991 -862 -1957 -828
rect -1957 -862 -1948 -828
rect -2000 -868 -1948 -862
rect -1654 -2022 -1602 -1970
rect -828 -789 -776 -737
rect 1235 1492 1287 1544
rect 4386 -79 4438 -27
rect -417 -1048 -365 -996
rect -296 -1106 -244 -1097
rect -296 -1140 -287 -1106
rect -287 -1140 -253 -1106
rect -253 -1140 -244 -1106
rect -296 -1149 -244 -1140
rect 4368 -343 4420 -291
rect 1336 -824 1388 -807
rect 1336 -858 1337 -824
rect 1337 -858 1371 -824
rect 1371 -858 1388 -824
rect 1336 -859 1388 -858
rect 1917 -855 1969 -803
rect 1430 -1102 1482 -1050
rect -825 -2097 -773 -2045
rect -446 -2447 -394 -2395
rect -54 -2023 -2 -1971
rect 996 -2068 1048 -2016
<< metal2 >>
rect 1620 2234 3482 2238
rect 5065 2234 5267 2292
rect 1620 2175 5267 2234
rect -7106 1875 -6904 2003
rect -2634 1879 -2562 1888
rect -7106 1874 -5382 1875
rect -2634 1874 -2622 1879
rect -7106 1827 -2622 1874
rect -2570 1827 -2562 1879
rect -7106 1825 -2562 1827
rect -6929 1823 -2562 1825
rect -5699 1822 -2562 1823
rect -2634 1816 -2562 1822
rect -2628 1764 -2556 1773
rect -7113 1760 -6911 1762
rect -7113 1758 -5391 1760
rect -2628 1758 -2616 1764
rect -7113 1712 -2616 1758
rect -2564 1712 -2556 1764
rect -7113 1708 -2556 1712
rect -7113 1584 -6911 1708
rect -5706 1706 -2556 1708
rect -2628 1701 -2556 1706
rect -1537 1702 -1460 1715
rect -1537 1646 -1526 1702
rect -1470 1646 -1460 1702
rect -1537 1630 -1460 1646
rect -5592 1588 -5448 1626
rect -5592 1532 -5549 1588
rect -5493 1532 -5448 1588
rect -5592 1496 -5448 1532
rect -3934 1588 -3790 1626
rect -3934 1532 -3891 1588
rect -3835 1532 -3790 1588
rect -3934 1496 -3790 1532
rect 1222 1546 1299 1559
rect 1222 1490 1233 1546
rect 1289 1490 1299 1546
rect 1222 1474 1299 1490
rect -3302 261 -3230 284
rect -5384 243 -5309 255
rect -5384 191 -5378 243
rect -5326 232 -5309 243
rect -4964 247 -4900 253
rect -4964 232 -4958 247
rect -5326 202 -4958 232
rect -5326 191 -5309 202
rect -5384 182 -5309 191
rect -4964 195 -4958 202
rect -4906 232 -4900 247
rect -3302 232 -3292 261
rect -4906 209 -3292 232
rect -3240 209 -3230 261
rect -4906 202 -3230 209
rect -4906 195 -4900 202
rect -3302 197 -3230 202
rect -4964 189 -4900 195
rect -5274 44 -5130 82
rect -5274 -12 -5231 44
rect -5175 -12 -5130 44
rect -5274 -48 -5130 -12
rect -3616 44 -3472 82
rect -3616 -12 -3573 44
rect -3517 -12 -3472 44
rect -3616 -48 -3472 -12
rect -7102 -125 -6900 -67
rect -7102 -167 -5503 -125
rect -7102 -245 -6900 -167
rect -7112 -536 -6910 -449
rect -7112 -567 -5711 -536
rect -7112 -627 -6910 -567
rect -5758 -821 -5711 -567
rect -5565 -619 -5503 -167
rect -2237 -492 -2174 -484
rect -2237 -544 -2232 -492
rect -2180 -508 -2174 -492
rect -1866 -492 -1802 -481
rect -1866 -508 -1859 -492
rect -2180 -544 -1859 -508
rect -1807 -544 -1802 -492
rect -2237 -550 -1802 -544
rect -1775 -612 -1711 -601
rect -5565 -620 -2200 -619
rect -1775 -620 -1768 -612
rect -5565 -660 -1768 -620
rect -5397 -661 -1768 -660
rect -1775 -664 -1768 -661
rect -1716 -664 -1711 -612
rect -1775 -670 -1711 -664
rect 1620 -692 1659 2175
rect 3307 2171 5267 2175
rect 5065 2114 5267 2171
rect 4339 -23 4485 12
rect 993 -722 1659 -692
rect 2297 -25 4485 -23
rect 2297 -78 4385 -25
rect -3218 -730 -3154 -724
rect -3218 -782 -3212 -730
rect -3160 -745 -3154 -730
rect -834 -737 -770 -731
rect -834 -745 -828 -737
rect -3160 -778 -828 -745
rect -3160 -782 -3154 -778
rect -3218 -788 -3154 -782
rect -834 -789 -828 -778
rect -776 -748 -770 -737
rect 993 -748 1027 -722
rect -776 -778 1027 -748
rect -776 -789 -770 -778
rect -834 -795 -770 -789
rect -2012 -816 -1939 -806
rect -5758 -822 -3975 -821
rect -5758 -823 -2435 -822
rect -2012 -823 -2000 -816
rect -5758 -852 -2000 -823
rect -5546 -853 -2000 -852
rect -5396 -854 -2000 -853
rect -2012 -868 -2000 -854
rect -1948 -868 -1939 -816
rect -2012 -875 -1939 -868
rect 1323 -807 1394 -801
rect 1323 -859 1336 -807
rect 1388 -815 1394 -807
rect 1911 -803 1975 -797
rect 1911 -815 1917 -803
rect 1388 -845 1917 -815
rect 1388 -859 1394 -845
rect 1323 -873 1394 -859
rect 1911 -855 1917 -845
rect 1969 -855 1975 -803
rect 1911 -861 1975 -855
rect -4988 -889 -4924 -883
rect -4988 -941 -4982 -889
rect -4930 -904 -4924 -889
rect 1332 -904 1378 -873
rect -4930 -934 1378 -904
rect 1422 -883 1496 -874
rect -4930 -941 -4924 -934
rect -4988 -947 -4924 -941
rect 1422 -939 1430 -883
rect 1486 -939 1496 -883
rect 1422 -943 1496 -939
rect 1422 -944 1494 -943
rect -7114 -1002 -6912 -986
rect -423 -996 -359 -990
rect -7114 -1003 -849 -1002
rect -423 -1003 -417 -996
rect -7114 -1032 -417 -1003
rect -7114 -1164 -6912 -1032
rect -5264 -1033 -417 -1032
rect -423 -1048 -417 -1033
rect -365 -1048 -359 -996
rect -423 -1054 -359 -1048
rect 1421 -1050 1494 -944
rect -308 -1097 -232 -1088
rect -5584 -1111 -728 -1110
rect -308 -1111 -296 -1097
rect -5584 -1144 -296 -1111
rect -7117 -1590 -6915 -1521
rect -5584 -1590 -5529 -1144
rect -5244 -1145 -296 -1144
rect -308 -1149 -296 -1145
rect -244 -1149 -232 -1097
rect 1421 -1102 1430 -1050
rect 1482 -1102 1494 -1050
rect 1421 -1105 1494 -1102
rect 1421 -1106 1490 -1105
rect -308 -1160 -232 -1149
rect -7117 -1637 -5529 -1590
rect -7117 -1699 -6915 -1637
rect -1665 -1968 -1596 -1961
rect -60 -1968 5 -1964
rect -1665 -1970 5 -1968
rect -1665 -2022 -1654 -1970
rect -1602 -1971 5 -1970
rect -1602 -2002 -54 -1971
rect -1602 -2022 -1596 -2002
rect -61 -2006 -54 -2002
rect -1665 -2029 -1596 -2022
rect -60 -2023 -54 -2006
rect -2 -2023 5 -1971
rect -60 -2030 5 -2023
rect 990 -2016 1054 -2010
rect 990 -2026 996 -2016
rect -838 -2043 -761 -2030
rect -7117 -2150 -6915 -2078
rect -838 -2099 -827 -2043
rect -771 -2099 -761 -2043
rect 989 -2056 996 -2026
rect 990 -2068 996 -2056
rect 1048 -2068 1054 -2016
rect 990 -2074 1054 -2068
rect -838 -2115 -761 -2099
rect -7117 -2151 612 -2150
rect 999 -2151 1045 -2074
rect -7117 -2197 1044 -2151
rect -7117 -2256 -6915 -2197
rect -5246 -2198 1044 -2197
rect -452 -2395 -388 -2389
rect -452 -2447 -446 -2395
rect -394 -2412 -388 -2395
rect 2297 -2412 2331 -78
rect 4339 -81 4385 -78
rect 4441 -81 4485 -25
rect 4339 -118 4485 -81
rect 4340 -119 4484 -118
rect 4318 -282 4470 -248
rect 4925 -282 5127 -215
rect 4318 -289 5127 -282
rect 4318 -345 4366 -289
rect 4422 -345 5127 -289
rect 4318 -391 4470 -345
rect 4925 -393 5127 -345
rect -394 -2446 2331 -2412
rect -394 -2447 -388 -2446
rect -452 -2453 -388 -2447
<< via2 >>
rect -1526 1700 -1470 1702
rect -1526 1648 -1524 1700
rect -1524 1648 -1472 1700
rect -1472 1648 -1470 1700
rect -1526 1646 -1470 1648
rect -5549 1586 -5493 1588
rect -5549 1534 -5546 1586
rect -5546 1534 -5494 1586
rect -5494 1534 -5493 1586
rect -5549 1532 -5493 1534
rect -3891 1586 -3835 1588
rect -3891 1534 -3888 1586
rect -3888 1534 -3836 1586
rect -3836 1534 -3835 1586
rect -3891 1532 -3835 1534
rect 1233 1544 1289 1546
rect 1233 1492 1235 1544
rect 1235 1492 1287 1544
rect 1287 1492 1289 1544
rect 1233 1490 1289 1492
rect -5231 42 -5175 44
rect -5231 -10 -5228 42
rect -5228 -10 -5176 42
rect -5176 -10 -5175 42
rect -5231 -12 -5175 -10
rect -3573 42 -3517 44
rect -3573 -10 -3570 42
rect -3570 -10 -3518 42
rect -3518 -10 -3517 42
rect -3573 -12 -3517 -10
rect 4385 -27 4441 -25
rect 1430 -939 1486 -883
rect -827 -2045 -771 -2043
rect -827 -2097 -825 -2045
rect -825 -2097 -773 -2045
rect -773 -2097 -771 -2045
rect -827 -2099 -771 -2097
rect 4385 -79 4386 -27
rect 4386 -79 4438 -27
rect 4438 -79 4441 -27
rect 4385 -81 4441 -79
rect 4366 -291 4422 -289
rect 4366 -343 4368 -291
rect 4368 -343 4420 -291
rect 4420 -343 4422 -291
rect 4366 -345 4422 -343
<< metal3 >>
rect -1537 1702 -1460 1715
rect -1537 1646 -1526 1702
rect -1470 1646 -1460 1702
rect -1537 1630 -1460 1646
rect -5592 1592 -5450 1624
rect -5592 1528 -5554 1592
rect -5490 1528 -5450 1592
rect -5592 1496 -5450 1528
rect -3934 1592 -3792 1624
rect -3934 1528 -3896 1592
rect -3832 1528 -3792 1592
rect -3934 1496 -3792 1528
rect -5274 48 -5132 80
rect -5274 -16 -5236 48
rect -5172 -16 -5132 48
rect -5274 -48 -5132 -16
rect -3616 48 -3474 80
rect -3616 -16 -3578 48
rect -3514 -16 -3474 48
rect -3616 -48 -3474 -16
rect -1534 -2031 -1462 1630
rect 1222 1546 1299 1559
rect 1222 1490 1233 1546
rect 1289 1490 1299 1546
rect 1222 1474 1299 1490
rect 1230 -831 1293 1474
rect 4342 -21 4484 11
rect 4342 -85 4382 -21
rect 4446 -85 4484 -21
rect 4342 -117 4484 -85
rect 4318 -285 4470 -248
rect 4318 -349 4362 -285
rect 4426 -349 4470 -285
rect 4318 -391 4470 -349
rect 1230 -883 1496 -831
rect 1230 -894 1430 -883
rect 1422 -939 1430 -894
rect 1486 -939 1496 -883
rect 1422 -944 1496 -939
rect -838 -2031 -761 -2030
rect -1534 -2043 -761 -2031
rect -1534 -2099 -827 -2043
rect -771 -2099 -761 -2043
rect -1534 -2112 -761 -2099
rect -838 -2115 -761 -2112
<< via3 >>
rect -5554 1588 -5490 1592
rect -5554 1532 -5549 1588
rect -5549 1532 -5493 1588
rect -5493 1532 -5490 1588
rect -5554 1528 -5490 1532
rect -3896 1588 -3832 1592
rect -3896 1532 -3891 1588
rect -3891 1532 -3835 1588
rect -3835 1532 -3832 1588
rect -3896 1528 -3832 1532
rect -5236 44 -5172 48
rect -5236 -12 -5231 44
rect -5231 -12 -5175 44
rect -5175 -12 -5172 44
rect -5236 -16 -5172 -12
rect -3578 44 -3514 48
rect -3578 -12 -3573 44
rect -3573 -12 -3517 44
rect -3517 -12 -3514 44
rect -3578 -16 -3514 -12
rect 4382 -25 4446 -21
rect 4382 -81 4385 -25
rect 4385 -81 4441 -25
rect 4441 -81 4446 -25
rect 4382 -85 4446 -81
rect 4362 -289 4426 -285
rect 4362 -345 4366 -289
rect 4366 -345 4422 -289
rect 4422 -345 4426 -289
rect 4362 -349 4426 -345
<< metal4 >>
rect -5594 1592 -5448 1626
rect -5594 1528 -5554 1592
rect -5490 1528 -5448 1592
rect -5594 1496 -5448 1528
rect -3936 1592 -3790 1626
rect -3936 1528 -3896 1592
rect -3832 1528 -3790 1592
rect -3936 1496 -3790 1528
rect -5539 1259 -5476 1496
rect -5540 844 -5476 1259
rect -3880 981 -3817 1496
rect -3878 932 -3817 981
rect -5234 82 -5174 456
rect -3576 82 -3516 626
rect 4359 83 4465 1075
rect -5276 48 -5130 82
rect -5276 -16 -5236 48
rect -5172 -16 -5130 48
rect -5276 -48 -5130 -16
rect -3618 48 -3472 82
rect -3618 -16 -3578 48
rect -3514 -16 -3472 48
rect 4360 11 4466 83
rect -3618 -48 -3472 -16
rect 4340 -21 4486 11
rect -5218 -60 -5158 -48
rect -3560 -60 -3500 -48
rect 4340 -85 4382 -21
rect 4446 -85 4486 -21
rect 4340 -119 4486 -85
rect 4318 -285 4470 -248
rect 4318 -349 4362 -285
rect 4426 -349 4470 -285
rect 4318 -391 4470 -349
rect 4350 -690 4435 -391
rect 2884 -2586 4206 -1531
rect 4354 -2073 4430 -690
use res20_046K  res20_046K_0
timestamp 1669522153
transform 1 0 -4718 0 1 145
box -300 0 72 1528
use res20_046K  res20_046K_1
timestamp 1669522153
transform 1 0 -3060 0 1 39
box -300 0 72 1528
use sky130_fd_pr__cap_mim_m3_1_2TJQJA  sky130_fd_pr__cap_mim_m3_1_2TJQJA_0
timestamp 1669522153
transform 1 0 -3849 0 1 818
box -356 -306 355 306
use sky130_fd_pr__cap_mim_m3_1_2TJQJA  sky130_fd_pr__cap_mim_m3_1_2TJQJA_1
timestamp 1669522153
transform 1 0 -5510 0 1 715
box -356 -306 355 306
use sky130_fd_pr__cap_mim_m3_1_UJT6R3  sky130_fd_pr__cap_mim_m3_1_UJT6R3_0
timestamp 1669522153
transform 1 0 3614 0 1 1014
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_UJT6R3  sky130_fd_pr__cap_mim_m3_1_UJT6R3_1
timestamp 1669522153
transform 1 0 3595 0 1 -1301
box -850 -800 849 800
use sky130_fd_pr__nfet_01v8_4LH4MW  sky130_fd_pr__nfet_01v8_4LH4MW_0
timestamp 1669522153
transform 1 0 -1036 0 1 -1486
box -173 -326 173 369
use sky130_fd_pr__nfet_01v8_DDE7UB  sky130_fd_pr__nfet_01v8_DDE7UB_0
timestamp 1669522153
transform 1 0 -1750 0 1 -1537
box -144 -357 144 357
use sky130_fd_pr__nfet_01v8_PW4FSF  sky130_fd_pr__nfet_01v8_PW4FSF_0
timestamp 1669522153
transform 1 0 1140 0 1 -1486
box -114 -388 114 388
use sky130_fd_pr__nfet_01v8_PW4FSF  sky130_fd_pr__nfet_01v8_PW4FSF_1
timestamp 1669522153
transform 1 0 529 0 1 -1489
box -114 -388 114 388
use sky130_fd_pr__nfet_01v8_PW4FSF  sky130_fd_pr__nfet_01v8_PW4FSF_2
timestamp 1669522153
transform 1 0 411 0 1 -1489
box -114 -388 114 388
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_0
timestamp 1669522153
transform 1 0 -505 0 1 -1516
box -114 -357 114 357
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_1
timestamp 1669522153
transform 1 0 1022 0 1 -1517
box -114 -357 114 357
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_2
timestamp 1669522153
transform 1 0 904 0 1 -1517
box -114 -357 114 357
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_3
timestamp 1669522153
transform 1 0 -1325 0 1 -1520
box -114 -357 114 357
use sky130_fd_pr__nfet_01v8_QSQEJU  sky130_fd_pr__nfet_01v8_QSQEJU_0
timestamp 1669522153
transform 1 0 -121 0 1 -1454
box -144 -357 144 357
use sky130_fd_pr__nfet_01v8_QSSMMX  sky130_fd_pr__nfet_01v8_QSSMMX_0
timestamp 1669522153
transform 1 0 -2434 0 1 -1601
box -114 -357 114 357
use sky130_fd_pr__nfet_01v8_VXZ4X9  sky130_fd_pr__nfet_01v8_VXZ4X9_0
timestamp 1669522153
transform 1 0 1576 0 1 -1703
box -114 -657 114 657
use sky130_fd_pr__nfet_01v8_VXZ4X9  sky130_fd_pr__nfet_01v8_VXZ4X9_1
timestamp 1669522153
transform 1 0 1458 0 1 -1703
box -114 -657 114 657
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_0
timestamp 1669522153
transform 1 0 1818 0 1 -1401
box -114 -357 114 372
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_1
timestamp 1669522153
transform 1 0 145 0 1 -1454
box -114 -357 114 372
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_2
timestamp 1669522153
transform 1 0 27 0 1 -1454
box -114 -357 114 372
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_3
timestamp 1669522153
transform 1 0 -269 0 1 -1454
box -114 -357 114 372
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_4
timestamp 1669522153
transform 1 0 -387 0 1 -1454
box -114 -357 114 372
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_5
timestamp 1669522153
transform 1 0 -2316 0 1 -1601
box -114 -357 114 372
use sky130_fd_pr__nfet_01v8_ZG8UN4  sky130_fd_pr__nfet_01v8_ZG8UN4_0
timestamp 1669522153
transform 1 0 -800 0 1 -1517
box -173 -357 173 398
use sky130_fd_pr__pfet_01v8_3AH94A  sky130_fd_pr__pfet_01v8_3AH94A_0
timestamp 1669522153
transform 1 0 -1744 0 1 525
box -124 -1024 124 1058
use sky130_fd_pr__pfet_01v8_BGAJ3C  sky130_fd_pr__pfet_01v8_BGAJ3C_0
timestamp 1669522153
transform 1 0 -2160 0 1 567
box -124 -1058 124 1024
use sky130_fd_pr__pfet_01v8_BGN7SB  sky130_fd_pr__pfet_01v8_BGN7SB_0
timestamp 1669522153
transform 1 0 -930 0 1 556
box -183 -1058 183 1024
use sky130_fd_pr__pfet_01v8_DLEZW3  sky130_fd_pr__pfet_01v8_DLEZW3_0
timestamp 1669522153
transform 1 0 -2278 0 1 567
box -124 -1058 124 1024
use sky130_fd_pr__pfet_01v8_FHN7S9  sky130_fd_pr__pfet_01v8_FHN7S9_0
timestamp 1669522153
transform 1 0 990 0 1 424
box -183 -1024 183 1058
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_0
timestamp 1669522153
transform 1 0 -269 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_1
timestamp 1669522153
transform 1 0 -387 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_2
timestamp 1669522153
transform 1 0 -505 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_3
timestamp 1669522153
transform 1 0 -623 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_4
timestamp 1669522153
transform 1 0 452 0 1 478
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_5
timestamp 1669522153
transform 1 0 334 0 1 478
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_6
timestamp 1669522153
transform 1 0 682 0 1 472
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_XLJZXD  sky130_fd_pr__pfet_01v8_XLJZXD_0
timestamp 1669522153
transform 1 0 -1325 0 1 579
box -124 -1084 124 1118
use sky130_fd_pr__pfet_01v8_ZF98YR  sky130_fd_pr__pfet_01v8_ZF98YR_0
timestamp 1669522153
transform 1 0 27 0 1 -7
box -184 -544 184 578
<< labels >>
rlabel locali s -2612 -2948 2008 -2688 4 GND
port 1 nsew
rlabel locali s -2216 2018 1290 2144 4 VDD
port 2 nsew
rlabel metal2 s -7086 1611 -6936 1738 4 Vabp
port 3 nsew
rlabel metal2 s -7080 1844 -6935 1987 4 Vabn
port 4 nsew
rlabel metal2 s 5089 2133 5240 2275 4 Vop
port 5 nsew
rlabel metal2 s 4948 -367 5103 -236 4 Von
port 6 nsew
rlabel metal2 s -7085 -1145 -6943 -1015 4 Vip
port 7 nsew
rlabel metal2 s -7090 -2230 -6948 -2100 4 Vin
port 8 nsew
rlabel metal2 s -7075 -218 -6925 -88 4 Vbp
port 9 nsew
rlabel metal2 s -7093 -1680 -6944 -1550 4 Vbiasn
port 10 nsew
rlabel metal2 s -7086 -599 -6932 -465 4 Vcm
port 11 nsew
<< end >>
