magic
tech sky130A
magscale 1 2
timestamp 1668984253
<< psubdiff >>
rect -4250 20507 -4226 20810
rect -3655 20507 -3631 20810
rect 12184 20657 12208 20783
rect 12765 20657 12789 20783
rect -4290 20340 -4266 20507
rect -4260 -962 -4236 -522
rect -3567 -632 -3543 -522
rect 12147 -632 12171 -474
rect -3567 -962 -3543 -799
rect 12147 -863 12171 -799
rect 12837 -863 12861 -474
<< psubdiffcont >>
rect -4226 20507 -3655 20810
rect 12208 20657 12765 20783
rect 12234 20507 12718 20657
rect -4266 20340 12718 20507
rect -4170 -522 -3686 20340
rect 12234 -474 12718 20340
rect -4236 -632 -3567 -522
rect 12171 -632 12837 -474
rect -4236 -799 12837 -632
rect -4236 -962 -3567 -799
rect 12171 -863 12837 -799
<< poly >>
rect 2953 20233 5250 20235
rect 2892 20190 5250 20233
rect 2892 20179 2965 20190
rect 3120 20180 5250 20190
rect 2892 20143 2958 20179
rect 5219 20104 5250 20180
rect 5219 20057 5388 20104
rect 8189 20102 8255 20113
rect 8189 20068 8205 20102
rect 8239 20068 8255 20102
rect 8189 20052 8255 20068
<< polycont >>
rect 8205 20068 8239 20102
<< locali >>
rect -4242 20507 -4226 20810
rect -3655 20507 -3639 20810
rect 12192 20657 12208 20783
rect 12765 20657 12781 20783
rect -4282 20340 -4266 20507
rect 8189 20142 8480 20147
rect 8189 20102 8423 20142
rect 8189 20068 8205 20102
rect 8239 20084 8423 20102
rect 8476 20084 8480 20142
rect 8239 20079 8480 20084
rect 8239 20068 8255 20079
rect 8189 20065 8255 20068
rect -2534 760 -2500 920
rect -2298 760 -2264 919
rect -2062 760 -2028 919
rect -1826 760 -1792 919
rect -1590 760 -1556 919
rect -1354 760 -1320 921
rect -2535 756 -1320 760
rect -2535 729 -1316 756
rect 253 729 287 869
rect -2535 722 287 729
rect -1350 710 287 722
rect 489 710 523 869
rect 725 710 759 870
rect 961 710 995 870
rect 1197 710 1231 869
rect 1433 710 1467 871
rect 1669 710 1703 870
rect 1905 710 1939 872
rect 2141 710 2175 870
rect 2377 710 2411 871
rect 2613 710 2647 870
rect 2849 710 2883 870
rect 3085 710 3119 871
rect -1350 687 3119 710
rect 253 681 3119 687
rect 253 676 3118 681
rect 5432 680 5466 839
rect 5668 680 5702 839
rect 5904 680 5938 840
rect 6140 680 6174 840
rect 6376 680 6410 839
rect 6612 680 6646 841
rect 6848 680 6882 840
rect 7084 680 7118 842
rect 7320 680 7354 840
rect 7556 680 7590 841
rect 7792 680 7826 840
rect 8028 680 8062 840
rect 8264 740 8298 841
rect 10072 754 10106 914
rect 10308 754 10342 913
rect 10544 754 10578 913
rect 10780 754 10814 913
rect 11016 754 11050 913
rect 11252 754 11286 915
rect 10071 740 11286 754
rect 8264 733 11286 740
rect 8264 716 11284 733
rect 8264 680 10108 716
rect 5432 646 10108 680
rect 8264 645 10108 646
rect 4416 -141 4485 -129
rect 4416 -175 4430 -141
rect 4468 -175 4485 -141
rect 4416 -181 4485 -175
rect -4252 -962 -4236 -522
rect -3567 -632 -3551 -522
rect 4424 -632 4473 -181
rect 12155 -632 12171 -474
rect -3567 -962 -3551 -799
rect 4404 -958 4479 -799
rect 12155 -863 12171 -799
rect 12837 -863 12853 -474
rect 4162 -1382 4716 -958
<< viali >>
rect 8205 20068 8239 20102
rect 8423 20084 8476 20142
rect -2475 12944 -2441 12978
rect 4430 -175 4468 -141
<< metal1 >>
rect 1013 21023 1290 21034
rect 1013 20867 1033 21023
rect 1277 20867 1290 21023
rect 1013 20756 1290 20867
rect 914 20735 1290 20756
rect 7388 21007 7665 21018
rect 7388 20851 7408 21007
rect 7652 20851 7665 21007
rect 7388 20775 7665 20851
rect 914 20668 1193 20735
rect 7388 20687 7758 20775
rect 1055 20266 1193 20668
rect 134 20185 1310 20266
rect 7406 20254 7545 20687
rect 5901 20243 6521 20245
rect 7093 20243 7713 20254
rect 5314 20193 7713 20243
rect -5344 12983 -5276 13020
rect -5344 12981 -4228 12983
rect -2526 12981 -2425 12984
rect -5344 12978 -2425 12981
rect -5344 12944 -2475 12978
rect -2441 12944 -2425 12978
rect -5344 12941 -2425 12944
rect -5344 12940 -4228 12941
rect -5344 12910 -5276 12940
rect -2526 12938 -2425 12941
rect -2416 671 -2382 12894
rect -2180 671 -2146 12894
rect -1944 671 -1910 12894
rect -1708 671 -1674 12894
rect -1472 671 -1438 12894
rect -2416 642 -1438 671
rect -2416 641 -1439 642
rect -2180 639 -2146 641
rect -1676 434 -1639 641
rect 135 519 169 20185
rect 5314 20184 7123 20193
rect 5314 20182 5934 20184
rect 6503 20182 7123 20184
rect 5314 20157 5349 20182
rect 15446 20160 15862 20368
rect 371 519 405 20046
rect 607 519 641 20046
rect 843 519 877 20046
rect 1079 519 1113 20046
rect 1315 519 1349 20046
rect 1551 519 1585 20046
rect 1787 519 1821 20046
rect 2023 519 2057 20046
rect 2259 519 2293 20046
rect 2495 519 2529 20046
rect 2731 519 2765 20046
rect 2967 519 3001 20046
rect 5314 554 5348 20157
rect 12132 20155 15862 20160
rect 8412 20142 15862 20155
rect 8189 20102 8255 20117
rect 8189 20068 8205 20102
rect 8239 20068 8255 20102
rect 8189 20062 8255 20068
rect 8412 20084 8423 20142
rect 8476 20084 15862 20142
rect 8412 20072 15862 20084
rect 8412 20067 12157 20072
rect 5550 554 5584 20015
rect 5786 554 5820 20015
rect 6022 554 6056 20015
rect 6258 554 6292 20015
rect 6494 554 6528 20015
rect 6730 554 6764 20015
rect 6966 554 7000 20015
rect 7202 554 7236 20015
rect 7438 554 7472 20015
rect 7674 554 7708 20015
rect 7910 554 7944 20015
rect 8146 554 8180 20015
rect 15446 19928 15862 20072
rect 10125 13103 11384 13131
rect 10115 13058 11384 13103
rect 10115 12932 10178 13058
rect 11322 12974 11383 13058
rect 13040 12974 13108 13008
rect 11322 12956 13108 12974
rect 11330 12933 13108 12956
rect 13040 12898 13108 12933
rect 10190 657 10224 12888
rect 10426 657 10460 12888
rect 10662 657 10696 12888
rect 10898 657 10932 12888
rect 11134 657 11168 12888
rect 10189 623 11169 657
rect 135 485 3001 519
rect 5311 494 8182 554
rect 135 478 169 485
rect 371 479 405 485
rect 607 484 641 485
rect 1079 483 1113 485
rect 1315 484 1349 485
rect 1551 480 1585 485
rect 1787 481 1821 485
rect 2023 480 2057 485
rect 2259 482 2293 485
rect 2731 482 2765 485
rect 2967 481 3001 485
rect 10371 437 10416 623
rect 10371 436 10415 437
rect 9410 435 10415 436
rect 3876 434 10415 435
rect -1676 413 10415 434
rect -1668 400 10415 413
rect -1668 399 3884 400
rect 4420 -129 4476 400
rect 4416 -141 4485 -129
rect 4416 -175 4430 -141
rect 4468 -175 4485 -141
rect 4416 -181 4485 -175
<< via1 >>
rect 1033 20867 1277 21023
rect 7408 20851 7652 21007
<< metal2 >>
rect 992 21436 1310 21504
rect 992 21272 1035 21436
rect 1267 21272 1310 21436
rect 992 21023 1310 21272
rect 992 20867 1033 21023
rect 1277 20867 1310 21023
rect 992 20842 1310 20867
rect 7367 21420 7685 21488
rect 7367 21256 7410 21420
rect 7642 21256 7685 21420
rect 7367 21007 7685 21256
rect 7367 20851 7408 21007
rect 7652 20851 7685 21007
rect 7367 20826 7685 20851
<< via2 >>
rect 1035 21272 1267 21436
rect 7410 21256 7642 21420
<< metal3 >>
rect 957 22082 1336 22151
rect 957 21866 1009 22082
rect 1276 21866 1336 22082
rect 957 21436 1336 21866
rect 957 21272 1035 21436
rect 1267 21272 1336 21436
rect 957 21177 1336 21272
rect 7332 22066 7711 22135
rect 7332 21850 7384 22066
rect 7651 21850 7711 22066
rect 7332 21420 7711 21850
rect 7332 21256 7410 21420
rect 7642 21256 7711 21420
rect 7332 21161 7711 21256
<< via3 >>
rect 1009 21866 1276 22082
rect 7384 21850 7651 22066
<< metal4 >>
rect 914 22711 1362 22746
rect 914 22453 957 22711
rect 1328 22453 1362 22711
rect 914 22082 1362 22453
rect 914 21866 1009 22082
rect 1276 21866 1362 22082
rect 914 21737 1362 21866
rect 7289 22695 7737 22730
rect 7289 22437 7332 22695
rect 7703 22437 7737 22695
rect 7289 22066 7737 22437
rect 7289 21850 7384 22066
rect 7651 21850 7737 22066
rect 7289 21721 7737 21850
rect 10578 21446 11584 21506
rect 15656 21446 16374 21738
rect 9684 21408 16374 21446
rect -1858 21200 16374 21408
rect -1858 21020 9928 21200
rect 15656 21038 16374 21200
rect -2732 20974 9928 21020
rect -1858 20972 9928 20974
<< via4 >>
rect 957 22453 1328 22711
rect 7332 22437 7703 22695
<< metal5 >>
rect 462 23894 1256 23908
rect 2126 23894 2844 24076
rect 462 23536 2844 23894
rect 462 22908 1388 23536
rect 2126 23376 2844 23536
rect 5472 23910 6190 24016
rect 6820 23914 8416 24392
rect 6816 23910 8416 23914
rect 5472 23552 8416 23910
rect 5472 23316 6190 23552
rect 6816 23550 8416 23552
rect 6820 23098 8416 23550
rect 888 22711 1388 22908
rect 7262 22762 7763 23098
rect 888 22453 957 22711
rect 1328 22453 1388 22711
rect 888 22375 1388 22453
rect 7263 22695 7763 22762
rect 7263 22437 7332 22695
rect 7703 22437 7763 22695
rect 7263 22359 7763 22437
use sky130_fd_pr__nfet_01v8_MWCSZB  XM2
timestamp 1668922623
transform 1 0 10679 0 1 6900
box -645 -6088 645 6088
use sky130_fd_pr__nfet_01v8_TXCS3D  XM4
timestamp 1668922623
transform 1 0 6806 0 1 10426
box -1530 -9688 1530 9688
use ind_PA  ind_PA_0
timestamp 1668922623
transform 1 0 7180 0 -1 21188
box 1200 -12000 11600 -300
use ind_PA  ind_PA_1
timestamp 1668922623
transform -1 0 1668 0 -1 20710
box 1200 -12000 11600 -300
use sky130_fd_pr__nfet_01v8_MWCSZB  sky130_fd_pr__nfet_01v8_MWCSZB_0
timestamp 1668922623
transform 1 0 -1927 0 1 6906
box -645 -6088 645 6088
use sky130_fd_pr__nfet_01v8_TXCS3D  sky130_fd_pr__nfet_01v8_TXCS3D_0
timestamp 1668922623
transform 1 0 1627 0 1 10457
box -1530 -9688 1530 9688
<< labels >>
rlabel metal5 2126 23376 2844 24076 1 Vx
port 1 n
rlabel metal5 5472 23316 6190 24016 1 Vy
port 2 n
rlabel metal4 15656 21038 16374 21738 1 VDD
port 3 n
rlabel locali 4162 -1382 4716 -958 1 GND
port 4 n
rlabel metal1 15446 19928 15862 20368 1 Vb
port 5 n
rlabel metal1 13040 12898 13108 13008 1 Vina
port 6 n
rlabel metal1 -5344 12910 -5276 13020 1 Vin
port 7 n
<< end >>
