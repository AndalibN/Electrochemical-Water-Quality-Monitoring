magic
tech sky130A
magscale 1 2
timestamp 1668702877
<< error_p >>
rect -324 6989 -266 6995
rect -206 6989 -148 6995
rect -88 6989 -30 6995
rect 30 6989 88 6995
rect 148 6989 206 6995
rect 266 6989 324 6995
rect -324 6955 -312 6989
rect -206 6955 -194 6989
rect -88 6955 -76 6989
rect 30 6955 42 6989
rect 148 6955 160 6989
rect 266 6955 278 6989
rect -324 6949 -266 6955
rect -206 6949 -148 6955
rect -88 6949 -30 6955
rect 30 6949 88 6955
rect 148 6949 206 6955
rect 266 6949 324 6955
rect -324 -6955 -266 -6949
rect -206 -6955 -148 -6949
rect -88 -6955 -30 -6949
rect 30 -6955 88 -6949
rect 148 -6955 206 -6949
rect 266 -6955 324 -6949
rect -324 -6989 -312 -6955
rect -206 -6989 -194 -6955
rect -88 -6989 -76 -6955
rect 30 -6989 42 -6955
rect 148 -6989 160 -6955
rect 266 -6989 278 -6955
rect -324 -6995 -266 -6989
rect -206 -6995 -148 -6989
rect -88 -6995 -30 -6989
rect 30 -6995 88 -6989
rect 148 -6995 206 -6989
rect 266 -6995 324 -6989
<< nmos >>
rect -325 -6917 -265 6917
rect -207 -6917 -147 6917
rect -89 -6917 -29 6917
rect 29 -6917 89 6917
rect 147 -6917 207 6917
rect 265 -6917 325 6917
<< ndiff >>
rect -383 6905 -325 6917
rect -383 -6905 -371 6905
rect -337 -6905 -325 6905
rect -383 -6917 -325 -6905
rect -265 6905 -207 6917
rect -265 -6905 -253 6905
rect -219 -6905 -207 6905
rect -265 -6917 -207 -6905
rect -147 6905 -89 6917
rect -147 -6905 -135 6905
rect -101 -6905 -89 6905
rect -147 -6917 -89 -6905
rect -29 6905 29 6917
rect -29 -6905 -17 6905
rect 17 -6905 29 6905
rect -29 -6917 29 -6905
rect 89 6905 147 6917
rect 89 -6905 101 6905
rect 135 -6905 147 6905
rect 89 -6917 147 -6905
rect 207 6905 265 6917
rect 207 -6905 219 6905
rect 253 -6905 265 6905
rect 207 -6917 265 -6905
rect 325 6905 383 6917
rect 325 -6905 337 6905
rect 371 -6905 383 6905
rect 325 -6917 383 -6905
<< ndiffc >>
rect -371 -6905 -337 6905
rect -253 -6905 -219 6905
rect -135 -6905 -101 6905
rect -17 -6905 17 6905
rect 101 -6905 135 6905
rect 219 -6905 253 6905
rect 337 -6905 371 6905
<< poly >>
rect -328 6989 -262 7005
rect -328 6955 -312 6989
rect -278 6955 -262 6989
rect -328 6939 -262 6955
rect -210 6989 -144 7005
rect -210 6955 -194 6989
rect -160 6955 -144 6989
rect -210 6939 -144 6955
rect -92 6989 -26 7005
rect -92 6955 -76 6989
rect -42 6955 -26 6989
rect -92 6939 -26 6955
rect 26 6989 92 7005
rect 26 6955 42 6989
rect 76 6955 92 6989
rect 26 6939 92 6955
rect 144 6989 210 7005
rect 144 6955 160 6989
rect 194 6955 210 6989
rect 144 6939 210 6955
rect 262 6989 328 7005
rect 262 6955 278 6989
rect 312 6955 328 6989
rect 262 6939 328 6955
rect -325 6917 -265 6939
rect -207 6917 -147 6939
rect -89 6917 -29 6939
rect 29 6917 89 6939
rect 147 6917 207 6939
rect 265 6917 325 6939
rect -325 -6939 -265 -6917
rect -207 -6939 -147 -6917
rect -89 -6939 -29 -6917
rect 29 -6939 89 -6917
rect 147 -6939 207 -6917
rect 265 -6939 325 -6917
rect -328 -6955 -262 -6939
rect -328 -6989 -312 -6955
rect -278 -6989 -262 -6955
rect -328 -7005 -262 -6989
rect -210 -6955 -144 -6939
rect -210 -6989 -194 -6955
rect -160 -6989 -144 -6955
rect -210 -7005 -144 -6989
rect -92 -6955 -26 -6939
rect -92 -6989 -76 -6955
rect -42 -6989 -26 -6955
rect -92 -7005 -26 -6989
rect 26 -6955 92 -6939
rect 26 -6989 42 -6955
rect 76 -6989 92 -6955
rect 26 -7005 92 -6989
rect 144 -6955 210 -6939
rect 144 -6989 160 -6955
rect 194 -6989 210 -6955
rect 144 -7005 210 -6989
rect 262 -6955 328 -6939
rect 262 -6989 278 -6955
rect 312 -6989 328 -6955
rect 262 -7005 328 -6989
<< polycont >>
rect -312 6955 -278 6989
rect -194 6955 -160 6989
rect -76 6955 -42 6989
rect 42 6955 76 6989
rect 160 6955 194 6989
rect 278 6955 312 6989
rect -312 -6989 -278 -6955
rect -194 -6989 -160 -6955
rect -76 -6989 -42 -6955
rect 42 -6989 76 -6955
rect 160 -6989 194 -6955
rect 278 -6989 312 -6955
<< locali >>
rect -328 6955 -312 6989
rect -278 6955 -262 6989
rect -210 6955 -194 6989
rect -160 6955 -144 6989
rect -92 6955 -76 6989
rect -42 6955 -26 6989
rect 26 6955 42 6989
rect 76 6955 92 6989
rect 144 6955 160 6989
rect 194 6955 210 6989
rect 262 6955 278 6989
rect 312 6955 328 6989
rect -371 6905 -337 6921
rect -371 -6921 -337 -6905
rect -253 6905 -219 6921
rect -253 -6921 -219 -6905
rect -135 6905 -101 6921
rect -135 -6921 -101 -6905
rect -17 6905 17 6921
rect -17 -6921 17 -6905
rect 101 6905 135 6921
rect 101 -6921 135 -6905
rect 219 6905 253 6921
rect 219 -6921 253 -6905
rect 337 6905 371 6921
rect 337 -6921 371 -6905
rect -328 -6989 -312 -6955
rect -278 -6989 -262 -6955
rect -210 -6989 -194 -6955
rect -160 -6989 -144 -6955
rect -92 -6989 -76 -6955
rect -42 -6989 -26 -6955
rect 26 -6989 42 -6955
rect 76 -6989 92 -6955
rect 144 -6989 160 -6955
rect 194 -6989 210 -6955
rect 262 -6989 278 -6955
rect 312 -6989 328 -6955
<< viali >>
rect -312 6955 -278 6989
rect -194 6955 -160 6989
rect -76 6955 -42 6989
rect 42 6955 76 6989
rect 160 6955 194 6989
rect 278 6955 312 6989
rect -371 -6905 -337 6905
rect -253 -6905 -219 6905
rect -135 -6905 -101 6905
rect -17 -6905 17 6905
rect 101 -6905 135 6905
rect 219 -6905 253 6905
rect 337 -6905 371 6905
rect -312 -6989 -278 -6955
rect -194 -6989 -160 -6955
rect -76 -6989 -42 -6955
rect 42 -6989 76 -6955
rect 160 -6989 194 -6955
rect 278 -6989 312 -6955
<< metal1 >>
rect -324 6989 -266 6995
rect -324 6955 -312 6989
rect -278 6955 -266 6989
rect -324 6949 -266 6955
rect -206 6989 -148 6995
rect -206 6955 -194 6989
rect -160 6955 -148 6989
rect -206 6949 -148 6955
rect -88 6989 -30 6995
rect -88 6955 -76 6989
rect -42 6955 -30 6989
rect -88 6949 -30 6955
rect 30 6989 88 6995
rect 30 6955 42 6989
rect 76 6955 88 6989
rect 30 6949 88 6955
rect 148 6989 206 6995
rect 148 6955 160 6989
rect 194 6955 206 6989
rect 148 6949 206 6955
rect 266 6989 324 6995
rect 266 6955 278 6989
rect 312 6955 324 6989
rect 266 6949 324 6955
rect -377 6905 -331 6917
rect -377 -6905 -371 6905
rect -337 -6905 -331 6905
rect -377 -6917 -331 -6905
rect -259 6905 -213 6917
rect -259 -6905 -253 6905
rect -219 -6905 -213 6905
rect -259 -6917 -213 -6905
rect -141 6905 -95 6917
rect -141 -6905 -135 6905
rect -101 -6905 -95 6905
rect -141 -6917 -95 -6905
rect -23 6905 23 6917
rect -23 -6905 -17 6905
rect 17 -6905 23 6905
rect -23 -6917 23 -6905
rect 95 6905 141 6917
rect 95 -6905 101 6905
rect 135 -6905 141 6905
rect 95 -6917 141 -6905
rect 213 6905 259 6917
rect 213 -6905 219 6905
rect 253 -6905 259 6905
rect 213 -6917 259 -6905
rect 331 6905 377 6917
rect 331 -6905 337 6905
rect 371 -6905 377 6905
rect 331 -6917 377 -6905
rect -324 -6955 -266 -6949
rect -324 -6989 -312 -6955
rect -278 -6989 -266 -6955
rect -324 -6995 -266 -6989
rect -206 -6955 -148 -6949
rect -206 -6989 -194 -6955
rect -160 -6989 -148 -6955
rect -206 -6995 -148 -6989
rect -88 -6955 -30 -6949
rect -88 -6989 -76 -6955
rect -42 -6989 -30 -6955
rect -88 -6995 -30 -6989
rect 30 -6955 88 -6949
rect 30 -6989 42 -6955
rect 76 -6989 88 -6955
rect 30 -6995 88 -6989
rect 148 -6955 206 -6949
rect 148 -6989 160 -6955
rect 194 -6989 206 -6955
rect 148 -6995 206 -6989
rect 266 -6955 324 -6949
rect 266 -6989 278 -6955
rect 312 -6989 324 -6955
rect 266 -6995 324 -6989
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 69.17 l 0.3 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
