magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect 142 2556 200 2562
rect 142 2522 154 2556
rect 142 2516 200 2522
<< pwell >>
rect -283 -2506 283 2506
<< nmos >>
rect -199 -2480 -143 2480
rect -85 -2480 -29 2480
rect 29 -2480 85 2480
rect 143 -2480 199 2480
<< ndiff >>
rect -257 2465 -199 2480
rect -257 2431 -245 2465
rect -211 2431 -199 2465
rect -257 2397 -199 2431
rect -257 2363 -245 2397
rect -211 2363 -199 2397
rect -257 2329 -199 2363
rect -257 2295 -245 2329
rect -211 2295 -199 2329
rect -257 2261 -199 2295
rect -257 2227 -245 2261
rect -211 2227 -199 2261
rect -257 2193 -199 2227
rect -257 2159 -245 2193
rect -211 2159 -199 2193
rect -257 2125 -199 2159
rect -257 2091 -245 2125
rect -211 2091 -199 2125
rect -257 2057 -199 2091
rect -257 2023 -245 2057
rect -211 2023 -199 2057
rect -257 1989 -199 2023
rect -257 1955 -245 1989
rect -211 1955 -199 1989
rect -257 1921 -199 1955
rect -257 1887 -245 1921
rect -211 1887 -199 1921
rect -257 1853 -199 1887
rect -257 1819 -245 1853
rect -211 1819 -199 1853
rect -257 1785 -199 1819
rect -257 1751 -245 1785
rect -211 1751 -199 1785
rect -257 1717 -199 1751
rect -257 1683 -245 1717
rect -211 1683 -199 1717
rect -257 1649 -199 1683
rect -257 1615 -245 1649
rect -211 1615 -199 1649
rect -257 1581 -199 1615
rect -257 1547 -245 1581
rect -211 1547 -199 1581
rect -257 1513 -199 1547
rect -257 1479 -245 1513
rect -211 1479 -199 1513
rect -257 1445 -199 1479
rect -257 1411 -245 1445
rect -211 1411 -199 1445
rect -257 1377 -199 1411
rect -257 1343 -245 1377
rect -211 1343 -199 1377
rect -257 1309 -199 1343
rect -257 1275 -245 1309
rect -211 1275 -199 1309
rect -257 1241 -199 1275
rect -257 1207 -245 1241
rect -211 1207 -199 1241
rect -257 1173 -199 1207
rect -257 1139 -245 1173
rect -211 1139 -199 1173
rect -257 1105 -199 1139
rect -257 1071 -245 1105
rect -211 1071 -199 1105
rect -257 1037 -199 1071
rect -257 1003 -245 1037
rect -211 1003 -199 1037
rect -257 969 -199 1003
rect -257 935 -245 969
rect -211 935 -199 969
rect -257 901 -199 935
rect -257 867 -245 901
rect -211 867 -199 901
rect -257 833 -199 867
rect -257 799 -245 833
rect -211 799 -199 833
rect -257 765 -199 799
rect -257 731 -245 765
rect -211 731 -199 765
rect -257 697 -199 731
rect -257 663 -245 697
rect -211 663 -199 697
rect -257 629 -199 663
rect -257 595 -245 629
rect -211 595 -199 629
rect -257 561 -199 595
rect -257 527 -245 561
rect -211 527 -199 561
rect -257 493 -199 527
rect -257 459 -245 493
rect -211 459 -199 493
rect -257 425 -199 459
rect -257 391 -245 425
rect -211 391 -199 425
rect -257 357 -199 391
rect -257 323 -245 357
rect -211 323 -199 357
rect -257 289 -199 323
rect -257 255 -245 289
rect -211 255 -199 289
rect -257 221 -199 255
rect -257 187 -245 221
rect -211 187 -199 221
rect -257 153 -199 187
rect -257 119 -245 153
rect -211 119 -199 153
rect -257 85 -199 119
rect -257 51 -245 85
rect -211 51 -199 85
rect -257 17 -199 51
rect -257 -17 -245 17
rect -211 -17 -199 17
rect -257 -51 -199 -17
rect -257 -85 -245 -51
rect -211 -85 -199 -51
rect -257 -119 -199 -85
rect -257 -153 -245 -119
rect -211 -153 -199 -119
rect -257 -187 -199 -153
rect -257 -221 -245 -187
rect -211 -221 -199 -187
rect -257 -255 -199 -221
rect -257 -289 -245 -255
rect -211 -289 -199 -255
rect -257 -323 -199 -289
rect -257 -357 -245 -323
rect -211 -357 -199 -323
rect -257 -391 -199 -357
rect -257 -425 -245 -391
rect -211 -425 -199 -391
rect -257 -459 -199 -425
rect -257 -493 -245 -459
rect -211 -493 -199 -459
rect -257 -527 -199 -493
rect -257 -561 -245 -527
rect -211 -561 -199 -527
rect -257 -595 -199 -561
rect -257 -629 -245 -595
rect -211 -629 -199 -595
rect -257 -663 -199 -629
rect -257 -697 -245 -663
rect -211 -697 -199 -663
rect -257 -731 -199 -697
rect -257 -765 -245 -731
rect -211 -765 -199 -731
rect -257 -799 -199 -765
rect -257 -833 -245 -799
rect -211 -833 -199 -799
rect -257 -867 -199 -833
rect -257 -901 -245 -867
rect -211 -901 -199 -867
rect -257 -935 -199 -901
rect -257 -969 -245 -935
rect -211 -969 -199 -935
rect -257 -1003 -199 -969
rect -257 -1037 -245 -1003
rect -211 -1037 -199 -1003
rect -257 -1071 -199 -1037
rect -257 -1105 -245 -1071
rect -211 -1105 -199 -1071
rect -257 -1139 -199 -1105
rect -257 -1173 -245 -1139
rect -211 -1173 -199 -1139
rect -257 -1207 -199 -1173
rect -257 -1241 -245 -1207
rect -211 -1241 -199 -1207
rect -257 -1275 -199 -1241
rect -257 -1309 -245 -1275
rect -211 -1309 -199 -1275
rect -257 -1343 -199 -1309
rect -257 -1377 -245 -1343
rect -211 -1377 -199 -1343
rect -257 -1411 -199 -1377
rect -257 -1445 -245 -1411
rect -211 -1445 -199 -1411
rect -257 -1479 -199 -1445
rect -257 -1513 -245 -1479
rect -211 -1513 -199 -1479
rect -257 -1547 -199 -1513
rect -257 -1581 -245 -1547
rect -211 -1581 -199 -1547
rect -257 -1615 -199 -1581
rect -257 -1649 -245 -1615
rect -211 -1649 -199 -1615
rect -257 -1683 -199 -1649
rect -257 -1717 -245 -1683
rect -211 -1717 -199 -1683
rect -257 -1751 -199 -1717
rect -257 -1785 -245 -1751
rect -211 -1785 -199 -1751
rect -257 -1819 -199 -1785
rect -257 -1853 -245 -1819
rect -211 -1853 -199 -1819
rect -257 -1887 -199 -1853
rect -257 -1921 -245 -1887
rect -211 -1921 -199 -1887
rect -257 -1955 -199 -1921
rect -257 -1989 -245 -1955
rect -211 -1989 -199 -1955
rect -257 -2023 -199 -1989
rect -257 -2057 -245 -2023
rect -211 -2057 -199 -2023
rect -257 -2091 -199 -2057
rect -257 -2125 -245 -2091
rect -211 -2125 -199 -2091
rect -257 -2159 -199 -2125
rect -257 -2193 -245 -2159
rect -211 -2193 -199 -2159
rect -257 -2227 -199 -2193
rect -257 -2261 -245 -2227
rect -211 -2261 -199 -2227
rect -257 -2295 -199 -2261
rect -257 -2329 -245 -2295
rect -211 -2329 -199 -2295
rect -257 -2363 -199 -2329
rect -257 -2397 -245 -2363
rect -211 -2397 -199 -2363
rect -257 -2431 -199 -2397
rect -257 -2465 -245 -2431
rect -211 -2465 -199 -2431
rect -257 -2480 -199 -2465
rect -143 2465 -85 2480
rect -143 2431 -131 2465
rect -97 2431 -85 2465
rect -143 2397 -85 2431
rect -143 2363 -131 2397
rect -97 2363 -85 2397
rect -143 2329 -85 2363
rect -143 2295 -131 2329
rect -97 2295 -85 2329
rect -143 2261 -85 2295
rect -143 2227 -131 2261
rect -97 2227 -85 2261
rect -143 2193 -85 2227
rect -143 2159 -131 2193
rect -97 2159 -85 2193
rect -143 2125 -85 2159
rect -143 2091 -131 2125
rect -97 2091 -85 2125
rect -143 2057 -85 2091
rect -143 2023 -131 2057
rect -97 2023 -85 2057
rect -143 1989 -85 2023
rect -143 1955 -131 1989
rect -97 1955 -85 1989
rect -143 1921 -85 1955
rect -143 1887 -131 1921
rect -97 1887 -85 1921
rect -143 1853 -85 1887
rect -143 1819 -131 1853
rect -97 1819 -85 1853
rect -143 1785 -85 1819
rect -143 1751 -131 1785
rect -97 1751 -85 1785
rect -143 1717 -85 1751
rect -143 1683 -131 1717
rect -97 1683 -85 1717
rect -143 1649 -85 1683
rect -143 1615 -131 1649
rect -97 1615 -85 1649
rect -143 1581 -85 1615
rect -143 1547 -131 1581
rect -97 1547 -85 1581
rect -143 1513 -85 1547
rect -143 1479 -131 1513
rect -97 1479 -85 1513
rect -143 1445 -85 1479
rect -143 1411 -131 1445
rect -97 1411 -85 1445
rect -143 1377 -85 1411
rect -143 1343 -131 1377
rect -97 1343 -85 1377
rect -143 1309 -85 1343
rect -143 1275 -131 1309
rect -97 1275 -85 1309
rect -143 1241 -85 1275
rect -143 1207 -131 1241
rect -97 1207 -85 1241
rect -143 1173 -85 1207
rect -143 1139 -131 1173
rect -97 1139 -85 1173
rect -143 1105 -85 1139
rect -143 1071 -131 1105
rect -97 1071 -85 1105
rect -143 1037 -85 1071
rect -143 1003 -131 1037
rect -97 1003 -85 1037
rect -143 969 -85 1003
rect -143 935 -131 969
rect -97 935 -85 969
rect -143 901 -85 935
rect -143 867 -131 901
rect -97 867 -85 901
rect -143 833 -85 867
rect -143 799 -131 833
rect -97 799 -85 833
rect -143 765 -85 799
rect -143 731 -131 765
rect -97 731 -85 765
rect -143 697 -85 731
rect -143 663 -131 697
rect -97 663 -85 697
rect -143 629 -85 663
rect -143 595 -131 629
rect -97 595 -85 629
rect -143 561 -85 595
rect -143 527 -131 561
rect -97 527 -85 561
rect -143 493 -85 527
rect -143 459 -131 493
rect -97 459 -85 493
rect -143 425 -85 459
rect -143 391 -131 425
rect -97 391 -85 425
rect -143 357 -85 391
rect -143 323 -131 357
rect -97 323 -85 357
rect -143 289 -85 323
rect -143 255 -131 289
rect -97 255 -85 289
rect -143 221 -85 255
rect -143 187 -131 221
rect -97 187 -85 221
rect -143 153 -85 187
rect -143 119 -131 153
rect -97 119 -85 153
rect -143 85 -85 119
rect -143 51 -131 85
rect -97 51 -85 85
rect -143 17 -85 51
rect -143 -17 -131 17
rect -97 -17 -85 17
rect -143 -51 -85 -17
rect -143 -85 -131 -51
rect -97 -85 -85 -51
rect -143 -119 -85 -85
rect -143 -153 -131 -119
rect -97 -153 -85 -119
rect -143 -187 -85 -153
rect -143 -221 -131 -187
rect -97 -221 -85 -187
rect -143 -255 -85 -221
rect -143 -289 -131 -255
rect -97 -289 -85 -255
rect -143 -323 -85 -289
rect -143 -357 -131 -323
rect -97 -357 -85 -323
rect -143 -391 -85 -357
rect -143 -425 -131 -391
rect -97 -425 -85 -391
rect -143 -459 -85 -425
rect -143 -493 -131 -459
rect -97 -493 -85 -459
rect -143 -527 -85 -493
rect -143 -561 -131 -527
rect -97 -561 -85 -527
rect -143 -595 -85 -561
rect -143 -629 -131 -595
rect -97 -629 -85 -595
rect -143 -663 -85 -629
rect -143 -697 -131 -663
rect -97 -697 -85 -663
rect -143 -731 -85 -697
rect -143 -765 -131 -731
rect -97 -765 -85 -731
rect -143 -799 -85 -765
rect -143 -833 -131 -799
rect -97 -833 -85 -799
rect -143 -867 -85 -833
rect -143 -901 -131 -867
rect -97 -901 -85 -867
rect -143 -935 -85 -901
rect -143 -969 -131 -935
rect -97 -969 -85 -935
rect -143 -1003 -85 -969
rect -143 -1037 -131 -1003
rect -97 -1037 -85 -1003
rect -143 -1071 -85 -1037
rect -143 -1105 -131 -1071
rect -97 -1105 -85 -1071
rect -143 -1139 -85 -1105
rect -143 -1173 -131 -1139
rect -97 -1173 -85 -1139
rect -143 -1207 -85 -1173
rect -143 -1241 -131 -1207
rect -97 -1241 -85 -1207
rect -143 -1275 -85 -1241
rect -143 -1309 -131 -1275
rect -97 -1309 -85 -1275
rect -143 -1343 -85 -1309
rect -143 -1377 -131 -1343
rect -97 -1377 -85 -1343
rect -143 -1411 -85 -1377
rect -143 -1445 -131 -1411
rect -97 -1445 -85 -1411
rect -143 -1479 -85 -1445
rect -143 -1513 -131 -1479
rect -97 -1513 -85 -1479
rect -143 -1547 -85 -1513
rect -143 -1581 -131 -1547
rect -97 -1581 -85 -1547
rect -143 -1615 -85 -1581
rect -143 -1649 -131 -1615
rect -97 -1649 -85 -1615
rect -143 -1683 -85 -1649
rect -143 -1717 -131 -1683
rect -97 -1717 -85 -1683
rect -143 -1751 -85 -1717
rect -143 -1785 -131 -1751
rect -97 -1785 -85 -1751
rect -143 -1819 -85 -1785
rect -143 -1853 -131 -1819
rect -97 -1853 -85 -1819
rect -143 -1887 -85 -1853
rect -143 -1921 -131 -1887
rect -97 -1921 -85 -1887
rect -143 -1955 -85 -1921
rect -143 -1989 -131 -1955
rect -97 -1989 -85 -1955
rect -143 -2023 -85 -1989
rect -143 -2057 -131 -2023
rect -97 -2057 -85 -2023
rect -143 -2091 -85 -2057
rect -143 -2125 -131 -2091
rect -97 -2125 -85 -2091
rect -143 -2159 -85 -2125
rect -143 -2193 -131 -2159
rect -97 -2193 -85 -2159
rect -143 -2227 -85 -2193
rect -143 -2261 -131 -2227
rect -97 -2261 -85 -2227
rect -143 -2295 -85 -2261
rect -143 -2329 -131 -2295
rect -97 -2329 -85 -2295
rect -143 -2363 -85 -2329
rect -143 -2397 -131 -2363
rect -97 -2397 -85 -2363
rect -143 -2431 -85 -2397
rect -143 -2465 -131 -2431
rect -97 -2465 -85 -2431
rect -143 -2480 -85 -2465
rect -29 2465 29 2480
rect -29 2431 -17 2465
rect 17 2431 29 2465
rect -29 2397 29 2431
rect -29 2363 -17 2397
rect 17 2363 29 2397
rect -29 2329 29 2363
rect -29 2295 -17 2329
rect 17 2295 29 2329
rect -29 2261 29 2295
rect -29 2227 -17 2261
rect 17 2227 29 2261
rect -29 2193 29 2227
rect -29 2159 -17 2193
rect 17 2159 29 2193
rect -29 2125 29 2159
rect -29 2091 -17 2125
rect 17 2091 29 2125
rect -29 2057 29 2091
rect -29 2023 -17 2057
rect 17 2023 29 2057
rect -29 1989 29 2023
rect -29 1955 -17 1989
rect 17 1955 29 1989
rect -29 1921 29 1955
rect -29 1887 -17 1921
rect 17 1887 29 1921
rect -29 1853 29 1887
rect -29 1819 -17 1853
rect 17 1819 29 1853
rect -29 1785 29 1819
rect -29 1751 -17 1785
rect 17 1751 29 1785
rect -29 1717 29 1751
rect -29 1683 -17 1717
rect 17 1683 29 1717
rect -29 1649 29 1683
rect -29 1615 -17 1649
rect 17 1615 29 1649
rect -29 1581 29 1615
rect -29 1547 -17 1581
rect 17 1547 29 1581
rect -29 1513 29 1547
rect -29 1479 -17 1513
rect 17 1479 29 1513
rect -29 1445 29 1479
rect -29 1411 -17 1445
rect 17 1411 29 1445
rect -29 1377 29 1411
rect -29 1343 -17 1377
rect 17 1343 29 1377
rect -29 1309 29 1343
rect -29 1275 -17 1309
rect 17 1275 29 1309
rect -29 1241 29 1275
rect -29 1207 -17 1241
rect 17 1207 29 1241
rect -29 1173 29 1207
rect -29 1139 -17 1173
rect 17 1139 29 1173
rect -29 1105 29 1139
rect -29 1071 -17 1105
rect 17 1071 29 1105
rect -29 1037 29 1071
rect -29 1003 -17 1037
rect 17 1003 29 1037
rect -29 969 29 1003
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1003 29 -969
rect -29 -1037 -17 -1003
rect 17 -1037 29 -1003
rect -29 -1071 29 -1037
rect -29 -1105 -17 -1071
rect 17 -1105 29 -1071
rect -29 -1139 29 -1105
rect -29 -1173 -17 -1139
rect 17 -1173 29 -1139
rect -29 -1207 29 -1173
rect -29 -1241 -17 -1207
rect 17 -1241 29 -1207
rect -29 -1275 29 -1241
rect -29 -1309 -17 -1275
rect 17 -1309 29 -1275
rect -29 -1343 29 -1309
rect -29 -1377 -17 -1343
rect 17 -1377 29 -1343
rect -29 -1411 29 -1377
rect -29 -1445 -17 -1411
rect 17 -1445 29 -1411
rect -29 -1479 29 -1445
rect -29 -1513 -17 -1479
rect 17 -1513 29 -1479
rect -29 -1547 29 -1513
rect -29 -1581 -17 -1547
rect 17 -1581 29 -1547
rect -29 -1615 29 -1581
rect -29 -1649 -17 -1615
rect 17 -1649 29 -1615
rect -29 -1683 29 -1649
rect -29 -1717 -17 -1683
rect 17 -1717 29 -1683
rect -29 -1751 29 -1717
rect -29 -1785 -17 -1751
rect 17 -1785 29 -1751
rect -29 -1819 29 -1785
rect -29 -1853 -17 -1819
rect 17 -1853 29 -1819
rect -29 -1887 29 -1853
rect -29 -1921 -17 -1887
rect 17 -1921 29 -1887
rect -29 -1955 29 -1921
rect -29 -1989 -17 -1955
rect 17 -1989 29 -1955
rect -29 -2023 29 -1989
rect -29 -2057 -17 -2023
rect 17 -2057 29 -2023
rect -29 -2091 29 -2057
rect -29 -2125 -17 -2091
rect 17 -2125 29 -2091
rect -29 -2159 29 -2125
rect -29 -2193 -17 -2159
rect 17 -2193 29 -2159
rect -29 -2227 29 -2193
rect -29 -2261 -17 -2227
rect 17 -2261 29 -2227
rect -29 -2295 29 -2261
rect -29 -2329 -17 -2295
rect 17 -2329 29 -2295
rect -29 -2363 29 -2329
rect -29 -2397 -17 -2363
rect 17 -2397 29 -2363
rect -29 -2431 29 -2397
rect -29 -2465 -17 -2431
rect 17 -2465 29 -2431
rect -29 -2480 29 -2465
rect 85 2465 143 2480
rect 85 2431 97 2465
rect 131 2431 143 2465
rect 85 2397 143 2431
rect 85 2363 97 2397
rect 131 2363 143 2397
rect 85 2329 143 2363
rect 85 2295 97 2329
rect 131 2295 143 2329
rect 85 2261 143 2295
rect 85 2227 97 2261
rect 131 2227 143 2261
rect 85 2193 143 2227
rect 85 2159 97 2193
rect 131 2159 143 2193
rect 85 2125 143 2159
rect 85 2091 97 2125
rect 131 2091 143 2125
rect 85 2057 143 2091
rect 85 2023 97 2057
rect 131 2023 143 2057
rect 85 1989 143 2023
rect 85 1955 97 1989
rect 131 1955 143 1989
rect 85 1921 143 1955
rect 85 1887 97 1921
rect 131 1887 143 1921
rect 85 1853 143 1887
rect 85 1819 97 1853
rect 131 1819 143 1853
rect 85 1785 143 1819
rect 85 1751 97 1785
rect 131 1751 143 1785
rect 85 1717 143 1751
rect 85 1683 97 1717
rect 131 1683 143 1717
rect 85 1649 143 1683
rect 85 1615 97 1649
rect 131 1615 143 1649
rect 85 1581 143 1615
rect 85 1547 97 1581
rect 131 1547 143 1581
rect 85 1513 143 1547
rect 85 1479 97 1513
rect 131 1479 143 1513
rect 85 1445 143 1479
rect 85 1411 97 1445
rect 131 1411 143 1445
rect 85 1377 143 1411
rect 85 1343 97 1377
rect 131 1343 143 1377
rect 85 1309 143 1343
rect 85 1275 97 1309
rect 131 1275 143 1309
rect 85 1241 143 1275
rect 85 1207 97 1241
rect 131 1207 143 1241
rect 85 1173 143 1207
rect 85 1139 97 1173
rect 131 1139 143 1173
rect 85 1105 143 1139
rect 85 1071 97 1105
rect 131 1071 143 1105
rect 85 1037 143 1071
rect 85 1003 97 1037
rect 131 1003 143 1037
rect 85 969 143 1003
rect 85 935 97 969
rect 131 935 143 969
rect 85 901 143 935
rect 85 867 97 901
rect 131 867 143 901
rect 85 833 143 867
rect 85 799 97 833
rect 131 799 143 833
rect 85 765 143 799
rect 85 731 97 765
rect 131 731 143 765
rect 85 697 143 731
rect 85 663 97 697
rect 131 663 143 697
rect 85 629 143 663
rect 85 595 97 629
rect 131 595 143 629
rect 85 561 143 595
rect 85 527 97 561
rect 131 527 143 561
rect 85 493 143 527
rect 85 459 97 493
rect 131 459 143 493
rect 85 425 143 459
rect 85 391 97 425
rect 131 391 143 425
rect 85 357 143 391
rect 85 323 97 357
rect 131 323 143 357
rect 85 289 143 323
rect 85 255 97 289
rect 131 255 143 289
rect 85 221 143 255
rect 85 187 97 221
rect 131 187 143 221
rect 85 153 143 187
rect 85 119 97 153
rect 131 119 143 153
rect 85 85 143 119
rect 85 51 97 85
rect 131 51 143 85
rect 85 17 143 51
rect 85 -17 97 17
rect 131 -17 143 17
rect 85 -51 143 -17
rect 85 -85 97 -51
rect 131 -85 143 -51
rect 85 -119 143 -85
rect 85 -153 97 -119
rect 131 -153 143 -119
rect 85 -187 143 -153
rect 85 -221 97 -187
rect 131 -221 143 -187
rect 85 -255 143 -221
rect 85 -289 97 -255
rect 131 -289 143 -255
rect 85 -323 143 -289
rect 85 -357 97 -323
rect 131 -357 143 -323
rect 85 -391 143 -357
rect 85 -425 97 -391
rect 131 -425 143 -391
rect 85 -459 143 -425
rect 85 -493 97 -459
rect 131 -493 143 -459
rect 85 -527 143 -493
rect 85 -561 97 -527
rect 131 -561 143 -527
rect 85 -595 143 -561
rect 85 -629 97 -595
rect 131 -629 143 -595
rect 85 -663 143 -629
rect 85 -697 97 -663
rect 131 -697 143 -663
rect 85 -731 143 -697
rect 85 -765 97 -731
rect 131 -765 143 -731
rect 85 -799 143 -765
rect 85 -833 97 -799
rect 131 -833 143 -799
rect 85 -867 143 -833
rect 85 -901 97 -867
rect 131 -901 143 -867
rect 85 -935 143 -901
rect 85 -969 97 -935
rect 131 -969 143 -935
rect 85 -1003 143 -969
rect 85 -1037 97 -1003
rect 131 -1037 143 -1003
rect 85 -1071 143 -1037
rect 85 -1105 97 -1071
rect 131 -1105 143 -1071
rect 85 -1139 143 -1105
rect 85 -1173 97 -1139
rect 131 -1173 143 -1139
rect 85 -1207 143 -1173
rect 85 -1241 97 -1207
rect 131 -1241 143 -1207
rect 85 -1275 143 -1241
rect 85 -1309 97 -1275
rect 131 -1309 143 -1275
rect 85 -1343 143 -1309
rect 85 -1377 97 -1343
rect 131 -1377 143 -1343
rect 85 -1411 143 -1377
rect 85 -1445 97 -1411
rect 131 -1445 143 -1411
rect 85 -1479 143 -1445
rect 85 -1513 97 -1479
rect 131 -1513 143 -1479
rect 85 -1547 143 -1513
rect 85 -1581 97 -1547
rect 131 -1581 143 -1547
rect 85 -1615 143 -1581
rect 85 -1649 97 -1615
rect 131 -1649 143 -1615
rect 85 -1683 143 -1649
rect 85 -1717 97 -1683
rect 131 -1717 143 -1683
rect 85 -1751 143 -1717
rect 85 -1785 97 -1751
rect 131 -1785 143 -1751
rect 85 -1819 143 -1785
rect 85 -1853 97 -1819
rect 131 -1853 143 -1819
rect 85 -1887 143 -1853
rect 85 -1921 97 -1887
rect 131 -1921 143 -1887
rect 85 -1955 143 -1921
rect 85 -1989 97 -1955
rect 131 -1989 143 -1955
rect 85 -2023 143 -1989
rect 85 -2057 97 -2023
rect 131 -2057 143 -2023
rect 85 -2091 143 -2057
rect 85 -2125 97 -2091
rect 131 -2125 143 -2091
rect 85 -2159 143 -2125
rect 85 -2193 97 -2159
rect 131 -2193 143 -2159
rect 85 -2227 143 -2193
rect 85 -2261 97 -2227
rect 131 -2261 143 -2227
rect 85 -2295 143 -2261
rect 85 -2329 97 -2295
rect 131 -2329 143 -2295
rect 85 -2363 143 -2329
rect 85 -2397 97 -2363
rect 131 -2397 143 -2363
rect 85 -2431 143 -2397
rect 85 -2465 97 -2431
rect 131 -2465 143 -2431
rect 85 -2480 143 -2465
rect 199 2465 257 2480
rect 199 2431 211 2465
rect 245 2431 257 2465
rect 199 2397 257 2431
rect 199 2363 211 2397
rect 245 2363 257 2397
rect 199 2329 257 2363
rect 199 2295 211 2329
rect 245 2295 257 2329
rect 199 2261 257 2295
rect 199 2227 211 2261
rect 245 2227 257 2261
rect 199 2193 257 2227
rect 199 2159 211 2193
rect 245 2159 257 2193
rect 199 2125 257 2159
rect 199 2091 211 2125
rect 245 2091 257 2125
rect 199 2057 257 2091
rect 199 2023 211 2057
rect 245 2023 257 2057
rect 199 1989 257 2023
rect 199 1955 211 1989
rect 245 1955 257 1989
rect 199 1921 257 1955
rect 199 1887 211 1921
rect 245 1887 257 1921
rect 199 1853 257 1887
rect 199 1819 211 1853
rect 245 1819 257 1853
rect 199 1785 257 1819
rect 199 1751 211 1785
rect 245 1751 257 1785
rect 199 1717 257 1751
rect 199 1683 211 1717
rect 245 1683 257 1717
rect 199 1649 257 1683
rect 199 1615 211 1649
rect 245 1615 257 1649
rect 199 1581 257 1615
rect 199 1547 211 1581
rect 245 1547 257 1581
rect 199 1513 257 1547
rect 199 1479 211 1513
rect 245 1479 257 1513
rect 199 1445 257 1479
rect 199 1411 211 1445
rect 245 1411 257 1445
rect 199 1377 257 1411
rect 199 1343 211 1377
rect 245 1343 257 1377
rect 199 1309 257 1343
rect 199 1275 211 1309
rect 245 1275 257 1309
rect 199 1241 257 1275
rect 199 1207 211 1241
rect 245 1207 257 1241
rect 199 1173 257 1207
rect 199 1139 211 1173
rect 245 1139 257 1173
rect 199 1105 257 1139
rect 199 1071 211 1105
rect 245 1071 257 1105
rect 199 1037 257 1071
rect 199 1003 211 1037
rect 245 1003 257 1037
rect 199 969 257 1003
rect 199 935 211 969
rect 245 935 257 969
rect 199 901 257 935
rect 199 867 211 901
rect 245 867 257 901
rect 199 833 257 867
rect 199 799 211 833
rect 245 799 257 833
rect 199 765 257 799
rect 199 731 211 765
rect 245 731 257 765
rect 199 697 257 731
rect 199 663 211 697
rect 245 663 257 697
rect 199 629 257 663
rect 199 595 211 629
rect 245 595 257 629
rect 199 561 257 595
rect 199 527 211 561
rect 245 527 257 561
rect 199 493 257 527
rect 199 459 211 493
rect 245 459 257 493
rect 199 425 257 459
rect 199 391 211 425
rect 245 391 257 425
rect 199 357 257 391
rect 199 323 211 357
rect 245 323 257 357
rect 199 289 257 323
rect 199 255 211 289
rect 245 255 257 289
rect 199 221 257 255
rect 199 187 211 221
rect 245 187 257 221
rect 199 153 257 187
rect 199 119 211 153
rect 245 119 257 153
rect 199 85 257 119
rect 199 51 211 85
rect 245 51 257 85
rect 199 17 257 51
rect 199 -17 211 17
rect 245 -17 257 17
rect 199 -51 257 -17
rect 199 -85 211 -51
rect 245 -85 257 -51
rect 199 -119 257 -85
rect 199 -153 211 -119
rect 245 -153 257 -119
rect 199 -187 257 -153
rect 199 -221 211 -187
rect 245 -221 257 -187
rect 199 -255 257 -221
rect 199 -289 211 -255
rect 245 -289 257 -255
rect 199 -323 257 -289
rect 199 -357 211 -323
rect 245 -357 257 -323
rect 199 -391 257 -357
rect 199 -425 211 -391
rect 245 -425 257 -391
rect 199 -459 257 -425
rect 199 -493 211 -459
rect 245 -493 257 -459
rect 199 -527 257 -493
rect 199 -561 211 -527
rect 245 -561 257 -527
rect 199 -595 257 -561
rect 199 -629 211 -595
rect 245 -629 257 -595
rect 199 -663 257 -629
rect 199 -697 211 -663
rect 245 -697 257 -663
rect 199 -731 257 -697
rect 199 -765 211 -731
rect 245 -765 257 -731
rect 199 -799 257 -765
rect 199 -833 211 -799
rect 245 -833 257 -799
rect 199 -867 257 -833
rect 199 -901 211 -867
rect 245 -901 257 -867
rect 199 -935 257 -901
rect 199 -969 211 -935
rect 245 -969 257 -935
rect 199 -1003 257 -969
rect 199 -1037 211 -1003
rect 245 -1037 257 -1003
rect 199 -1071 257 -1037
rect 199 -1105 211 -1071
rect 245 -1105 257 -1071
rect 199 -1139 257 -1105
rect 199 -1173 211 -1139
rect 245 -1173 257 -1139
rect 199 -1207 257 -1173
rect 199 -1241 211 -1207
rect 245 -1241 257 -1207
rect 199 -1275 257 -1241
rect 199 -1309 211 -1275
rect 245 -1309 257 -1275
rect 199 -1343 257 -1309
rect 199 -1377 211 -1343
rect 245 -1377 257 -1343
rect 199 -1411 257 -1377
rect 199 -1445 211 -1411
rect 245 -1445 257 -1411
rect 199 -1479 257 -1445
rect 199 -1513 211 -1479
rect 245 -1513 257 -1479
rect 199 -1547 257 -1513
rect 199 -1581 211 -1547
rect 245 -1581 257 -1547
rect 199 -1615 257 -1581
rect 199 -1649 211 -1615
rect 245 -1649 257 -1615
rect 199 -1683 257 -1649
rect 199 -1717 211 -1683
rect 245 -1717 257 -1683
rect 199 -1751 257 -1717
rect 199 -1785 211 -1751
rect 245 -1785 257 -1751
rect 199 -1819 257 -1785
rect 199 -1853 211 -1819
rect 245 -1853 257 -1819
rect 199 -1887 257 -1853
rect 199 -1921 211 -1887
rect 245 -1921 257 -1887
rect 199 -1955 257 -1921
rect 199 -1989 211 -1955
rect 245 -1989 257 -1955
rect 199 -2023 257 -1989
rect 199 -2057 211 -2023
rect 245 -2057 257 -2023
rect 199 -2091 257 -2057
rect 199 -2125 211 -2091
rect 245 -2125 257 -2091
rect 199 -2159 257 -2125
rect 199 -2193 211 -2159
rect 245 -2193 257 -2159
rect 199 -2227 257 -2193
rect 199 -2261 211 -2227
rect 245 -2261 257 -2227
rect 199 -2295 257 -2261
rect 199 -2329 211 -2295
rect 245 -2329 257 -2295
rect 199 -2363 257 -2329
rect 199 -2397 211 -2363
rect 245 -2397 257 -2363
rect 199 -2431 257 -2397
rect 199 -2465 211 -2431
rect 245 -2465 257 -2431
rect 199 -2480 257 -2465
<< ndiffc >>
rect -245 2431 -211 2465
rect -245 2363 -211 2397
rect -245 2295 -211 2329
rect -245 2227 -211 2261
rect -245 2159 -211 2193
rect -245 2091 -211 2125
rect -245 2023 -211 2057
rect -245 1955 -211 1989
rect -245 1887 -211 1921
rect -245 1819 -211 1853
rect -245 1751 -211 1785
rect -245 1683 -211 1717
rect -245 1615 -211 1649
rect -245 1547 -211 1581
rect -245 1479 -211 1513
rect -245 1411 -211 1445
rect -245 1343 -211 1377
rect -245 1275 -211 1309
rect -245 1207 -211 1241
rect -245 1139 -211 1173
rect -245 1071 -211 1105
rect -245 1003 -211 1037
rect -245 935 -211 969
rect -245 867 -211 901
rect -245 799 -211 833
rect -245 731 -211 765
rect -245 663 -211 697
rect -245 595 -211 629
rect -245 527 -211 561
rect -245 459 -211 493
rect -245 391 -211 425
rect -245 323 -211 357
rect -245 255 -211 289
rect -245 187 -211 221
rect -245 119 -211 153
rect -245 51 -211 85
rect -245 -17 -211 17
rect -245 -85 -211 -51
rect -245 -153 -211 -119
rect -245 -221 -211 -187
rect -245 -289 -211 -255
rect -245 -357 -211 -323
rect -245 -425 -211 -391
rect -245 -493 -211 -459
rect -245 -561 -211 -527
rect -245 -629 -211 -595
rect -245 -697 -211 -663
rect -245 -765 -211 -731
rect -245 -833 -211 -799
rect -245 -901 -211 -867
rect -245 -969 -211 -935
rect -245 -1037 -211 -1003
rect -245 -1105 -211 -1071
rect -245 -1173 -211 -1139
rect -245 -1241 -211 -1207
rect -245 -1309 -211 -1275
rect -245 -1377 -211 -1343
rect -245 -1445 -211 -1411
rect -245 -1513 -211 -1479
rect -245 -1581 -211 -1547
rect -245 -1649 -211 -1615
rect -245 -1717 -211 -1683
rect -245 -1785 -211 -1751
rect -245 -1853 -211 -1819
rect -245 -1921 -211 -1887
rect -245 -1989 -211 -1955
rect -245 -2057 -211 -2023
rect -245 -2125 -211 -2091
rect -245 -2193 -211 -2159
rect -245 -2261 -211 -2227
rect -245 -2329 -211 -2295
rect -245 -2397 -211 -2363
rect -245 -2465 -211 -2431
rect -131 2431 -97 2465
rect -131 2363 -97 2397
rect -131 2295 -97 2329
rect -131 2227 -97 2261
rect -131 2159 -97 2193
rect -131 2091 -97 2125
rect -131 2023 -97 2057
rect -131 1955 -97 1989
rect -131 1887 -97 1921
rect -131 1819 -97 1853
rect -131 1751 -97 1785
rect -131 1683 -97 1717
rect -131 1615 -97 1649
rect -131 1547 -97 1581
rect -131 1479 -97 1513
rect -131 1411 -97 1445
rect -131 1343 -97 1377
rect -131 1275 -97 1309
rect -131 1207 -97 1241
rect -131 1139 -97 1173
rect -131 1071 -97 1105
rect -131 1003 -97 1037
rect -131 935 -97 969
rect -131 867 -97 901
rect -131 799 -97 833
rect -131 731 -97 765
rect -131 663 -97 697
rect -131 595 -97 629
rect -131 527 -97 561
rect -131 459 -97 493
rect -131 391 -97 425
rect -131 323 -97 357
rect -131 255 -97 289
rect -131 187 -97 221
rect -131 119 -97 153
rect -131 51 -97 85
rect -131 -17 -97 17
rect -131 -85 -97 -51
rect -131 -153 -97 -119
rect -131 -221 -97 -187
rect -131 -289 -97 -255
rect -131 -357 -97 -323
rect -131 -425 -97 -391
rect -131 -493 -97 -459
rect -131 -561 -97 -527
rect -131 -629 -97 -595
rect -131 -697 -97 -663
rect -131 -765 -97 -731
rect -131 -833 -97 -799
rect -131 -901 -97 -867
rect -131 -969 -97 -935
rect -131 -1037 -97 -1003
rect -131 -1105 -97 -1071
rect -131 -1173 -97 -1139
rect -131 -1241 -97 -1207
rect -131 -1309 -97 -1275
rect -131 -1377 -97 -1343
rect -131 -1445 -97 -1411
rect -131 -1513 -97 -1479
rect -131 -1581 -97 -1547
rect -131 -1649 -97 -1615
rect -131 -1717 -97 -1683
rect -131 -1785 -97 -1751
rect -131 -1853 -97 -1819
rect -131 -1921 -97 -1887
rect -131 -1989 -97 -1955
rect -131 -2057 -97 -2023
rect -131 -2125 -97 -2091
rect -131 -2193 -97 -2159
rect -131 -2261 -97 -2227
rect -131 -2329 -97 -2295
rect -131 -2397 -97 -2363
rect -131 -2465 -97 -2431
rect -17 2431 17 2465
rect -17 2363 17 2397
rect -17 2295 17 2329
rect -17 2227 17 2261
rect -17 2159 17 2193
rect -17 2091 17 2125
rect -17 2023 17 2057
rect -17 1955 17 1989
rect -17 1887 17 1921
rect -17 1819 17 1853
rect -17 1751 17 1785
rect -17 1683 17 1717
rect -17 1615 17 1649
rect -17 1547 17 1581
rect -17 1479 17 1513
rect -17 1411 17 1445
rect -17 1343 17 1377
rect -17 1275 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1173
rect -17 1071 17 1105
rect -17 1003 17 1037
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect -17 -1037 17 -1003
rect -17 -1105 17 -1071
rect -17 -1173 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1275
rect -17 -1377 17 -1343
rect -17 -1445 17 -1411
rect -17 -1513 17 -1479
rect -17 -1581 17 -1547
rect -17 -1649 17 -1615
rect -17 -1717 17 -1683
rect -17 -1785 17 -1751
rect -17 -1853 17 -1819
rect -17 -1921 17 -1887
rect -17 -1989 17 -1955
rect -17 -2057 17 -2023
rect -17 -2125 17 -2091
rect -17 -2193 17 -2159
rect -17 -2261 17 -2227
rect -17 -2329 17 -2295
rect -17 -2397 17 -2363
rect -17 -2465 17 -2431
rect 97 2431 131 2465
rect 97 2363 131 2397
rect 97 2295 131 2329
rect 97 2227 131 2261
rect 97 2159 131 2193
rect 97 2091 131 2125
rect 97 2023 131 2057
rect 97 1955 131 1989
rect 97 1887 131 1921
rect 97 1819 131 1853
rect 97 1751 131 1785
rect 97 1683 131 1717
rect 97 1615 131 1649
rect 97 1547 131 1581
rect 97 1479 131 1513
rect 97 1411 131 1445
rect 97 1343 131 1377
rect 97 1275 131 1309
rect 97 1207 131 1241
rect 97 1139 131 1173
rect 97 1071 131 1105
rect 97 1003 131 1037
rect 97 935 131 969
rect 97 867 131 901
rect 97 799 131 833
rect 97 731 131 765
rect 97 663 131 697
rect 97 595 131 629
rect 97 527 131 561
rect 97 459 131 493
rect 97 391 131 425
rect 97 323 131 357
rect 97 255 131 289
rect 97 187 131 221
rect 97 119 131 153
rect 97 51 131 85
rect 97 -17 131 17
rect 97 -85 131 -51
rect 97 -153 131 -119
rect 97 -221 131 -187
rect 97 -289 131 -255
rect 97 -357 131 -323
rect 97 -425 131 -391
rect 97 -493 131 -459
rect 97 -561 131 -527
rect 97 -629 131 -595
rect 97 -697 131 -663
rect 97 -765 131 -731
rect 97 -833 131 -799
rect 97 -901 131 -867
rect 97 -969 131 -935
rect 97 -1037 131 -1003
rect 97 -1105 131 -1071
rect 97 -1173 131 -1139
rect 97 -1241 131 -1207
rect 97 -1309 131 -1275
rect 97 -1377 131 -1343
rect 97 -1445 131 -1411
rect 97 -1513 131 -1479
rect 97 -1581 131 -1547
rect 97 -1649 131 -1615
rect 97 -1717 131 -1683
rect 97 -1785 131 -1751
rect 97 -1853 131 -1819
rect 97 -1921 131 -1887
rect 97 -1989 131 -1955
rect 97 -2057 131 -2023
rect 97 -2125 131 -2091
rect 97 -2193 131 -2159
rect 97 -2261 131 -2227
rect 97 -2329 131 -2295
rect 97 -2397 131 -2363
rect 97 -2465 131 -2431
rect 211 2431 245 2465
rect 211 2363 245 2397
rect 211 2295 245 2329
rect 211 2227 245 2261
rect 211 2159 245 2193
rect 211 2091 245 2125
rect 211 2023 245 2057
rect 211 1955 245 1989
rect 211 1887 245 1921
rect 211 1819 245 1853
rect 211 1751 245 1785
rect 211 1683 245 1717
rect 211 1615 245 1649
rect 211 1547 245 1581
rect 211 1479 245 1513
rect 211 1411 245 1445
rect 211 1343 245 1377
rect 211 1275 245 1309
rect 211 1207 245 1241
rect 211 1139 245 1173
rect 211 1071 245 1105
rect 211 1003 245 1037
rect 211 935 245 969
rect 211 867 245 901
rect 211 799 245 833
rect 211 731 245 765
rect 211 663 245 697
rect 211 595 245 629
rect 211 527 245 561
rect 211 459 245 493
rect 211 391 245 425
rect 211 323 245 357
rect 211 255 245 289
rect 211 187 245 221
rect 211 119 245 153
rect 211 51 245 85
rect 211 -17 245 17
rect 211 -85 245 -51
rect 211 -153 245 -119
rect 211 -221 245 -187
rect 211 -289 245 -255
rect 211 -357 245 -323
rect 211 -425 245 -391
rect 211 -493 245 -459
rect 211 -561 245 -527
rect 211 -629 245 -595
rect 211 -697 245 -663
rect 211 -765 245 -731
rect 211 -833 245 -799
rect 211 -901 245 -867
rect 211 -969 245 -935
rect 211 -1037 245 -1003
rect 211 -1105 245 -1071
rect 211 -1173 245 -1139
rect 211 -1241 245 -1207
rect 211 -1309 245 -1275
rect 211 -1377 245 -1343
rect 211 -1445 245 -1411
rect 211 -1513 245 -1479
rect 211 -1581 245 -1547
rect 211 -1649 245 -1615
rect 211 -1717 245 -1683
rect 211 -1785 245 -1751
rect 211 -1853 245 -1819
rect 211 -1921 245 -1887
rect 211 -1989 245 -1955
rect 211 -2057 245 -2023
rect 211 -2125 245 -2091
rect 211 -2193 245 -2159
rect 211 -2261 245 -2227
rect 211 -2329 245 -2295
rect 211 -2397 245 -2363
rect 211 -2465 245 -2431
<< poly >>
rect -204 2502 -138 2568
rect -90 2510 90 2568
rect -90 2502 -24 2510
rect 24 2502 90 2510
rect 138 2556 204 2568
rect 138 2522 154 2556
rect 188 2522 204 2556
rect 138 2502 204 2522
rect -199 2480 -143 2502
rect -85 2480 -29 2502
rect 29 2480 85 2502
rect 143 2480 199 2502
rect -199 -2502 -143 -2480
rect -85 -2502 -29 -2480
rect 29 -2502 85 -2480
rect 143 -2502 199 -2480
rect -204 -2504 -138 -2502
rect -90 -2504 -24 -2502
rect -204 -2568 -24 -2504
rect 24 -2510 90 -2502
rect 138 -2510 204 -2502
rect 24 -2568 204 -2510
<< polycont >>
rect 154 2522 188 2556
<< locali >>
rect 138 2522 154 2556
rect 188 2522 204 2556
rect -245 2465 -211 2484
rect -245 2397 -211 2431
rect -245 2329 -211 2359
rect -245 2261 -211 2287
rect -245 2193 -211 2215
rect -245 2125 -211 2143
rect -245 2057 -211 2071
rect -245 1989 -211 1999
rect -245 1921 -211 1927
rect -245 1853 -211 1855
rect -245 1817 -211 1819
rect -245 1745 -211 1751
rect -245 1673 -211 1683
rect -245 1601 -211 1615
rect -245 1529 -211 1547
rect -245 1457 -211 1479
rect -245 1385 -211 1411
rect -245 1313 -211 1343
rect -245 1241 -211 1275
rect -245 1173 -211 1207
rect -245 1105 -211 1135
rect -245 1037 -211 1063
rect -245 969 -211 991
rect -245 901 -211 919
rect -245 833 -211 847
rect -245 765 -211 775
rect -245 697 -211 703
rect -245 629 -211 631
rect -245 593 -211 595
rect -245 521 -211 527
rect -245 449 -211 459
rect -245 377 -211 391
rect -245 305 -211 323
rect -245 233 -211 255
rect -245 161 -211 187
rect -245 89 -211 119
rect -245 17 -211 51
rect -245 -51 -211 -17
rect -245 -119 -211 -89
rect -245 -187 -211 -161
rect -245 -255 -211 -233
rect -245 -323 -211 -305
rect -245 -391 -211 -377
rect -245 -459 -211 -449
rect -245 -527 -211 -521
rect -245 -595 -211 -593
rect -245 -631 -211 -629
rect -245 -703 -211 -697
rect -245 -775 -211 -765
rect -245 -847 -211 -833
rect -245 -919 -211 -901
rect -245 -991 -211 -969
rect -245 -1063 -211 -1037
rect -245 -1135 -211 -1105
rect -245 -1207 -211 -1173
rect -245 -1275 -211 -1241
rect -245 -1343 -211 -1313
rect -245 -1411 -211 -1385
rect -245 -1479 -211 -1457
rect -245 -1547 -211 -1529
rect -245 -1615 -211 -1601
rect -245 -1683 -211 -1673
rect -245 -1751 -211 -1745
rect -245 -1819 -211 -1817
rect -245 -1855 -211 -1853
rect -245 -1927 -211 -1921
rect -245 -1999 -211 -1989
rect -245 -2071 -211 -2057
rect -245 -2143 -211 -2125
rect -245 -2215 -211 -2193
rect -245 -2287 -211 -2261
rect -245 -2359 -211 -2329
rect -245 -2431 -211 -2397
rect -245 -2484 -211 -2465
rect -131 2465 -97 2484
rect -131 2397 -97 2431
rect -131 2329 -97 2359
rect -131 2261 -97 2287
rect -131 2193 -97 2215
rect -131 2125 -97 2143
rect -131 2057 -97 2071
rect -131 1989 -97 1999
rect -131 1921 -97 1927
rect -131 1853 -97 1855
rect -131 1817 -97 1819
rect -131 1745 -97 1751
rect -131 1673 -97 1683
rect -131 1601 -97 1615
rect -131 1529 -97 1547
rect -131 1457 -97 1479
rect -131 1385 -97 1411
rect -131 1313 -97 1343
rect -131 1241 -97 1275
rect -131 1173 -97 1207
rect -131 1105 -97 1135
rect -131 1037 -97 1063
rect -131 969 -97 991
rect -131 901 -97 919
rect -131 833 -97 847
rect -131 765 -97 775
rect -131 697 -97 703
rect -131 629 -97 631
rect -131 593 -97 595
rect -131 521 -97 527
rect -131 449 -97 459
rect -131 377 -97 391
rect -131 305 -97 323
rect -131 233 -97 255
rect -131 161 -97 187
rect -131 89 -97 119
rect -131 17 -97 51
rect -131 -51 -97 -17
rect -131 -119 -97 -89
rect -131 -187 -97 -161
rect -131 -255 -97 -233
rect -131 -323 -97 -305
rect -131 -391 -97 -377
rect -131 -459 -97 -449
rect -131 -527 -97 -521
rect -131 -595 -97 -593
rect -131 -631 -97 -629
rect -131 -703 -97 -697
rect -131 -775 -97 -765
rect -131 -847 -97 -833
rect -131 -919 -97 -901
rect -131 -991 -97 -969
rect -131 -1063 -97 -1037
rect -131 -1135 -97 -1105
rect -131 -1207 -97 -1173
rect -131 -1275 -97 -1241
rect -131 -1343 -97 -1313
rect -131 -1411 -97 -1385
rect -131 -1479 -97 -1457
rect -131 -1547 -97 -1529
rect -131 -1615 -97 -1601
rect -131 -1683 -97 -1673
rect -131 -1751 -97 -1745
rect -131 -1819 -97 -1817
rect -131 -1855 -97 -1853
rect -131 -1927 -97 -1921
rect -131 -1999 -97 -1989
rect -131 -2071 -97 -2057
rect -131 -2143 -97 -2125
rect -131 -2215 -97 -2193
rect -131 -2287 -97 -2261
rect -131 -2359 -97 -2329
rect -131 -2431 -97 -2397
rect -131 -2484 -97 -2465
rect -17 2465 17 2484
rect -17 2397 17 2431
rect -17 2329 17 2359
rect -17 2261 17 2287
rect -17 2193 17 2215
rect -17 2125 17 2143
rect -17 2057 17 2071
rect -17 1989 17 1999
rect -17 1921 17 1927
rect -17 1853 17 1855
rect -17 1817 17 1819
rect -17 1745 17 1751
rect -17 1673 17 1683
rect -17 1601 17 1615
rect -17 1529 17 1547
rect -17 1457 17 1479
rect -17 1385 17 1411
rect -17 1313 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1135
rect -17 1037 17 1063
rect -17 969 17 991
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -991 17 -969
rect -17 -1063 17 -1037
rect -17 -1135 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1313
rect -17 -1411 17 -1385
rect -17 -1479 17 -1457
rect -17 -1547 17 -1529
rect -17 -1615 17 -1601
rect -17 -1683 17 -1673
rect -17 -1751 17 -1745
rect -17 -1819 17 -1817
rect -17 -1855 17 -1853
rect -17 -1927 17 -1921
rect -17 -1999 17 -1989
rect -17 -2071 17 -2057
rect -17 -2143 17 -2125
rect -17 -2215 17 -2193
rect -17 -2287 17 -2261
rect -17 -2359 17 -2329
rect -17 -2431 17 -2397
rect -17 -2484 17 -2465
rect 97 2465 131 2484
rect 97 2397 131 2431
rect 97 2329 131 2359
rect 97 2261 131 2287
rect 97 2193 131 2215
rect 97 2125 131 2143
rect 97 2057 131 2071
rect 97 1989 131 1999
rect 97 1921 131 1927
rect 97 1853 131 1855
rect 97 1817 131 1819
rect 97 1745 131 1751
rect 97 1673 131 1683
rect 97 1601 131 1615
rect 97 1529 131 1547
rect 97 1457 131 1479
rect 97 1385 131 1411
rect 97 1313 131 1343
rect 97 1241 131 1275
rect 97 1173 131 1207
rect 97 1105 131 1135
rect 97 1037 131 1063
rect 97 969 131 991
rect 97 901 131 919
rect 97 833 131 847
rect 97 765 131 775
rect 97 697 131 703
rect 97 629 131 631
rect 97 593 131 595
rect 97 521 131 527
rect 97 449 131 459
rect 97 377 131 391
rect 97 305 131 323
rect 97 233 131 255
rect 97 161 131 187
rect 97 89 131 119
rect 97 17 131 51
rect 97 -51 131 -17
rect 97 -119 131 -89
rect 97 -187 131 -161
rect 97 -255 131 -233
rect 97 -323 131 -305
rect 97 -391 131 -377
rect 97 -459 131 -449
rect 97 -527 131 -521
rect 97 -595 131 -593
rect 97 -631 131 -629
rect 97 -703 131 -697
rect 97 -775 131 -765
rect 97 -847 131 -833
rect 97 -919 131 -901
rect 97 -991 131 -969
rect 97 -1063 131 -1037
rect 97 -1135 131 -1105
rect 97 -1207 131 -1173
rect 97 -1275 131 -1241
rect 97 -1343 131 -1313
rect 97 -1411 131 -1385
rect 97 -1479 131 -1457
rect 97 -1547 131 -1529
rect 97 -1615 131 -1601
rect 97 -1683 131 -1673
rect 97 -1751 131 -1745
rect 97 -1819 131 -1817
rect 97 -1855 131 -1853
rect 97 -1927 131 -1921
rect 97 -1999 131 -1989
rect 97 -2071 131 -2057
rect 97 -2143 131 -2125
rect 97 -2215 131 -2193
rect 97 -2287 131 -2261
rect 97 -2359 131 -2329
rect 97 -2431 131 -2397
rect 97 -2484 131 -2465
rect 211 2465 245 2484
rect 211 2397 245 2431
rect 211 2329 245 2359
rect 211 2261 245 2287
rect 211 2193 245 2215
rect 211 2125 245 2143
rect 211 2057 245 2071
rect 211 1989 245 1999
rect 211 1921 245 1927
rect 211 1853 245 1855
rect 211 1817 245 1819
rect 211 1745 245 1751
rect 211 1673 245 1683
rect 211 1601 245 1615
rect 211 1529 245 1547
rect 211 1457 245 1479
rect 211 1385 245 1411
rect 211 1313 245 1343
rect 211 1241 245 1275
rect 211 1173 245 1207
rect 211 1105 245 1135
rect 211 1037 245 1063
rect 211 969 245 991
rect 211 901 245 919
rect 211 833 245 847
rect 211 765 245 775
rect 211 697 245 703
rect 211 629 245 631
rect 211 593 245 595
rect 211 521 245 527
rect 211 449 245 459
rect 211 377 245 391
rect 211 305 245 323
rect 211 233 245 255
rect 211 161 245 187
rect 211 89 245 119
rect 211 17 245 51
rect 211 -51 245 -17
rect 211 -119 245 -89
rect 211 -187 245 -161
rect 211 -255 245 -233
rect 211 -323 245 -305
rect 211 -391 245 -377
rect 211 -459 245 -449
rect 211 -527 245 -521
rect 211 -595 245 -593
rect 211 -631 245 -629
rect 211 -703 245 -697
rect 211 -775 245 -765
rect 211 -847 245 -833
rect 211 -919 245 -901
rect 211 -991 245 -969
rect 211 -1063 245 -1037
rect 211 -1135 245 -1105
rect 211 -1207 245 -1173
rect 211 -1275 245 -1241
rect 211 -1343 245 -1313
rect 211 -1411 245 -1385
rect 211 -1479 245 -1457
rect 211 -1547 245 -1529
rect 211 -1615 245 -1601
rect 211 -1683 245 -1673
rect 211 -1751 245 -1745
rect 211 -1819 245 -1817
rect 211 -1855 245 -1853
rect 211 -1927 245 -1921
rect 211 -1999 245 -1989
rect 211 -2071 245 -2057
rect 211 -2143 245 -2125
rect 211 -2215 245 -2193
rect 211 -2287 245 -2261
rect 211 -2359 245 -2329
rect 211 -2431 245 -2397
rect 211 -2484 245 -2465
<< viali >>
rect 154 2522 188 2556
rect -245 2431 -211 2465
rect -245 2363 -211 2393
rect -245 2359 -211 2363
rect -245 2295 -211 2321
rect -245 2287 -211 2295
rect -245 2227 -211 2249
rect -245 2215 -211 2227
rect -245 2159 -211 2177
rect -245 2143 -211 2159
rect -245 2091 -211 2105
rect -245 2071 -211 2091
rect -245 2023 -211 2033
rect -245 1999 -211 2023
rect -245 1955 -211 1961
rect -245 1927 -211 1955
rect -245 1887 -211 1889
rect -245 1855 -211 1887
rect -245 1785 -211 1817
rect -245 1783 -211 1785
rect -245 1717 -211 1745
rect -245 1711 -211 1717
rect -245 1649 -211 1673
rect -245 1639 -211 1649
rect -245 1581 -211 1601
rect -245 1567 -211 1581
rect -245 1513 -211 1529
rect -245 1495 -211 1513
rect -245 1445 -211 1457
rect -245 1423 -211 1445
rect -245 1377 -211 1385
rect -245 1351 -211 1377
rect -245 1309 -211 1313
rect -245 1279 -211 1309
rect -245 1207 -211 1241
rect -245 1139 -211 1169
rect -245 1135 -211 1139
rect -245 1071 -211 1097
rect -245 1063 -211 1071
rect -245 1003 -211 1025
rect -245 991 -211 1003
rect -245 935 -211 953
rect -245 919 -211 935
rect -245 867 -211 881
rect -245 847 -211 867
rect -245 799 -211 809
rect -245 775 -211 799
rect -245 731 -211 737
rect -245 703 -211 731
rect -245 663 -211 665
rect -245 631 -211 663
rect -245 561 -211 593
rect -245 559 -211 561
rect -245 493 -211 521
rect -245 487 -211 493
rect -245 425 -211 449
rect -245 415 -211 425
rect -245 357 -211 377
rect -245 343 -211 357
rect -245 289 -211 305
rect -245 271 -211 289
rect -245 221 -211 233
rect -245 199 -211 221
rect -245 153 -211 161
rect -245 127 -211 153
rect -245 85 -211 89
rect -245 55 -211 85
rect -245 -17 -211 17
rect -245 -85 -211 -55
rect -245 -89 -211 -85
rect -245 -153 -211 -127
rect -245 -161 -211 -153
rect -245 -221 -211 -199
rect -245 -233 -211 -221
rect -245 -289 -211 -271
rect -245 -305 -211 -289
rect -245 -357 -211 -343
rect -245 -377 -211 -357
rect -245 -425 -211 -415
rect -245 -449 -211 -425
rect -245 -493 -211 -487
rect -245 -521 -211 -493
rect -245 -561 -211 -559
rect -245 -593 -211 -561
rect -245 -663 -211 -631
rect -245 -665 -211 -663
rect -245 -731 -211 -703
rect -245 -737 -211 -731
rect -245 -799 -211 -775
rect -245 -809 -211 -799
rect -245 -867 -211 -847
rect -245 -881 -211 -867
rect -245 -935 -211 -919
rect -245 -953 -211 -935
rect -245 -1003 -211 -991
rect -245 -1025 -211 -1003
rect -245 -1071 -211 -1063
rect -245 -1097 -211 -1071
rect -245 -1139 -211 -1135
rect -245 -1169 -211 -1139
rect -245 -1241 -211 -1207
rect -245 -1309 -211 -1279
rect -245 -1313 -211 -1309
rect -245 -1377 -211 -1351
rect -245 -1385 -211 -1377
rect -245 -1445 -211 -1423
rect -245 -1457 -211 -1445
rect -245 -1513 -211 -1495
rect -245 -1529 -211 -1513
rect -245 -1581 -211 -1567
rect -245 -1601 -211 -1581
rect -245 -1649 -211 -1639
rect -245 -1673 -211 -1649
rect -245 -1717 -211 -1711
rect -245 -1745 -211 -1717
rect -245 -1785 -211 -1783
rect -245 -1817 -211 -1785
rect -245 -1887 -211 -1855
rect -245 -1889 -211 -1887
rect -245 -1955 -211 -1927
rect -245 -1961 -211 -1955
rect -245 -2023 -211 -1999
rect -245 -2033 -211 -2023
rect -245 -2091 -211 -2071
rect -245 -2105 -211 -2091
rect -245 -2159 -211 -2143
rect -245 -2177 -211 -2159
rect -245 -2227 -211 -2215
rect -245 -2249 -211 -2227
rect -245 -2295 -211 -2287
rect -245 -2321 -211 -2295
rect -245 -2363 -211 -2359
rect -245 -2393 -211 -2363
rect -245 -2465 -211 -2431
rect -131 2431 -97 2465
rect -131 2363 -97 2393
rect -131 2359 -97 2363
rect -131 2295 -97 2321
rect -131 2287 -97 2295
rect -131 2227 -97 2249
rect -131 2215 -97 2227
rect -131 2159 -97 2177
rect -131 2143 -97 2159
rect -131 2091 -97 2105
rect -131 2071 -97 2091
rect -131 2023 -97 2033
rect -131 1999 -97 2023
rect -131 1955 -97 1961
rect -131 1927 -97 1955
rect -131 1887 -97 1889
rect -131 1855 -97 1887
rect -131 1785 -97 1817
rect -131 1783 -97 1785
rect -131 1717 -97 1745
rect -131 1711 -97 1717
rect -131 1649 -97 1673
rect -131 1639 -97 1649
rect -131 1581 -97 1601
rect -131 1567 -97 1581
rect -131 1513 -97 1529
rect -131 1495 -97 1513
rect -131 1445 -97 1457
rect -131 1423 -97 1445
rect -131 1377 -97 1385
rect -131 1351 -97 1377
rect -131 1309 -97 1313
rect -131 1279 -97 1309
rect -131 1207 -97 1241
rect -131 1139 -97 1169
rect -131 1135 -97 1139
rect -131 1071 -97 1097
rect -131 1063 -97 1071
rect -131 1003 -97 1025
rect -131 991 -97 1003
rect -131 935 -97 953
rect -131 919 -97 935
rect -131 867 -97 881
rect -131 847 -97 867
rect -131 799 -97 809
rect -131 775 -97 799
rect -131 731 -97 737
rect -131 703 -97 731
rect -131 663 -97 665
rect -131 631 -97 663
rect -131 561 -97 593
rect -131 559 -97 561
rect -131 493 -97 521
rect -131 487 -97 493
rect -131 425 -97 449
rect -131 415 -97 425
rect -131 357 -97 377
rect -131 343 -97 357
rect -131 289 -97 305
rect -131 271 -97 289
rect -131 221 -97 233
rect -131 199 -97 221
rect -131 153 -97 161
rect -131 127 -97 153
rect -131 85 -97 89
rect -131 55 -97 85
rect -131 -17 -97 17
rect -131 -85 -97 -55
rect -131 -89 -97 -85
rect -131 -153 -97 -127
rect -131 -161 -97 -153
rect -131 -221 -97 -199
rect -131 -233 -97 -221
rect -131 -289 -97 -271
rect -131 -305 -97 -289
rect -131 -357 -97 -343
rect -131 -377 -97 -357
rect -131 -425 -97 -415
rect -131 -449 -97 -425
rect -131 -493 -97 -487
rect -131 -521 -97 -493
rect -131 -561 -97 -559
rect -131 -593 -97 -561
rect -131 -663 -97 -631
rect -131 -665 -97 -663
rect -131 -731 -97 -703
rect -131 -737 -97 -731
rect -131 -799 -97 -775
rect -131 -809 -97 -799
rect -131 -867 -97 -847
rect -131 -881 -97 -867
rect -131 -935 -97 -919
rect -131 -953 -97 -935
rect -131 -1003 -97 -991
rect -131 -1025 -97 -1003
rect -131 -1071 -97 -1063
rect -131 -1097 -97 -1071
rect -131 -1139 -97 -1135
rect -131 -1169 -97 -1139
rect -131 -1241 -97 -1207
rect -131 -1309 -97 -1279
rect -131 -1313 -97 -1309
rect -131 -1377 -97 -1351
rect -131 -1385 -97 -1377
rect -131 -1445 -97 -1423
rect -131 -1457 -97 -1445
rect -131 -1513 -97 -1495
rect -131 -1529 -97 -1513
rect -131 -1581 -97 -1567
rect -131 -1601 -97 -1581
rect -131 -1649 -97 -1639
rect -131 -1673 -97 -1649
rect -131 -1717 -97 -1711
rect -131 -1745 -97 -1717
rect -131 -1785 -97 -1783
rect -131 -1817 -97 -1785
rect -131 -1887 -97 -1855
rect -131 -1889 -97 -1887
rect -131 -1955 -97 -1927
rect -131 -1961 -97 -1955
rect -131 -2023 -97 -1999
rect -131 -2033 -97 -2023
rect -131 -2091 -97 -2071
rect -131 -2105 -97 -2091
rect -131 -2159 -97 -2143
rect -131 -2177 -97 -2159
rect -131 -2227 -97 -2215
rect -131 -2249 -97 -2227
rect -131 -2295 -97 -2287
rect -131 -2321 -97 -2295
rect -131 -2363 -97 -2359
rect -131 -2393 -97 -2363
rect -131 -2465 -97 -2431
rect -17 2431 17 2465
rect -17 2363 17 2393
rect -17 2359 17 2363
rect -17 2295 17 2321
rect -17 2287 17 2295
rect -17 2227 17 2249
rect -17 2215 17 2227
rect -17 2159 17 2177
rect -17 2143 17 2159
rect -17 2091 17 2105
rect -17 2071 17 2091
rect -17 2023 17 2033
rect -17 1999 17 2023
rect -17 1955 17 1961
rect -17 1927 17 1955
rect -17 1887 17 1889
rect -17 1855 17 1887
rect -17 1785 17 1817
rect -17 1783 17 1785
rect -17 1717 17 1745
rect -17 1711 17 1717
rect -17 1649 17 1673
rect -17 1639 17 1649
rect -17 1581 17 1601
rect -17 1567 17 1581
rect -17 1513 17 1529
rect -17 1495 17 1513
rect -17 1445 17 1457
rect -17 1423 17 1445
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect -17 -1445 17 -1423
rect -17 -1457 17 -1445
rect -17 -1513 17 -1495
rect -17 -1529 17 -1513
rect -17 -1581 17 -1567
rect -17 -1601 17 -1581
rect -17 -1649 17 -1639
rect -17 -1673 17 -1649
rect -17 -1717 17 -1711
rect -17 -1745 17 -1717
rect -17 -1785 17 -1783
rect -17 -1817 17 -1785
rect -17 -1887 17 -1855
rect -17 -1889 17 -1887
rect -17 -1955 17 -1927
rect -17 -1961 17 -1955
rect -17 -2023 17 -1999
rect -17 -2033 17 -2023
rect -17 -2091 17 -2071
rect -17 -2105 17 -2091
rect -17 -2159 17 -2143
rect -17 -2177 17 -2159
rect -17 -2227 17 -2215
rect -17 -2249 17 -2227
rect -17 -2295 17 -2287
rect -17 -2321 17 -2295
rect -17 -2363 17 -2359
rect -17 -2393 17 -2363
rect -17 -2465 17 -2431
rect 97 2431 131 2465
rect 97 2363 131 2393
rect 97 2359 131 2363
rect 97 2295 131 2321
rect 97 2287 131 2295
rect 97 2227 131 2249
rect 97 2215 131 2227
rect 97 2159 131 2177
rect 97 2143 131 2159
rect 97 2091 131 2105
rect 97 2071 131 2091
rect 97 2023 131 2033
rect 97 1999 131 2023
rect 97 1955 131 1961
rect 97 1927 131 1955
rect 97 1887 131 1889
rect 97 1855 131 1887
rect 97 1785 131 1817
rect 97 1783 131 1785
rect 97 1717 131 1745
rect 97 1711 131 1717
rect 97 1649 131 1673
rect 97 1639 131 1649
rect 97 1581 131 1601
rect 97 1567 131 1581
rect 97 1513 131 1529
rect 97 1495 131 1513
rect 97 1445 131 1457
rect 97 1423 131 1445
rect 97 1377 131 1385
rect 97 1351 131 1377
rect 97 1309 131 1313
rect 97 1279 131 1309
rect 97 1207 131 1241
rect 97 1139 131 1169
rect 97 1135 131 1139
rect 97 1071 131 1097
rect 97 1063 131 1071
rect 97 1003 131 1025
rect 97 991 131 1003
rect 97 935 131 953
rect 97 919 131 935
rect 97 867 131 881
rect 97 847 131 867
rect 97 799 131 809
rect 97 775 131 799
rect 97 731 131 737
rect 97 703 131 731
rect 97 663 131 665
rect 97 631 131 663
rect 97 561 131 593
rect 97 559 131 561
rect 97 493 131 521
rect 97 487 131 493
rect 97 425 131 449
rect 97 415 131 425
rect 97 357 131 377
rect 97 343 131 357
rect 97 289 131 305
rect 97 271 131 289
rect 97 221 131 233
rect 97 199 131 221
rect 97 153 131 161
rect 97 127 131 153
rect 97 85 131 89
rect 97 55 131 85
rect 97 -17 131 17
rect 97 -85 131 -55
rect 97 -89 131 -85
rect 97 -153 131 -127
rect 97 -161 131 -153
rect 97 -221 131 -199
rect 97 -233 131 -221
rect 97 -289 131 -271
rect 97 -305 131 -289
rect 97 -357 131 -343
rect 97 -377 131 -357
rect 97 -425 131 -415
rect 97 -449 131 -425
rect 97 -493 131 -487
rect 97 -521 131 -493
rect 97 -561 131 -559
rect 97 -593 131 -561
rect 97 -663 131 -631
rect 97 -665 131 -663
rect 97 -731 131 -703
rect 97 -737 131 -731
rect 97 -799 131 -775
rect 97 -809 131 -799
rect 97 -867 131 -847
rect 97 -881 131 -867
rect 97 -935 131 -919
rect 97 -953 131 -935
rect 97 -1003 131 -991
rect 97 -1025 131 -1003
rect 97 -1071 131 -1063
rect 97 -1097 131 -1071
rect 97 -1139 131 -1135
rect 97 -1169 131 -1139
rect 97 -1241 131 -1207
rect 97 -1309 131 -1279
rect 97 -1313 131 -1309
rect 97 -1377 131 -1351
rect 97 -1385 131 -1377
rect 97 -1445 131 -1423
rect 97 -1457 131 -1445
rect 97 -1513 131 -1495
rect 97 -1529 131 -1513
rect 97 -1581 131 -1567
rect 97 -1601 131 -1581
rect 97 -1649 131 -1639
rect 97 -1673 131 -1649
rect 97 -1717 131 -1711
rect 97 -1745 131 -1717
rect 97 -1785 131 -1783
rect 97 -1817 131 -1785
rect 97 -1887 131 -1855
rect 97 -1889 131 -1887
rect 97 -1955 131 -1927
rect 97 -1961 131 -1955
rect 97 -2023 131 -1999
rect 97 -2033 131 -2023
rect 97 -2091 131 -2071
rect 97 -2105 131 -2091
rect 97 -2159 131 -2143
rect 97 -2177 131 -2159
rect 97 -2227 131 -2215
rect 97 -2249 131 -2227
rect 97 -2295 131 -2287
rect 97 -2321 131 -2295
rect 97 -2363 131 -2359
rect 97 -2393 131 -2363
rect 97 -2465 131 -2431
rect 211 2431 245 2465
rect 211 2363 245 2393
rect 211 2359 245 2363
rect 211 2295 245 2321
rect 211 2287 245 2295
rect 211 2227 245 2249
rect 211 2215 245 2227
rect 211 2159 245 2177
rect 211 2143 245 2159
rect 211 2091 245 2105
rect 211 2071 245 2091
rect 211 2023 245 2033
rect 211 1999 245 2023
rect 211 1955 245 1961
rect 211 1927 245 1955
rect 211 1887 245 1889
rect 211 1855 245 1887
rect 211 1785 245 1817
rect 211 1783 245 1785
rect 211 1717 245 1745
rect 211 1711 245 1717
rect 211 1649 245 1673
rect 211 1639 245 1649
rect 211 1581 245 1601
rect 211 1567 245 1581
rect 211 1513 245 1529
rect 211 1495 245 1513
rect 211 1445 245 1457
rect 211 1423 245 1445
rect 211 1377 245 1385
rect 211 1351 245 1377
rect 211 1309 245 1313
rect 211 1279 245 1309
rect 211 1207 245 1241
rect 211 1139 245 1169
rect 211 1135 245 1139
rect 211 1071 245 1097
rect 211 1063 245 1071
rect 211 1003 245 1025
rect 211 991 245 1003
rect 211 935 245 953
rect 211 919 245 935
rect 211 867 245 881
rect 211 847 245 867
rect 211 799 245 809
rect 211 775 245 799
rect 211 731 245 737
rect 211 703 245 731
rect 211 663 245 665
rect 211 631 245 663
rect 211 561 245 593
rect 211 559 245 561
rect 211 493 245 521
rect 211 487 245 493
rect 211 425 245 449
rect 211 415 245 425
rect 211 357 245 377
rect 211 343 245 357
rect 211 289 245 305
rect 211 271 245 289
rect 211 221 245 233
rect 211 199 245 221
rect 211 153 245 161
rect 211 127 245 153
rect 211 85 245 89
rect 211 55 245 85
rect 211 -17 245 17
rect 211 -85 245 -55
rect 211 -89 245 -85
rect 211 -153 245 -127
rect 211 -161 245 -153
rect 211 -221 245 -199
rect 211 -233 245 -221
rect 211 -289 245 -271
rect 211 -305 245 -289
rect 211 -357 245 -343
rect 211 -377 245 -357
rect 211 -425 245 -415
rect 211 -449 245 -425
rect 211 -493 245 -487
rect 211 -521 245 -493
rect 211 -561 245 -559
rect 211 -593 245 -561
rect 211 -663 245 -631
rect 211 -665 245 -663
rect 211 -731 245 -703
rect 211 -737 245 -731
rect 211 -799 245 -775
rect 211 -809 245 -799
rect 211 -867 245 -847
rect 211 -881 245 -867
rect 211 -935 245 -919
rect 211 -953 245 -935
rect 211 -1003 245 -991
rect 211 -1025 245 -1003
rect 211 -1071 245 -1063
rect 211 -1097 245 -1071
rect 211 -1139 245 -1135
rect 211 -1169 245 -1139
rect 211 -1241 245 -1207
rect 211 -1309 245 -1279
rect 211 -1313 245 -1309
rect 211 -1377 245 -1351
rect 211 -1385 245 -1377
rect 211 -1445 245 -1423
rect 211 -1457 245 -1445
rect 211 -1513 245 -1495
rect 211 -1529 245 -1513
rect 211 -1581 245 -1567
rect 211 -1601 245 -1581
rect 211 -1649 245 -1639
rect 211 -1673 245 -1649
rect 211 -1717 245 -1711
rect 211 -1745 245 -1717
rect 211 -1785 245 -1783
rect 211 -1817 245 -1785
rect 211 -1887 245 -1855
rect 211 -1889 245 -1887
rect 211 -1955 245 -1927
rect 211 -1961 245 -1955
rect 211 -2023 245 -1999
rect 211 -2033 245 -2023
rect 211 -2091 245 -2071
rect 211 -2105 245 -2091
rect 211 -2159 245 -2143
rect 211 -2177 245 -2159
rect 211 -2227 245 -2215
rect 211 -2249 245 -2227
rect 211 -2295 245 -2287
rect 211 -2321 245 -2295
rect 211 -2363 245 -2359
rect 211 -2393 245 -2363
rect 211 -2465 245 -2431
<< metal1 >>
rect 142 2556 200 2562
rect 142 2522 154 2556
rect 188 2522 200 2556
rect 142 2516 200 2522
rect -251 2465 -205 2480
rect -251 2431 -245 2465
rect -211 2431 -205 2465
rect -251 2393 -205 2431
rect -251 2359 -245 2393
rect -211 2359 -205 2393
rect -251 2321 -205 2359
rect -251 2287 -245 2321
rect -211 2287 -205 2321
rect -251 2249 -205 2287
rect -251 2215 -245 2249
rect -211 2215 -205 2249
rect -251 2177 -205 2215
rect -251 2143 -245 2177
rect -211 2143 -205 2177
rect -251 2105 -205 2143
rect -251 2071 -245 2105
rect -211 2071 -205 2105
rect -251 2033 -205 2071
rect -251 1999 -245 2033
rect -211 1999 -205 2033
rect -251 1961 -205 1999
rect -251 1927 -245 1961
rect -211 1927 -205 1961
rect -251 1889 -205 1927
rect -251 1855 -245 1889
rect -211 1855 -205 1889
rect -251 1817 -205 1855
rect -251 1783 -245 1817
rect -211 1783 -205 1817
rect -251 1745 -205 1783
rect -251 1711 -245 1745
rect -211 1711 -205 1745
rect -251 1673 -205 1711
rect -251 1639 -245 1673
rect -211 1639 -205 1673
rect -251 1601 -205 1639
rect -251 1567 -245 1601
rect -211 1567 -205 1601
rect -251 1529 -205 1567
rect -251 1495 -245 1529
rect -211 1495 -205 1529
rect -251 1457 -205 1495
rect -251 1423 -245 1457
rect -211 1423 -205 1457
rect -251 1385 -205 1423
rect -251 1351 -245 1385
rect -211 1351 -205 1385
rect -251 1313 -205 1351
rect -251 1279 -245 1313
rect -211 1279 -205 1313
rect -251 1241 -205 1279
rect -251 1207 -245 1241
rect -211 1207 -205 1241
rect -251 1169 -205 1207
rect -251 1135 -245 1169
rect -211 1135 -205 1169
rect -251 1097 -205 1135
rect -251 1063 -245 1097
rect -211 1063 -205 1097
rect -251 1025 -205 1063
rect -251 991 -245 1025
rect -211 991 -205 1025
rect -251 953 -205 991
rect -251 919 -245 953
rect -211 919 -205 953
rect -251 881 -205 919
rect -251 847 -245 881
rect -211 847 -205 881
rect -251 809 -205 847
rect -251 775 -245 809
rect -211 775 -205 809
rect -251 737 -205 775
rect -251 703 -245 737
rect -211 703 -205 737
rect -251 665 -205 703
rect -251 631 -245 665
rect -211 631 -205 665
rect -251 593 -205 631
rect -251 559 -245 593
rect -211 559 -205 593
rect -251 521 -205 559
rect -251 487 -245 521
rect -211 487 -205 521
rect -251 449 -205 487
rect -251 415 -245 449
rect -211 415 -205 449
rect -251 377 -205 415
rect -251 343 -245 377
rect -211 343 -205 377
rect -251 305 -205 343
rect -251 271 -245 305
rect -211 271 -205 305
rect -251 233 -205 271
rect -251 199 -245 233
rect -211 199 -205 233
rect -251 161 -205 199
rect -251 127 -245 161
rect -211 127 -205 161
rect -251 89 -205 127
rect -251 55 -245 89
rect -211 55 -205 89
rect -251 17 -205 55
rect -251 -17 -245 17
rect -211 -17 -205 17
rect -251 -55 -205 -17
rect -251 -89 -245 -55
rect -211 -89 -205 -55
rect -251 -127 -205 -89
rect -251 -161 -245 -127
rect -211 -161 -205 -127
rect -251 -199 -205 -161
rect -251 -233 -245 -199
rect -211 -233 -205 -199
rect -251 -271 -205 -233
rect -251 -305 -245 -271
rect -211 -305 -205 -271
rect -251 -343 -205 -305
rect -251 -377 -245 -343
rect -211 -377 -205 -343
rect -251 -415 -205 -377
rect -251 -449 -245 -415
rect -211 -449 -205 -415
rect -251 -487 -205 -449
rect -251 -521 -245 -487
rect -211 -521 -205 -487
rect -251 -559 -205 -521
rect -251 -593 -245 -559
rect -211 -593 -205 -559
rect -251 -631 -205 -593
rect -251 -665 -245 -631
rect -211 -665 -205 -631
rect -251 -703 -205 -665
rect -251 -737 -245 -703
rect -211 -737 -205 -703
rect -251 -775 -205 -737
rect -251 -809 -245 -775
rect -211 -809 -205 -775
rect -251 -847 -205 -809
rect -251 -881 -245 -847
rect -211 -881 -205 -847
rect -251 -919 -205 -881
rect -251 -953 -245 -919
rect -211 -953 -205 -919
rect -251 -991 -205 -953
rect -251 -1025 -245 -991
rect -211 -1025 -205 -991
rect -251 -1063 -205 -1025
rect -251 -1097 -245 -1063
rect -211 -1097 -205 -1063
rect -251 -1135 -205 -1097
rect -251 -1169 -245 -1135
rect -211 -1169 -205 -1135
rect -251 -1207 -205 -1169
rect -251 -1241 -245 -1207
rect -211 -1241 -205 -1207
rect -251 -1279 -205 -1241
rect -251 -1313 -245 -1279
rect -211 -1313 -205 -1279
rect -251 -1351 -205 -1313
rect -251 -1385 -245 -1351
rect -211 -1385 -205 -1351
rect -251 -1423 -205 -1385
rect -251 -1457 -245 -1423
rect -211 -1457 -205 -1423
rect -251 -1495 -205 -1457
rect -251 -1529 -245 -1495
rect -211 -1529 -205 -1495
rect -251 -1567 -205 -1529
rect -251 -1601 -245 -1567
rect -211 -1601 -205 -1567
rect -251 -1639 -205 -1601
rect -251 -1673 -245 -1639
rect -211 -1673 -205 -1639
rect -251 -1711 -205 -1673
rect -251 -1745 -245 -1711
rect -211 -1745 -205 -1711
rect -251 -1783 -205 -1745
rect -251 -1817 -245 -1783
rect -211 -1817 -205 -1783
rect -251 -1855 -205 -1817
rect -251 -1889 -245 -1855
rect -211 -1889 -205 -1855
rect -251 -1927 -205 -1889
rect -251 -1961 -245 -1927
rect -211 -1961 -205 -1927
rect -251 -1999 -205 -1961
rect -251 -2033 -245 -1999
rect -211 -2033 -205 -1999
rect -251 -2071 -205 -2033
rect -251 -2105 -245 -2071
rect -211 -2105 -205 -2071
rect -251 -2143 -205 -2105
rect -251 -2177 -245 -2143
rect -211 -2177 -205 -2143
rect -251 -2215 -205 -2177
rect -251 -2249 -245 -2215
rect -211 -2249 -205 -2215
rect -251 -2287 -205 -2249
rect -251 -2321 -245 -2287
rect -211 -2321 -205 -2287
rect -251 -2359 -205 -2321
rect -251 -2393 -245 -2359
rect -211 -2393 -205 -2359
rect -251 -2431 -205 -2393
rect -251 -2465 -245 -2431
rect -211 -2465 -205 -2431
rect -251 -2480 -205 -2465
rect -137 2465 -91 2480
rect -137 2431 -131 2465
rect -97 2431 -91 2465
rect -137 2393 -91 2431
rect -137 2359 -131 2393
rect -97 2359 -91 2393
rect -137 2321 -91 2359
rect -137 2287 -131 2321
rect -97 2287 -91 2321
rect -137 2249 -91 2287
rect -137 2215 -131 2249
rect -97 2215 -91 2249
rect -137 2177 -91 2215
rect -137 2143 -131 2177
rect -97 2143 -91 2177
rect -137 2105 -91 2143
rect -137 2071 -131 2105
rect -97 2071 -91 2105
rect -137 2033 -91 2071
rect -137 1999 -131 2033
rect -97 1999 -91 2033
rect -137 1961 -91 1999
rect -137 1927 -131 1961
rect -97 1927 -91 1961
rect -137 1889 -91 1927
rect -137 1855 -131 1889
rect -97 1855 -91 1889
rect -137 1817 -91 1855
rect -137 1783 -131 1817
rect -97 1783 -91 1817
rect -137 1745 -91 1783
rect -137 1711 -131 1745
rect -97 1711 -91 1745
rect -137 1673 -91 1711
rect -137 1639 -131 1673
rect -97 1639 -91 1673
rect -137 1601 -91 1639
rect -137 1567 -131 1601
rect -97 1567 -91 1601
rect -137 1529 -91 1567
rect -137 1495 -131 1529
rect -97 1495 -91 1529
rect -137 1457 -91 1495
rect -137 1423 -131 1457
rect -97 1423 -91 1457
rect -137 1385 -91 1423
rect -137 1351 -131 1385
rect -97 1351 -91 1385
rect -137 1313 -91 1351
rect -137 1279 -131 1313
rect -97 1279 -91 1313
rect -137 1241 -91 1279
rect -137 1207 -131 1241
rect -97 1207 -91 1241
rect -137 1169 -91 1207
rect -137 1135 -131 1169
rect -97 1135 -91 1169
rect -137 1097 -91 1135
rect -137 1063 -131 1097
rect -97 1063 -91 1097
rect -137 1025 -91 1063
rect -137 991 -131 1025
rect -97 991 -91 1025
rect -137 953 -91 991
rect -137 919 -131 953
rect -97 919 -91 953
rect -137 881 -91 919
rect -137 847 -131 881
rect -97 847 -91 881
rect -137 809 -91 847
rect -137 775 -131 809
rect -97 775 -91 809
rect -137 737 -91 775
rect -137 703 -131 737
rect -97 703 -91 737
rect -137 665 -91 703
rect -137 631 -131 665
rect -97 631 -91 665
rect -137 593 -91 631
rect -137 559 -131 593
rect -97 559 -91 593
rect -137 521 -91 559
rect -137 487 -131 521
rect -97 487 -91 521
rect -137 449 -91 487
rect -137 415 -131 449
rect -97 415 -91 449
rect -137 377 -91 415
rect -137 343 -131 377
rect -97 343 -91 377
rect -137 305 -91 343
rect -137 271 -131 305
rect -97 271 -91 305
rect -137 233 -91 271
rect -137 199 -131 233
rect -97 199 -91 233
rect -137 161 -91 199
rect -137 127 -131 161
rect -97 127 -91 161
rect -137 89 -91 127
rect -137 55 -131 89
rect -97 55 -91 89
rect -137 17 -91 55
rect -137 -17 -131 17
rect -97 -17 -91 17
rect -137 -55 -91 -17
rect -137 -89 -131 -55
rect -97 -89 -91 -55
rect -137 -127 -91 -89
rect -137 -161 -131 -127
rect -97 -161 -91 -127
rect -137 -199 -91 -161
rect -137 -233 -131 -199
rect -97 -233 -91 -199
rect -137 -271 -91 -233
rect -137 -305 -131 -271
rect -97 -305 -91 -271
rect -137 -343 -91 -305
rect -137 -377 -131 -343
rect -97 -377 -91 -343
rect -137 -415 -91 -377
rect -137 -449 -131 -415
rect -97 -449 -91 -415
rect -137 -487 -91 -449
rect -137 -521 -131 -487
rect -97 -521 -91 -487
rect -137 -559 -91 -521
rect -137 -593 -131 -559
rect -97 -593 -91 -559
rect -137 -631 -91 -593
rect -137 -665 -131 -631
rect -97 -665 -91 -631
rect -137 -703 -91 -665
rect -137 -737 -131 -703
rect -97 -737 -91 -703
rect -137 -775 -91 -737
rect -137 -809 -131 -775
rect -97 -809 -91 -775
rect -137 -847 -91 -809
rect -137 -881 -131 -847
rect -97 -881 -91 -847
rect -137 -919 -91 -881
rect -137 -953 -131 -919
rect -97 -953 -91 -919
rect -137 -991 -91 -953
rect -137 -1025 -131 -991
rect -97 -1025 -91 -991
rect -137 -1063 -91 -1025
rect -137 -1097 -131 -1063
rect -97 -1097 -91 -1063
rect -137 -1135 -91 -1097
rect -137 -1169 -131 -1135
rect -97 -1169 -91 -1135
rect -137 -1207 -91 -1169
rect -137 -1241 -131 -1207
rect -97 -1241 -91 -1207
rect -137 -1279 -91 -1241
rect -137 -1313 -131 -1279
rect -97 -1313 -91 -1279
rect -137 -1351 -91 -1313
rect -137 -1385 -131 -1351
rect -97 -1385 -91 -1351
rect -137 -1423 -91 -1385
rect -137 -1457 -131 -1423
rect -97 -1457 -91 -1423
rect -137 -1495 -91 -1457
rect -137 -1529 -131 -1495
rect -97 -1529 -91 -1495
rect -137 -1567 -91 -1529
rect -137 -1601 -131 -1567
rect -97 -1601 -91 -1567
rect -137 -1639 -91 -1601
rect -137 -1673 -131 -1639
rect -97 -1673 -91 -1639
rect -137 -1711 -91 -1673
rect -137 -1745 -131 -1711
rect -97 -1745 -91 -1711
rect -137 -1783 -91 -1745
rect -137 -1817 -131 -1783
rect -97 -1817 -91 -1783
rect -137 -1855 -91 -1817
rect -137 -1889 -131 -1855
rect -97 -1889 -91 -1855
rect -137 -1927 -91 -1889
rect -137 -1961 -131 -1927
rect -97 -1961 -91 -1927
rect -137 -1999 -91 -1961
rect -137 -2033 -131 -1999
rect -97 -2033 -91 -1999
rect -137 -2071 -91 -2033
rect -137 -2105 -131 -2071
rect -97 -2105 -91 -2071
rect -137 -2143 -91 -2105
rect -137 -2177 -131 -2143
rect -97 -2177 -91 -2143
rect -137 -2215 -91 -2177
rect -137 -2249 -131 -2215
rect -97 -2249 -91 -2215
rect -137 -2287 -91 -2249
rect -137 -2321 -131 -2287
rect -97 -2321 -91 -2287
rect -137 -2359 -91 -2321
rect -137 -2393 -131 -2359
rect -97 -2393 -91 -2359
rect -137 -2431 -91 -2393
rect -137 -2465 -131 -2431
rect -97 -2465 -91 -2431
rect -137 -2480 -91 -2465
rect -23 2465 23 2480
rect -23 2431 -17 2465
rect 17 2431 23 2465
rect -23 2393 23 2431
rect -23 2359 -17 2393
rect 17 2359 23 2393
rect -23 2321 23 2359
rect -23 2287 -17 2321
rect 17 2287 23 2321
rect -23 2249 23 2287
rect -23 2215 -17 2249
rect 17 2215 23 2249
rect -23 2177 23 2215
rect -23 2143 -17 2177
rect 17 2143 23 2177
rect -23 2105 23 2143
rect -23 2071 -17 2105
rect 17 2071 23 2105
rect -23 2033 23 2071
rect -23 1999 -17 2033
rect 17 1999 23 2033
rect -23 1961 23 1999
rect -23 1927 -17 1961
rect 17 1927 23 1961
rect -23 1889 23 1927
rect -23 1855 -17 1889
rect 17 1855 23 1889
rect -23 1817 23 1855
rect -23 1783 -17 1817
rect 17 1783 23 1817
rect -23 1745 23 1783
rect -23 1711 -17 1745
rect 17 1711 23 1745
rect -23 1673 23 1711
rect -23 1639 -17 1673
rect 17 1639 23 1673
rect -23 1601 23 1639
rect -23 1567 -17 1601
rect 17 1567 23 1601
rect -23 1529 23 1567
rect -23 1495 -17 1529
rect 17 1495 23 1529
rect -23 1457 23 1495
rect -23 1423 -17 1457
rect 17 1423 23 1457
rect -23 1385 23 1423
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1423 23 -1385
rect -23 -1457 -17 -1423
rect 17 -1457 23 -1423
rect -23 -1495 23 -1457
rect -23 -1529 -17 -1495
rect 17 -1529 23 -1495
rect -23 -1567 23 -1529
rect -23 -1601 -17 -1567
rect 17 -1601 23 -1567
rect -23 -1639 23 -1601
rect -23 -1673 -17 -1639
rect 17 -1673 23 -1639
rect -23 -1711 23 -1673
rect -23 -1745 -17 -1711
rect 17 -1745 23 -1711
rect -23 -1783 23 -1745
rect -23 -1817 -17 -1783
rect 17 -1817 23 -1783
rect -23 -1855 23 -1817
rect -23 -1889 -17 -1855
rect 17 -1889 23 -1855
rect -23 -1927 23 -1889
rect -23 -1961 -17 -1927
rect 17 -1961 23 -1927
rect -23 -1999 23 -1961
rect -23 -2033 -17 -1999
rect 17 -2033 23 -1999
rect -23 -2071 23 -2033
rect -23 -2105 -17 -2071
rect 17 -2105 23 -2071
rect -23 -2143 23 -2105
rect -23 -2177 -17 -2143
rect 17 -2177 23 -2143
rect -23 -2215 23 -2177
rect -23 -2249 -17 -2215
rect 17 -2249 23 -2215
rect -23 -2287 23 -2249
rect -23 -2321 -17 -2287
rect 17 -2321 23 -2287
rect -23 -2359 23 -2321
rect -23 -2393 -17 -2359
rect 17 -2393 23 -2359
rect -23 -2431 23 -2393
rect -23 -2465 -17 -2431
rect 17 -2465 23 -2431
rect -23 -2480 23 -2465
rect 91 2465 137 2480
rect 91 2431 97 2465
rect 131 2431 137 2465
rect 91 2393 137 2431
rect 91 2359 97 2393
rect 131 2359 137 2393
rect 91 2321 137 2359
rect 91 2287 97 2321
rect 131 2287 137 2321
rect 91 2249 137 2287
rect 91 2215 97 2249
rect 131 2215 137 2249
rect 91 2177 137 2215
rect 91 2143 97 2177
rect 131 2143 137 2177
rect 91 2105 137 2143
rect 91 2071 97 2105
rect 131 2071 137 2105
rect 91 2033 137 2071
rect 91 1999 97 2033
rect 131 1999 137 2033
rect 91 1961 137 1999
rect 91 1927 97 1961
rect 131 1927 137 1961
rect 91 1889 137 1927
rect 91 1855 97 1889
rect 131 1855 137 1889
rect 91 1817 137 1855
rect 91 1783 97 1817
rect 131 1783 137 1817
rect 91 1745 137 1783
rect 91 1711 97 1745
rect 131 1711 137 1745
rect 91 1673 137 1711
rect 91 1639 97 1673
rect 131 1639 137 1673
rect 91 1601 137 1639
rect 91 1567 97 1601
rect 131 1567 137 1601
rect 91 1529 137 1567
rect 91 1495 97 1529
rect 131 1495 137 1529
rect 91 1457 137 1495
rect 91 1423 97 1457
rect 131 1423 137 1457
rect 91 1385 137 1423
rect 91 1351 97 1385
rect 131 1351 137 1385
rect 91 1313 137 1351
rect 91 1279 97 1313
rect 131 1279 137 1313
rect 91 1241 137 1279
rect 91 1207 97 1241
rect 131 1207 137 1241
rect 91 1169 137 1207
rect 91 1135 97 1169
rect 131 1135 137 1169
rect 91 1097 137 1135
rect 91 1063 97 1097
rect 131 1063 137 1097
rect 91 1025 137 1063
rect 91 991 97 1025
rect 131 991 137 1025
rect 91 953 137 991
rect 91 919 97 953
rect 131 919 137 953
rect 91 881 137 919
rect 91 847 97 881
rect 131 847 137 881
rect 91 809 137 847
rect 91 775 97 809
rect 131 775 137 809
rect 91 737 137 775
rect 91 703 97 737
rect 131 703 137 737
rect 91 665 137 703
rect 91 631 97 665
rect 131 631 137 665
rect 91 593 137 631
rect 91 559 97 593
rect 131 559 137 593
rect 91 521 137 559
rect 91 487 97 521
rect 131 487 137 521
rect 91 449 137 487
rect 91 415 97 449
rect 131 415 137 449
rect 91 377 137 415
rect 91 343 97 377
rect 131 343 137 377
rect 91 305 137 343
rect 91 271 97 305
rect 131 271 137 305
rect 91 233 137 271
rect 91 199 97 233
rect 131 199 137 233
rect 91 161 137 199
rect 91 127 97 161
rect 131 127 137 161
rect 91 89 137 127
rect 91 55 97 89
rect 131 55 137 89
rect 91 17 137 55
rect 91 -17 97 17
rect 131 -17 137 17
rect 91 -55 137 -17
rect 91 -89 97 -55
rect 131 -89 137 -55
rect 91 -127 137 -89
rect 91 -161 97 -127
rect 131 -161 137 -127
rect 91 -199 137 -161
rect 91 -233 97 -199
rect 131 -233 137 -199
rect 91 -271 137 -233
rect 91 -305 97 -271
rect 131 -305 137 -271
rect 91 -343 137 -305
rect 91 -377 97 -343
rect 131 -377 137 -343
rect 91 -415 137 -377
rect 91 -449 97 -415
rect 131 -449 137 -415
rect 91 -487 137 -449
rect 91 -521 97 -487
rect 131 -521 137 -487
rect 91 -559 137 -521
rect 91 -593 97 -559
rect 131 -593 137 -559
rect 91 -631 137 -593
rect 91 -665 97 -631
rect 131 -665 137 -631
rect 91 -703 137 -665
rect 91 -737 97 -703
rect 131 -737 137 -703
rect 91 -775 137 -737
rect 91 -809 97 -775
rect 131 -809 137 -775
rect 91 -847 137 -809
rect 91 -881 97 -847
rect 131 -881 137 -847
rect 91 -919 137 -881
rect 91 -953 97 -919
rect 131 -953 137 -919
rect 91 -991 137 -953
rect 91 -1025 97 -991
rect 131 -1025 137 -991
rect 91 -1063 137 -1025
rect 91 -1097 97 -1063
rect 131 -1097 137 -1063
rect 91 -1135 137 -1097
rect 91 -1169 97 -1135
rect 131 -1169 137 -1135
rect 91 -1207 137 -1169
rect 91 -1241 97 -1207
rect 131 -1241 137 -1207
rect 91 -1279 137 -1241
rect 91 -1313 97 -1279
rect 131 -1313 137 -1279
rect 91 -1351 137 -1313
rect 91 -1385 97 -1351
rect 131 -1385 137 -1351
rect 91 -1423 137 -1385
rect 91 -1457 97 -1423
rect 131 -1457 137 -1423
rect 91 -1495 137 -1457
rect 91 -1529 97 -1495
rect 131 -1529 137 -1495
rect 91 -1567 137 -1529
rect 91 -1601 97 -1567
rect 131 -1601 137 -1567
rect 91 -1639 137 -1601
rect 91 -1673 97 -1639
rect 131 -1673 137 -1639
rect 91 -1711 137 -1673
rect 91 -1745 97 -1711
rect 131 -1745 137 -1711
rect 91 -1783 137 -1745
rect 91 -1817 97 -1783
rect 131 -1817 137 -1783
rect 91 -1855 137 -1817
rect 91 -1889 97 -1855
rect 131 -1889 137 -1855
rect 91 -1927 137 -1889
rect 91 -1961 97 -1927
rect 131 -1961 137 -1927
rect 91 -1999 137 -1961
rect 91 -2033 97 -1999
rect 131 -2033 137 -1999
rect 91 -2071 137 -2033
rect 91 -2105 97 -2071
rect 131 -2105 137 -2071
rect 91 -2143 137 -2105
rect 91 -2177 97 -2143
rect 131 -2177 137 -2143
rect 91 -2215 137 -2177
rect 91 -2249 97 -2215
rect 131 -2249 137 -2215
rect 91 -2287 137 -2249
rect 91 -2321 97 -2287
rect 131 -2321 137 -2287
rect 91 -2359 137 -2321
rect 91 -2393 97 -2359
rect 131 -2393 137 -2359
rect 91 -2431 137 -2393
rect 91 -2465 97 -2431
rect 131 -2465 137 -2431
rect 91 -2480 137 -2465
rect 205 2465 251 2480
rect 205 2431 211 2465
rect 245 2431 251 2465
rect 205 2393 251 2431
rect 205 2359 211 2393
rect 245 2359 251 2393
rect 205 2321 251 2359
rect 205 2287 211 2321
rect 245 2287 251 2321
rect 205 2249 251 2287
rect 205 2215 211 2249
rect 245 2215 251 2249
rect 205 2177 251 2215
rect 205 2143 211 2177
rect 245 2143 251 2177
rect 205 2105 251 2143
rect 205 2071 211 2105
rect 245 2071 251 2105
rect 205 2033 251 2071
rect 205 1999 211 2033
rect 245 1999 251 2033
rect 205 1961 251 1999
rect 205 1927 211 1961
rect 245 1927 251 1961
rect 205 1889 251 1927
rect 205 1855 211 1889
rect 245 1855 251 1889
rect 205 1817 251 1855
rect 205 1783 211 1817
rect 245 1783 251 1817
rect 205 1745 251 1783
rect 205 1711 211 1745
rect 245 1711 251 1745
rect 205 1673 251 1711
rect 205 1639 211 1673
rect 245 1639 251 1673
rect 205 1601 251 1639
rect 205 1567 211 1601
rect 245 1567 251 1601
rect 205 1529 251 1567
rect 205 1495 211 1529
rect 245 1495 251 1529
rect 205 1457 251 1495
rect 205 1423 211 1457
rect 245 1423 251 1457
rect 205 1385 251 1423
rect 205 1351 211 1385
rect 245 1351 251 1385
rect 205 1313 251 1351
rect 205 1279 211 1313
rect 245 1279 251 1313
rect 205 1241 251 1279
rect 205 1207 211 1241
rect 245 1207 251 1241
rect 205 1169 251 1207
rect 205 1135 211 1169
rect 245 1135 251 1169
rect 205 1097 251 1135
rect 205 1063 211 1097
rect 245 1063 251 1097
rect 205 1025 251 1063
rect 205 991 211 1025
rect 245 991 251 1025
rect 205 953 251 991
rect 205 919 211 953
rect 245 919 251 953
rect 205 881 251 919
rect 205 847 211 881
rect 245 847 251 881
rect 205 809 251 847
rect 205 775 211 809
rect 245 775 251 809
rect 205 737 251 775
rect 205 703 211 737
rect 245 703 251 737
rect 205 665 251 703
rect 205 631 211 665
rect 245 631 251 665
rect 205 593 251 631
rect 205 559 211 593
rect 245 559 251 593
rect 205 521 251 559
rect 205 487 211 521
rect 245 487 251 521
rect 205 449 251 487
rect 205 415 211 449
rect 245 415 251 449
rect 205 377 251 415
rect 205 343 211 377
rect 245 343 251 377
rect 205 305 251 343
rect 205 271 211 305
rect 245 271 251 305
rect 205 233 251 271
rect 205 199 211 233
rect 245 199 251 233
rect 205 161 251 199
rect 205 127 211 161
rect 245 127 251 161
rect 205 89 251 127
rect 205 55 211 89
rect 245 55 251 89
rect 205 17 251 55
rect 205 -17 211 17
rect 245 -17 251 17
rect 205 -55 251 -17
rect 205 -89 211 -55
rect 245 -89 251 -55
rect 205 -127 251 -89
rect 205 -161 211 -127
rect 245 -161 251 -127
rect 205 -199 251 -161
rect 205 -233 211 -199
rect 245 -233 251 -199
rect 205 -271 251 -233
rect 205 -305 211 -271
rect 245 -305 251 -271
rect 205 -343 251 -305
rect 205 -377 211 -343
rect 245 -377 251 -343
rect 205 -415 251 -377
rect 205 -449 211 -415
rect 245 -449 251 -415
rect 205 -487 251 -449
rect 205 -521 211 -487
rect 245 -521 251 -487
rect 205 -559 251 -521
rect 205 -593 211 -559
rect 245 -593 251 -559
rect 205 -631 251 -593
rect 205 -665 211 -631
rect 245 -665 251 -631
rect 205 -703 251 -665
rect 205 -737 211 -703
rect 245 -737 251 -703
rect 205 -775 251 -737
rect 205 -809 211 -775
rect 245 -809 251 -775
rect 205 -847 251 -809
rect 205 -881 211 -847
rect 245 -881 251 -847
rect 205 -919 251 -881
rect 205 -953 211 -919
rect 245 -953 251 -919
rect 205 -991 251 -953
rect 205 -1025 211 -991
rect 245 -1025 251 -991
rect 205 -1063 251 -1025
rect 205 -1097 211 -1063
rect 245 -1097 251 -1063
rect 205 -1135 251 -1097
rect 205 -1169 211 -1135
rect 245 -1169 251 -1135
rect 205 -1207 251 -1169
rect 205 -1241 211 -1207
rect 245 -1241 251 -1207
rect 205 -1279 251 -1241
rect 205 -1313 211 -1279
rect 245 -1313 251 -1279
rect 205 -1351 251 -1313
rect 205 -1385 211 -1351
rect 245 -1385 251 -1351
rect 205 -1423 251 -1385
rect 205 -1457 211 -1423
rect 245 -1457 251 -1423
rect 205 -1495 251 -1457
rect 205 -1529 211 -1495
rect 245 -1529 251 -1495
rect 205 -1567 251 -1529
rect 205 -1601 211 -1567
rect 245 -1601 251 -1567
rect 205 -1639 251 -1601
rect 205 -1673 211 -1639
rect 245 -1673 251 -1639
rect 205 -1711 251 -1673
rect 205 -1745 211 -1711
rect 245 -1745 251 -1711
rect 205 -1783 251 -1745
rect 205 -1817 211 -1783
rect 245 -1817 251 -1783
rect 205 -1855 251 -1817
rect 205 -1889 211 -1855
rect 245 -1889 251 -1855
rect 205 -1927 251 -1889
rect 205 -1961 211 -1927
rect 245 -1961 251 -1927
rect 205 -1999 251 -1961
rect 205 -2033 211 -1999
rect 245 -2033 251 -1999
rect 205 -2071 251 -2033
rect 205 -2105 211 -2071
rect 245 -2105 251 -2071
rect 205 -2143 251 -2105
rect 205 -2177 211 -2143
rect 245 -2177 251 -2143
rect 205 -2215 251 -2177
rect 205 -2249 211 -2215
rect 245 -2249 251 -2215
rect 205 -2287 251 -2249
rect 205 -2321 211 -2287
rect 245 -2321 251 -2287
rect 205 -2359 251 -2321
rect 205 -2393 211 -2359
rect 245 -2393 251 -2359
rect 205 -2431 251 -2393
rect 205 -2465 211 -2431
rect 245 -2465 251 -2431
rect 205 -2480 251 -2465
<< end >>
