magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nwell >>
rect -381 -2600 381 2600
<< pmos >>
rect -287 -2500 -187 2500
rect -129 -2500 -29 2500
rect 29 -2500 129 2500
rect 187 -2500 287 2500
<< pdiff >>
rect -345 2488 -287 2500
rect -345 -2488 -333 2488
rect -299 -2488 -287 2488
rect -345 -2500 -287 -2488
rect -187 2488 -129 2500
rect -187 -2488 -175 2488
rect -141 -2488 -129 2488
rect -187 -2500 -129 -2488
rect -29 2488 29 2500
rect -29 -2488 -17 2488
rect 17 -2488 29 2488
rect -29 -2500 29 -2488
rect 129 2488 187 2500
rect 129 -2488 141 2488
rect 175 -2488 187 2488
rect 129 -2500 187 -2488
rect 287 2488 345 2500
rect 287 -2488 299 2488
rect 333 -2488 345 2488
rect 287 -2500 345 -2488
<< pdiffc >>
rect -333 -2488 -299 2488
rect -175 -2488 -141 2488
rect -17 -2488 17 2488
rect 141 -2488 175 2488
rect 299 -2488 333 2488
<< poly >>
rect -287 2581 -187 2597
rect -287 2547 -271 2581
rect -203 2547 -187 2581
rect -287 2500 -187 2547
rect -129 2581 -29 2597
rect -129 2547 -113 2581
rect -45 2547 -29 2581
rect -129 2500 -29 2547
rect 29 2581 129 2597
rect 29 2547 45 2581
rect 113 2547 129 2581
rect 29 2500 129 2547
rect 187 2581 287 2597
rect 187 2547 203 2581
rect 271 2547 287 2581
rect 187 2500 287 2547
rect -287 -2547 -187 -2500
rect -287 -2581 -271 -2547
rect -203 -2581 -187 -2547
rect -287 -2597 -187 -2581
rect -129 -2547 -29 -2500
rect -129 -2581 -113 -2547
rect -45 -2581 -29 -2547
rect -129 -2597 -29 -2581
rect 29 -2547 129 -2500
rect 29 -2581 45 -2547
rect 113 -2581 129 -2547
rect 29 -2597 129 -2581
rect 187 -2547 287 -2500
rect 187 -2581 203 -2547
rect 271 -2581 287 -2547
rect 187 -2597 287 -2581
<< polycont >>
rect -271 2547 -203 2581
rect -113 2547 -45 2581
rect 45 2547 113 2581
rect 203 2547 271 2581
rect -271 -2581 -203 -2547
rect -113 -2581 -45 -2547
rect 45 -2581 113 -2547
rect 203 -2581 271 -2547
<< locali >>
rect -287 2547 -271 2581
rect -203 2547 -187 2581
rect -129 2547 -113 2581
rect -45 2547 -29 2581
rect 29 2547 45 2581
rect 113 2547 129 2581
rect 187 2547 203 2581
rect 271 2547 287 2581
rect -333 2488 -299 2504
rect -333 -2504 -299 -2488
rect -175 2488 -141 2504
rect -175 -2504 -141 -2488
rect -17 2488 17 2504
rect -17 -2504 17 -2488
rect 141 2488 175 2504
rect 141 -2504 175 -2488
rect 299 2488 333 2504
rect 299 -2504 333 -2488
rect -287 -2581 -271 -2547
rect -203 -2581 -187 -2547
rect -129 -2581 -113 -2547
rect -45 -2581 -29 -2547
rect 29 -2581 45 -2547
rect 113 -2581 129 -2547
rect 187 -2581 203 -2547
rect 271 -2581 287 -2547
<< viali >>
rect -271 2547 -203 2581
rect -113 2547 -45 2581
rect 45 2547 113 2581
rect 203 2547 271 2581
rect -333 -2488 -299 2488
rect -175 -2488 -141 2488
rect -17 -2488 17 2488
rect 141 -2488 175 2488
rect 299 -2488 333 2488
rect -271 -2581 -203 -2547
rect -113 -2581 -45 -2547
rect 45 -2581 113 -2547
rect 203 -2581 271 -2547
<< metal1 >>
rect -283 2581 -191 2587
rect -283 2547 -271 2581
rect -203 2547 -191 2581
rect -283 2541 -191 2547
rect -125 2581 -33 2587
rect -125 2547 -113 2581
rect -45 2547 -33 2581
rect -125 2541 -33 2547
rect 33 2581 125 2587
rect 33 2547 45 2581
rect 113 2547 125 2581
rect 33 2541 125 2547
rect 191 2581 283 2587
rect 191 2547 203 2581
rect 271 2547 283 2581
rect 191 2541 283 2547
rect -339 2488 -293 2500
rect -339 -2488 -333 2488
rect -299 -2488 -293 2488
rect -339 -2500 -293 -2488
rect -181 2488 -135 2500
rect -181 -2488 -175 2488
rect -141 -2488 -135 2488
rect -181 -2500 -135 -2488
rect -23 2488 23 2500
rect -23 -2488 -17 2488
rect 17 -2488 23 2488
rect -23 -2500 23 -2488
rect 135 2488 181 2500
rect 135 -2488 141 2488
rect 175 -2488 181 2488
rect 135 -2500 181 -2488
rect 293 2488 339 2500
rect 293 -2488 299 2488
rect 333 -2488 339 2488
rect 293 -2500 339 -2488
rect -283 -2547 -191 -2541
rect -283 -2581 -271 -2547
rect -203 -2581 -191 -2547
rect -283 -2587 -191 -2581
rect -125 -2547 -33 -2541
rect -125 -2581 -113 -2547
rect -45 -2581 -33 -2547
rect -125 -2587 -33 -2581
rect 33 -2547 125 -2541
rect 33 -2581 45 -2547
rect 113 -2581 125 -2547
rect 33 -2587 125 -2581
rect 191 -2547 283 -2541
rect 191 -2581 203 -2547
rect 271 -2581 283 -2547
rect 191 -2587 283 -2581
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 25 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
