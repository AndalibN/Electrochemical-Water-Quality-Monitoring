magic
tech sky130A
magscale 1 2
timestamp 1666200384
<< error_p >>
rect -213 18 213 236
<< nwell >>
rect -213 18 213 518
rect -213 -518 213 -18
<< pmos >>
rect -119 118 -29 418
rect 29 118 119 418
rect -119 -418 -29 -118
rect 29 -418 119 -118
<< pdiff >>
rect -177 406 -119 418
rect -177 130 -165 406
rect -131 130 -119 406
rect -177 118 -119 130
rect -29 406 29 418
rect -29 130 -17 406
rect 17 130 29 406
rect -29 118 29 130
rect 119 406 177 418
rect 119 130 131 406
rect 165 130 177 406
rect 119 118 177 130
rect -177 -130 -119 -118
rect -177 -406 -165 -130
rect -131 -406 -119 -130
rect -177 -418 -119 -406
rect -29 -130 29 -118
rect -29 -406 -17 -130
rect 17 -406 29 -130
rect -29 -418 29 -406
rect 119 -130 177 -118
rect 119 -406 131 -130
rect 165 -406 177 -130
rect 119 -418 177 -406
<< pdiffc >>
rect -165 130 -131 406
rect -17 130 17 406
rect 131 130 165 406
rect -165 -406 -131 -130
rect -17 -406 17 -130
rect 131 -406 165 -130
<< poly >>
rect -119 499 -29 515
rect -119 465 -103 499
rect -45 465 -29 499
rect -119 418 -29 465
rect 29 499 119 515
rect 29 465 45 499
rect 103 465 119 499
rect 29 418 119 465
rect -119 71 -29 118
rect -119 37 -103 71
rect -45 37 -29 71
rect -119 21 -29 37
rect 29 71 119 118
rect 29 37 45 71
rect 103 37 119 71
rect 29 21 119 37
rect -119 -37 -29 -21
rect -119 -71 -103 -37
rect -45 -71 -29 -37
rect -119 -118 -29 -71
rect 29 -37 119 -21
rect 29 -71 45 -37
rect 103 -71 119 -37
rect 29 -118 119 -71
rect -119 -465 -29 -418
rect -119 -499 -103 -465
rect -45 -499 -29 -465
rect -119 -515 -29 -499
rect 29 -465 119 -418
rect 29 -499 45 -465
rect 103 -499 119 -465
rect 29 -515 119 -499
<< polycont >>
rect -103 465 -45 499
rect 45 465 103 499
rect -103 37 -45 71
rect 45 37 103 71
rect -103 -71 -45 -37
rect 45 -71 103 -37
rect -103 -499 -45 -465
rect 45 -499 103 -465
<< locali >>
rect -119 465 -103 499
rect -45 465 -29 499
rect 29 465 45 499
rect 103 465 119 499
rect -165 406 -131 422
rect -165 114 -131 130
rect -17 406 17 422
rect -17 114 17 130
rect 131 406 165 422
rect 131 114 165 130
rect -119 37 -103 71
rect -45 37 -29 71
rect 29 37 45 71
rect 103 37 119 71
rect -119 -71 -103 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 103 -71 119 -37
rect -165 -130 -131 -114
rect -165 -422 -131 -406
rect -17 -130 17 -114
rect -17 -422 17 -406
rect 131 -130 165 -114
rect 131 -422 165 -406
rect -119 -499 -103 -465
rect -45 -499 -29 -465
rect 29 -499 45 -465
rect 103 -499 119 -465
<< viali >>
rect -103 465 -45 499
rect 45 465 103 499
rect -165 130 -131 406
rect -17 130 17 406
rect 131 130 165 406
rect -103 37 -45 71
rect 45 37 103 71
rect -103 -71 -45 -37
rect 45 -71 103 -37
rect -165 -406 -131 -130
rect -17 -406 17 -130
rect 131 -406 165 -130
rect -103 -499 -45 -465
rect 45 -499 103 -465
<< metal1 >>
rect -115 499 -33 505
rect -115 465 -103 499
rect -45 465 -33 499
rect -115 459 -33 465
rect 33 499 115 505
rect 33 465 45 499
rect 103 465 115 499
rect 33 459 115 465
rect -171 406 -125 418
rect -171 130 -165 406
rect -131 130 -125 406
rect -171 118 -125 130
rect -23 406 23 418
rect -23 130 -17 406
rect 17 130 23 406
rect -23 118 23 130
rect 125 406 171 418
rect 125 130 131 406
rect 165 130 171 406
rect 125 118 171 130
rect -115 71 -33 77
rect -115 37 -103 71
rect -45 37 -33 71
rect -115 31 -33 37
rect 33 71 115 77
rect 33 37 45 71
rect 103 37 115 71
rect 33 31 115 37
rect -115 -37 -33 -31
rect -115 -71 -103 -37
rect -45 -71 -33 -37
rect -115 -77 -33 -71
rect 33 -37 115 -31
rect 33 -71 45 -37
rect 103 -71 115 -37
rect 33 -77 115 -71
rect -171 -130 -125 -118
rect -171 -406 -165 -130
rect -131 -406 -125 -130
rect -171 -418 -125 -406
rect -23 -130 23 -118
rect -23 -406 -17 -130
rect 17 -406 23 -130
rect -23 -418 23 -406
rect 125 -130 171 -118
rect 125 -406 131 -130
rect 165 -406 171 -130
rect 125 -418 171 -406
rect -115 -465 -33 -459
rect -115 -499 -103 -465
rect -45 -499 -33 -465
rect -115 -505 -33 -499
rect 33 -465 115 -459
rect 33 -499 45 -465
rect 103 -499 115 -465
rect 33 -505 115 -499
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.45 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
