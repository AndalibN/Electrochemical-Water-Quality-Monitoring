magic
tech sky130A
magscale 1 2
timestamp 1666625676
<< xpolycontact >>
rect -15776 5200 -15706 5632
rect -15776 -5632 -15706 -5200
rect -15458 5200 -15388 5632
rect -15458 -5632 -15388 -5200
rect -15140 5200 -15070 5632
rect -15140 -5632 -15070 -5200
rect -14822 5200 -14752 5632
rect -14822 -5632 -14752 -5200
rect -14504 5200 -14434 5632
rect -14504 -5632 -14434 -5200
rect -14186 5200 -14116 5632
rect -14186 -5632 -14116 -5200
rect -13868 5200 -13798 5632
rect -13868 -5632 -13798 -5200
rect -13550 5200 -13480 5632
rect -13550 -5632 -13480 -5200
rect -13232 5200 -13162 5632
rect -13232 -5632 -13162 -5200
rect -12914 5200 -12844 5632
rect -12914 -5632 -12844 -5200
rect -12596 5200 -12526 5632
rect -12596 -5632 -12526 -5200
rect -12278 5200 -12208 5632
rect -12278 -5632 -12208 -5200
rect -11960 5200 -11890 5632
rect -11960 -5632 -11890 -5200
rect -11642 5200 -11572 5632
rect -11642 -5632 -11572 -5200
rect -11324 5200 -11254 5632
rect -11324 -5632 -11254 -5200
rect -11006 5200 -10936 5632
rect -11006 -5632 -10936 -5200
rect -10688 5200 -10618 5632
rect -10688 -5632 -10618 -5200
rect -10370 5200 -10300 5632
rect -10370 -5632 -10300 -5200
rect -10052 5200 -9982 5632
rect -10052 -5632 -9982 -5200
rect -9734 5200 -9664 5632
rect -9734 -5632 -9664 -5200
rect -9416 5200 -9346 5632
rect -9416 -5632 -9346 -5200
rect -9098 5200 -9028 5632
rect -9098 -5632 -9028 -5200
rect -8780 5200 -8710 5632
rect -8780 -5632 -8710 -5200
rect -8462 5200 -8392 5632
rect -8462 -5632 -8392 -5200
rect -8144 5200 -8074 5632
rect -8144 -5632 -8074 -5200
rect -7826 5200 -7756 5632
rect -7826 -5632 -7756 -5200
rect -7508 5200 -7438 5632
rect -7508 -5632 -7438 -5200
rect -7190 5200 -7120 5632
rect -7190 -5632 -7120 -5200
rect -6872 5200 -6802 5632
rect -6872 -5632 -6802 -5200
rect -6554 5200 -6484 5632
rect -6554 -5632 -6484 -5200
rect -6236 5200 -6166 5632
rect -6236 -5632 -6166 -5200
rect -5918 5200 -5848 5632
rect -5918 -5632 -5848 -5200
rect -5600 5200 -5530 5632
rect -5600 -5632 -5530 -5200
rect -5282 5200 -5212 5632
rect -5282 -5632 -5212 -5200
rect -4964 5200 -4894 5632
rect -4964 -5632 -4894 -5200
rect -4646 5200 -4576 5632
rect -4646 -5632 -4576 -5200
rect -4328 5200 -4258 5632
rect -4328 -5632 -4258 -5200
rect -4010 5200 -3940 5632
rect -4010 -5632 -3940 -5200
rect -3692 5200 -3622 5632
rect -3692 -5632 -3622 -5200
rect -3374 5200 -3304 5632
rect -3374 -5632 -3304 -5200
rect -3056 5200 -2986 5632
rect -3056 -5632 -2986 -5200
rect -2738 5200 -2668 5632
rect -2738 -5632 -2668 -5200
rect -2420 5200 -2350 5632
rect -2420 -5632 -2350 -5200
rect -2102 5200 -2032 5632
rect -2102 -5632 -2032 -5200
rect -1784 5200 -1714 5632
rect -1784 -5632 -1714 -5200
rect -1466 5200 -1396 5632
rect -1466 -5632 -1396 -5200
rect -1148 5200 -1078 5632
rect -1148 -5632 -1078 -5200
rect -830 5200 -760 5632
rect -830 -5632 -760 -5200
rect -512 5200 -442 5632
rect -512 -5632 -442 -5200
rect -194 5200 -124 5632
rect -194 -5632 -124 -5200
rect 124 5200 194 5632
rect 124 -5632 194 -5200
rect 442 5200 512 5632
rect 442 -5632 512 -5200
rect 760 5200 830 5632
rect 760 -5632 830 -5200
rect 1078 5200 1148 5632
rect 1078 -5632 1148 -5200
rect 1396 5200 1466 5632
rect 1396 -5632 1466 -5200
rect 1714 5200 1784 5632
rect 1714 -5632 1784 -5200
rect 2032 5200 2102 5632
rect 2032 -5632 2102 -5200
rect 2350 5200 2420 5632
rect 2350 -5632 2420 -5200
rect 2668 5200 2738 5632
rect 2668 -5632 2738 -5200
rect 2986 5200 3056 5632
rect 2986 -5632 3056 -5200
rect 3304 5200 3374 5632
rect 3304 -5632 3374 -5200
rect 3622 5200 3692 5632
rect 3622 -5632 3692 -5200
rect 3940 5200 4010 5632
rect 3940 -5632 4010 -5200
rect 4258 5200 4328 5632
rect 4258 -5632 4328 -5200
rect 4576 5200 4646 5632
rect 4576 -5632 4646 -5200
rect 4894 5200 4964 5632
rect 4894 -5632 4964 -5200
rect 5212 5200 5282 5632
rect 5212 -5632 5282 -5200
rect 5530 5200 5600 5632
rect 5530 -5632 5600 -5200
rect 5848 5200 5918 5632
rect 5848 -5632 5918 -5200
rect 6166 5200 6236 5632
rect 6166 -5632 6236 -5200
rect 6484 5200 6554 5632
rect 6484 -5632 6554 -5200
rect 6802 5200 6872 5632
rect 6802 -5632 6872 -5200
rect 7120 5200 7190 5632
rect 7120 -5632 7190 -5200
rect 7438 5200 7508 5632
rect 7438 -5632 7508 -5200
rect 7756 5200 7826 5632
rect 7756 -5632 7826 -5200
rect 8074 5200 8144 5632
rect 8074 -5632 8144 -5200
rect 8392 5200 8462 5632
rect 8392 -5632 8462 -5200
rect 8710 5200 8780 5632
rect 8710 -5632 8780 -5200
rect 9028 5200 9098 5632
rect 9028 -5632 9098 -5200
rect 9346 5200 9416 5632
rect 9346 -5632 9416 -5200
rect 9664 5200 9734 5632
rect 9664 -5632 9734 -5200
rect 9982 5200 10052 5632
rect 9982 -5632 10052 -5200
rect 10300 5200 10370 5632
rect 10300 -5632 10370 -5200
rect 10618 5200 10688 5632
rect 10618 -5632 10688 -5200
rect 10936 5200 11006 5632
rect 10936 -5632 11006 -5200
rect 11254 5200 11324 5632
rect 11254 -5632 11324 -5200
rect 11572 5200 11642 5632
rect 11572 -5632 11642 -5200
rect 11890 5200 11960 5632
rect 11890 -5632 11960 -5200
rect 12208 5200 12278 5632
rect 12208 -5632 12278 -5200
rect 12526 5200 12596 5632
rect 12526 -5632 12596 -5200
rect 12844 5200 12914 5632
rect 12844 -5632 12914 -5200
rect 13162 5200 13232 5632
rect 13162 -5632 13232 -5200
rect 13480 5200 13550 5632
rect 13480 -5632 13550 -5200
rect 13798 5200 13868 5632
rect 13798 -5632 13868 -5200
rect 14116 5200 14186 5632
rect 14116 -5632 14186 -5200
rect 14434 5200 14504 5632
rect 14434 -5632 14504 -5200
rect 14752 5200 14822 5632
rect 14752 -5632 14822 -5200
rect 15070 5200 15140 5632
rect 15070 -5632 15140 -5200
rect 15388 5200 15458 5632
rect 15388 -5632 15458 -5200
rect 15706 5200 15776 5632
rect 15706 -5632 15776 -5200
<< xpolyres >>
rect -15776 -5200 -15706 5200
rect -15458 -5200 -15388 5200
rect -15140 -5200 -15070 5200
rect -14822 -5200 -14752 5200
rect -14504 -5200 -14434 5200
rect -14186 -5200 -14116 5200
rect -13868 -5200 -13798 5200
rect -13550 -5200 -13480 5200
rect -13232 -5200 -13162 5200
rect -12914 -5200 -12844 5200
rect -12596 -5200 -12526 5200
rect -12278 -5200 -12208 5200
rect -11960 -5200 -11890 5200
rect -11642 -5200 -11572 5200
rect -11324 -5200 -11254 5200
rect -11006 -5200 -10936 5200
rect -10688 -5200 -10618 5200
rect -10370 -5200 -10300 5200
rect -10052 -5200 -9982 5200
rect -9734 -5200 -9664 5200
rect -9416 -5200 -9346 5200
rect -9098 -5200 -9028 5200
rect -8780 -5200 -8710 5200
rect -8462 -5200 -8392 5200
rect -8144 -5200 -8074 5200
rect -7826 -5200 -7756 5200
rect -7508 -5200 -7438 5200
rect -7190 -5200 -7120 5200
rect -6872 -5200 -6802 5200
rect -6554 -5200 -6484 5200
rect -6236 -5200 -6166 5200
rect -5918 -5200 -5848 5200
rect -5600 -5200 -5530 5200
rect -5282 -5200 -5212 5200
rect -4964 -5200 -4894 5200
rect -4646 -5200 -4576 5200
rect -4328 -5200 -4258 5200
rect -4010 -5200 -3940 5200
rect -3692 -5200 -3622 5200
rect -3374 -5200 -3304 5200
rect -3056 -5200 -2986 5200
rect -2738 -5200 -2668 5200
rect -2420 -5200 -2350 5200
rect -2102 -5200 -2032 5200
rect -1784 -5200 -1714 5200
rect -1466 -5200 -1396 5200
rect -1148 -5200 -1078 5200
rect -830 -5200 -760 5200
rect -512 -5200 -442 5200
rect -194 -5200 -124 5200
rect 124 -5200 194 5200
rect 442 -5200 512 5200
rect 760 -5200 830 5200
rect 1078 -5200 1148 5200
rect 1396 -5200 1466 5200
rect 1714 -5200 1784 5200
rect 2032 -5200 2102 5200
rect 2350 -5200 2420 5200
rect 2668 -5200 2738 5200
rect 2986 -5200 3056 5200
rect 3304 -5200 3374 5200
rect 3622 -5200 3692 5200
rect 3940 -5200 4010 5200
rect 4258 -5200 4328 5200
rect 4576 -5200 4646 5200
rect 4894 -5200 4964 5200
rect 5212 -5200 5282 5200
rect 5530 -5200 5600 5200
rect 5848 -5200 5918 5200
rect 6166 -5200 6236 5200
rect 6484 -5200 6554 5200
rect 6802 -5200 6872 5200
rect 7120 -5200 7190 5200
rect 7438 -5200 7508 5200
rect 7756 -5200 7826 5200
rect 8074 -5200 8144 5200
rect 8392 -5200 8462 5200
rect 8710 -5200 8780 5200
rect 9028 -5200 9098 5200
rect 9346 -5200 9416 5200
rect 9664 -5200 9734 5200
rect 9982 -5200 10052 5200
rect 10300 -5200 10370 5200
rect 10618 -5200 10688 5200
rect 10936 -5200 11006 5200
rect 11254 -5200 11324 5200
rect 11572 -5200 11642 5200
rect 11890 -5200 11960 5200
rect 12208 -5200 12278 5200
rect 12526 -5200 12596 5200
rect 12844 -5200 12914 5200
rect 13162 -5200 13232 5200
rect 13480 -5200 13550 5200
rect 13798 -5200 13868 5200
rect 14116 -5200 14186 5200
rect 14434 -5200 14504 5200
rect 14752 -5200 14822 5200
rect 15070 -5200 15140 5200
rect 15388 -5200 15458 5200
rect 15706 -5200 15776 5200
<< viali >>
rect -15760 5217 -15722 5614
rect -15442 5217 -15404 5614
rect -15124 5217 -15086 5614
rect -14806 5217 -14768 5614
rect -14488 5217 -14450 5614
rect -14170 5217 -14132 5614
rect -13852 5217 -13814 5614
rect -13534 5217 -13496 5614
rect -13216 5217 -13178 5614
rect -12898 5217 -12860 5614
rect -12580 5217 -12542 5614
rect -12262 5217 -12224 5614
rect -11944 5217 -11906 5614
rect -11626 5217 -11588 5614
rect -11308 5217 -11270 5614
rect -10990 5217 -10952 5614
rect -10672 5217 -10634 5614
rect -10354 5217 -10316 5614
rect -10036 5217 -9998 5614
rect -9718 5217 -9680 5614
rect -9400 5217 -9362 5614
rect -9082 5217 -9044 5614
rect -8764 5217 -8726 5614
rect -8446 5217 -8408 5614
rect -8128 5217 -8090 5614
rect -7810 5217 -7772 5614
rect -7492 5217 -7454 5614
rect -7174 5217 -7136 5614
rect -6856 5217 -6818 5614
rect -6538 5217 -6500 5614
rect -6220 5217 -6182 5614
rect -5902 5217 -5864 5614
rect -5584 5217 -5546 5614
rect -5266 5217 -5228 5614
rect -4948 5217 -4910 5614
rect -4630 5217 -4592 5614
rect -4312 5217 -4274 5614
rect -3994 5217 -3956 5614
rect -3676 5217 -3638 5614
rect -3358 5217 -3320 5614
rect -3040 5217 -3002 5614
rect -2722 5217 -2684 5614
rect -2404 5217 -2366 5614
rect -2086 5217 -2048 5614
rect -1768 5217 -1730 5614
rect -1450 5217 -1412 5614
rect -1132 5217 -1094 5614
rect -814 5217 -776 5614
rect -496 5217 -458 5614
rect -178 5217 -140 5614
rect 140 5217 178 5614
rect 458 5217 496 5614
rect 776 5217 814 5614
rect 1094 5217 1132 5614
rect 1412 5217 1450 5614
rect 1730 5217 1768 5614
rect 2048 5217 2086 5614
rect 2366 5217 2404 5614
rect 2684 5217 2722 5614
rect 3002 5217 3040 5614
rect 3320 5217 3358 5614
rect 3638 5217 3676 5614
rect 3956 5217 3994 5614
rect 4274 5217 4312 5614
rect 4592 5217 4630 5614
rect 4910 5217 4948 5614
rect 5228 5217 5266 5614
rect 5546 5217 5584 5614
rect 5864 5217 5902 5614
rect 6182 5217 6220 5614
rect 6500 5217 6538 5614
rect 6818 5217 6856 5614
rect 7136 5217 7174 5614
rect 7454 5217 7492 5614
rect 7772 5217 7810 5614
rect 8090 5217 8128 5614
rect 8408 5217 8446 5614
rect 8726 5217 8764 5614
rect 9044 5217 9082 5614
rect 9362 5217 9400 5614
rect 9680 5217 9718 5614
rect 9998 5217 10036 5614
rect 10316 5217 10354 5614
rect 10634 5217 10672 5614
rect 10952 5217 10990 5614
rect 11270 5217 11308 5614
rect 11588 5217 11626 5614
rect 11906 5217 11944 5614
rect 12224 5217 12262 5614
rect 12542 5217 12580 5614
rect 12860 5217 12898 5614
rect 13178 5217 13216 5614
rect 13496 5217 13534 5614
rect 13814 5217 13852 5614
rect 14132 5217 14170 5614
rect 14450 5217 14488 5614
rect 14768 5217 14806 5614
rect 15086 5217 15124 5614
rect 15404 5217 15442 5614
rect 15722 5217 15760 5614
rect -15760 -5614 -15722 -5217
rect -15442 -5614 -15404 -5217
rect -15124 -5614 -15086 -5217
rect -14806 -5614 -14768 -5217
rect -14488 -5614 -14450 -5217
rect -14170 -5614 -14132 -5217
rect -13852 -5614 -13814 -5217
rect -13534 -5614 -13496 -5217
rect -13216 -5614 -13178 -5217
rect -12898 -5614 -12860 -5217
rect -12580 -5614 -12542 -5217
rect -12262 -5614 -12224 -5217
rect -11944 -5614 -11906 -5217
rect -11626 -5614 -11588 -5217
rect -11308 -5614 -11270 -5217
rect -10990 -5614 -10952 -5217
rect -10672 -5614 -10634 -5217
rect -10354 -5614 -10316 -5217
rect -10036 -5614 -9998 -5217
rect -9718 -5614 -9680 -5217
rect -9400 -5614 -9362 -5217
rect -9082 -5614 -9044 -5217
rect -8764 -5614 -8726 -5217
rect -8446 -5614 -8408 -5217
rect -8128 -5614 -8090 -5217
rect -7810 -5614 -7772 -5217
rect -7492 -5614 -7454 -5217
rect -7174 -5614 -7136 -5217
rect -6856 -5614 -6818 -5217
rect -6538 -5614 -6500 -5217
rect -6220 -5614 -6182 -5217
rect -5902 -5614 -5864 -5217
rect -5584 -5614 -5546 -5217
rect -5266 -5614 -5228 -5217
rect -4948 -5614 -4910 -5217
rect -4630 -5614 -4592 -5217
rect -4312 -5614 -4274 -5217
rect -3994 -5614 -3956 -5217
rect -3676 -5614 -3638 -5217
rect -3358 -5614 -3320 -5217
rect -3040 -5614 -3002 -5217
rect -2722 -5614 -2684 -5217
rect -2404 -5614 -2366 -5217
rect -2086 -5614 -2048 -5217
rect -1768 -5614 -1730 -5217
rect -1450 -5614 -1412 -5217
rect -1132 -5614 -1094 -5217
rect -814 -5614 -776 -5217
rect -496 -5614 -458 -5217
rect -178 -5614 -140 -5217
rect 140 -5614 178 -5217
rect 458 -5614 496 -5217
rect 776 -5614 814 -5217
rect 1094 -5614 1132 -5217
rect 1412 -5614 1450 -5217
rect 1730 -5614 1768 -5217
rect 2048 -5614 2086 -5217
rect 2366 -5614 2404 -5217
rect 2684 -5614 2722 -5217
rect 3002 -5614 3040 -5217
rect 3320 -5614 3358 -5217
rect 3638 -5614 3676 -5217
rect 3956 -5614 3994 -5217
rect 4274 -5614 4312 -5217
rect 4592 -5614 4630 -5217
rect 4910 -5614 4948 -5217
rect 5228 -5614 5266 -5217
rect 5546 -5614 5584 -5217
rect 5864 -5614 5902 -5217
rect 6182 -5614 6220 -5217
rect 6500 -5614 6538 -5217
rect 6818 -5614 6856 -5217
rect 7136 -5614 7174 -5217
rect 7454 -5614 7492 -5217
rect 7772 -5614 7810 -5217
rect 8090 -5614 8128 -5217
rect 8408 -5614 8446 -5217
rect 8726 -5614 8764 -5217
rect 9044 -5614 9082 -5217
rect 9362 -5614 9400 -5217
rect 9680 -5614 9718 -5217
rect 9998 -5614 10036 -5217
rect 10316 -5614 10354 -5217
rect 10634 -5614 10672 -5217
rect 10952 -5614 10990 -5217
rect 11270 -5614 11308 -5217
rect 11588 -5614 11626 -5217
rect 11906 -5614 11944 -5217
rect 12224 -5614 12262 -5217
rect 12542 -5614 12580 -5217
rect 12860 -5614 12898 -5217
rect 13178 -5614 13216 -5217
rect 13496 -5614 13534 -5217
rect 13814 -5614 13852 -5217
rect 14132 -5614 14170 -5217
rect 14450 -5614 14488 -5217
rect 14768 -5614 14806 -5217
rect 15086 -5614 15124 -5217
rect 15404 -5614 15442 -5217
rect 15722 -5614 15760 -5217
<< metal1 >>
rect -15766 5614 -15716 5626
rect -15766 5217 -15760 5614
rect -15722 5217 -15716 5614
rect -15766 5205 -15716 5217
rect -15448 5614 -15398 5626
rect -15448 5217 -15442 5614
rect -15404 5217 -15398 5614
rect -15448 5205 -15398 5217
rect -15130 5614 -15080 5626
rect -15130 5217 -15124 5614
rect -15086 5217 -15080 5614
rect -15130 5205 -15080 5217
rect -14812 5614 -14762 5626
rect -14812 5217 -14806 5614
rect -14768 5217 -14762 5614
rect -14812 5205 -14762 5217
rect -14494 5614 -14444 5626
rect -14494 5217 -14488 5614
rect -14450 5217 -14444 5614
rect -14494 5205 -14444 5217
rect -14176 5614 -14126 5626
rect -14176 5217 -14170 5614
rect -14132 5217 -14126 5614
rect -14176 5205 -14126 5217
rect -13858 5614 -13808 5626
rect -13858 5217 -13852 5614
rect -13814 5217 -13808 5614
rect -13858 5205 -13808 5217
rect -13540 5614 -13490 5626
rect -13540 5217 -13534 5614
rect -13496 5217 -13490 5614
rect -13540 5205 -13490 5217
rect -13222 5614 -13172 5626
rect -13222 5217 -13216 5614
rect -13178 5217 -13172 5614
rect -13222 5205 -13172 5217
rect -12904 5614 -12854 5626
rect -12904 5217 -12898 5614
rect -12860 5217 -12854 5614
rect -12904 5205 -12854 5217
rect -12586 5614 -12536 5626
rect -12586 5217 -12580 5614
rect -12542 5217 -12536 5614
rect -12586 5205 -12536 5217
rect -12268 5614 -12218 5626
rect -12268 5217 -12262 5614
rect -12224 5217 -12218 5614
rect -12268 5205 -12218 5217
rect -11950 5614 -11900 5626
rect -11950 5217 -11944 5614
rect -11906 5217 -11900 5614
rect -11950 5205 -11900 5217
rect -11632 5614 -11582 5626
rect -11632 5217 -11626 5614
rect -11588 5217 -11582 5614
rect -11632 5205 -11582 5217
rect -11314 5614 -11264 5626
rect -11314 5217 -11308 5614
rect -11270 5217 -11264 5614
rect -11314 5205 -11264 5217
rect -10996 5614 -10946 5626
rect -10996 5217 -10990 5614
rect -10952 5217 -10946 5614
rect -10996 5205 -10946 5217
rect -10678 5614 -10628 5626
rect -10678 5217 -10672 5614
rect -10634 5217 -10628 5614
rect -10678 5205 -10628 5217
rect -10360 5614 -10310 5626
rect -10360 5217 -10354 5614
rect -10316 5217 -10310 5614
rect -10360 5205 -10310 5217
rect -10042 5614 -9992 5626
rect -10042 5217 -10036 5614
rect -9998 5217 -9992 5614
rect -10042 5205 -9992 5217
rect -9724 5614 -9674 5626
rect -9724 5217 -9718 5614
rect -9680 5217 -9674 5614
rect -9724 5205 -9674 5217
rect -9406 5614 -9356 5626
rect -9406 5217 -9400 5614
rect -9362 5217 -9356 5614
rect -9406 5205 -9356 5217
rect -9088 5614 -9038 5626
rect -9088 5217 -9082 5614
rect -9044 5217 -9038 5614
rect -9088 5205 -9038 5217
rect -8770 5614 -8720 5626
rect -8770 5217 -8764 5614
rect -8726 5217 -8720 5614
rect -8770 5205 -8720 5217
rect -8452 5614 -8402 5626
rect -8452 5217 -8446 5614
rect -8408 5217 -8402 5614
rect -8452 5205 -8402 5217
rect -8134 5614 -8084 5626
rect -8134 5217 -8128 5614
rect -8090 5217 -8084 5614
rect -8134 5205 -8084 5217
rect -7816 5614 -7766 5626
rect -7816 5217 -7810 5614
rect -7772 5217 -7766 5614
rect -7816 5205 -7766 5217
rect -7498 5614 -7448 5626
rect -7498 5217 -7492 5614
rect -7454 5217 -7448 5614
rect -7498 5205 -7448 5217
rect -7180 5614 -7130 5626
rect -7180 5217 -7174 5614
rect -7136 5217 -7130 5614
rect -7180 5205 -7130 5217
rect -6862 5614 -6812 5626
rect -6862 5217 -6856 5614
rect -6818 5217 -6812 5614
rect -6862 5205 -6812 5217
rect -6544 5614 -6494 5626
rect -6544 5217 -6538 5614
rect -6500 5217 -6494 5614
rect -6544 5205 -6494 5217
rect -6226 5614 -6176 5626
rect -6226 5217 -6220 5614
rect -6182 5217 -6176 5614
rect -6226 5205 -6176 5217
rect -5908 5614 -5858 5626
rect -5908 5217 -5902 5614
rect -5864 5217 -5858 5614
rect -5908 5205 -5858 5217
rect -5590 5614 -5540 5626
rect -5590 5217 -5584 5614
rect -5546 5217 -5540 5614
rect -5590 5205 -5540 5217
rect -5272 5614 -5222 5626
rect -5272 5217 -5266 5614
rect -5228 5217 -5222 5614
rect -5272 5205 -5222 5217
rect -4954 5614 -4904 5626
rect -4954 5217 -4948 5614
rect -4910 5217 -4904 5614
rect -4954 5205 -4904 5217
rect -4636 5614 -4586 5626
rect -4636 5217 -4630 5614
rect -4592 5217 -4586 5614
rect -4636 5205 -4586 5217
rect -4318 5614 -4268 5626
rect -4318 5217 -4312 5614
rect -4274 5217 -4268 5614
rect -4318 5205 -4268 5217
rect -4000 5614 -3950 5626
rect -4000 5217 -3994 5614
rect -3956 5217 -3950 5614
rect -4000 5205 -3950 5217
rect -3682 5614 -3632 5626
rect -3682 5217 -3676 5614
rect -3638 5217 -3632 5614
rect -3682 5205 -3632 5217
rect -3364 5614 -3314 5626
rect -3364 5217 -3358 5614
rect -3320 5217 -3314 5614
rect -3364 5205 -3314 5217
rect -3046 5614 -2996 5626
rect -3046 5217 -3040 5614
rect -3002 5217 -2996 5614
rect -3046 5205 -2996 5217
rect -2728 5614 -2678 5626
rect -2728 5217 -2722 5614
rect -2684 5217 -2678 5614
rect -2728 5205 -2678 5217
rect -2410 5614 -2360 5626
rect -2410 5217 -2404 5614
rect -2366 5217 -2360 5614
rect -2410 5205 -2360 5217
rect -2092 5614 -2042 5626
rect -2092 5217 -2086 5614
rect -2048 5217 -2042 5614
rect -2092 5205 -2042 5217
rect -1774 5614 -1724 5626
rect -1774 5217 -1768 5614
rect -1730 5217 -1724 5614
rect -1774 5205 -1724 5217
rect -1456 5614 -1406 5626
rect -1456 5217 -1450 5614
rect -1412 5217 -1406 5614
rect -1456 5205 -1406 5217
rect -1138 5614 -1088 5626
rect -1138 5217 -1132 5614
rect -1094 5217 -1088 5614
rect -1138 5205 -1088 5217
rect -820 5614 -770 5626
rect -820 5217 -814 5614
rect -776 5217 -770 5614
rect -820 5205 -770 5217
rect -502 5614 -452 5626
rect -502 5217 -496 5614
rect -458 5217 -452 5614
rect -502 5205 -452 5217
rect -184 5614 -134 5626
rect -184 5217 -178 5614
rect -140 5217 -134 5614
rect -184 5205 -134 5217
rect 134 5614 184 5626
rect 134 5217 140 5614
rect 178 5217 184 5614
rect 134 5205 184 5217
rect 452 5614 502 5626
rect 452 5217 458 5614
rect 496 5217 502 5614
rect 452 5205 502 5217
rect 770 5614 820 5626
rect 770 5217 776 5614
rect 814 5217 820 5614
rect 770 5205 820 5217
rect 1088 5614 1138 5626
rect 1088 5217 1094 5614
rect 1132 5217 1138 5614
rect 1088 5205 1138 5217
rect 1406 5614 1456 5626
rect 1406 5217 1412 5614
rect 1450 5217 1456 5614
rect 1406 5205 1456 5217
rect 1724 5614 1774 5626
rect 1724 5217 1730 5614
rect 1768 5217 1774 5614
rect 1724 5205 1774 5217
rect 2042 5614 2092 5626
rect 2042 5217 2048 5614
rect 2086 5217 2092 5614
rect 2042 5205 2092 5217
rect 2360 5614 2410 5626
rect 2360 5217 2366 5614
rect 2404 5217 2410 5614
rect 2360 5205 2410 5217
rect 2678 5614 2728 5626
rect 2678 5217 2684 5614
rect 2722 5217 2728 5614
rect 2678 5205 2728 5217
rect 2996 5614 3046 5626
rect 2996 5217 3002 5614
rect 3040 5217 3046 5614
rect 2996 5205 3046 5217
rect 3314 5614 3364 5626
rect 3314 5217 3320 5614
rect 3358 5217 3364 5614
rect 3314 5205 3364 5217
rect 3632 5614 3682 5626
rect 3632 5217 3638 5614
rect 3676 5217 3682 5614
rect 3632 5205 3682 5217
rect 3950 5614 4000 5626
rect 3950 5217 3956 5614
rect 3994 5217 4000 5614
rect 3950 5205 4000 5217
rect 4268 5614 4318 5626
rect 4268 5217 4274 5614
rect 4312 5217 4318 5614
rect 4268 5205 4318 5217
rect 4586 5614 4636 5626
rect 4586 5217 4592 5614
rect 4630 5217 4636 5614
rect 4586 5205 4636 5217
rect 4904 5614 4954 5626
rect 4904 5217 4910 5614
rect 4948 5217 4954 5614
rect 4904 5205 4954 5217
rect 5222 5614 5272 5626
rect 5222 5217 5228 5614
rect 5266 5217 5272 5614
rect 5222 5205 5272 5217
rect 5540 5614 5590 5626
rect 5540 5217 5546 5614
rect 5584 5217 5590 5614
rect 5540 5205 5590 5217
rect 5858 5614 5908 5626
rect 5858 5217 5864 5614
rect 5902 5217 5908 5614
rect 5858 5205 5908 5217
rect 6176 5614 6226 5626
rect 6176 5217 6182 5614
rect 6220 5217 6226 5614
rect 6176 5205 6226 5217
rect 6494 5614 6544 5626
rect 6494 5217 6500 5614
rect 6538 5217 6544 5614
rect 6494 5205 6544 5217
rect 6812 5614 6862 5626
rect 6812 5217 6818 5614
rect 6856 5217 6862 5614
rect 6812 5205 6862 5217
rect 7130 5614 7180 5626
rect 7130 5217 7136 5614
rect 7174 5217 7180 5614
rect 7130 5205 7180 5217
rect 7448 5614 7498 5626
rect 7448 5217 7454 5614
rect 7492 5217 7498 5614
rect 7448 5205 7498 5217
rect 7766 5614 7816 5626
rect 7766 5217 7772 5614
rect 7810 5217 7816 5614
rect 7766 5205 7816 5217
rect 8084 5614 8134 5626
rect 8084 5217 8090 5614
rect 8128 5217 8134 5614
rect 8084 5205 8134 5217
rect 8402 5614 8452 5626
rect 8402 5217 8408 5614
rect 8446 5217 8452 5614
rect 8402 5205 8452 5217
rect 8720 5614 8770 5626
rect 8720 5217 8726 5614
rect 8764 5217 8770 5614
rect 8720 5205 8770 5217
rect 9038 5614 9088 5626
rect 9038 5217 9044 5614
rect 9082 5217 9088 5614
rect 9038 5205 9088 5217
rect 9356 5614 9406 5626
rect 9356 5217 9362 5614
rect 9400 5217 9406 5614
rect 9356 5205 9406 5217
rect 9674 5614 9724 5626
rect 9674 5217 9680 5614
rect 9718 5217 9724 5614
rect 9674 5205 9724 5217
rect 9992 5614 10042 5626
rect 9992 5217 9998 5614
rect 10036 5217 10042 5614
rect 9992 5205 10042 5217
rect 10310 5614 10360 5626
rect 10310 5217 10316 5614
rect 10354 5217 10360 5614
rect 10310 5205 10360 5217
rect 10628 5614 10678 5626
rect 10628 5217 10634 5614
rect 10672 5217 10678 5614
rect 10628 5205 10678 5217
rect 10946 5614 10996 5626
rect 10946 5217 10952 5614
rect 10990 5217 10996 5614
rect 10946 5205 10996 5217
rect 11264 5614 11314 5626
rect 11264 5217 11270 5614
rect 11308 5217 11314 5614
rect 11264 5205 11314 5217
rect 11582 5614 11632 5626
rect 11582 5217 11588 5614
rect 11626 5217 11632 5614
rect 11582 5205 11632 5217
rect 11900 5614 11950 5626
rect 11900 5217 11906 5614
rect 11944 5217 11950 5614
rect 11900 5205 11950 5217
rect 12218 5614 12268 5626
rect 12218 5217 12224 5614
rect 12262 5217 12268 5614
rect 12218 5205 12268 5217
rect 12536 5614 12586 5626
rect 12536 5217 12542 5614
rect 12580 5217 12586 5614
rect 12536 5205 12586 5217
rect 12854 5614 12904 5626
rect 12854 5217 12860 5614
rect 12898 5217 12904 5614
rect 12854 5205 12904 5217
rect 13172 5614 13222 5626
rect 13172 5217 13178 5614
rect 13216 5217 13222 5614
rect 13172 5205 13222 5217
rect 13490 5614 13540 5626
rect 13490 5217 13496 5614
rect 13534 5217 13540 5614
rect 13490 5205 13540 5217
rect 13808 5614 13858 5626
rect 13808 5217 13814 5614
rect 13852 5217 13858 5614
rect 13808 5205 13858 5217
rect 14126 5614 14176 5626
rect 14126 5217 14132 5614
rect 14170 5217 14176 5614
rect 14126 5205 14176 5217
rect 14444 5614 14494 5626
rect 14444 5217 14450 5614
rect 14488 5217 14494 5614
rect 14444 5205 14494 5217
rect 14762 5614 14812 5626
rect 14762 5217 14768 5614
rect 14806 5217 14812 5614
rect 14762 5205 14812 5217
rect 15080 5614 15130 5626
rect 15080 5217 15086 5614
rect 15124 5217 15130 5614
rect 15080 5205 15130 5217
rect 15398 5614 15448 5626
rect 15398 5217 15404 5614
rect 15442 5217 15448 5614
rect 15398 5205 15448 5217
rect 15716 5614 15766 5626
rect 15716 5217 15722 5614
rect 15760 5217 15766 5614
rect 15716 5205 15766 5217
rect -15766 -5217 -15716 -5205
rect -15766 -5614 -15760 -5217
rect -15722 -5614 -15716 -5217
rect -15766 -5626 -15716 -5614
rect -15448 -5217 -15398 -5205
rect -15448 -5614 -15442 -5217
rect -15404 -5614 -15398 -5217
rect -15448 -5626 -15398 -5614
rect -15130 -5217 -15080 -5205
rect -15130 -5614 -15124 -5217
rect -15086 -5614 -15080 -5217
rect -15130 -5626 -15080 -5614
rect -14812 -5217 -14762 -5205
rect -14812 -5614 -14806 -5217
rect -14768 -5614 -14762 -5217
rect -14812 -5626 -14762 -5614
rect -14494 -5217 -14444 -5205
rect -14494 -5614 -14488 -5217
rect -14450 -5614 -14444 -5217
rect -14494 -5626 -14444 -5614
rect -14176 -5217 -14126 -5205
rect -14176 -5614 -14170 -5217
rect -14132 -5614 -14126 -5217
rect -14176 -5626 -14126 -5614
rect -13858 -5217 -13808 -5205
rect -13858 -5614 -13852 -5217
rect -13814 -5614 -13808 -5217
rect -13858 -5626 -13808 -5614
rect -13540 -5217 -13490 -5205
rect -13540 -5614 -13534 -5217
rect -13496 -5614 -13490 -5217
rect -13540 -5626 -13490 -5614
rect -13222 -5217 -13172 -5205
rect -13222 -5614 -13216 -5217
rect -13178 -5614 -13172 -5217
rect -13222 -5626 -13172 -5614
rect -12904 -5217 -12854 -5205
rect -12904 -5614 -12898 -5217
rect -12860 -5614 -12854 -5217
rect -12904 -5626 -12854 -5614
rect -12586 -5217 -12536 -5205
rect -12586 -5614 -12580 -5217
rect -12542 -5614 -12536 -5217
rect -12586 -5626 -12536 -5614
rect -12268 -5217 -12218 -5205
rect -12268 -5614 -12262 -5217
rect -12224 -5614 -12218 -5217
rect -12268 -5626 -12218 -5614
rect -11950 -5217 -11900 -5205
rect -11950 -5614 -11944 -5217
rect -11906 -5614 -11900 -5217
rect -11950 -5626 -11900 -5614
rect -11632 -5217 -11582 -5205
rect -11632 -5614 -11626 -5217
rect -11588 -5614 -11582 -5217
rect -11632 -5626 -11582 -5614
rect -11314 -5217 -11264 -5205
rect -11314 -5614 -11308 -5217
rect -11270 -5614 -11264 -5217
rect -11314 -5626 -11264 -5614
rect -10996 -5217 -10946 -5205
rect -10996 -5614 -10990 -5217
rect -10952 -5614 -10946 -5217
rect -10996 -5626 -10946 -5614
rect -10678 -5217 -10628 -5205
rect -10678 -5614 -10672 -5217
rect -10634 -5614 -10628 -5217
rect -10678 -5626 -10628 -5614
rect -10360 -5217 -10310 -5205
rect -10360 -5614 -10354 -5217
rect -10316 -5614 -10310 -5217
rect -10360 -5626 -10310 -5614
rect -10042 -5217 -9992 -5205
rect -10042 -5614 -10036 -5217
rect -9998 -5614 -9992 -5217
rect -10042 -5626 -9992 -5614
rect -9724 -5217 -9674 -5205
rect -9724 -5614 -9718 -5217
rect -9680 -5614 -9674 -5217
rect -9724 -5626 -9674 -5614
rect -9406 -5217 -9356 -5205
rect -9406 -5614 -9400 -5217
rect -9362 -5614 -9356 -5217
rect -9406 -5626 -9356 -5614
rect -9088 -5217 -9038 -5205
rect -9088 -5614 -9082 -5217
rect -9044 -5614 -9038 -5217
rect -9088 -5626 -9038 -5614
rect -8770 -5217 -8720 -5205
rect -8770 -5614 -8764 -5217
rect -8726 -5614 -8720 -5217
rect -8770 -5626 -8720 -5614
rect -8452 -5217 -8402 -5205
rect -8452 -5614 -8446 -5217
rect -8408 -5614 -8402 -5217
rect -8452 -5626 -8402 -5614
rect -8134 -5217 -8084 -5205
rect -8134 -5614 -8128 -5217
rect -8090 -5614 -8084 -5217
rect -8134 -5626 -8084 -5614
rect -7816 -5217 -7766 -5205
rect -7816 -5614 -7810 -5217
rect -7772 -5614 -7766 -5217
rect -7816 -5626 -7766 -5614
rect -7498 -5217 -7448 -5205
rect -7498 -5614 -7492 -5217
rect -7454 -5614 -7448 -5217
rect -7498 -5626 -7448 -5614
rect -7180 -5217 -7130 -5205
rect -7180 -5614 -7174 -5217
rect -7136 -5614 -7130 -5217
rect -7180 -5626 -7130 -5614
rect -6862 -5217 -6812 -5205
rect -6862 -5614 -6856 -5217
rect -6818 -5614 -6812 -5217
rect -6862 -5626 -6812 -5614
rect -6544 -5217 -6494 -5205
rect -6544 -5614 -6538 -5217
rect -6500 -5614 -6494 -5217
rect -6544 -5626 -6494 -5614
rect -6226 -5217 -6176 -5205
rect -6226 -5614 -6220 -5217
rect -6182 -5614 -6176 -5217
rect -6226 -5626 -6176 -5614
rect -5908 -5217 -5858 -5205
rect -5908 -5614 -5902 -5217
rect -5864 -5614 -5858 -5217
rect -5908 -5626 -5858 -5614
rect -5590 -5217 -5540 -5205
rect -5590 -5614 -5584 -5217
rect -5546 -5614 -5540 -5217
rect -5590 -5626 -5540 -5614
rect -5272 -5217 -5222 -5205
rect -5272 -5614 -5266 -5217
rect -5228 -5614 -5222 -5217
rect -5272 -5626 -5222 -5614
rect -4954 -5217 -4904 -5205
rect -4954 -5614 -4948 -5217
rect -4910 -5614 -4904 -5217
rect -4954 -5626 -4904 -5614
rect -4636 -5217 -4586 -5205
rect -4636 -5614 -4630 -5217
rect -4592 -5614 -4586 -5217
rect -4636 -5626 -4586 -5614
rect -4318 -5217 -4268 -5205
rect -4318 -5614 -4312 -5217
rect -4274 -5614 -4268 -5217
rect -4318 -5626 -4268 -5614
rect -4000 -5217 -3950 -5205
rect -4000 -5614 -3994 -5217
rect -3956 -5614 -3950 -5217
rect -4000 -5626 -3950 -5614
rect -3682 -5217 -3632 -5205
rect -3682 -5614 -3676 -5217
rect -3638 -5614 -3632 -5217
rect -3682 -5626 -3632 -5614
rect -3364 -5217 -3314 -5205
rect -3364 -5614 -3358 -5217
rect -3320 -5614 -3314 -5217
rect -3364 -5626 -3314 -5614
rect -3046 -5217 -2996 -5205
rect -3046 -5614 -3040 -5217
rect -3002 -5614 -2996 -5217
rect -3046 -5626 -2996 -5614
rect -2728 -5217 -2678 -5205
rect -2728 -5614 -2722 -5217
rect -2684 -5614 -2678 -5217
rect -2728 -5626 -2678 -5614
rect -2410 -5217 -2360 -5205
rect -2410 -5614 -2404 -5217
rect -2366 -5614 -2360 -5217
rect -2410 -5626 -2360 -5614
rect -2092 -5217 -2042 -5205
rect -2092 -5614 -2086 -5217
rect -2048 -5614 -2042 -5217
rect -2092 -5626 -2042 -5614
rect -1774 -5217 -1724 -5205
rect -1774 -5614 -1768 -5217
rect -1730 -5614 -1724 -5217
rect -1774 -5626 -1724 -5614
rect -1456 -5217 -1406 -5205
rect -1456 -5614 -1450 -5217
rect -1412 -5614 -1406 -5217
rect -1456 -5626 -1406 -5614
rect -1138 -5217 -1088 -5205
rect -1138 -5614 -1132 -5217
rect -1094 -5614 -1088 -5217
rect -1138 -5626 -1088 -5614
rect -820 -5217 -770 -5205
rect -820 -5614 -814 -5217
rect -776 -5614 -770 -5217
rect -820 -5626 -770 -5614
rect -502 -5217 -452 -5205
rect -502 -5614 -496 -5217
rect -458 -5614 -452 -5217
rect -502 -5626 -452 -5614
rect -184 -5217 -134 -5205
rect -184 -5614 -178 -5217
rect -140 -5614 -134 -5217
rect -184 -5626 -134 -5614
rect 134 -5217 184 -5205
rect 134 -5614 140 -5217
rect 178 -5614 184 -5217
rect 134 -5626 184 -5614
rect 452 -5217 502 -5205
rect 452 -5614 458 -5217
rect 496 -5614 502 -5217
rect 452 -5626 502 -5614
rect 770 -5217 820 -5205
rect 770 -5614 776 -5217
rect 814 -5614 820 -5217
rect 770 -5626 820 -5614
rect 1088 -5217 1138 -5205
rect 1088 -5614 1094 -5217
rect 1132 -5614 1138 -5217
rect 1088 -5626 1138 -5614
rect 1406 -5217 1456 -5205
rect 1406 -5614 1412 -5217
rect 1450 -5614 1456 -5217
rect 1406 -5626 1456 -5614
rect 1724 -5217 1774 -5205
rect 1724 -5614 1730 -5217
rect 1768 -5614 1774 -5217
rect 1724 -5626 1774 -5614
rect 2042 -5217 2092 -5205
rect 2042 -5614 2048 -5217
rect 2086 -5614 2092 -5217
rect 2042 -5626 2092 -5614
rect 2360 -5217 2410 -5205
rect 2360 -5614 2366 -5217
rect 2404 -5614 2410 -5217
rect 2360 -5626 2410 -5614
rect 2678 -5217 2728 -5205
rect 2678 -5614 2684 -5217
rect 2722 -5614 2728 -5217
rect 2678 -5626 2728 -5614
rect 2996 -5217 3046 -5205
rect 2996 -5614 3002 -5217
rect 3040 -5614 3046 -5217
rect 2996 -5626 3046 -5614
rect 3314 -5217 3364 -5205
rect 3314 -5614 3320 -5217
rect 3358 -5614 3364 -5217
rect 3314 -5626 3364 -5614
rect 3632 -5217 3682 -5205
rect 3632 -5614 3638 -5217
rect 3676 -5614 3682 -5217
rect 3632 -5626 3682 -5614
rect 3950 -5217 4000 -5205
rect 3950 -5614 3956 -5217
rect 3994 -5614 4000 -5217
rect 3950 -5626 4000 -5614
rect 4268 -5217 4318 -5205
rect 4268 -5614 4274 -5217
rect 4312 -5614 4318 -5217
rect 4268 -5626 4318 -5614
rect 4586 -5217 4636 -5205
rect 4586 -5614 4592 -5217
rect 4630 -5614 4636 -5217
rect 4586 -5626 4636 -5614
rect 4904 -5217 4954 -5205
rect 4904 -5614 4910 -5217
rect 4948 -5614 4954 -5217
rect 4904 -5626 4954 -5614
rect 5222 -5217 5272 -5205
rect 5222 -5614 5228 -5217
rect 5266 -5614 5272 -5217
rect 5222 -5626 5272 -5614
rect 5540 -5217 5590 -5205
rect 5540 -5614 5546 -5217
rect 5584 -5614 5590 -5217
rect 5540 -5626 5590 -5614
rect 5858 -5217 5908 -5205
rect 5858 -5614 5864 -5217
rect 5902 -5614 5908 -5217
rect 5858 -5626 5908 -5614
rect 6176 -5217 6226 -5205
rect 6176 -5614 6182 -5217
rect 6220 -5614 6226 -5217
rect 6176 -5626 6226 -5614
rect 6494 -5217 6544 -5205
rect 6494 -5614 6500 -5217
rect 6538 -5614 6544 -5217
rect 6494 -5626 6544 -5614
rect 6812 -5217 6862 -5205
rect 6812 -5614 6818 -5217
rect 6856 -5614 6862 -5217
rect 6812 -5626 6862 -5614
rect 7130 -5217 7180 -5205
rect 7130 -5614 7136 -5217
rect 7174 -5614 7180 -5217
rect 7130 -5626 7180 -5614
rect 7448 -5217 7498 -5205
rect 7448 -5614 7454 -5217
rect 7492 -5614 7498 -5217
rect 7448 -5626 7498 -5614
rect 7766 -5217 7816 -5205
rect 7766 -5614 7772 -5217
rect 7810 -5614 7816 -5217
rect 7766 -5626 7816 -5614
rect 8084 -5217 8134 -5205
rect 8084 -5614 8090 -5217
rect 8128 -5614 8134 -5217
rect 8084 -5626 8134 -5614
rect 8402 -5217 8452 -5205
rect 8402 -5614 8408 -5217
rect 8446 -5614 8452 -5217
rect 8402 -5626 8452 -5614
rect 8720 -5217 8770 -5205
rect 8720 -5614 8726 -5217
rect 8764 -5614 8770 -5217
rect 8720 -5626 8770 -5614
rect 9038 -5217 9088 -5205
rect 9038 -5614 9044 -5217
rect 9082 -5614 9088 -5217
rect 9038 -5626 9088 -5614
rect 9356 -5217 9406 -5205
rect 9356 -5614 9362 -5217
rect 9400 -5614 9406 -5217
rect 9356 -5626 9406 -5614
rect 9674 -5217 9724 -5205
rect 9674 -5614 9680 -5217
rect 9718 -5614 9724 -5217
rect 9674 -5626 9724 -5614
rect 9992 -5217 10042 -5205
rect 9992 -5614 9998 -5217
rect 10036 -5614 10042 -5217
rect 9992 -5626 10042 -5614
rect 10310 -5217 10360 -5205
rect 10310 -5614 10316 -5217
rect 10354 -5614 10360 -5217
rect 10310 -5626 10360 -5614
rect 10628 -5217 10678 -5205
rect 10628 -5614 10634 -5217
rect 10672 -5614 10678 -5217
rect 10628 -5626 10678 -5614
rect 10946 -5217 10996 -5205
rect 10946 -5614 10952 -5217
rect 10990 -5614 10996 -5217
rect 10946 -5626 10996 -5614
rect 11264 -5217 11314 -5205
rect 11264 -5614 11270 -5217
rect 11308 -5614 11314 -5217
rect 11264 -5626 11314 -5614
rect 11582 -5217 11632 -5205
rect 11582 -5614 11588 -5217
rect 11626 -5614 11632 -5217
rect 11582 -5626 11632 -5614
rect 11900 -5217 11950 -5205
rect 11900 -5614 11906 -5217
rect 11944 -5614 11950 -5217
rect 11900 -5626 11950 -5614
rect 12218 -5217 12268 -5205
rect 12218 -5614 12224 -5217
rect 12262 -5614 12268 -5217
rect 12218 -5626 12268 -5614
rect 12536 -5217 12586 -5205
rect 12536 -5614 12542 -5217
rect 12580 -5614 12586 -5217
rect 12536 -5626 12586 -5614
rect 12854 -5217 12904 -5205
rect 12854 -5614 12860 -5217
rect 12898 -5614 12904 -5217
rect 12854 -5626 12904 -5614
rect 13172 -5217 13222 -5205
rect 13172 -5614 13178 -5217
rect 13216 -5614 13222 -5217
rect 13172 -5626 13222 -5614
rect 13490 -5217 13540 -5205
rect 13490 -5614 13496 -5217
rect 13534 -5614 13540 -5217
rect 13490 -5626 13540 -5614
rect 13808 -5217 13858 -5205
rect 13808 -5614 13814 -5217
rect 13852 -5614 13858 -5217
rect 13808 -5626 13858 -5614
rect 14126 -5217 14176 -5205
rect 14126 -5614 14132 -5217
rect 14170 -5614 14176 -5217
rect 14126 -5626 14176 -5614
rect 14444 -5217 14494 -5205
rect 14444 -5614 14450 -5217
rect 14488 -5614 14494 -5217
rect 14444 -5626 14494 -5614
rect 14762 -5217 14812 -5205
rect 14762 -5614 14768 -5217
rect 14806 -5614 14812 -5217
rect 14762 -5626 14812 -5614
rect 15080 -5217 15130 -5205
rect 15080 -5614 15086 -5217
rect 15124 -5614 15130 -5217
rect 15080 -5626 15130 -5614
rect 15398 -5217 15448 -5205
rect 15398 -5614 15404 -5217
rect 15442 -5614 15448 -5217
rect 15398 -5626 15448 -5614
rect 15716 -5217 15766 -5205
rect 15716 -5614 15722 -5217
rect 15760 -5614 15766 -5217
rect 15716 -5626 15766 -5614
<< res0p35 >>
rect -15778 -5202 -15704 5202
rect -15460 -5202 -15386 5202
rect -15142 -5202 -15068 5202
rect -14824 -5202 -14750 5202
rect -14506 -5202 -14432 5202
rect -14188 -5202 -14114 5202
rect -13870 -5202 -13796 5202
rect -13552 -5202 -13478 5202
rect -13234 -5202 -13160 5202
rect -12916 -5202 -12842 5202
rect -12598 -5202 -12524 5202
rect -12280 -5202 -12206 5202
rect -11962 -5202 -11888 5202
rect -11644 -5202 -11570 5202
rect -11326 -5202 -11252 5202
rect -11008 -5202 -10934 5202
rect -10690 -5202 -10616 5202
rect -10372 -5202 -10298 5202
rect -10054 -5202 -9980 5202
rect -9736 -5202 -9662 5202
rect -9418 -5202 -9344 5202
rect -9100 -5202 -9026 5202
rect -8782 -5202 -8708 5202
rect -8464 -5202 -8390 5202
rect -8146 -5202 -8072 5202
rect -7828 -5202 -7754 5202
rect -7510 -5202 -7436 5202
rect -7192 -5202 -7118 5202
rect -6874 -5202 -6800 5202
rect -6556 -5202 -6482 5202
rect -6238 -5202 -6164 5202
rect -5920 -5202 -5846 5202
rect -5602 -5202 -5528 5202
rect -5284 -5202 -5210 5202
rect -4966 -5202 -4892 5202
rect -4648 -5202 -4574 5202
rect -4330 -5202 -4256 5202
rect -4012 -5202 -3938 5202
rect -3694 -5202 -3620 5202
rect -3376 -5202 -3302 5202
rect -3058 -5202 -2984 5202
rect -2740 -5202 -2666 5202
rect -2422 -5202 -2348 5202
rect -2104 -5202 -2030 5202
rect -1786 -5202 -1712 5202
rect -1468 -5202 -1394 5202
rect -1150 -5202 -1076 5202
rect -832 -5202 -758 5202
rect -514 -5202 -440 5202
rect -196 -5202 -122 5202
rect 122 -5202 196 5202
rect 440 -5202 514 5202
rect 758 -5202 832 5202
rect 1076 -5202 1150 5202
rect 1394 -5202 1468 5202
rect 1712 -5202 1786 5202
rect 2030 -5202 2104 5202
rect 2348 -5202 2422 5202
rect 2666 -5202 2740 5202
rect 2984 -5202 3058 5202
rect 3302 -5202 3376 5202
rect 3620 -5202 3694 5202
rect 3938 -5202 4012 5202
rect 4256 -5202 4330 5202
rect 4574 -5202 4648 5202
rect 4892 -5202 4966 5202
rect 5210 -5202 5284 5202
rect 5528 -5202 5602 5202
rect 5846 -5202 5920 5202
rect 6164 -5202 6238 5202
rect 6482 -5202 6556 5202
rect 6800 -5202 6874 5202
rect 7118 -5202 7192 5202
rect 7436 -5202 7510 5202
rect 7754 -5202 7828 5202
rect 8072 -5202 8146 5202
rect 8390 -5202 8464 5202
rect 8708 -5202 8782 5202
rect 9026 -5202 9100 5202
rect 9344 -5202 9418 5202
rect 9662 -5202 9736 5202
rect 9980 -5202 10054 5202
rect 10298 -5202 10372 5202
rect 10616 -5202 10690 5202
rect 10934 -5202 11008 5202
rect 11252 -5202 11326 5202
rect 11570 -5202 11644 5202
rect 11888 -5202 11962 5202
rect 12206 -5202 12280 5202
rect 12524 -5202 12598 5202
rect 12842 -5202 12916 5202
rect 13160 -5202 13234 5202
rect 13478 -5202 13552 5202
rect 13796 -5202 13870 5202
rect 14114 -5202 14188 5202
rect 14432 -5202 14506 5202
rect 14750 -5202 14824 5202
rect 15068 -5202 15142 5202
rect 15386 -5202 15460 5202
rect 15704 -5202 15778 5202
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 52 m 1 nx 100 wmin 0.350 lmin 0.50 rho 2000 val 298.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
