magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -144 -1064 144 1098
<< pmos >>
rect -50 -964 50 1036
<< pdiff >>
rect -108 1005 -50 1036
rect -108 971 -96 1005
rect -62 971 -50 1005
rect -108 937 -50 971
rect -108 903 -96 937
rect -62 903 -50 937
rect -108 869 -50 903
rect -108 835 -96 869
rect -62 835 -50 869
rect -108 801 -50 835
rect -108 767 -96 801
rect -62 767 -50 801
rect -108 733 -50 767
rect -108 699 -96 733
rect -62 699 -50 733
rect -108 665 -50 699
rect -108 631 -96 665
rect -62 631 -50 665
rect -108 597 -50 631
rect -108 563 -96 597
rect -62 563 -50 597
rect -108 529 -50 563
rect -108 495 -96 529
rect -62 495 -50 529
rect -108 461 -50 495
rect -108 427 -96 461
rect -62 427 -50 461
rect -108 393 -50 427
rect -108 359 -96 393
rect -62 359 -50 393
rect -108 325 -50 359
rect -108 291 -96 325
rect -62 291 -50 325
rect -108 257 -50 291
rect -108 223 -96 257
rect -62 223 -50 257
rect -108 189 -50 223
rect -108 155 -96 189
rect -62 155 -50 189
rect -108 121 -50 155
rect -108 87 -96 121
rect -62 87 -50 121
rect -108 53 -50 87
rect -108 19 -96 53
rect -62 19 -50 53
rect -108 -15 -50 19
rect -108 -49 -96 -15
rect -62 -49 -50 -15
rect -108 -83 -50 -49
rect -108 -117 -96 -83
rect -62 -117 -50 -83
rect -108 -151 -50 -117
rect -108 -185 -96 -151
rect -62 -185 -50 -151
rect -108 -219 -50 -185
rect -108 -253 -96 -219
rect -62 -253 -50 -219
rect -108 -287 -50 -253
rect -108 -321 -96 -287
rect -62 -321 -50 -287
rect -108 -355 -50 -321
rect -108 -389 -96 -355
rect -62 -389 -50 -355
rect -108 -423 -50 -389
rect -108 -457 -96 -423
rect -62 -457 -50 -423
rect -108 -491 -50 -457
rect -108 -525 -96 -491
rect -62 -525 -50 -491
rect -108 -559 -50 -525
rect -108 -593 -96 -559
rect -62 -593 -50 -559
rect -108 -627 -50 -593
rect -108 -661 -96 -627
rect -62 -661 -50 -627
rect -108 -695 -50 -661
rect -108 -729 -96 -695
rect -62 -729 -50 -695
rect -108 -763 -50 -729
rect -108 -797 -96 -763
rect -62 -797 -50 -763
rect -108 -831 -50 -797
rect -108 -865 -96 -831
rect -62 -865 -50 -831
rect -108 -899 -50 -865
rect -108 -933 -96 -899
rect -62 -933 -50 -899
rect -108 -964 -50 -933
rect 50 1005 108 1036
rect 50 971 62 1005
rect 96 971 108 1005
rect 50 937 108 971
rect 50 903 62 937
rect 96 903 108 937
rect 50 869 108 903
rect 50 835 62 869
rect 96 835 108 869
rect 50 801 108 835
rect 50 767 62 801
rect 96 767 108 801
rect 50 733 108 767
rect 50 699 62 733
rect 96 699 108 733
rect 50 665 108 699
rect 50 631 62 665
rect 96 631 108 665
rect 50 597 108 631
rect 50 563 62 597
rect 96 563 108 597
rect 50 529 108 563
rect 50 495 62 529
rect 96 495 108 529
rect 50 461 108 495
rect 50 427 62 461
rect 96 427 108 461
rect 50 393 108 427
rect 50 359 62 393
rect 96 359 108 393
rect 50 325 108 359
rect 50 291 62 325
rect 96 291 108 325
rect 50 257 108 291
rect 50 223 62 257
rect 96 223 108 257
rect 50 189 108 223
rect 50 155 62 189
rect 96 155 108 189
rect 50 121 108 155
rect 50 87 62 121
rect 96 87 108 121
rect 50 53 108 87
rect 50 19 62 53
rect 96 19 108 53
rect 50 -15 108 19
rect 50 -49 62 -15
rect 96 -49 108 -15
rect 50 -83 108 -49
rect 50 -117 62 -83
rect 96 -117 108 -83
rect 50 -151 108 -117
rect 50 -185 62 -151
rect 96 -185 108 -151
rect 50 -219 108 -185
rect 50 -253 62 -219
rect 96 -253 108 -219
rect 50 -287 108 -253
rect 50 -321 62 -287
rect 96 -321 108 -287
rect 50 -355 108 -321
rect 50 -389 62 -355
rect 96 -389 108 -355
rect 50 -423 108 -389
rect 50 -457 62 -423
rect 96 -457 108 -423
rect 50 -491 108 -457
rect 50 -525 62 -491
rect 96 -525 108 -491
rect 50 -559 108 -525
rect 50 -593 62 -559
rect 96 -593 108 -559
rect 50 -627 108 -593
rect 50 -661 62 -627
rect 96 -661 108 -627
rect 50 -695 108 -661
rect 50 -729 62 -695
rect 96 -729 108 -695
rect 50 -763 108 -729
rect 50 -797 62 -763
rect 96 -797 108 -763
rect 50 -831 108 -797
rect 50 -865 62 -831
rect 96 -865 108 -831
rect 50 -899 108 -865
rect 50 -933 62 -899
rect 96 -933 108 -899
rect 50 -964 108 -933
<< pdiffc >>
rect -96 971 -62 1005
rect -96 903 -62 937
rect -96 835 -62 869
rect -96 767 -62 801
rect -96 699 -62 733
rect -96 631 -62 665
rect -96 563 -62 597
rect -96 495 -62 529
rect -96 427 -62 461
rect -96 359 -62 393
rect -96 291 -62 325
rect -96 223 -62 257
rect -96 155 -62 189
rect -96 87 -62 121
rect -96 19 -62 53
rect -96 -49 -62 -15
rect -96 -117 -62 -83
rect -96 -185 -62 -151
rect -96 -253 -62 -219
rect -96 -321 -62 -287
rect -96 -389 -62 -355
rect -96 -457 -62 -423
rect -96 -525 -62 -491
rect -96 -593 -62 -559
rect -96 -661 -62 -627
rect -96 -729 -62 -695
rect -96 -797 -62 -763
rect -96 -865 -62 -831
rect -96 -933 -62 -899
rect 62 971 96 1005
rect 62 903 96 937
rect 62 835 96 869
rect 62 767 96 801
rect 62 699 96 733
rect 62 631 96 665
rect 62 563 96 597
rect 62 495 96 529
rect 62 427 96 461
rect 62 359 96 393
rect 62 291 96 325
rect 62 223 96 257
rect 62 155 96 189
rect 62 87 96 121
rect 62 19 96 53
rect 62 -49 96 -15
rect 62 -117 96 -83
rect 62 -185 96 -151
rect 62 -253 96 -219
rect 62 -321 96 -287
rect 62 -389 96 -355
rect 62 -457 96 -423
rect 62 -525 96 -491
rect 62 -593 96 -559
rect 62 -661 96 -627
rect 62 -729 96 -695
rect 62 -797 96 -763
rect 62 -865 96 -831
rect 62 -933 96 -899
<< poly >>
rect -50 1036 50 1062
rect -50 -1011 50 -964
rect -50 -1045 -17 -1011
rect 17 -1045 50 -1011
rect -50 -1061 50 -1045
<< polycont >>
rect -17 -1045 17 -1011
<< locali >>
rect -96 1005 -62 1040
rect -96 937 -62 955
rect -96 869 -62 883
rect -96 801 -62 811
rect -96 733 -62 739
rect -96 665 -62 667
rect -96 629 -62 631
rect -96 557 -62 563
rect -96 485 -62 495
rect -96 413 -62 427
rect -96 341 -62 359
rect -96 269 -62 291
rect -96 197 -62 223
rect -96 125 -62 155
rect -96 53 -62 87
rect -96 -15 -62 19
rect -96 -83 -62 -53
rect -96 -151 -62 -125
rect -96 -219 -62 -197
rect -96 -287 -62 -269
rect -96 -355 -62 -341
rect -96 -423 -62 -413
rect -96 -491 -62 -485
rect -96 -559 -62 -557
rect -96 -595 -62 -593
rect -96 -667 -62 -661
rect -96 -739 -62 -729
rect -96 -811 -62 -797
rect -96 -883 -62 -865
rect -96 -968 -62 -933
rect 62 1005 96 1040
rect 62 937 96 955
rect 62 869 96 883
rect 62 801 96 811
rect 62 733 96 739
rect 62 665 96 667
rect 62 629 96 631
rect 62 557 96 563
rect 62 485 96 495
rect 62 413 96 427
rect 62 341 96 359
rect 62 269 96 291
rect 62 197 96 223
rect 62 125 96 155
rect 62 53 96 87
rect 62 -15 96 19
rect 62 -83 96 -53
rect 62 -151 96 -125
rect 62 -219 96 -197
rect 62 -287 96 -269
rect 62 -355 96 -341
rect 62 -423 96 -413
rect 62 -491 96 -485
rect 62 -559 96 -557
rect 62 -595 96 -593
rect 62 -667 96 -661
rect 62 -739 96 -729
rect 62 -811 96 -797
rect 62 -883 96 -865
rect 62 -968 96 -933
rect -50 -1045 -17 -1011
rect 17 -1045 50 -1011
<< viali >>
rect -96 971 -62 989
rect -96 955 -62 971
rect -96 903 -62 917
rect -96 883 -62 903
rect -96 835 -62 845
rect -96 811 -62 835
rect -96 767 -62 773
rect -96 739 -62 767
rect -96 699 -62 701
rect -96 667 -62 699
rect -96 597 -62 629
rect -96 595 -62 597
rect -96 529 -62 557
rect -96 523 -62 529
rect -96 461 -62 485
rect -96 451 -62 461
rect -96 393 -62 413
rect -96 379 -62 393
rect -96 325 -62 341
rect -96 307 -62 325
rect -96 257 -62 269
rect -96 235 -62 257
rect -96 189 -62 197
rect -96 163 -62 189
rect -96 121 -62 125
rect -96 91 -62 121
rect -96 19 -62 53
rect -96 -49 -62 -19
rect -96 -53 -62 -49
rect -96 -117 -62 -91
rect -96 -125 -62 -117
rect -96 -185 -62 -163
rect -96 -197 -62 -185
rect -96 -253 -62 -235
rect -96 -269 -62 -253
rect -96 -321 -62 -307
rect -96 -341 -62 -321
rect -96 -389 -62 -379
rect -96 -413 -62 -389
rect -96 -457 -62 -451
rect -96 -485 -62 -457
rect -96 -525 -62 -523
rect -96 -557 -62 -525
rect -96 -627 -62 -595
rect -96 -629 -62 -627
rect -96 -695 -62 -667
rect -96 -701 -62 -695
rect -96 -763 -62 -739
rect -96 -773 -62 -763
rect -96 -831 -62 -811
rect -96 -845 -62 -831
rect -96 -899 -62 -883
rect -96 -917 -62 -899
rect 62 971 96 989
rect 62 955 96 971
rect 62 903 96 917
rect 62 883 96 903
rect 62 835 96 845
rect 62 811 96 835
rect 62 767 96 773
rect 62 739 96 767
rect 62 699 96 701
rect 62 667 96 699
rect 62 597 96 629
rect 62 595 96 597
rect 62 529 96 557
rect 62 523 96 529
rect 62 461 96 485
rect 62 451 96 461
rect 62 393 96 413
rect 62 379 96 393
rect 62 325 96 341
rect 62 307 96 325
rect 62 257 96 269
rect 62 235 96 257
rect 62 189 96 197
rect 62 163 96 189
rect 62 121 96 125
rect 62 91 96 121
rect 62 19 96 53
rect 62 -49 96 -19
rect 62 -53 96 -49
rect 62 -117 96 -91
rect 62 -125 96 -117
rect 62 -185 96 -163
rect 62 -197 96 -185
rect 62 -253 96 -235
rect 62 -269 96 -253
rect 62 -321 96 -307
rect 62 -341 96 -321
rect 62 -389 96 -379
rect 62 -413 96 -389
rect 62 -457 96 -451
rect 62 -485 96 -457
rect 62 -525 96 -523
rect 62 -557 96 -525
rect 62 -627 96 -595
rect 62 -629 96 -627
rect 62 -695 96 -667
rect 62 -701 96 -695
rect 62 -763 96 -739
rect 62 -773 96 -763
rect 62 -831 96 -811
rect 62 -845 96 -831
rect 62 -899 96 -883
rect 62 -917 96 -899
rect -17 -1045 17 -1011
<< metal1 >>
rect -102 989 -56 1036
rect -102 955 -96 989
rect -62 955 -56 989
rect -102 917 -56 955
rect -102 883 -96 917
rect -62 883 -56 917
rect -102 845 -56 883
rect -102 811 -96 845
rect -62 811 -56 845
rect -102 773 -56 811
rect -102 739 -96 773
rect -62 739 -56 773
rect -102 701 -56 739
rect -102 667 -96 701
rect -62 667 -56 701
rect -102 629 -56 667
rect -102 595 -96 629
rect -62 595 -56 629
rect -102 557 -56 595
rect -102 523 -96 557
rect -62 523 -56 557
rect -102 485 -56 523
rect -102 451 -96 485
rect -62 451 -56 485
rect -102 413 -56 451
rect -102 379 -96 413
rect -62 379 -56 413
rect -102 341 -56 379
rect -102 307 -96 341
rect -62 307 -56 341
rect -102 269 -56 307
rect -102 235 -96 269
rect -62 235 -56 269
rect -102 197 -56 235
rect -102 163 -96 197
rect -62 163 -56 197
rect -102 125 -56 163
rect -102 91 -96 125
rect -62 91 -56 125
rect -102 53 -56 91
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -91 -56 -53
rect -102 -125 -96 -91
rect -62 -125 -56 -91
rect -102 -163 -56 -125
rect -102 -197 -96 -163
rect -62 -197 -56 -163
rect -102 -235 -56 -197
rect -102 -269 -96 -235
rect -62 -269 -56 -235
rect -102 -307 -56 -269
rect -102 -341 -96 -307
rect -62 -341 -56 -307
rect -102 -379 -56 -341
rect -102 -413 -96 -379
rect -62 -413 -56 -379
rect -102 -451 -56 -413
rect -102 -485 -96 -451
rect -62 -485 -56 -451
rect -102 -523 -56 -485
rect -102 -557 -96 -523
rect -62 -557 -56 -523
rect -102 -595 -56 -557
rect -102 -629 -96 -595
rect -62 -629 -56 -595
rect -102 -667 -56 -629
rect -102 -701 -96 -667
rect -62 -701 -56 -667
rect -102 -739 -56 -701
rect -102 -773 -96 -739
rect -62 -773 -56 -739
rect -102 -811 -56 -773
rect -102 -845 -96 -811
rect -62 -845 -56 -811
rect -102 -883 -56 -845
rect -102 -917 -96 -883
rect -62 -917 -56 -883
rect -102 -964 -56 -917
rect 56 989 102 1036
rect 56 955 62 989
rect 96 955 102 989
rect 56 917 102 955
rect 56 883 62 917
rect 96 883 102 917
rect 56 845 102 883
rect 56 811 62 845
rect 96 811 102 845
rect 56 773 102 811
rect 56 739 62 773
rect 96 739 102 773
rect 56 701 102 739
rect 56 667 62 701
rect 96 667 102 701
rect 56 629 102 667
rect 56 595 62 629
rect 96 595 102 629
rect 56 557 102 595
rect 56 523 62 557
rect 96 523 102 557
rect 56 485 102 523
rect 56 451 62 485
rect 96 451 102 485
rect 56 413 102 451
rect 56 379 62 413
rect 96 379 102 413
rect 56 341 102 379
rect 56 307 62 341
rect 96 307 102 341
rect 56 269 102 307
rect 56 235 62 269
rect 96 235 102 269
rect 56 197 102 235
rect 56 163 62 197
rect 96 163 102 197
rect 56 125 102 163
rect 56 91 62 125
rect 96 91 102 125
rect 56 53 102 91
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -91 102 -53
rect 56 -125 62 -91
rect 96 -125 102 -91
rect 56 -163 102 -125
rect 56 -197 62 -163
rect 96 -197 102 -163
rect 56 -235 102 -197
rect 56 -269 62 -235
rect 96 -269 102 -235
rect 56 -307 102 -269
rect 56 -341 62 -307
rect 96 -341 102 -307
rect 56 -379 102 -341
rect 56 -413 62 -379
rect 96 -413 102 -379
rect 56 -451 102 -413
rect 56 -485 62 -451
rect 96 -485 102 -451
rect 56 -523 102 -485
rect 56 -557 62 -523
rect 96 -557 102 -523
rect 56 -595 102 -557
rect 56 -629 62 -595
rect 96 -629 102 -595
rect 56 -667 102 -629
rect 56 -701 62 -667
rect 96 -701 102 -667
rect 56 -739 102 -701
rect 56 -773 62 -739
rect 96 -773 102 -739
rect 56 -811 102 -773
rect 56 -845 62 -811
rect 96 -845 102 -811
rect 56 -883 102 -845
rect 56 -917 62 -883
rect 96 -917 102 -883
rect 56 -964 102 -917
rect -46 -1011 46 -1005
rect -46 -1045 -17 -1011
rect 17 -1045 46 -1011
rect -46 -1051 46 -1045
<< end >>
