magic
tech sky130A
magscale 1 2
timestamp 1667443905
<< nwell >>
rect -194 -800 194 800
<< pmos >>
rect -100 -700 100 700
<< pdiff >>
rect -158 688 -100 700
rect -158 -688 -146 688
rect -112 -688 -100 688
rect -158 -700 -100 -688
rect 100 688 158 700
rect 100 -688 112 688
rect 146 -688 158 688
rect 100 -700 158 -688
<< pdiffc >>
rect -146 -688 -112 688
rect 112 -688 146 688
<< poly >>
rect -100 781 100 797
rect -100 747 -84 781
rect 84 747 100 781
rect -100 700 100 747
rect -100 -747 100 -700
rect -100 -781 -84 -747
rect 84 -781 100 -747
rect -100 -797 100 -781
<< polycont >>
rect -84 747 84 781
rect -84 -781 84 -747
<< locali >>
rect -100 747 -84 781
rect 84 747 100 781
rect -146 688 -112 704
rect -146 -704 -112 -688
rect 112 688 146 704
rect 112 -704 146 -688
rect -100 -781 -84 -747
rect 84 -781 100 -747
<< viali >>
rect -84 747 84 781
rect -146 -688 -112 688
rect 112 -688 146 688
rect -84 -781 84 -747
<< metal1 >>
rect -96 781 96 787
rect -96 747 -84 781
rect 84 747 96 781
rect -96 741 96 747
rect -152 688 -106 700
rect -152 -688 -146 688
rect -112 -688 -106 688
rect -152 -700 -106 -688
rect 106 688 152 700
rect 106 -688 112 688
rect 146 -688 152 688
rect 106 -700 152 -688
rect -96 -747 96 -741
rect -96 -781 -84 -747
rect 84 -781 96 -747
rect -96 -787 96 -781
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
