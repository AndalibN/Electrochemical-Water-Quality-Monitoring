magic
tech sky130A
magscale 1 2
timestamp 1668227999
<< metal3 >>
rect -1009 922 -10 950
rect -1009 78 -94 922
rect -30 78 -10 922
rect -1009 50 -10 78
rect 70 922 1069 950
rect 70 78 985 922
rect 1049 78 1069 922
rect 70 50 1069 78
rect -1009 -78 -10 -50
rect -1009 -922 -94 -78
rect -30 -922 -10 -78
rect -1009 -950 -10 -922
rect 70 -78 1069 -50
rect 70 -922 985 -78
rect 1049 -922 1069 -78
rect 70 -950 1069 -922
<< via3 >>
rect -94 78 -30 922
rect 985 78 1049 922
rect -94 -922 -30 -78
rect 985 -922 1049 -78
<< mimcap >>
rect -909 810 -209 850
rect -909 190 -869 810
rect -249 190 -209 810
rect -909 150 -209 190
rect 170 810 870 850
rect 170 190 210 810
rect 830 190 870 810
rect 170 150 870 190
rect -909 -190 -209 -150
rect -909 -810 -869 -190
rect -249 -810 -209 -190
rect -909 -850 -209 -810
rect 170 -190 870 -150
rect 170 -810 210 -190
rect 830 -810 870 -190
rect 170 -850 870 -810
<< mimcapcontact >>
rect -869 190 -249 810
rect 210 190 830 810
rect -869 -810 -249 -190
rect 210 -810 830 -190
<< metal4 >>
rect -611 811 -507 1000
rect -141 938 -37 1000
rect -141 922 -14 938
rect -870 810 -248 811
rect -870 190 -869 810
rect -249 190 -248 810
rect -870 189 -248 190
rect -611 -189 -507 189
rect -141 78 -94 922
rect -30 78 -14 922
rect 468 811 572 1000
rect 938 938 1042 1000
rect 938 922 1065 938
rect 209 810 831 811
rect 209 190 210 810
rect 830 190 831 810
rect 209 189 831 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -870 -190 -248 -189
rect -870 -810 -869 -190
rect -249 -810 -248 -190
rect -870 -811 -248 -810
rect -611 -1000 -507 -811
rect -141 -922 -94 -78
rect -30 -922 -14 -78
rect 468 -189 572 189
rect 938 78 985 922
rect 1049 78 1065 922
rect 938 62 1065 78
rect 938 -62 1042 62
rect 938 -78 1065 -62
rect 209 -190 831 -189
rect 209 -810 210 -190
rect 830 -810 831 -190
rect 209 -811 831 -810
rect -141 -938 -14 -922
rect -141 -1000 -37 -938
rect 468 -1000 572 -811
rect 938 -922 985 -78
rect 1049 -922 1065 -78
rect 938 -938 1065 -922
rect 938 -1000 1042 -938
<< properties >>
string FIXED_BBOX 10 50 910 950
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.5 l 3.5 val 27.16 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
