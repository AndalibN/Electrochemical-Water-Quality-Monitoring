magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -345 -1498 323 1464
<< pmos >>
rect -251 -1436 -51 1364
rect 7 -1436 207 1364
<< pdiff >>
rect -309 1341 -251 1364
rect -309 1307 -297 1341
rect -263 1307 -251 1341
rect -309 1273 -251 1307
rect -309 1239 -297 1273
rect -263 1239 -251 1273
rect -309 1205 -251 1239
rect -309 1171 -297 1205
rect -263 1171 -251 1205
rect -309 1137 -251 1171
rect -309 1103 -297 1137
rect -263 1103 -251 1137
rect -309 1069 -251 1103
rect -309 1035 -297 1069
rect -263 1035 -251 1069
rect -309 1001 -251 1035
rect -309 967 -297 1001
rect -263 967 -251 1001
rect -309 933 -251 967
rect -309 899 -297 933
rect -263 899 -251 933
rect -309 865 -251 899
rect -309 831 -297 865
rect -263 831 -251 865
rect -309 797 -251 831
rect -309 763 -297 797
rect -263 763 -251 797
rect -309 729 -251 763
rect -309 695 -297 729
rect -263 695 -251 729
rect -309 661 -251 695
rect -309 627 -297 661
rect -263 627 -251 661
rect -309 593 -251 627
rect -309 559 -297 593
rect -263 559 -251 593
rect -309 525 -251 559
rect -309 491 -297 525
rect -263 491 -251 525
rect -309 457 -251 491
rect -309 423 -297 457
rect -263 423 -251 457
rect -309 389 -251 423
rect -309 355 -297 389
rect -263 355 -251 389
rect -309 321 -251 355
rect -309 287 -297 321
rect -263 287 -251 321
rect -309 253 -251 287
rect -309 219 -297 253
rect -263 219 -251 253
rect -309 185 -251 219
rect -309 151 -297 185
rect -263 151 -251 185
rect -309 117 -251 151
rect -309 83 -297 117
rect -263 83 -251 117
rect -309 49 -251 83
rect -309 15 -297 49
rect -263 15 -251 49
rect -309 -19 -251 15
rect -309 -53 -297 -19
rect -263 -53 -251 -19
rect -309 -87 -251 -53
rect -309 -121 -297 -87
rect -263 -121 -251 -87
rect -309 -155 -251 -121
rect -309 -189 -297 -155
rect -263 -189 -251 -155
rect -309 -223 -251 -189
rect -309 -257 -297 -223
rect -263 -257 -251 -223
rect -309 -291 -251 -257
rect -309 -325 -297 -291
rect -263 -325 -251 -291
rect -309 -359 -251 -325
rect -309 -393 -297 -359
rect -263 -393 -251 -359
rect -309 -427 -251 -393
rect -309 -461 -297 -427
rect -263 -461 -251 -427
rect -309 -495 -251 -461
rect -309 -529 -297 -495
rect -263 -529 -251 -495
rect -309 -563 -251 -529
rect -309 -597 -297 -563
rect -263 -597 -251 -563
rect -309 -631 -251 -597
rect -309 -665 -297 -631
rect -263 -665 -251 -631
rect -309 -699 -251 -665
rect -309 -733 -297 -699
rect -263 -733 -251 -699
rect -309 -767 -251 -733
rect -309 -801 -297 -767
rect -263 -801 -251 -767
rect -309 -835 -251 -801
rect -309 -869 -297 -835
rect -263 -869 -251 -835
rect -309 -903 -251 -869
rect -309 -937 -297 -903
rect -263 -937 -251 -903
rect -309 -971 -251 -937
rect -309 -1005 -297 -971
rect -263 -1005 -251 -971
rect -309 -1039 -251 -1005
rect -309 -1073 -297 -1039
rect -263 -1073 -251 -1039
rect -309 -1107 -251 -1073
rect -309 -1141 -297 -1107
rect -263 -1141 -251 -1107
rect -309 -1175 -251 -1141
rect -309 -1209 -297 -1175
rect -263 -1209 -251 -1175
rect -309 -1243 -251 -1209
rect -309 -1277 -297 -1243
rect -263 -1277 -251 -1243
rect -309 -1311 -251 -1277
rect -309 -1345 -297 -1311
rect -263 -1345 -251 -1311
rect -309 -1379 -251 -1345
rect -309 -1413 -297 -1379
rect -263 -1413 -251 -1379
rect -309 -1436 -251 -1413
rect -51 1341 7 1364
rect -51 1307 -39 1341
rect -5 1307 7 1341
rect -51 1273 7 1307
rect -51 1239 -39 1273
rect -5 1239 7 1273
rect -51 1205 7 1239
rect -51 1171 -39 1205
rect -5 1171 7 1205
rect -51 1137 7 1171
rect -51 1103 -39 1137
rect -5 1103 7 1137
rect -51 1069 7 1103
rect -51 1035 -39 1069
rect -5 1035 7 1069
rect -51 1001 7 1035
rect -51 967 -39 1001
rect -5 967 7 1001
rect -51 933 7 967
rect -51 899 -39 933
rect -5 899 7 933
rect -51 865 7 899
rect -51 831 -39 865
rect -5 831 7 865
rect -51 797 7 831
rect -51 763 -39 797
rect -5 763 7 797
rect -51 729 7 763
rect -51 695 -39 729
rect -5 695 7 729
rect -51 661 7 695
rect -51 627 -39 661
rect -5 627 7 661
rect -51 593 7 627
rect -51 559 -39 593
rect -5 559 7 593
rect -51 525 7 559
rect -51 491 -39 525
rect -5 491 7 525
rect -51 457 7 491
rect -51 423 -39 457
rect -5 423 7 457
rect -51 389 7 423
rect -51 355 -39 389
rect -5 355 7 389
rect -51 321 7 355
rect -51 287 -39 321
rect -5 287 7 321
rect -51 253 7 287
rect -51 219 -39 253
rect -5 219 7 253
rect -51 185 7 219
rect -51 151 -39 185
rect -5 151 7 185
rect -51 117 7 151
rect -51 83 -39 117
rect -5 83 7 117
rect -51 49 7 83
rect -51 15 -39 49
rect -5 15 7 49
rect -51 -19 7 15
rect -51 -53 -39 -19
rect -5 -53 7 -19
rect -51 -87 7 -53
rect -51 -121 -39 -87
rect -5 -121 7 -87
rect -51 -155 7 -121
rect -51 -189 -39 -155
rect -5 -189 7 -155
rect -51 -223 7 -189
rect -51 -257 -39 -223
rect -5 -257 7 -223
rect -51 -291 7 -257
rect -51 -325 -39 -291
rect -5 -325 7 -291
rect -51 -359 7 -325
rect -51 -393 -39 -359
rect -5 -393 7 -359
rect -51 -427 7 -393
rect -51 -461 -39 -427
rect -5 -461 7 -427
rect -51 -495 7 -461
rect -51 -529 -39 -495
rect -5 -529 7 -495
rect -51 -563 7 -529
rect -51 -597 -39 -563
rect -5 -597 7 -563
rect -51 -631 7 -597
rect -51 -665 -39 -631
rect -5 -665 7 -631
rect -51 -699 7 -665
rect -51 -733 -39 -699
rect -5 -733 7 -699
rect -51 -767 7 -733
rect -51 -801 -39 -767
rect -5 -801 7 -767
rect -51 -835 7 -801
rect -51 -869 -39 -835
rect -5 -869 7 -835
rect -51 -903 7 -869
rect -51 -937 -39 -903
rect -5 -937 7 -903
rect -51 -971 7 -937
rect -51 -1005 -39 -971
rect -5 -1005 7 -971
rect -51 -1039 7 -1005
rect -51 -1073 -39 -1039
rect -5 -1073 7 -1039
rect -51 -1107 7 -1073
rect -51 -1141 -39 -1107
rect -5 -1141 7 -1107
rect -51 -1175 7 -1141
rect -51 -1209 -39 -1175
rect -5 -1209 7 -1175
rect -51 -1243 7 -1209
rect -51 -1277 -39 -1243
rect -5 -1277 7 -1243
rect -51 -1311 7 -1277
rect -51 -1345 -39 -1311
rect -5 -1345 7 -1311
rect -51 -1379 7 -1345
rect -51 -1413 -39 -1379
rect -5 -1413 7 -1379
rect -51 -1436 7 -1413
rect 207 1341 287 1364
rect 207 1307 230 1341
rect 264 1307 287 1341
rect 207 1273 287 1307
rect 207 1239 230 1273
rect 264 1239 287 1273
rect 207 1205 287 1239
rect 207 1171 230 1205
rect 264 1171 287 1205
rect 207 1137 287 1171
rect 207 1103 230 1137
rect 264 1103 287 1137
rect 207 1069 287 1103
rect 207 1035 230 1069
rect 264 1035 287 1069
rect 207 1001 287 1035
rect 207 967 230 1001
rect 264 967 287 1001
rect 207 933 287 967
rect 207 899 230 933
rect 264 899 287 933
rect 207 865 287 899
rect 207 831 230 865
rect 264 831 287 865
rect 207 797 287 831
rect 207 763 230 797
rect 264 763 287 797
rect 207 729 287 763
rect 207 695 230 729
rect 264 695 287 729
rect 207 661 287 695
rect 207 627 230 661
rect 264 627 287 661
rect 207 593 287 627
rect 207 559 230 593
rect 264 559 287 593
rect 207 525 287 559
rect 207 491 230 525
rect 264 491 287 525
rect 207 457 287 491
rect 207 423 230 457
rect 264 423 287 457
rect 207 389 287 423
rect 207 355 230 389
rect 264 355 287 389
rect 207 321 287 355
rect 207 287 230 321
rect 264 287 287 321
rect 207 253 287 287
rect 207 219 230 253
rect 264 219 287 253
rect 207 185 287 219
rect 207 151 230 185
rect 264 151 287 185
rect 207 117 287 151
rect 207 83 230 117
rect 264 83 287 117
rect 207 49 287 83
rect 207 15 230 49
rect 264 15 287 49
rect 207 -19 287 15
rect 207 -53 230 -19
rect 264 -53 287 -19
rect 207 -87 287 -53
rect 207 -121 230 -87
rect 264 -121 287 -87
rect 207 -155 287 -121
rect 207 -189 230 -155
rect 264 -189 287 -155
rect 207 -223 287 -189
rect 207 -257 230 -223
rect 264 -257 287 -223
rect 207 -291 287 -257
rect 207 -325 230 -291
rect 264 -325 287 -291
rect 207 -359 287 -325
rect 207 -393 230 -359
rect 264 -393 287 -359
rect 207 -427 287 -393
rect 207 -461 230 -427
rect 264 -461 287 -427
rect 207 -495 287 -461
rect 207 -529 230 -495
rect 264 -529 287 -495
rect 207 -563 287 -529
rect 207 -597 230 -563
rect 264 -597 287 -563
rect 207 -631 287 -597
rect 207 -665 230 -631
rect 264 -665 287 -631
rect 207 -699 287 -665
rect 207 -733 230 -699
rect 264 -733 287 -699
rect 207 -767 287 -733
rect 207 -801 230 -767
rect 264 -801 287 -767
rect 207 -835 287 -801
rect 207 -869 230 -835
rect 264 -869 287 -835
rect 207 -903 287 -869
rect 207 -937 230 -903
rect 264 -937 287 -903
rect 207 -971 287 -937
rect 207 -1005 230 -971
rect 264 -1005 287 -971
rect 207 -1039 287 -1005
rect 207 -1073 230 -1039
rect 264 -1073 287 -1039
rect 207 -1107 287 -1073
rect 207 -1141 230 -1107
rect 264 -1141 287 -1107
rect 207 -1175 287 -1141
rect 207 -1209 230 -1175
rect 264 -1209 287 -1175
rect 207 -1243 287 -1209
rect 207 -1277 230 -1243
rect 264 -1277 287 -1243
rect 207 -1311 287 -1277
rect 207 -1345 230 -1311
rect 264 -1345 287 -1311
rect 207 -1379 287 -1345
rect 207 -1413 230 -1379
rect 264 -1413 287 -1379
rect 207 -1436 287 -1413
<< pdiffc >>
rect -297 1307 -263 1341
rect -297 1239 -263 1273
rect -297 1171 -263 1205
rect -297 1103 -263 1137
rect -297 1035 -263 1069
rect -297 967 -263 1001
rect -297 899 -263 933
rect -297 831 -263 865
rect -297 763 -263 797
rect -297 695 -263 729
rect -297 627 -263 661
rect -297 559 -263 593
rect -297 491 -263 525
rect -297 423 -263 457
rect -297 355 -263 389
rect -297 287 -263 321
rect -297 219 -263 253
rect -297 151 -263 185
rect -297 83 -263 117
rect -297 15 -263 49
rect -297 -53 -263 -19
rect -297 -121 -263 -87
rect -297 -189 -263 -155
rect -297 -257 -263 -223
rect -297 -325 -263 -291
rect -297 -393 -263 -359
rect -297 -461 -263 -427
rect -297 -529 -263 -495
rect -297 -597 -263 -563
rect -297 -665 -263 -631
rect -297 -733 -263 -699
rect -297 -801 -263 -767
rect -297 -869 -263 -835
rect -297 -937 -263 -903
rect -297 -1005 -263 -971
rect -297 -1073 -263 -1039
rect -297 -1141 -263 -1107
rect -297 -1209 -263 -1175
rect -297 -1277 -263 -1243
rect -297 -1345 -263 -1311
rect -297 -1413 -263 -1379
rect -39 1307 -5 1341
rect -39 1239 -5 1273
rect -39 1171 -5 1205
rect -39 1103 -5 1137
rect -39 1035 -5 1069
rect -39 967 -5 1001
rect -39 899 -5 933
rect -39 831 -5 865
rect -39 763 -5 797
rect -39 695 -5 729
rect -39 627 -5 661
rect -39 559 -5 593
rect -39 491 -5 525
rect -39 423 -5 457
rect -39 355 -5 389
rect -39 287 -5 321
rect -39 219 -5 253
rect -39 151 -5 185
rect -39 83 -5 117
rect -39 15 -5 49
rect -39 -53 -5 -19
rect -39 -121 -5 -87
rect -39 -189 -5 -155
rect -39 -257 -5 -223
rect -39 -325 -5 -291
rect -39 -393 -5 -359
rect -39 -461 -5 -427
rect -39 -529 -5 -495
rect -39 -597 -5 -563
rect -39 -665 -5 -631
rect -39 -733 -5 -699
rect -39 -801 -5 -767
rect -39 -869 -5 -835
rect -39 -937 -5 -903
rect -39 -1005 -5 -971
rect -39 -1073 -5 -1039
rect -39 -1141 -5 -1107
rect -39 -1209 -5 -1175
rect -39 -1277 -5 -1243
rect -39 -1345 -5 -1311
rect -39 -1413 -5 -1379
rect 230 1307 264 1341
rect 230 1239 264 1273
rect 230 1171 264 1205
rect 230 1103 264 1137
rect 230 1035 264 1069
rect 230 967 264 1001
rect 230 899 264 933
rect 230 831 264 865
rect 230 763 264 797
rect 230 695 264 729
rect 230 627 264 661
rect 230 559 264 593
rect 230 491 264 525
rect 230 423 264 457
rect 230 355 264 389
rect 230 287 264 321
rect 230 219 264 253
rect 230 151 264 185
rect 230 83 264 117
rect 230 15 264 49
rect 230 -53 264 -19
rect 230 -121 264 -87
rect 230 -189 264 -155
rect 230 -257 264 -223
rect 230 -325 264 -291
rect 230 -393 264 -359
rect 230 -461 264 -427
rect 230 -529 264 -495
rect 230 -597 264 -563
rect 230 -665 264 -631
rect 230 -733 264 -699
rect 230 -801 264 -767
rect 230 -869 264 -835
rect 230 -937 264 -903
rect 230 -1005 264 -971
rect 230 -1073 264 -1039
rect 230 -1141 264 -1107
rect 230 -1209 264 -1175
rect 230 -1277 264 -1243
rect 230 -1345 264 -1311
rect 230 -1413 264 -1379
<< poly >>
rect -251 1445 -51 1461
rect -251 1411 -202 1445
rect -168 1411 -134 1445
rect -100 1411 -51 1445
rect -251 1364 -51 1411
rect 7 1364 207 1461
rect -251 -1451 -51 -1436
rect 7 -1451 207 -1436
rect -251 -1491 207 -1451
<< polycont >>
rect -202 1411 -168 1445
rect -134 1411 -100 1445
<< locali >>
rect -251 1411 -204 1445
rect -168 1411 -134 1445
rect -98 1411 -51 1445
rect -297 1349 -263 1368
rect -297 1277 -263 1307
rect -297 1205 -263 1239
rect -297 1137 -263 1171
rect -297 1069 -263 1099
rect -297 1001 -263 1027
rect -297 933 -263 955
rect -297 865 -263 883
rect -297 797 -263 811
rect -297 729 -263 739
rect -297 661 -263 667
rect -297 593 -263 595
rect -297 557 -263 559
rect -297 485 -263 491
rect -297 413 -263 423
rect -297 341 -263 355
rect -297 269 -263 287
rect -297 197 -263 219
rect -297 125 -263 151
rect -297 53 -263 83
rect -297 -19 -263 15
rect -297 -87 -263 -53
rect -297 -155 -263 -125
rect -297 -223 -263 -197
rect -297 -291 -263 -269
rect -297 -359 -263 -341
rect -297 -427 -263 -413
rect -297 -495 -263 -485
rect -297 -563 -263 -557
rect -297 -631 -263 -629
rect -297 -667 -263 -665
rect -297 -739 -263 -733
rect -297 -811 -263 -801
rect -297 -883 -263 -869
rect -297 -955 -263 -937
rect -297 -1027 -263 -1005
rect -297 -1099 -263 -1073
rect -297 -1171 -263 -1141
rect -297 -1243 -263 -1209
rect -297 -1311 -263 -1277
rect -297 -1379 -263 -1349
rect -297 -1440 -263 -1421
rect -39 1349 -5 1368
rect -39 1277 -5 1307
rect -39 1205 -5 1239
rect -39 1137 -5 1171
rect -39 1069 -5 1099
rect -39 1001 -5 1027
rect -39 933 -5 955
rect -39 865 -5 883
rect -39 797 -5 811
rect -39 729 -5 739
rect -39 661 -5 667
rect -39 593 -5 595
rect -39 557 -5 559
rect -39 485 -5 491
rect -39 413 -5 423
rect -39 341 -5 355
rect -39 269 -5 287
rect -39 197 -5 219
rect -39 125 -5 151
rect -39 53 -5 83
rect -39 -19 -5 15
rect -39 -87 -5 -53
rect -39 -155 -5 -125
rect -39 -223 -5 -197
rect -39 -291 -5 -269
rect -39 -359 -5 -341
rect -39 -427 -5 -413
rect -39 -495 -5 -485
rect -39 -563 -5 -557
rect -39 -631 -5 -629
rect -39 -667 -5 -665
rect -39 -739 -5 -733
rect -39 -811 -5 -801
rect -39 -883 -5 -869
rect -39 -955 -5 -937
rect -39 -1027 -5 -1005
rect -39 -1099 -5 -1073
rect -39 -1171 -5 -1141
rect -39 -1243 -5 -1209
rect -39 -1311 -5 -1277
rect -39 -1379 -5 -1349
rect -39 -1440 -5 -1421
rect 230 1349 264 1368
rect 230 1277 264 1307
rect 230 1205 264 1239
rect 230 1137 264 1171
rect 230 1069 264 1099
rect 230 1001 264 1027
rect 230 933 264 955
rect 230 865 264 883
rect 230 797 264 811
rect 230 729 264 739
rect 230 661 264 667
rect 230 593 264 595
rect 230 557 264 559
rect 230 485 264 491
rect 230 413 264 423
rect 230 341 264 355
rect 230 269 264 287
rect 230 197 264 219
rect 230 125 264 151
rect 230 53 264 83
rect 230 -19 264 15
rect 230 -87 264 -53
rect 230 -155 264 -125
rect 230 -223 264 -197
rect 230 -291 264 -269
rect 230 -359 264 -341
rect 230 -427 264 -413
rect 230 -495 264 -485
rect 230 -563 264 -557
rect 230 -631 264 -629
rect 230 -667 264 -665
rect 230 -739 264 -733
rect 230 -811 264 -801
rect 230 -883 264 -869
rect 230 -955 264 -937
rect 230 -1027 264 -1005
rect 230 -1099 264 -1073
rect 230 -1171 264 -1141
rect 230 -1243 264 -1209
rect 230 -1311 264 -1277
rect 230 -1379 264 -1349
rect 230 -1440 264 -1421
<< viali >>
rect -204 1411 -202 1445
rect -202 1411 -170 1445
rect -132 1411 -100 1445
rect -100 1411 -98 1445
rect -297 1341 -263 1349
rect -297 1315 -263 1341
rect -297 1273 -263 1277
rect -297 1243 -263 1273
rect -297 1171 -263 1205
rect -297 1103 -263 1133
rect -297 1099 -263 1103
rect -297 1035 -263 1061
rect -297 1027 -263 1035
rect -297 967 -263 989
rect -297 955 -263 967
rect -297 899 -263 917
rect -297 883 -263 899
rect -297 831 -263 845
rect -297 811 -263 831
rect -297 763 -263 773
rect -297 739 -263 763
rect -297 695 -263 701
rect -297 667 -263 695
rect -297 627 -263 629
rect -297 595 -263 627
rect -297 525 -263 557
rect -297 523 -263 525
rect -297 457 -263 485
rect -297 451 -263 457
rect -297 389 -263 413
rect -297 379 -263 389
rect -297 321 -263 341
rect -297 307 -263 321
rect -297 253 -263 269
rect -297 235 -263 253
rect -297 185 -263 197
rect -297 163 -263 185
rect -297 117 -263 125
rect -297 91 -263 117
rect -297 49 -263 53
rect -297 19 -263 49
rect -297 -53 -263 -19
rect -297 -121 -263 -91
rect -297 -125 -263 -121
rect -297 -189 -263 -163
rect -297 -197 -263 -189
rect -297 -257 -263 -235
rect -297 -269 -263 -257
rect -297 -325 -263 -307
rect -297 -341 -263 -325
rect -297 -393 -263 -379
rect -297 -413 -263 -393
rect -297 -461 -263 -451
rect -297 -485 -263 -461
rect -297 -529 -263 -523
rect -297 -557 -263 -529
rect -297 -597 -263 -595
rect -297 -629 -263 -597
rect -297 -699 -263 -667
rect -297 -701 -263 -699
rect -297 -767 -263 -739
rect -297 -773 -263 -767
rect -297 -835 -263 -811
rect -297 -845 -263 -835
rect -297 -903 -263 -883
rect -297 -917 -263 -903
rect -297 -971 -263 -955
rect -297 -989 -263 -971
rect -297 -1039 -263 -1027
rect -297 -1061 -263 -1039
rect -297 -1107 -263 -1099
rect -297 -1133 -263 -1107
rect -297 -1175 -263 -1171
rect -297 -1205 -263 -1175
rect -297 -1277 -263 -1243
rect -297 -1345 -263 -1315
rect -297 -1349 -263 -1345
rect -297 -1413 -263 -1387
rect -297 -1421 -263 -1413
rect -39 1341 -5 1349
rect -39 1315 -5 1341
rect -39 1273 -5 1277
rect -39 1243 -5 1273
rect -39 1171 -5 1205
rect -39 1103 -5 1133
rect -39 1099 -5 1103
rect -39 1035 -5 1061
rect -39 1027 -5 1035
rect -39 967 -5 989
rect -39 955 -5 967
rect -39 899 -5 917
rect -39 883 -5 899
rect -39 831 -5 845
rect -39 811 -5 831
rect -39 763 -5 773
rect -39 739 -5 763
rect -39 695 -5 701
rect -39 667 -5 695
rect -39 627 -5 629
rect -39 595 -5 627
rect -39 525 -5 557
rect -39 523 -5 525
rect -39 457 -5 485
rect -39 451 -5 457
rect -39 389 -5 413
rect -39 379 -5 389
rect -39 321 -5 341
rect -39 307 -5 321
rect -39 253 -5 269
rect -39 235 -5 253
rect -39 185 -5 197
rect -39 163 -5 185
rect -39 117 -5 125
rect -39 91 -5 117
rect -39 49 -5 53
rect -39 19 -5 49
rect -39 -53 -5 -19
rect -39 -121 -5 -91
rect -39 -125 -5 -121
rect -39 -189 -5 -163
rect -39 -197 -5 -189
rect -39 -257 -5 -235
rect -39 -269 -5 -257
rect -39 -325 -5 -307
rect -39 -341 -5 -325
rect -39 -393 -5 -379
rect -39 -413 -5 -393
rect -39 -461 -5 -451
rect -39 -485 -5 -461
rect -39 -529 -5 -523
rect -39 -557 -5 -529
rect -39 -597 -5 -595
rect -39 -629 -5 -597
rect -39 -699 -5 -667
rect -39 -701 -5 -699
rect -39 -767 -5 -739
rect -39 -773 -5 -767
rect -39 -835 -5 -811
rect -39 -845 -5 -835
rect -39 -903 -5 -883
rect -39 -917 -5 -903
rect -39 -971 -5 -955
rect -39 -989 -5 -971
rect -39 -1039 -5 -1027
rect -39 -1061 -5 -1039
rect -39 -1107 -5 -1099
rect -39 -1133 -5 -1107
rect -39 -1175 -5 -1171
rect -39 -1205 -5 -1175
rect -39 -1277 -5 -1243
rect -39 -1345 -5 -1315
rect -39 -1349 -5 -1345
rect -39 -1413 -5 -1387
rect -39 -1421 -5 -1413
rect 230 1341 264 1349
rect 230 1315 264 1341
rect 230 1273 264 1277
rect 230 1243 264 1273
rect 230 1171 264 1205
rect 230 1103 264 1133
rect 230 1099 264 1103
rect 230 1035 264 1061
rect 230 1027 264 1035
rect 230 967 264 989
rect 230 955 264 967
rect 230 899 264 917
rect 230 883 264 899
rect 230 831 264 845
rect 230 811 264 831
rect 230 763 264 773
rect 230 739 264 763
rect 230 695 264 701
rect 230 667 264 695
rect 230 627 264 629
rect 230 595 264 627
rect 230 525 264 557
rect 230 523 264 525
rect 230 457 264 485
rect 230 451 264 457
rect 230 389 264 413
rect 230 379 264 389
rect 230 321 264 341
rect 230 307 264 321
rect 230 253 264 269
rect 230 235 264 253
rect 230 185 264 197
rect 230 163 264 185
rect 230 117 264 125
rect 230 91 264 117
rect 230 49 264 53
rect 230 19 264 49
rect 230 -53 264 -19
rect 230 -121 264 -91
rect 230 -125 264 -121
rect 230 -189 264 -163
rect 230 -197 264 -189
rect 230 -257 264 -235
rect 230 -269 264 -257
rect 230 -325 264 -307
rect 230 -341 264 -325
rect 230 -393 264 -379
rect 230 -413 264 -393
rect 230 -461 264 -451
rect 230 -485 264 -461
rect 230 -529 264 -523
rect 230 -557 264 -529
rect 230 -597 264 -595
rect 230 -629 264 -597
rect 230 -699 264 -667
rect 230 -701 264 -699
rect 230 -767 264 -739
rect 230 -773 264 -767
rect 230 -835 264 -811
rect 230 -845 264 -835
rect 230 -903 264 -883
rect 230 -917 264 -903
rect 230 -971 264 -955
rect 230 -989 264 -971
rect 230 -1039 264 -1027
rect 230 -1061 264 -1039
rect 230 -1107 264 -1099
rect 230 -1133 264 -1107
rect 230 -1175 264 -1171
rect 230 -1205 264 -1175
rect 230 -1277 264 -1243
rect 230 -1345 264 -1315
rect 230 -1349 264 -1345
rect 230 -1413 264 -1387
rect 230 -1421 264 -1413
<< metal1 >>
rect -247 1445 -55 1451
rect -247 1411 -204 1445
rect -170 1411 -132 1445
rect -98 1411 -55 1445
rect -247 1405 -55 1411
rect -303 1349 -257 1364
rect -303 1315 -297 1349
rect -263 1315 -257 1349
rect -303 1277 -257 1315
rect -303 1243 -297 1277
rect -263 1243 -257 1277
rect -303 1205 -257 1243
rect -303 1171 -297 1205
rect -263 1171 -257 1205
rect -303 1133 -257 1171
rect -303 1099 -297 1133
rect -263 1099 -257 1133
rect -303 1061 -257 1099
rect -303 1027 -297 1061
rect -263 1027 -257 1061
rect -303 989 -257 1027
rect -303 955 -297 989
rect -263 955 -257 989
rect -303 917 -257 955
rect -303 883 -297 917
rect -263 883 -257 917
rect -303 845 -257 883
rect -303 811 -297 845
rect -263 811 -257 845
rect -303 773 -257 811
rect -303 739 -297 773
rect -263 739 -257 773
rect -303 701 -257 739
rect -303 667 -297 701
rect -263 667 -257 701
rect -303 629 -257 667
rect -303 595 -297 629
rect -263 595 -257 629
rect -303 557 -257 595
rect -303 523 -297 557
rect -263 523 -257 557
rect -303 485 -257 523
rect -303 451 -297 485
rect -263 451 -257 485
rect -303 413 -257 451
rect -303 379 -297 413
rect -263 379 -257 413
rect -303 341 -257 379
rect -303 307 -297 341
rect -263 307 -257 341
rect -303 269 -257 307
rect -303 235 -297 269
rect -263 235 -257 269
rect -303 197 -257 235
rect -303 163 -297 197
rect -263 163 -257 197
rect -303 125 -257 163
rect -303 91 -297 125
rect -263 91 -257 125
rect -303 53 -257 91
rect -303 19 -297 53
rect -263 19 -257 53
rect -303 -19 -257 19
rect -303 -53 -297 -19
rect -263 -53 -257 -19
rect -303 -91 -257 -53
rect -303 -125 -297 -91
rect -263 -125 -257 -91
rect -303 -163 -257 -125
rect -303 -197 -297 -163
rect -263 -197 -257 -163
rect -303 -235 -257 -197
rect -303 -269 -297 -235
rect -263 -269 -257 -235
rect -303 -307 -257 -269
rect -303 -341 -297 -307
rect -263 -341 -257 -307
rect -303 -379 -257 -341
rect -303 -413 -297 -379
rect -263 -413 -257 -379
rect -303 -451 -257 -413
rect -303 -485 -297 -451
rect -263 -485 -257 -451
rect -303 -523 -257 -485
rect -303 -557 -297 -523
rect -263 -557 -257 -523
rect -303 -595 -257 -557
rect -303 -629 -297 -595
rect -263 -629 -257 -595
rect -303 -667 -257 -629
rect -303 -701 -297 -667
rect -263 -701 -257 -667
rect -303 -739 -257 -701
rect -303 -773 -297 -739
rect -263 -773 -257 -739
rect -303 -811 -257 -773
rect -303 -845 -297 -811
rect -263 -845 -257 -811
rect -303 -883 -257 -845
rect -303 -917 -297 -883
rect -263 -917 -257 -883
rect -303 -955 -257 -917
rect -303 -989 -297 -955
rect -263 -989 -257 -955
rect -303 -1027 -257 -989
rect -303 -1061 -297 -1027
rect -263 -1061 -257 -1027
rect -303 -1099 -257 -1061
rect -303 -1133 -297 -1099
rect -263 -1133 -257 -1099
rect -303 -1171 -257 -1133
rect -303 -1205 -297 -1171
rect -263 -1205 -257 -1171
rect -303 -1243 -257 -1205
rect -303 -1277 -297 -1243
rect -263 -1277 -257 -1243
rect -303 -1315 -257 -1277
rect -303 -1349 -297 -1315
rect -263 -1349 -257 -1315
rect -303 -1387 -257 -1349
rect -303 -1421 -297 -1387
rect -263 -1421 -257 -1387
rect -303 -1436 -257 -1421
rect -45 1349 1 1364
rect -45 1315 -39 1349
rect -5 1315 1 1349
rect -45 1277 1 1315
rect -45 1243 -39 1277
rect -5 1243 1 1277
rect -45 1205 1 1243
rect -45 1171 -39 1205
rect -5 1171 1 1205
rect -45 1133 1 1171
rect -45 1099 -39 1133
rect -5 1099 1 1133
rect -45 1061 1 1099
rect -45 1027 -39 1061
rect -5 1027 1 1061
rect -45 989 1 1027
rect -45 955 -39 989
rect -5 955 1 989
rect -45 917 1 955
rect -45 883 -39 917
rect -5 883 1 917
rect -45 845 1 883
rect -45 811 -39 845
rect -5 811 1 845
rect -45 773 1 811
rect -45 739 -39 773
rect -5 739 1 773
rect -45 701 1 739
rect -45 667 -39 701
rect -5 667 1 701
rect -45 629 1 667
rect -45 595 -39 629
rect -5 595 1 629
rect -45 557 1 595
rect -45 523 -39 557
rect -5 523 1 557
rect -45 485 1 523
rect -45 451 -39 485
rect -5 451 1 485
rect -45 413 1 451
rect -45 379 -39 413
rect -5 379 1 413
rect -45 341 1 379
rect -45 307 -39 341
rect -5 307 1 341
rect -45 269 1 307
rect -45 235 -39 269
rect -5 235 1 269
rect -45 197 1 235
rect -45 163 -39 197
rect -5 163 1 197
rect -45 125 1 163
rect -45 91 -39 125
rect -5 91 1 125
rect -45 53 1 91
rect -45 19 -39 53
rect -5 19 1 53
rect -45 -19 1 19
rect -45 -53 -39 -19
rect -5 -53 1 -19
rect -45 -91 1 -53
rect -45 -125 -39 -91
rect -5 -125 1 -91
rect -45 -163 1 -125
rect -45 -197 -39 -163
rect -5 -197 1 -163
rect -45 -235 1 -197
rect -45 -269 -39 -235
rect -5 -269 1 -235
rect -45 -307 1 -269
rect -45 -341 -39 -307
rect -5 -341 1 -307
rect -45 -379 1 -341
rect -45 -413 -39 -379
rect -5 -413 1 -379
rect -45 -451 1 -413
rect -45 -485 -39 -451
rect -5 -485 1 -451
rect -45 -523 1 -485
rect -45 -557 -39 -523
rect -5 -557 1 -523
rect -45 -595 1 -557
rect -45 -629 -39 -595
rect -5 -629 1 -595
rect -45 -667 1 -629
rect -45 -701 -39 -667
rect -5 -701 1 -667
rect -45 -739 1 -701
rect -45 -773 -39 -739
rect -5 -773 1 -739
rect -45 -811 1 -773
rect -45 -845 -39 -811
rect -5 -845 1 -811
rect -45 -883 1 -845
rect -45 -917 -39 -883
rect -5 -917 1 -883
rect -45 -955 1 -917
rect -45 -989 -39 -955
rect -5 -989 1 -955
rect -45 -1027 1 -989
rect -45 -1061 -39 -1027
rect -5 -1061 1 -1027
rect -45 -1099 1 -1061
rect -45 -1133 -39 -1099
rect -5 -1133 1 -1099
rect -45 -1171 1 -1133
rect -45 -1205 -39 -1171
rect -5 -1205 1 -1171
rect -45 -1243 1 -1205
rect -45 -1277 -39 -1243
rect -5 -1277 1 -1243
rect -45 -1315 1 -1277
rect -45 -1349 -39 -1315
rect -5 -1349 1 -1315
rect -45 -1387 1 -1349
rect -45 -1421 -39 -1387
rect -5 -1421 1 -1387
rect -45 -1436 1 -1421
rect 224 1349 270 1364
rect 224 1315 230 1349
rect 264 1315 270 1349
rect 224 1277 270 1315
rect 224 1243 230 1277
rect 264 1243 270 1277
rect 224 1205 270 1243
rect 224 1171 230 1205
rect 264 1171 270 1205
rect 224 1133 270 1171
rect 224 1099 230 1133
rect 264 1099 270 1133
rect 224 1061 270 1099
rect 224 1027 230 1061
rect 264 1027 270 1061
rect 224 989 270 1027
rect 224 955 230 989
rect 264 955 270 989
rect 224 917 270 955
rect 224 883 230 917
rect 264 883 270 917
rect 224 845 270 883
rect 224 811 230 845
rect 264 811 270 845
rect 224 773 270 811
rect 224 739 230 773
rect 264 739 270 773
rect 224 701 270 739
rect 224 667 230 701
rect 264 667 270 701
rect 224 629 270 667
rect 224 595 230 629
rect 264 595 270 629
rect 224 557 270 595
rect 224 523 230 557
rect 264 523 270 557
rect 224 485 270 523
rect 224 451 230 485
rect 264 451 270 485
rect 224 413 270 451
rect 224 379 230 413
rect 264 379 270 413
rect 224 341 270 379
rect 224 307 230 341
rect 264 307 270 341
rect 224 269 270 307
rect 224 235 230 269
rect 264 235 270 269
rect 224 197 270 235
rect 224 163 230 197
rect 264 163 270 197
rect 224 125 270 163
rect 224 91 230 125
rect 264 91 270 125
rect 224 53 270 91
rect 224 19 230 53
rect 264 19 270 53
rect 224 -19 270 19
rect 224 -53 230 -19
rect 264 -53 270 -19
rect 224 -91 270 -53
rect 224 -125 230 -91
rect 264 -125 270 -91
rect 224 -163 270 -125
rect 224 -197 230 -163
rect 264 -197 270 -163
rect 224 -235 270 -197
rect 224 -269 230 -235
rect 264 -269 270 -235
rect 224 -307 270 -269
rect 224 -341 230 -307
rect 264 -341 270 -307
rect 224 -379 270 -341
rect 224 -413 230 -379
rect 264 -413 270 -379
rect 224 -451 270 -413
rect 224 -485 230 -451
rect 264 -485 270 -451
rect 224 -523 270 -485
rect 224 -557 230 -523
rect 264 -557 270 -523
rect 224 -595 270 -557
rect 224 -629 230 -595
rect 264 -629 270 -595
rect 224 -667 270 -629
rect 224 -701 230 -667
rect 264 -701 270 -667
rect 224 -739 270 -701
rect 224 -773 230 -739
rect 264 -773 270 -739
rect 224 -811 270 -773
rect 224 -845 230 -811
rect 264 -845 270 -811
rect 224 -883 270 -845
rect 224 -917 230 -883
rect 264 -917 270 -883
rect 224 -955 270 -917
rect 224 -989 230 -955
rect 264 -989 270 -955
rect 224 -1027 270 -989
rect 224 -1061 230 -1027
rect 264 -1061 270 -1027
rect 224 -1099 270 -1061
rect 224 -1133 230 -1099
rect 264 -1133 270 -1099
rect 224 -1171 270 -1133
rect 224 -1205 230 -1171
rect 264 -1205 270 -1171
rect 224 -1243 270 -1205
rect 224 -1277 230 -1243
rect 264 -1277 270 -1243
rect 224 -1315 270 -1277
rect 224 -1349 230 -1315
rect 264 -1349 270 -1315
rect 224 -1387 270 -1349
rect 224 -1421 230 -1387
rect 264 -1421 270 -1387
rect 224 -1436 270 -1421
<< end >>
