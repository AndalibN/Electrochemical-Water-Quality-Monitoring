magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -2088 1892 -1089 1950
rect -2088 1828 -1173 1892
rect -1109 1828 -1089 1892
rect -2088 1812 -1089 1828
rect -2088 1748 -1173 1812
rect -1109 1748 -1089 1812
rect -2088 1732 -1089 1748
rect -2088 1668 -1173 1732
rect -1109 1668 -1089 1732
rect -2088 1652 -1089 1668
rect -2088 1588 -1173 1652
rect -1109 1588 -1089 1652
rect -2088 1572 -1089 1588
rect -2088 1508 -1173 1572
rect -1109 1508 -1089 1572
rect -2088 1492 -1089 1508
rect -2088 1428 -1173 1492
rect -1109 1428 -1089 1492
rect -2088 1412 -1089 1428
rect -2088 1348 -1173 1412
rect -1109 1348 -1089 1412
rect -2088 1332 -1089 1348
rect -2088 1268 -1173 1332
rect -1109 1268 -1089 1332
rect -2088 1252 -1089 1268
rect -2088 1188 -1173 1252
rect -1109 1188 -1089 1252
rect -2088 1172 -1089 1188
rect -2088 1108 -1173 1172
rect -1109 1108 -1089 1172
rect -2088 1050 -1089 1108
rect -1009 1892 -10 1950
rect -1009 1828 -94 1892
rect -30 1828 -10 1892
rect -1009 1812 -10 1828
rect -1009 1748 -94 1812
rect -30 1748 -10 1812
rect -1009 1732 -10 1748
rect -1009 1668 -94 1732
rect -30 1668 -10 1732
rect -1009 1652 -10 1668
rect -1009 1588 -94 1652
rect -30 1588 -10 1652
rect -1009 1572 -10 1588
rect -1009 1508 -94 1572
rect -30 1508 -10 1572
rect -1009 1492 -10 1508
rect -1009 1428 -94 1492
rect -30 1428 -10 1492
rect -1009 1412 -10 1428
rect -1009 1348 -94 1412
rect -30 1348 -10 1412
rect -1009 1332 -10 1348
rect -1009 1268 -94 1332
rect -30 1268 -10 1332
rect -1009 1252 -10 1268
rect -1009 1188 -94 1252
rect -30 1188 -10 1252
rect -1009 1172 -10 1188
rect -1009 1108 -94 1172
rect -30 1108 -10 1172
rect -1009 1050 -10 1108
rect 74 1892 1073 1950
rect 74 1828 989 1892
rect 1053 1828 1073 1892
rect 74 1812 1073 1828
rect 74 1748 989 1812
rect 1053 1748 1073 1812
rect 74 1732 1073 1748
rect 74 1668 989 1732
rect 1053 1668 1073 1732
rect 74 1652 1073 1668
rect 74 1588 989 1652
rect 1053 1588 1073 1652
rect 74 1572 1073 1588
rect 74 1508 989 1572
rect 1053 1508 1073 1572
rect 74 1492 1073 1508
rect 74 1428 989 1492
rect 1053 1428 1073 1492
rect 74 1412 1073 1428
rect 74 1348 989 1412
rect 1053 1348 1073 1412
rect 74 1332 1073 1348
rect 74 1268 989 1332
rect 1053 1268 1073 1332
rect 74 1252 1073 1268
rect 74 1188 989 1252
rect 1053 1188 1073 1252
rect 74 1172 1073 1188
rect 74 1108 989 1172
rect 1053 1108 1073 1172
rect 74 1050 1073 1108
rect 1153 1892 2152 1950
rect 1153 1828 2068 1892
rect 2132 1828 2152 1892
rect 1153 1812 2152 1828
rect 1153 1748 2068 1812
rect 2132 1748 2152 1812
rect 1153 1732 2152 1748
rect 1153 1668 2068 1732
rect 2132 1668 2152 1732
rect 1153 1652 2152 1668
rect 1153 1588 2068 1652
rect 2132 1588 2152 1652
rect 1153 1572 2152 1588
rect 1153 1508 2068 1572
rect 2132 1508 2152 1572
rect 1153 1492 2152 1508
rect 1153 1428 2068 1492
rect 2132 1428 2152 1492
rect 1153 1412 2152 1428
rect 1153 1348 2068 1412
rect 2132 1348 2152 1412
rect 1153 1332 2152 1348
rect 1153 1268 2068 1332
rect 2132 1268 2152 1332
rect 1153 1252 2152 1268
rect 1153 1188 2068 1252
rect 2132 1188 2152 1252
rect 1153 1172 2152 1188
rect 1153 1108 2068 1172
rect 2132 1108 2152 1172
rect 1153 1050 2152 1108
rect -2088 892 -1089 950
rect -2088 828 -1173 892
rect -1109 828 -1089 892
rect -2088 812 -1089 828
rect -2088 748 -1173 812
rect -1109 748 -1089 812
rect -2088 732 -1089 748
rect -2088 668 -1173 732
rect -1109 668 -1089 732
rect -2088 652 -1089 668
rect -2088 588 -1173 652
rect -1109 588 -1089 652
rect -2088 572 -1089 588
rect -2088 508 -1173 572
rect -1109 508 -1089 572
rect -2088 492 -1089 508
rect -2088 428 -1173 492
rect -1109 428 -1089 492
rect -2088 412 -1089 428
rect -2088 348 -1173 412
rect -1109 348 -1089 412
rect -2088 332 -1089 348
rect -2088 268 -1173 332
rect -1109 268 -1089 332
rect -2088 252 -1089 268
rect -2088 188 -1173 252
rect -1109 188 -1089 252
rect -2088 172 -1089 188
rect -2088 108 -1173 172
rect -1109 108 -1089 172
rect -2088 50 -1089 108
rect -1009 892 -10 950
rect -1009 828 -94 892
rect -30 828 -10 892
rect -1009 812 -10 828
rect -1009 748 -94 812
rect -30 748 -10 812
rect -1009 732 -10 748
rect -1009 668 -94 732
rect -30 668 -10 732
rect -1009 652 -10 668
rect -1009 588 -94 652
rect -30 588 -10 652
rect -1009 572 -10 588
rect -1009 508 -94 572
rect -30 508 -10 572
rect -1009 492 -10 508
rect -1009 428 -94 492
rect -30 428 -10 492
rect -1009 412 -10 428
rect -1009 348 -94 412
rect -30 348 -10 412
rect -1009 332 -10 348
rect -1009 268 -94 332
rect -30 268 -10 332
rect -1009 252 -10 268
rect -1009 188 -94 252
rect -30 188 -10 252
rect -1009 172 -10 188
rect -1009 108 -94 172
rect -30 108 -10 172
rect -1009 50 -10 108
rect 74 892 1073 950
rect 74 828 989 892
rect 1053 828 1073 892
rect 74 812 1073 828
rect 74 748 989 812
rect 1053 748 1073 812
rect 74 732 1073 748
rect 74 668 989 732
rect 1053 668 1073 732
rect 74 652 1073 668
rect 74 588 989 652
rect 1053 588 1073 652
rect 74 572 1073 588
rect 74 508 989 572
rect 1053 508 1073 572
rect 74 492 1073 508
rect 74 428 989 492
rect 1053 428 1073 492
rect 74 412 1073 428
rect 74 348 989 412
rect 1053 348 1073 412
rect 74 332 1073 348
rect 74 268 989 332
rect 1053 268 1073 332
rect 74 252 1073 268
rect 74 188 989 252
rect 1053 188 1073 252
rect 74 172 1073 188
rect 74 108 989 172
rect 1053 108 1073 172
rect 74 50 1073 108
rect 1153 892 2152 950
rect 1153 828 2068 892
rect 2132 828 2152 892
rect 1153 812 2152 828
rect 1153 748 2068 812
rect 2132 748 2152 812
rect 1153 732 2152 748
rect 1153 668 2068 732
rect 2132 668 2152 732
rect 1153 652 2152 668
rect 1153 588 2068 652
rect 2132 588 2152 652
rect 1153 572 2152 588
rect 1153 508 2068 572
rect 2132 508 2152 572
rect 1153 492 2152 508
rect 1153 428 2068 492
rect 2132 428 2152 492
rect 1153 412 2152 428
rect 1153 348 2068 412
rect 2132 348 2152 412
rect 1153 332 2152 348
rect 1153 268 2068 332
rect 2132 268 2152 332
rect 1153 252 2152 268
rect 1153 188 2068 252
rect 2132 188 2152 252
rect 1153 172 2152 188
rect 1153 108 2068 172
rect 2132 108 2152 172
rect 1153 50 2152 108
rect -2088 -108 -1089 -50
rect -2088 -172 -1173 -108
rect -1109 -172 -1089 -108
rect -2088 -188 -1089 -172
rect -2088 -252 -1173 -188
rect -1109 -252 -1089 -188
rect -2088 -268 -1089 -252
rect -2088 -332 -1173 -268
rect -1109 -332 -1089 -268
rect -2088 -348 -1089 -332
rect -2088 -412 -1173 -348
rect -1109 -412 -1089 -348
rect -2088 -428 -1089 -412
rect -2088 -492 -1173 -428
rect -1109 -492 -1089 -428
rect -2088 -508 -1089 -492
rect -2088 -572 -1173 -508
rect -1109 -572 -1089 -508
rect -2088 -588 -1089 -572
rect -2088 -652 -1173 -588
rect -1109 -652 -1089 -588
rect -2088 -668 -1089 -652
rect -2088 -732 -1173 -668
rect -1109 -732 -1089 -668
rect -2088 -748 -1089 -732
rect -2088 -812 -1173 -748
rect -1109 -812 -1089 -748
rect -2088 -828 -1089 -812
rect -2088 -892 -1173 -828
rect -1109 -892 -1089 -828
rect -2088 -950 -1089 -892
rect -1009 -108 -10 -50
rect -1009 -172 -94 -108
rect -30 -172 -10 -108
rect -1009 -188 -10 -172
rect -1009 -252 -94 -188
rect -30 -252 -10 -188
rect -1009 -268 -10 -252
rect -1009 -332 -94 -268
rect -30 -332 -10 -268
rect -1009 -348 -10 -332
rect -1009 -412 -94 -348
rect -30 -412 -10 -348
rect -1009 -428 -10 -412
rect -1009 -492 -94 -428
rect -30 -492 -10 -428
rect -1009 -508 -10 -492
rect -1009 -572 -94 -508
rect -30 -572 -10 -508
rect -1009 -588 -10 -572
rect -1009 -652 -94 -588
rect -30 -652 -10 -588
rect -1009 -668 -10 -652
rect -1009 -732 -94 -668
rect -30 -732 -10 -668
rect -1009 -748 -10 -732
rect -1009 -812 -94 -748
rect -30 -812 -10 -748
rect -1009 -828 -10 -812
rect -1009 -892 -94 -828
rect -30 -892 -10 -828
rect -1009 -950 -10 -892
rect 74 -108 1073 -50
rect 74 -172 989 -108
rect 1053 -172 1073 -108
rect 74 -188 1073 -172
rect 74 -252 989 -188
rect 1053 -252 1073 -188
rect 74 -268 1073 -252
rect 74 -332 989 -268
rect 1053 -332 1073 -268
rect 74 -348 1073 -332
rect 74 -412 989 -348
rect 1053 -412 1073 -348
rect 74 -428 1073 -412
rect 74 -492 989 -428
rect 1053 -492 1073 -428
rect 74 -508 1073 -492
rect 74 -572 989 -508
rect 1053 -572 1073 -508
rect 74 -588 1073 -572
rect 74 -652 989 -588
rect 1053 -652 1073 -588
rect 74 -668 1073 -652
rect 74 -732 989 -668
rect 1053 -732 1073 -668
rect 74 -748 1073 -732
rect 74 -812 989 -748
rect 1053 -812 1073 -748
rect 74 -828 1073 -812
rect 74 -892 989 -828
rect 1053 -892 1073 -828
rect 74 -950 1073 -892
rect 1153 -108 2152 -50
rect 1153 -172 2068 -108
rect 2132 -172 2152 -108
rect 1153 -188 2152 -172
rect 1153 -252 2068 -188
rect 2132 -252 2152 -188
rect 1153 -268 2152 -252
rect 1153 -332 2068 -268
rect 2132 -332 2152 -268
rect 1153 -348 2152 -332
rect 1153 -412 2068 -348
rect 2132 -412 2152 -348
rect 1153 -428 2152 -412
rect 1153 -492 2068 -428
rect 2132 -492 2152 -428
rect 1153 -508 2152 -492
rect 1153 -572 2068 -508
rect 2132 -572 2152 -508
rect 1153 -588 2152 -572
rect 1153 -652 2068 -588
rect 2132 -652 2152 -588
rect 1153 -668 2152 -652
rect 1153 -732 2068 -668
rect 2132 -732 2152 -668
rect 1153 -748 2152 -732
rect 1153 -812 2068 -748
rect 2132 -812 2152 -748
rect 1153 -828 2152 -812
rect 1153 -892 2068 -828
rect 2132 -892 2152 -828
rect 1153 -950 2152 -892
rect -2088 -1108 -1089 -1050
rect -2088 -1172 -1173 -1108
rect -1109 -1172 -1089 -1108
rect -2088 -1188 -1089 -1172
rect -2088 -1252 -1173 -1188
rect -1109 -1252 -1089 -1188
rect -2088 -1268 -1089 -1252
rect -2088 -1332 -1173 -1268
rect -1109 -1332 -1089 -1268
rect -2088 -1348 -1089 -1332
rect -2088 -1412 -1173 -1348
rect -1109 -1412 -1089 -1348
rect -2088 -1428 -1089 -1412
rect -2088 -1492 -1173 -1428
rect -1109 -1492 -1089 -1428
rect -2088 -1508 -1089 -1492
rect -2088 -1572 -1173 -1508
rect -1109 -1572 -1089 -1508
rect -2088 -1588 -1089 -1572
rect -2088 -1652 -1173 -1588
rect -1109 -1652 -1089 -1588
rect -2088 -1668 -1089 -1652
rect -2088 -1732 -1173 -1668
rect -1109 -1732 -1089 -1668
rect -2088 -1748 -1089 -1732
rect -2088 -1812 -1173 -1748
rect -1109 -1812 -1089 -1748
rect -2088 -1828 -1089 -1812
rect -2088 -1892 -1173 -1828
rect -1109 -1892 -1089 -1828
rect -2088 -1950 -1089 -1892
rect -1009 -1108 -10 -1050
rect -1009 -1172 -94 -1108
rect -30 -1172 -10 -1108
rect -1009 -1188 -10 -1172
rect -1009 -1252 -94 -1188
rect -30 -1252 -10 -1188
rect -1009 -1268 -10 -1252
rect -1009 -1332 -94 -1268
rect -30 -1332 -10 -1268
rect -1009 -1348 -10 -1332
rect -1009 -1412 -94 -1348
rect -30 -1412 -10 -1348
rect -1009 -1428 -10 -1412
rect -1009 -1492 -94 -1428
rect -30 -1492 -10 -1428
rect -1009 -1508 -10 -1492
rect -1009 -1572 -94 -1508
rect -30 -1572 -10 -1508
rect -1009 -1588 -10 -1572
rect -1009 -1652 -94 -1588
rect -30 -1652 -10 -1588
rect -1009 -1668 -10 -1652
rect -1009 -1732 -94 -1668
rect -30 -1732 -10 -1668
rect -1009 -1748 -10 -1732
rect -1009 -1812 -94 -1748
rect -30 -1812 -10 -1748
rect -1009 -1828 -10 -1812
rect -1009 -1892 -94 -1828
rect -30 -1892 -10 -1828
rect -1009 -1950 -10 -1892
rect 74 -1108 1073 -1050
rect 74 -1172 989 -1108
rect 1053 -1172 1073 -1108
rect 74 -1188 1073 -1172
rect 74 -1252 989 -1188
rect 1053 -1252 1073 -1188
rect 74 -1268 1073 -1252
rect 74 -1332 989 -1268
rect 1053 -1332 1073 -1268
rect 74 -1348 1073 -1332
rect 74 -1412 989 -1348
rect 1053 -1412 1073 -1348
rect 74 -1428 1073 -1412
rect 74 -1492 989 -1428
rect 1053 -1492 1073 -1428
rect 74 -1508 1073 -1492
rect 74 -1572 989 -1508
rect 1053 -1572 1073 -1508
rect 74 -1588 1073 -1572
rect 74 -1652 989 -1588
rect 1053 -1652 1073 -1588
rect 74 -1668 1073 -1652
rect 74 -1732 989 -1668
rect 1053 -1732 1073 -1668
rect 74 -1748 1073 -1732
rect 74 -1812 989 -1748
rect 1053 -1812 1073 -1748
rect 74 -1828 1073 -1812
rect 74 -1892 989 -1828
rect 1053 -1892 1073 -1828
rect 74 -1949 1073 -1892
rect 1153 -1108 2152 -1050
rect 1153 -1172 2068 -1108
rect 2132 -1172 2152 -1108
rect 1153 -1188 2152 -1172
rect 1153 -1252 2068 -1188
rect 2132 -1252 2152 -1188
rect 1153 -1268 2152 -1252
rect 1153 -1332 2068 -1268
rect 2132 -1332 2152 -1268
rect 1153 -1348 2152 -1332
rect 1153 -1412 2068 -1348
rect 2132 -1412 2152 -1348
rect 1153 -1428 2152 -1412
rect 1153 -1492 2068 -1428
rect 2132 -1492 2152 -1428
rect 1153 -1508 2152 -1492
rect 1153 -1572 2068 -1508
rect 2132 -1572 2152 -1508
rect 1153 -1588 2152 -1572
rect 1153 -1652 2068 -1588
rect 2132 -1652 2152 -1588
rect 1153 -1668 2152 -1652
rect 1153 -1732 2068 -1668
rect 2132 -1732 2152 -1668
rect 1153 -1748 2152 -1732
rect 1153 -1812 2068 -1748
rect 2132 -1812 2152 -1748
rect 1153 -1828 2152 -1812
rect 1153 -1892 2068 -1828
rect 2132 -1892 2152 -1828
rect 1153 -1950 2152 -1892
<< via3 >>
rect -1173 1828 -1109 1892
rect -1173 1748 -1109 1812
rect -1173 1668 -1109 1732
rect -1173 1588 -1109 1652
rect -1173 1508 -1109 1572
rect -1173 1428 -1109 1492
rect -1173 1348 -1109 1412
rect -1173 1268 -1109 1332
rect -1173 1188 -1109 1252
rect -1173 1108 -1109 1172
rect -94 1828 -30 1892
rect -94 1748 -30 1812
rect -94 1668 -30 1732
rect -94 1588 -30 1652
rect -94 1508 -30 1572
rect -94 1428 -30 1492
rect -94 1348 -30 1412
rect -94 1268 -30 1332
rect -94 1188 -30 1252
rect -94 1108 -30 1172
rect 989 1828 1053 1892
rect 989 1748 1053 1812
rect 989 1668 1053 1732
rect 989 1588 1053 1652
rect 989 1508 1053 1572
rect 989 1428 1053 1492
rect 989 1348 1053 1412
rect 989 1268 1053 1332
rect 989 1188 1053 1252
rect 989 1108 1053 1172
rect 2068 1828 2132 1892
rect 2068 1748 2132 1812
rect 2068 1668 2132 1732
rect 2068 1588 2132 1652
rect 2068 1508 2132 1572
rect 2068 1428 2132 1492
rect 2068 1348 2132 1412
rect 2068 1268 2132 1332
rect 2068 1188 2132 1252
rect 2068 1108 2132 1172
rect -1173 828 -1109 892
rect -1173 748 -1109 812
rect -1173 668 -1109 732
rect -1173 588 -1109 652
rect -1173 508 -1109 572
rect -1173 428 -1109 492
rect -1173 348 -1109 412
rect -1173 268 -1109 332
rect -1173 188 -1109 252
rect -1173 108 -1109 172
rect -94 828 -30 892
rect -94 748 -30 812
rect -94 668 -30 732
rect -94 588 -30 652
rect -94 508 -30 572
rect -94 428 -30 492
rect -94 348 -30 412
rect -94 268 -30 332
rect -94 188 -30 252
rect -94 108 -30 172
rect 989 828 1053 892
rect 989 748 1053 812
rect 989 668 1053 732
rect 989 588 1053 652
rect 989 508 1053 572
rect 989 428 1053 492
rect 989 348 1053 412
rect 989 268 1053 332
rect 989 188 1053 252
rect 989 108 1053 172
rect 2068 828 2132 892
rect 2068 748 2132 812
rect 2068 668 2132 732
rect 2068 588 2132 652
rect 2068 508 2132 572
rect 2068 428 2132 492
rect 2068 348 2132 412
rect 2068 268 2132 332
rect 2068 188 2132 252
rect 2068 108 2132 172
rect -1173 -172 -1109 -108
rect -1173 -252 -1109 -188
rect -1173 -332 -1109 -268
rect -1173 -412 -1109 -348
rect -1173 -492 -1109 -428
rect -1173 -572 -1109 -508
rect -1173 -652 -1109 -588
rect -1173 -732 -1109 -668
rect -1173 -812 -1109 -748
rect -1173 -892 -1109 -828
rect -94 -172 -30 -108
rect -94 -252 -30 -188
rect -94 -332 -30 -268
rect -94 -412 -30 -348
rect -94 -492 -30 -428
rect -94 -572 -30 -508
rect -94 -652 -30 -588
rect -94 -732 -30 -668
rect -94 -812 -30 -748
rect -94 -892 -30 -828
rect 989 -172 1053 -108
rect 989 -252 1053 -188
rect 989 -332 1053 -268
rect 989 -412 1053 -348
rect 989 -492 1053 -428
rect 989 -572 1053 -508
rect 989 -652 1053 -588
rect 989 -732 1053 -668
rect 989 -812 1053 -748
rect 989 -892 1053 -828
rect 2068 -172 2132 -108
rect 2068 -252 2132 -188
rect 2068 -332 2132 -268
rect 2068 -412 2132 -348
rect 2068 -492 2132 -428
rect 2068 -572 2132 -508
rect 2068 -652 2132 -588
rect 2068 -732 2132 -668
rect 2068 -812 2132 -748
rect 2068 -892 2132 -828
rect -1173 -1172 -1109 -1108
rect -1173 -1252 -1109 -1188
rect -1173 -1332 -1109 -1268
rect -1173 -1412 -1109 -1348
rect -1173 -1492 -1109 -1428
rect -1173 -1572 -1109 -1508
rect -1173 -1652 -1109 -1588
rect -1173 -1732 -1109 -1668
rect -1173 -1812 -1109 -1748
rect -1173 -1892 -1109 -1828
rect -94 -1172 -30 -1108
rect -94 -1252 -30 -1188
rect -94 -1332 -30 -1268
rect -94 -1412 -30 -1348
rect -94 -1492 -30 -1428
rect -94 -1572 -30 -1508
rect -94 -1652 -30 -1588
rect -94 -1732 -30 -1668
rect -94 -1812 -30 -1748
rect -94 -1892 -30 -1828
rect 989 -1172 1053 -1108
rect 989 -1252 1053 -1188
rect 989 -1332 1053 -1268
rect 989 -1412 1053 -1348
rect 989 -1492 1053 -1428
rect 989 -1572 1053 -1508
rect 989 -1652 1053 -1588
rect 989 -1732 1053 -1668
rect 989 -1812 1053 -1748
rect 989 -1892 1053 -1828
rect 2068 -1172 2132 -1108
rect 2068 -1252 2132 -1188
rect 2068 -1332 2132 -1268
rect 2068 -1412 2132 -1348
rect 2068 -1492 2132 -1428
rect 2068 -1572 2132 -1508
rect 2068 -1652 2132 -1588
rect 2068 -1732 2132 -1668
rect 2068 -1812 2132 -1748
rect 2068 -1892 2132 -1828
<< mimcap >>
rect -1988 1772 -1288 1850
rect -1988 1228 -1910 1772
rect -1366 1228 -1288 1772
rect -1988 1150 -1288 1228
rect -909 1772 -209 1850
rect -909 1228 -831 1772
rect -287 1228 -209 1772
rect -909 1150 -209 1228
rect 174 1772 874 1850
rect 174 1228 252 1772
rect 796 1228 874 1772
rect 174 1150 874 1228
rect 1253 1772 1953 1850
rect 1253 1228 1331 1772
rect 1875 1228 1953 1772
rect 1253 1150 1953 1228
rect -1988 772 -1288 850
rect -1988 228 -1910 772
rect -1366 228 -1288 772
rect -1988 150 -1288 228
rect -909 772 -209 850
rect -909 228 -831 772
rect -287 228 -209 772
rect -909 150 -209 228
rect 174 772 874 850
rect 174 228 252 772
rect 796 228 874 772
rect 174 150 874 228
rect 1253 772 1953 850
rect 1253 228 1331 772
rect 1875 228 1953 772
rect 1253 150 1953 228
rect -1988 -228 -1288 -150
rect -1988 -772 -1910 -228
rect -1366 -772 -1288 -228
rect -1988 -850 -1288 -772
rect -909 -228 -209 -150
rect -909 -772 -831 -228
rect -287 -772 -209 -228
rect -909 -850 -209 -772
rect 174 -228 874 -150
rect 174 -772 252 -228
rect 796 -772 874 -228
rect 174 -850 874 -772
rect 1253 -228 1953 -150
rect 1253 -772 1331 -228
rect 1875 -772 1953 -228
rect 1253 -850 1953 -772
rect -1988 -1228 -1288 -1150
rect -1988 -1772 -1910 -1228
rect -1366 -1772 -1288 -1228
rect -1988 -1850 -1288 -1772
rect -909 -1228 -209 -1150
rect -909 -1772 -831 -1228
rect -287 -1772 -209 -1228
rect -909 -1850 -209 -1772
rect 174 -1228 874 -1150
rect 174 -1772 252 -1228
rect 796 -1772 874 -1228
rect 174 -1850 874 -1772
rect 1253 -1228 1953 -1150
rect 1253 -1772 1331 -1228
rect 1875 -1772 1953 -1228
rect 1253 -1850 1953 -1772
<< mimcapcontact >>
rect -1910 1228 -1366 1772
rect -831 1228 -287 1772
rect 252 1228 796 1772
rect 1331 1228 1875 1772
rect -1910 228 -1366 772
rect -831 228 -287 772
rect 252 228 796 772
rect 1331 228 1875 772
rect -1910 -772 -1366 -228
rect -831 -772 -287 -228
rect 252 -772 796 -228
rect 1331 -772 1875 -228
rect -1910 -1772 -1366 -1228
rect -831 -1772 -287 -1228
rect 252 -1772 796 -1228
rect 1331 -1772 1875 -1228
<< metal4 >>
rect -1949 1772 -1327 2000
rect -1949 1228 -1910 1772
rect -1366 1228 -1327 1772
rect -1949 772 -1327 1228
rect -1949 228 -1910 772
rect -1366 228 -1327 772
rect -1949 189 -1327 228
rect -1220 1892 -1093 2249
rect -1220 1828 -1173 1892
rect -1109 1828 -1093 1892
rect -1220 1812 -1093 1828
rect -1220 1748 -1173 1812
rect -1109 1748 -1093 1812
rect -1220 1732 -1093 1748
rect -1220 1668 -1173 1732
rect -1109 1668 -1093 1732
rect -1220 1652 -1093 1668
rect -1220 1588 -1173 1652
rect -1109 1588 -1093 1652
rect -1220 1572 -1093 1588
rect -1220 1508 -1173 1572
rect -1109 1508 -1093 1572
rect -1220 1492 -1093 1508
rect -1220 1428 -1173 1492
rect -1109 1428 -1093 1492
rect -1220 1412 -1093 1428
rect -1220 1348 -1173 1412
rect -1109 1348 -1093 1412
rect -1220 1332 -1093 1348
rect -1220 1268 -1173 1332
rect -1109 1268 -1093 1332
rect -1220 1252 -1093 1268
rect -1220 1188 -1173 1252
rect -1109 1188 -1093 1252
rect -1220 1172 -1093 1188
rect -1220 1108 -1173 1172
rect -1109 1108 -1093 1172
rect -1220 1062 -1093 1108
rect -870 1811 -249 2000
rect -141 1892 -14 2249
rect -141 1828 -94 1892
rect -30 1828 -14 1892
rect -141 1812 -14 1828
rect -870 1772 -248 1811
rect -870 1228 -831 1772
rect -287 1228 -248 1772
rect -1220 938 -1116 1062
rect -1220 892 -1093 938
rect -1220 828 -1173 892
rect -1109 828 -1093 892
rect -1220 812 -1093 828
rect -1220 748 -1173 812
rect -1109 748 -1093 812
rect -1220 732 -1093 748
rect -1220 668 -1173 732
rect -1109 668 -1093 732
rect -1220 652 -1093 668
rect -1220 588 -1173 652
rect -1109 588 -1093 652
rect -1220 572 -1093 588
rect -1220 508 -1173 572
rect -1109 508 -1093 572
rect -1220 492 -1093 508
rect -1220 428 -1173 492
rect -1109 428 -1093 492
rect -1220 412 -1093 428
rect -1220 348 -1173 412
rect -1109 348 -1093 412
rect -1220 332 -1093 348
rect -1220 268 -1173 332
rect -1109 268 -1093 332
rect -1220 252 -1093 268
rect -1946 -189 -1331 189
rect -1220 188 -1173 252
rect -1109 188 -1093 252
rect -870 772 -248 1228
rect -870 228 -831 772
rect -287 228 -248 772
rect -870 189 -248 228
rect -141 1748 -94 1812
rect -30 1748 -14 1812
rect -141 1732 -14 1748
rect -141 1668 -94 1732
rect -30 1668 -14 1732
rect -141 1652 -14 1668
rect -141 1588 -94 1652
rect -30 1588 -14 1652
rect -141 1572 -14 1588
rect -141 1508 -94 1572
rect -30 1508 -14 1572
rect -141 1492 -14 1508
rect -141 1428 -94 1492
rect -30 1428 -14 1492
rect -141 1412 -14 1428
rect -141 1348 -94 1412
rect -30 1348 -14 1412
rect -141 1332 -14 1348
rect -141 1268 -94 1332
rect -30 1268 -14 1332
rect -141 1252 -14 1268
rect -141 1188 -94 1252
rect -30 1188 -14 1252
rect -141 1172 -14 1188
rect -141 1108 -94 1172
rect -30 1108 -14 1172
rect -141 1062 -14 1108
rect 213 1772 835 2000
rect 213 1228 252 1772
rect 796 1228 835 1772
rect -141 938 -37 1062
rect -141 892 -14 938
rect -141 828 -94 892
rect -30 828 -14 892
rect -141 812 -14 828
rect -141 748 -94 812
rect -30 748 -14 812
rect -141 732 -14 748
rect -141 668 -94 732
rect -30 668 -14 732
rect -141 652 -14 668
rect -141 588 -94 652
rect -30 588 -14 652
rect -141 572 -14 588
rect -141 508 -94 572
rect -30 508 -14 572
rect -141 492 -14 508
rect -141 428 -94 492
rect -30 428 -14 492
rect -141 412 -14 428
rect -141 348 -94 412
rect -30 348 -14 412
rect -141 332 -14 348
rect -141 268 -94 332
rect -30 268 -14 332
rect -141 252 -14 268
rect -1220 172 -1093 188
rect -1220 108 -1173 172
rect -1109 108 -1093 172
rect -1220 62 -1093 108
rect -1220 -62 -1116 62
rect -1220 -108 -1093 -62
rect -1220 -172 -1173 -108
rect -1109 -172 -1093 -108
rect -1220 -188 -1093 -172
rect -1949 -228 -1327 -189
rect -1949 -772 -1910 -228
rect -1366 -772 -1327 -228
rect -1949 -811 -1327 -772
rect -1220 -252 -1173 -188
rect -1109 -252 -1093 -188
rect -864 -189 -252 189
rect -141 188 -94 252
rect -30 188 -14 252
rect -141 172 -14 188
rect -141 108 -94 172
rect -30 108 -14 172
rect -141 62 -14 108
rect 213 772 835 1228
rect 213 228 252 772
rect 796 228 835 772
rect -141 -62 -37 62
rect -141 -108 -14 -62
rect -141 -172 -94 -108
rect -30 -172 -14 -108
rect -141 -188 -14 -172
rect -1220 -268 -1093 -252
rect -1220 -332 -1173 -268
rect -1109 -332 -1093 -268
rect -1220 -348 -1093 -332
rect -1220 -412 -1173 -348
rect -1109 -412 -1093 -348
rect -1220 -428 -1093 -412
rect -1220 -492 -1173 -428
rect -1109 -492 -1093 -428
rect -1220 -508 -1093 -492
rect -1220 -572 -1173 -508
rect -1109 -572 -1093 -508
rect -1220 -588 -1093 -572
rect -1220 -652 -1173 -588
rect -1109 -652 -1093 -588
rect -1220 -668 -1093 -652
rect -1220 -732 -1173 -668
rect -1109 -732 -1093 -668
rect -1220 -748 -1093 -732
rect -1940 -1189 -1337 -811
rect -1220 -812 -1173 -748
rect -1109 -812 -1093 -748
rect -1220 -828 -1093 -812
rect -1220 -892 -1173 -828
rect -1109 -892 -1093 -828
rect -1220 -1108 -1093 -892
rect -1220 -1172 -1173 -1108
rect -1109 -1172 -1093 -1108
rect -1220 -1188 -1093 -1172
rect -1949 -1228 -1327 -1189
rect -1949 -1772 -1910 -1228
rect -1366 -1772 -1327 -1228
rect -1949 -1811 -1327 -1772
rect -1220 -1252 -1173 -1188
rect -1109 -1252 -1093 -1188
rect -1220 -1268 -1093 -1252
rect -1220 -1332 -1173 -1268
rect -1109 -1332 -1093 -1268
rect -1220 -1348 -1093 -1332
rect -1220 -1412 -1173 -1348
rect -1109 -1412 -1093 -1348
rect -1220 -1428 -1093 -1412
rect -1220 -1492 -1173 -1428
rect -1109 -1492 -1093 -1428
rect -1220 -1508 -1093 -1492
rect -1220 -1572 -1173 -1508
rect -1109 -1572 -1093 -1508
rect -1220 -1588 -1093 -1572
rect -1220 -1652 -1173 -1588
rect -1109 -1652 -1093 -1588
rect -1220 -1668 -1093 -1652
rect -1220 -1732 -1173 -1668
rect -1109 -1732 -1093 -1668
rect -1220 -1748 -1093 -1732
rect -1949 -2288 -1348 -1811
rect -1220 -1812 -1173 -1748
rect -1109 -1812 -1093 -1748
rect -870 -228 -248 -189
rect -870 -772 -831 -228
rect -287 -772 -248 -228
rect -870 -1228 -248 -772
rect -870 -1772 -831 -1228
rect -287 -1772 -248 -1228
rect -870 -1811 -248 -1772
rect -1220 -1828 -1093 -1812
rect -1220 -1892 -1173 -1828
rect -1109 -1892 -1093 -1828
rect -1220 -1938 -1093 -1892
rect -860 -2202 -248 -1811
rect -141 -252 -94 -188
rect -30 -252 -14 -188
rect -141 -268 -14 -252
rect -141 -332 -94 -268
rect -30 -332 -14 -268
rect -141 -348 -14 -332
rect -141 -412 -94 -348
rect -30 -412 -14 -348
rect -141 -428 -14 -412
rect -141 -492 -94 -428
rect -30 -492 -14 -428
rect -141 -508 -14 -492
rect -141 -572 -94 -508
rect -30 -572 -14 -508
rect -141 -588 -14 -572
rect -141 -652 -94 -588
rect -30 -652 -14 -588
rect -141 -668 -14 -652
rect -141 -732 -94 -668
rect -30 -732 -14 -668
rect -141 -748 -14 -732
rect -141 -812 -94 -748
rect -30 -812 -14 -748
rect -141 -828 -14 -812
rect -141 -892 -94 -828
rect -30 -892 -14 -828
rect -141 -1108 -14 -892
rect -141 -1172 -94 -1108
rect -30 -1172 -14 -1108
rect -141 -1188 -14 -1172
rect -141 -1252 -94 -1188
rect -30 -1252 -14 -1188
rect -141 -1268 -14 -1252
rect -141 -1332 -94 -1268
rect -30 -1332 -14 -1268
rect -141 -1348 -14 -1332
rect -141 -1412 -94 -1348
rect -30 -1412 -14 -1348
rect -141 -1428 -14 -1412
rect -141 -1492 -94 -1428
rect -30 -1492 -14 -1428
rect -141 -1508 -14 -1492
rect -141 -1572 -94 -1508
rect -30 -1572 -14 -1508
rect -141 -1588 -14 -1572
rect -141 -1652 -94 -1588
rect -30 -1652 -14 -1588
rect -141 -1668 -14 -1652
rect -141 -1732 -94 -1668
rect -30 -1732 -14 -1668
rect -141 -1748 -14 -1732
rect -141 -1812 -94 -1748
rect -30 -1812 -14 -1748
rect 213 -228 835 228
rect 213 -772 252 -228
rect 796 -772 835 -228
rect 213 -1228 835 -772
rect 213 -1772 252 -1228
rect 796 -1772 835 -1228
rect 213 -1811 835 -1772
rect 942 1892 1069 2249
rect 942 1828 989 1892
rect 1053 1828 1069 1892
rect 942 1812 1069 1828
rect 942 1748 989 1812
rect 1053 1748 1069 1812
rect 1293 1811 1913 2000
rect 2021 1892 2148 2249
rect 2021 1828 2068 1892
rect 2132 1828 2148 1892
rect 2021 1812 2148 1828
rect 942 1732 1069 1748
rect 942 1668 989 1732
rect 1053 1668 1069 1732
rect 942 1652 1069 1668
rect 942 1588 989 1652
rect 1053 1588 1069 1652
rect 942 1572 1069 1588
rect 942 1508 989 1572
rect 1053 1508 1069 1572
rect 942 1492 1069 1508
rect 942 1428 989 1492
rect 1053 1428 1069 1492
rect 942 1412 1069 1428
rect 942 1348 989 1412
rect 1053 1348 1069 1412
rect 942 1332 1069 1348
rect 942 1268 989 1332
rect 1053 1268 1069 1332
rect 942 1252 1069 1268
rect 942 1188 989 1252
rect 1053 1188 1069 1252
rect 1292 1772 1914 1811
rect 1292 1228 1331 1772
rect 1875 1228 1914 1772
rect 1292 1189 1914 1228
rect 2021 1748 2068 1812
rect 2132 1748 2148 1812
rect 2021 1732 2148 1748
rect 2021 1668 2068 1732
rect 2132 1668 2148 1732
rect 2021 1652 2148 1668
rect 2021 1588 2068 1652
rect 2132 1588 2148 1652
rect 2021 1572 2148 1588
rect 2021 1508 2068 1572
rect 2132 1508 2148 1572
rect 2021 1492 2148 1508
rect 2021 1428 2068 1492
rect 2132 1428 2148 1492
rect 2021 1412 2148 1428
rect 2021 1348 2068 1412
rect 2132 1348 2148 1412
rect 2021 1332 2148 1348
rect 2021 1268 2068 1332
rect 2132 1268 2148 1332
rect 2021 1252 2148 1268
rect 942 1172 1069 1188
rect 942 1108 989 1172
rect 1053 1108 1069 1172
rect 942 1062 1069 1108
rect 942 938 1046 1062
rect 942 892 1069 938
rect 942 828 989 892
rect 1053 828 1069 892
rect 942 812 1069 828
rect 942 748 989 812
rect 1053 748 1069 812
rect 1300 811 1907 1189
rect 2021 1188 2068 1252
rect 2132 1188 2148 1252
rect 2021 1172 2148 1188
rect 2021 1108 2068 1172
rect 2132 1108 2148 1172
rect 2021 1062 2148 1108
rect 2021 938 2125 1062
rect 2021 892 2148 938
rect 2021 828 2068 892
rect 2132 828 2148 892
rect 2021 812 2148 828
rect 942 732 1069 748
rect 942 668 989 732
rect 1053 668 1069 732
rect 942 652 1069 668
rect 942 588 989 652
rect 1053 588 1069 652
rect 942 572 1069 588
rect 942 508 989 572
rect 1053 508 1069 572
rect 942 492 1069 508
rect 942 428 989 492
rect 1053 428 1069 492
rect 942 412 1069 428
rect 942 348 989 412
rect 1053 348 1069 412
rect 942 332 1069 348
rect 942 268 989 332
rect 1053 268 1069 332
rect 942 252 1069 268
rect 942 188 989 252
rect 1053 188 1069 252
rect 942 172 1069 188
rect 942 108 989 172
rect 1053 108 1069 172
rect 942 62 1069 108
rect 1292 772 1914 811
rect 1292 228 1331 772
rect 1875 228 1914 772
rect 942 -62 1046 62
rect 942 -108 1069 -62
rect 942 -172 989 -108
rect 1053 -172 1069 -108
rect 942 -188 1069 -172
rect 942 -252 989 -188
rect 1053 -252 1069 -188
rect 942 -268 1069 -252
rect 942 -332 989 -268
rect 1053 -332 1069 -268
rect 942 -348 1069 -332
rect 942 -412 989 -348
rect 1053 -412 1069 -348
rect 942 -428 1069 -412
rect 942 -492 989 -428
rect 1053 -492 1069 -428
rect 942 -508 1069 -492
rect 942 -572 989 -508
rect 1053 -572 1069 -508
rect 942 -588 1069 -572
rect 942 -652 989 -588
rect 1053 -652 1069 -588
rect 942 -668 1069 -652
rect 942 -732 989 -668
rect 1053 -732 1069 -668
rect 942 -748 1069 -732
rect 942 -812 989 -748
rect 1053 -812 1069 -748
rect 942 -828 1069 -812
rect 942 -892 989 -828
rect 1053 -892 1069 -828
rect 942 -938 1069 -892
rect 1292 -228 1914 228
rect 1292 -772 1331 -228
rect 1875 -772 1914 -228
rect 942 -1062 1046 -938
rect 942 -1108 1069 -1062
rect 942 -1172 989 -1108
rect 1053 -1172 1069 -1108
rect 942 -1188 1069 -1172
rect 942 -1252 989 -1188
rect 1053 -1252 1069 -1188
rect 942 -1268 1069 -1252
rect 942 -1332 989 -1268
rect 1053 -1332 1069 -1268
rect 942 -1348 1069 -1332
rect 942 -1412 989 -1348
rect 1053 -1412 1069 -1348
rect 942 -1428 1069 -1412
rect 942 -1492 989 -1428
rect 1053 -1492 1069 -1428
rect 942 -1508 1069 -1492
rect 942 -1572 989 -1508
rect 1053 -1572 1069 -1508
rect 942 -1588 1069 -1572
rect 942 -1652 989 -1588
rect 1053 -1652 1069 -1588
rect 942 -1668 1069 -1652
rect 942 -1732 989 -1668
rect 1053 -1732 1069 -1668
rect 942 -1748 1069 -1732
rect -141 -1828 -14 -1812
rect -141 -1892 -94 -1828
rect -30 -1892 -14 -1828
rect -141 -1938 -14 -1892
rect 219 -2202 830 -1811
rect 942 -1812 989 -1748
rect 1053 -1812 1069 -1748
rect 942 -1828 1069 -1812
rect 942 -1892 989 -1828
rect 1053 -1892 1069 -1828
rect 942 -1938 1069 -1892
rect 1292 -1228 1914 -772
rect 1292 -1772 1331 -1228
rect 1875 -1772 1914 -1228
rect 1292 -1811 1914 -1772
rect 2021 748 2068 812
rect 2132 748 2148 812
rect 2021 732 2148 748
rect 2021 668 2068 732
rect 2132 668 2148 732
rect 2021 652 2148 668
rect 2021 588 2068 652
rect 2132 588 2148 652
rect 2021 572 2148 588
rect 2021 508 2068 572
rect 2132 508 2148 572
rect 2021 492 2148 508
rect 2021 428 2068 492
rect 2132 428 2148 492
rect 2021 412 2148 428
rect 2021 348 2068 412
rect 2132 348 2148 412
rect 2021 332 2148 348
rect 2021 268 2068 332
rect 2132 268 2148 332
rect 2021 252 2148 268
rect 2021 188 2068 252
rect 2132 188 2148 252
rect 2021 172 2148 188
rect 2021 108 2068 172
rect 2132 108 2148 172
rect 2021 62 2148 108
rect 2021 -62 2125 62
rect 2021 -108 2148 -62
rect 2021 -172 2068 -108
rect 2132 -172 2148 -108
rect 2021 -188 2148 -172
rect 2021 -252 2068 -188
rect 2132 -252 2148 -188
rect 2021 -268 2148 -252
rect 2021 -332 2068 -268
rect 2132 -332 2148 -268
rect 2021 -348 2148 -332
rect 2021 -412 2068 -348
rect 2132 -412 2148 -348
rect 2021 -428 2148 -412
rect 2021 -492 2068 -428
rect 2132 -492 2148 -428
rect 2021 -508 2148 -492
rect 2021 -572 2068 -508
rect 2132 -572 2148 -508
rect 2021 -588 2148 -572
rect 2021 -652 2068 -588
rect 2132 -652 2148 -588
rect 2021 -668 2148 -652
rect 2021 -732 2068 -668
rect 2132 -732 2148 -668
rect 2021 -748 2148 -732
rect 2021 -812 2068 -748
rect 2132 -812 2148 -748
rect 2021 -828 2148 -812
rect 2021 -892 2068 -828
rect 2132 -892 2148 -828
rect 2021 -938 2148 -892
rect 2021 -1062 2125 -938
rect 2021 -1108 2148 -1062
rect 2021 -1172 2068 -1108
rect 2132 -1172 2148 -1108
rect 2021 -1188 2148 -1172
rect 2021 -1252 2068 -1188
rect 2132 -1252 2148 -1188
rect 2021 -1268 2148 -1252
rect 2021 -1332 2068 -1268
rect 2132 -1332 2148 -1268
rect 2021 -1348 2148 -1332
rect 2021 -1412 2068 -1348
rect 2132 -1412 2148 -1348
rect 2021 -1428 2148 -1412
rect 2021 -1492 2068 -1428
rect 2132 -1492 2148 -1428
rect 2021 -1508 2148 -1492
rect 2021 -1572 2068 -1508
rect 2132 -1572 2148 -1508
rect 2021 -1588 2148 -1572
rect 2021 -1652 2068 -1588
rect 2132 -1652 2148 -1588
rect 2021 -1668 2148 -1652
rect 2021 -1732 2068 -1668
rect 2132 -1732 2148 -1668
rect 2021 -1748 2148 -1732
rect 1292 -2202 1900 -1811
rect 2021 -1812 2068 -1748
rect 2132 -1812 2148 -1748
rect 2021 -1828 2148 -1812
rect 2021 -1892 2068 -1828
rect 2132 -1892 2148 -1828
rect 2021 -1938 2148 -1892
<< properties >>
string FIXED_BBOX 1029 1050 1929 1950
<< end >>
