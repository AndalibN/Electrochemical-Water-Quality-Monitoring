magic
tech sky130A
timestamp 1669522153
<< metal4 >>
rect 1700 -2766 2200 -1703
rect 1700 -2884 1766 -2766
rect 1884 -2884 1966 -2766
rect 2084 -2884 2200 -2766
rect 1700 -2966 2200 -2884
rect 1700 -3084 1816 -2966
rect 1934 -3084 2016 -2966
rect 2134 -3084 2200 -2966
rect 1700 -3200 2200 -3084
<< via4 >>
rect 1766 -2884 1884 -2766
rect 1966 -2884 2084 -2766
rect 1816 -3084 1934 -2966
rect 2016 -3084 2134 -2966
<< metal5 >>
rect 600 -1600 5800 -1100
rect 900 -2400 5000 -1900
rect 900 -5500 1400 -2400
rect 1700 -2766 2200 -2700
rect 1700 -2884 1766 -2766
rect 1884 -2884 1966 -2766
rect 2084 -2884 2200 -2766
rect 1700 -2966 2200 -2884
rect 1700 -3084 1816 -2966
rect 1934 -3084 2016 -2966
rect 2134 -3084 2200 -2966
rect 1700 -4600 2200 -3084
rect 4500 -4600 5000 -2400
rect 1700 -5200 5000 -4600
rect 5300 -5500 5800 -1600
rect 900 -6000 5800 -5500
<< end >>
