magic
tech sky130A
timestamp 1668102987
<< error_p >>
rect -14 186 14 189
rect -14 169 -8 186
rect -14 166 14 169
rect -14 -169 14 -166
rect -14 -186 -8 -169
rect -14 -189 14 -186
<< nmos >>
rect -15 -150 15 150
<< ndiff >>
rect -44 144 -15 150
rect -44 -144 -38 144
rect -21 -144 -15 144
rect -44 -150 -15 -144
rect 15 144 44 150
rect 15 -144 21 144
rect 38 -144 44 144
rect 15 -150 44 -144
<< ndiffc >>
rect -38 -144 -21 144
rect 21 -144 38 144
<< poly >>
rect -16 186 16 194
rect -16 169 -8 186
rect 8 169 16 186
rect -16 161 16 169
rect -15 150 15 161
rect -15 -161 15 -150
rect -16 -169 16 -161
rect -16 -186 -8 -169
rect 8 -186 16 -169
rect -16 -194 16 -186
<< polycont >>
rect -8 169 8 186
rect -8 -186 8 -169
<< locali >>
rect -16 169 -8 186
rect 8 169 16 186
rect -38 144 -21 152
rect -38 -152 -21 -144
rect 21 144 38 152
rect 21 -152 38 -144
rect -16 -186 -8 -169
rect 8 -186 16 -169
<< viali >>
rect -8 169 8 186
rect -38 -144 -21 144
rect 21 -144 38 144
rect -8 -186 8 -169
<< metal1 >>
rect -14 186 14 189
rect -14 169 -8 186
rect 8 169 14 186
rect -14 166 14 169
rect -41 144 -18 150
rect -41 -144 -38 144
rect -21 -144 -18 144
rect -41 -150 -18 -144
rect 18 144 41 150
rect 18 -144 21 144
rect 38 -144 41 144
rect 18 -150 41 -144
rect -14 -169 14 -166
rect -14 -186 -8 -169
rect 8 -186 14 -169
rect -14 -189 14 -186
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
