magic
tech sky130A
timestamp 1669522153
<< metal4 >>
rect 2700 -3566 3200 3378
rect 2700 -3684 2766 -3566
rect 2884 -3684 2966 -3566
rect 3084 -3684 3200 -3566
rect 2700 -3766 3200 -3684
rect 2700 -3884 2816 -3766
rect 2934 -3884 3016 -3766
rect 3134 -3884 3200 -3766
rect 2700 -4000 3200 -3884
<< via4 >>
rect 2766 -3684 2884 -3566
rect 2966 -3684 3084 -3566
rect 2816 -3884 2934 -3766
rect 3016 -3884 3134 -3766
<< metal5 >>
rect -1600 800 12300 1300
rect -1300 0 11500 500
rect -1300 -11800 -800 0
rect -500 -800 10700 -300
rect -500 -11000 0 -800
rect 300 -1600 9900 -1100
rect 300 -10200 800 -1600
rect 1100 -2400 9100 -1900
rect 1100 -9400 1600 -2400
rect 1900 -3200 8300 -2700
rect 1900 -8600 2400 -3200
rect 2700 -3566 3200 -3500
rect 2700 -3684 2766 -3566
rect 2884 -3684 2966 -3566
rect 3084 -3684 3200 -3566
rect 2700 -3766 3200 -3684
rect 2700 -3884 2816 -3766
rect 2934 -3884 3016 -3766
rect 3134 -3884 3200 -3766
rect 2700 -7800 3200 -3884
rect 7800 -7800 8300 -3200
rect 2700 -8300 8300 -7800
rect 8600 -8600 9100 -2400
rect 1900 -9100 9100 -8600
rect 9400 -9400 9900 -1600
rect 1100 -9900 9900 -9400
rect 10200 -10200 10700 -800
rect 300 -10700 10700 -10200
rect 11000 -11000 11500 0
rect -500 -11500 11500 -11000
rect 11800 -11800 12300 800
rect -1300 -12300 12300 -11800
<< end >>
