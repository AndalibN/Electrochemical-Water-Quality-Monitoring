magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -2688 2502 -1389 2550
rect -2688 2438 -1473 2502
rect -1409 2438 -1389 2502
rect -2688 2422 -1389 2438
rect -2688 2358 -1473 2422
rect -1409 2358 -1389 2422
rect -2688 2342 -1389 2358
rect -2688 2278 -1473 2342
rect -1409 2278 -1389 2342
rect -2688 2262 -1389 2278
rect -2688 2198 -1473 2262
rect -1409 2198 -1389 2262
rect -2688 2182 -1389 2198
rect -2688 2118 -1473 2182
rect -1409 2118 -1389 2182
rect -2688 2102 -1389 2118
rect -2688 2038 -1473 2102
rect -1409 2038 -1389 2102
rect -2688 2022 -1389 2038
rect -2688 1958 -1473 2022
rect -1409 1958 -1389 2022
rect -2688 1942 -1389 1958
rect -2688 1878 -1473 1942
rect -1409 1878 -1389 1942
rect -2688 1862 -1389 1878
rect -2688 1798 -1473 1862
rect -1409 1798 -1389 1862
rect -2688 1782 -1389 1798
rect -2688 1718 -1473 1782
rect -1409 1718 -1389 1782
rect -2688 1702 -1389 1718
rect -2688 1638 -1473 1702
rect -1409 1638 -1389 1702
rect -2688 1622 -1389 1638
rect -2688 1558 -1473 1622
rect -1409 1558 -1389 1622
rect -2688 1542 -1389 1558
rect -2688 1478 -1473 1542
rect -1409 1478 -1389 1542
rect -2688 1462 -1389 1478
rect -2688 1398 -1473 1462
rect -1409 1398 -1389 1462
rect -2688 1350 -1389 1398
rect -1309 2502 -10 2550
rect -1309 2438 -94 2502
rect -30 2438 -10 2502
rect -1309 2422 -10 2438
rect -1309 2358 -94 2422
rect -30 2358 -10 2422
rect -1309 2342 -10 2358
rect -1309 2278 -94 2342
rect -30 2278 -10 2342
rect -1309 2262 -10 2278
rect -1309 2198 -94 2262
rect -30 2198 -10 2262
rect -1309 2182 -10 2198
rect -1309 2118 -94 2182
rect -30 2118 -10 2182
rect -1309 2102 -10 2118
rect -1309 2038 -94 2102
rect -30 2038 -10 2102
rect -1309 2022 -10 2038
rect -1309 1958 -94 2022
rect -30 1958 -10 2022
rect -1309 1942 -10 1958
rect -1309 1878 -94 1942
rect -30 1878 -10 1942
rect -1309 1862 -10 1878
rect -1309 1798 -94 1862
rect -30 1798 -10 1862
rect -1309 1782 -10 1798
rect -1309 1718 -94 1782
rect -30 1718 -10 1782
rect -1309 1702 -10 1718
rect -1309 1638 -94 1702
rect -30 1638 -10 1702
rect -1309 1622 -10 1638
rect -1309 1558 -94 1622
rect -30 1558 -10 1622
rect -1309 1542 -10 1558
rect -1309 1478 -94 1542
rect -30 1478 -10 1542
rect -1309 1462 -10 1478
rect -1309 1398 -94 1462
rect -30 1398 -10 1462
rect -1309 1350 -10 1398
rect 70 2502 1369 2550
rect 70 2438 1285 2502
rect 1349 2438 1369 2502
rect 70 2422 1369 2438
rect 70 2358 1285 2422
rect 1349 2358 1369 2422
rect 70 2342 1369 2358
rect 70 2278 1285 2342
rect 1349 2278 1369 2342
rect 70 2262 1369 2278
rect 70 2198 1285 2262
rect 1349 2198 1369 2262
rect 70 2182 1369 2198
rect 70 2118 1285 2182
rect 1349 2118 1369 2182
rect 70 2102 1369 2118
rect 70 2038 1285 2102
rect 1349 2038 1369 2102
rect 70 2022 1369 2038
rect 70 1958 1285 2022
rect 1349 1958 1369 2022
rect 70 1942 1369 1958
rect 70 1878 1285 1942
rect 1349 1878 1369 1942
rect 70 1862 1369 1878
rect 70 1798 1285 1862
rect 1349 1798 1369 1862
rect 70 1782 1369 1798
rect 70 1718 1285 1782
rect 1349 1718 1369 1782
rect 70 1702 1369 1718
rect 70 1638 1285 1702
rect 1349 1638 1369 1702
rect 70 1622 1369 1638
rect 70 1558 1285 1622
rect 1349 1558 1369 1622
rect 70 1542 1369 1558
rect 70 1478 1285 1542
rect 1349 1478 1369 1542
rect 70 1462 1369 1478
rect 70 1398 1285 1462
rect 1349 1398 1369 1462
rect 70 1350 1369 1398
rect 1449 2502 2748 2550
rect 1449 2438 2664 2502
rect 2728 2438 2748 2502
rect 1449 2422 2748 2438
rect 1449 2358 2664 2422
rect 2728 2358 2748 2422
rect 1449 2342 2748 2358
rect 1449 2278 2664 2342
rect 2728 2278 2748 2342
rect 1449 2262 2748 2278
rect 1449 2198 2664 2262
rect 2728 2198 2748 2262
rect 1449 2182 2748 2198
rect 1449 2118 2664 2182
rect 2728 2118 2748 2182
rect 1449 2102 2748 2118
rect 1449 2038 2664 2102
rect 2728 2038 2748 2102
rect 1449 2022 2748 2038
rect 1449 1958 2664 2022
rect 2728 1958 2748 2022
rect 1449 1942 2748 1958
rect 1449 1878 2664 1942
rect 2728 1878 2748 1942
rect 1449 1862 2748 1878
rect 1449 1798 2664 1862
rect 2728 1798 2748 1862
rect 1449 1782 2748 1798
rect 1449 1718 2664 1782
rect 2728 1718 2748 1782
rect 1449 1702 2748 1718
rect 1449 1638 2664 1702
rect 2728 1638 2748 1702
rect 1449 1622 2748 1638
rect 1449 1558 2664 1622
rect 2728 1558 2748 1622
rect 1449 1542 2748 1558
rect 1449 1478 2664 1542
rect 2728 1478 2748 1542
rect 1449 1462 2748 1478
rect 1449 1398 2664 1462
rect 2728 1398 2748 1462
rect 1449 1350 2748 1398
rect -2688 1202 -1389 1250
rect -2688 1138 -1473 1202
rect -1409 1138 -1389 1202
rect -2688 1122 -1389 1138
rect -2688 1058 -1473 1122
rect -1409 1058 -1389 1122
rect -2688 1042 -1389 1058
rect -2688 978 -1473 1042
rect -1409 978 -1389 1042
rect -2688 962 -1389 978
rect -2688 898 -1473 962
rect -1409 898 -1389 962
rect -2688 882 -1389 898
rect -2688 818 -1473 882
rect -1409 818 -1389 882
rect -2688 802 -1389 818
rect -2688 738 -1473 802
rect -1409 738 -1389 802
rect -2688 722 -1389 738
rect -2688 658 -1473 722
rect -1409 658 -1389 722
rect -2688 642 -1389 658
rect -2688 578 -1473 642
rect -1409 578 -1389 642
rect -2688 562 -1389 578
rect -2688 498 -1473 562
rect -1409 498 -1389 562
rect -2688 482 -1389 498
rect -2688 418 -1473 482
rect -1409 418 -1389 482
rect -2688 402 -1389 418
rect -2688 338 -1473 402
rect -1409 338 -1389 402
rect -2688 322 -1389 338
rect -2688 258 -1473 322
rect -1409 258 -1389 322
rect -2688 242 -1389 258
rect -2688 178 -1473 242
rect -1409 178 -1389 242
rect -2688 162 -1389 178
rect -2688 98 -1473 162
rect -1409 98 -1389 162
rect -2688 50 -1389 98
rect -1309 1202 -10 1250
rect -1309 1138 -94 1202
rect -30 1138 -10 1202
rect -1309 1122 -10 1138
rect -1309 1058 -94 1122
rect -30 1058 -10 1122
rect -1309 1042 -10 1058
rect -1309 978 -94 1042
rect -30 978 -10 1042
rect -1309 962 -10 978
rect -1309 898 -94 962
rect -30 898 -10 962
rect -1309 882 -10 898
rect -1309 818 -94 882
rect -30 818 -10 882
rect -1309 802 -10 818
rect -1309 738 -94 802
rect -30 738 -10 802
rect -1309 722 -10 738
rect -1309 658 -94 722
rect -30 658 -10 722
rect -1309 642 -10 658
rect -1309 578 -94 642
rect -30 578 -10 642
rect -1309 562 -10 578
rect -1309 498 -94 562
rect -30 498 -10 562
rect -1309 482 -10 498
rect -1309 418 -94 482
rect -30 418 -10 482
rect -1309 402 -10 418
rect -1309 338 -94 402
rect -30 338 -10 402
rect -1309 322 -10 338
rect -1309 258 -94 322
rect -30 258 -10 322
rect -1309 242 -10 258
rect -1309 178 -94 242
rect -30 178 -10 242
rect -1309 162 -10 178
rect -1309 98 -94 162
rect -30 98 -10 162
rect -1309 50 -10 98
rect 70 1202 1369 1250
rect 70 1138 1285 1202
rect 1349 1138 1369 1202
rect 70 1122 1369 1138
rect 70 1058 1285 1122
rect 1349 1058 1369 1122
rect 70 1042 1369 1058
rect 70 978 1285 1042
rect 1349 978 1369 1042
rect 70 962 1369 978
rect 70 898 1285 962
rect 1349 898 1369 962
rect 70 882 1369 898
rect 70 818 1285 882
rect 1349 818 1369 882
rect 70 802 1369 818
rect 70 738 1285 802
rect 1349 738 1369 802
rect 70 722 1369 738
rect 70 658 1285 722
rect 1349 658 1369 722
rect 70 642 1369 658
rect 70 578 1285 642
rect 1349 578 1369 642
rect 70 562 1369 578
rect 70 498 1285 562
rect 1349 498 1369 562
rect 70 482 1369 498
rect 70 418 1285 482
rect 1349 418 1369 482
rect 70 402 1369 418
rect 70 338 1285 402
rect 1349 338 1369 402
rect 70 322 1369 338
rect 70 258 1285 322
rect 1349 258 1369 322
rect 70 242 1369 258
rect 70 178 1285 242
rect 1349 178 1369 242
rect 70 162 1369 178
rect 70 98 1285 162
rect 1349 98 1369 162
rect 70 50 1369 98
rect 1449 1202 2748 1250
rect 1449 1138 2664 1202
rect 2728 1138 2748 1202
rect 1449 1122 2748 1138
rect 1449 1058 2664 1122
rect 2728 1058 2748 1122
rect 1449 1042 2748 1058
rect 1449 978 2664 1042
rect 2728 978 2748 1042
rect 1449 962 2748 978
rect 1449 898 2664 962
rect 2728 898 2748 962
rect 1449 882 2748 898
rect 1449 818 2664 882
rect 2728 818 2748 882
rect 1449 802 2748 818
rect 1449 738 2664 802
rect 2728 738 2748 802
rect 1449 722 2748 738
rect 1449 658 2664 722
rect 2728 658 2748 722
rect 1449 642 2748 658
rect 1449 578 2664 642
rect 2728 578 2748 642
rect 1449 562 2748 578
rect 1449 498 2664 562
rect 2728 498 2748 562
rect 1449 482 2748 498
rect 1449 418 2664 482
rect 2728 418 2748 482
rect 1449 402 2748 418
rect 1449 338 2664 402
rect 2728 338 2748 402
rect 1449 322 2748 338
rect 1449 258 2664 322
rect 2728 258 2748 322
rect 1449 242 2748 258
rect 1449 178 2664 242
rect 2728 178 2748 242
rect 1449 162 2748 178
rect 1449 98 2664 162
rect 2728 98 2748 162
rect 1449 50 2748 98
rect -2688 -98 -1389 -50
rect -2688 -162 -1473 -98
rect -1409 -162 -1389 -98
rect -2688 -178 -1389 -162
rect -2688 -242 -1473 -178
rect -1409 -242 -1389 -178
rect -2688 -258 -1389 -242
rect -2688 -322 -1473 -258
rect -1409 -322 -1389 -258
rect -2688 -338 -1389 -322
rect -2688 -402 -1473 -338
rect -1409 -402 -1389 -338
rect -2688 -418 -1389 -402
rect -2688 -482 -1473 -418
rect -1409 -482 -1389 -418
rect -2688 -498 -1389 -482
rect -2688 -562 -1473 -498
rect -1409 -562 -1389 -498
rect -2688 -578 -1389 -562
rect -2688 -642 -1473 -578
rect -1409 -642 -1389 -578
rect -2688 -658 -1389 -642
rect -2688 -722 -1473 -658
rect -1409 -722 -1389 -658
rect -2688 -738 -1389 -722
rect -2688 -802 -1473 -738
rect -1409 -802 -1389 -738
rect -2688 -818 -1389 -802
rect -2688 -882 -1473 -818
rect -1409 -882 -1389 -818
rect -2688 -898 -1389 -882
rect -2688 -962 -1473 -898
rect -1409 -962 -1389 -898
rect -2688 -978 -1389 -962
rect -2688 -1042 -1473 -978
rect -1409 -1042 -1389 -978
rect -2688 -1058 -1389 -1042
rect -2688 -1122 -1473 -1058
rect -1409 -1122 -1389 -1058
rect -2688 -1138 -1389 -1122
rect -2688 -1202 -1473 -1138
rect -1409 -1202 -1389 -1138
rect -2688 -1250 -1389 -1202
rect -1309 -98 -10 -50
rect -1309 -162 -94 -98
rect -30 -162 -10 -98
rect -1309 -178 -10 -162
rect -1309 -242 -94 -178
rect -30 -242 -10 -178
rect -1309 -258 -10 -242
rect -1309 -322 -94 -258
rect -30 -322 -10 -258
rect -1309 -338 -10 -322
rect -1309 -402 -94 -338
rect -30 -402 -10 -338
rect -1309 -418 -10 -402
rect -1309 -482 -94 -418
rect -30 -482 -10 -418
rect -1309 -498 -10 -482
rect -1309 -562 -94 -498
rect -30 -562 -10 -498
rect -1309 -578 -10 -562
rect -1309 -642 -94 -578
rect -30 -642 -10 -578
rect -1309 -658 -10 -642
rect -1309 -722 -94 -658
rect -30 -722 -10 -658
rect -1309 -738 -10 -722
rect -1309 -802 -94 -738
rect -30 -802 -10 -738
rect -1309 -818 -10 -802
rect -1309 -882 -94 -818
rect -30 -882 -10 -818
rect -1309 -898 -10 -882
rect -1309 -962 -94 -898
rect -30 -962 -10 -898
rect -1309 -978 -10 -962
rect -1309 -1042 -94 -978
rect -30 -1042 -10 -978
rect -1309 -1058 -10 -1042
rect -1309 -1122 -94 -1058
rect -30 -1122 -10 -1058
rect -1309 -1138 -10 -1122
rect -1309 -1202 -94 -1138
rect -30 -1202 -10 -1138
rect -1309 -1250 -10 -1202
rect 70 -98 1369 -50
rect 70 -162 1285 -98
rect 1349 -162 1369 -98
rect 70 -178 1369 -162
rect 70 -242 1285 -178
rect 1349 -242 1369 -178
rect 70 -258 1369 -242
rect 70 -322 1285 -258
rect 1349 -322 1369 -258
rect 70 -338 1369 -322
rect 70 -402 1285 -338
rect 1349 -402 1369 -338
rect 70 -418 1369 -402
rect 70 -482 1285 -418
rect 1349 -482 1369 -418
rect 70 -498 1369 -482
rect 70 -562 1285 -498
rect 1349 -562 1369 -498
rect 70 -578 1369 -562
rect 70 -642 1285 -578
rect 1349 -642 1369 -578
rect 70 -658 1369 -642
rect 70 -722 1285 -658
rect 1349 -722 1369 -658
rect 70 -738 1369 -722
rect 70 -802 1285 -738
rect 1349 -802 1369 -738
rect 70 -818 1369 -802
rect 70 -882 1285 -818
rect 1349 -882 1369 -818
rect 70 -898 1369 -882
rect 70 -962 1285 -898
rect 1349 -962 1369 -898
rect 70 -978 1369 -962
rect 70 -1042 1285 -978
rect 1349 -1042 1369 -978
rect 70 -1058 1369 -1042
rect 70 -1122 1285 -1058
rect 1349 -1122 1369 -1058
rect 70 -1138 1369 -1122
rect 70 -1202 1285 -1138
rect 1349 -1202 1369 -1138
rect 70 -1250 1369 -1202
rect 1449 -98 2748 -50
rect 1449 -162 2664 -98
rect 2728 -162 2748 -98
rect 1449 -178 2748 -162
rect 1449 -242 2664 -178
rect 2728 -242 2748 -178
rect 1449 -258 2748 -242
rect 1449 -322 2664 -258
rect 2728 -322 2748 -258
rect 1449 -338 2748 -322
rect 1449 -402 2664 -338
rect 2728 -402 2748 -338
rect 1449 -418 2748 -402
rect 1449 -482 2664 -418
rect 2728 -482 2748 -418
rect 1449 -498 2748 -482
rect 1449 -562 2664 -498
rect 2728 -562 2748 -498
rect 1449 -578 2748 -562
rect 1449 -642 2664 -578
rect 2728 -642 2748 -578
rect 1449 -658 2748 -642
rect 1449 -722 2664 -658
rect 2728 -722 2748 -658
rect 1449 -738 2748 -722
rect 1449 -802 2664 -738
rect 2728 -802 2748 -738
rect 1449 -818 2748 -802
rect 1449 -882 2664 -818
rect 2728 -882 2748 -818
rect 1449 -898 2748 -882
rect 1449 -962 2664 -898
rect 2728 -962 2748 -898
rect 1449 -978 2748 -962
rect 1449 -1042 2664 -978
rect 2728 -1042 2748 -978
rect 1449 -1058 2748 -1042
rect 1449 -1122 2664 -1058
rect 2728 -1122 2748 -1058
rect 1449 -1138 2748 -1122
rect 1449 -1202 2664 -1138
rect 2728 -1202 2748 -1138
rect 1449 -1250 2748 -1202
rect -2688 -1398 -1389 -1350
rect -2688 -1462 -1473 -1398
rect -1409 -1462 -1389 -1398
rect -2688 -1478 -1389 -1462
rect -2688 -1542 -1473 -1478
rect -1409 -1542 -1389 -1478
rect -2688 -1558 -1389 -1542
rect -2688 -1622 -1473 -1558
rect -1409 -1622 -1389 -1558
rect -2688 -1638 -1389 -1622
rect -2688 -1702 -1473 -1638
rect -1409 -1702 -1389 -1638
rect -2688 -1718 -1389 -1702
rect -2688 -1782 -1473 -1718
rect -1409 -1782 -1389 -1718
rect -2688 -1798 -1389 -1782
rect -2688 -1862 -1473 -1798
rect -1409 -1862 -1389 -1798
rect -2688 -1878 -1389 -1862
rect -2688 -1942 -1473 -1878
rect -1409 -1942 -1389 -1878
rect -2688 -1958 -1389 -1942
rect -2688 -2022 -1473 -1958
rect -1409 -2022 -1389 -1958
rect -2688 -2038 -1389 -2022
rect -2688 -2102 -1473 -2038
rect -1409 -2102 -1389 -2038
rect -2688 -2118 -1389 -2102
rect -2688 -2182 -1473 -2118
rect -1409 -2182 -1389 -2118
rect -2688 -2198 -1389 -2182
rect -2688 -2262 -1473 -2198
rect -1409 -2262 -1389 -2198
rect -2688 -2278 -1389 -2262
rect -2688 -2342 -1473 -2278
rect -1409 -2342 -1389 -2278
rect -2688 -2358 -1389 -2342
rect -2688 -2422 -1473 -2358
rect -1409 -2422 -1389 -2358
rect -2688 -2438 -1389 -2422
rect -2688 -2502 -1473 -2438
rect -1409 -2502 -1389 -2438
rect -2688 -2550 -1389 -2502
rect -1309 -1398 -10 -1350
rect -1309 -1462 -94 -1398
rect -30 -1462 -10 -1398
rect -1309 -1478 -10 -1462
rect -1309 -1542 -94 -1478
rect -30 -1542 -10 -1478
rect -1309 -1558 -10 -1542
rect -1309 -1622 -94 -1558
rect -30 -1622 -10 -1558
rect -1309 -1638 -10 -1622
rect -1309 -1702 -94 -1638
rect -30 -1702 -10 -1638
rect -1309 -1718 -10 -1702
rect -1309 -1782 -94 -1718
rect -30 -1782 -10 -1718
rect -1309 -1798 -10 -1782
rect -1309 -1862 -94 -1798
rect -30 -1862 -10 -1798
rect -1309 -1878 -10 -1862
rect -1309 -1942 -94 -1878
rect -30 -1942 -10 -1878
rect -1309 -1958 -10 -1942
rect -1309 -2022 -94 -1958
rect -30 -2022 -10 -1958
rect -1309 -2038 -10 -2022
rect -1309 -2102 -94 -2038
rect -30 -2102 -10 -2038
rect -1309 -2118 -10 -2102
rect -1309 -2182 -94 -2118
rect -30 -2182 -10 -2118
rect -1309 -2198 -10 -2182
rect -1309 -2262 -94 -2198
rect -30 -2262 -10 -2198
rect -1309 -2278 -10 -2262
rect -1309 -2342 -94 -2278
rect -30 -2342 -10 -2278
rect -1309 -2358 -10 -2342
rect -1309 -2422 -94 -2358
rect -30 -2422 -10 -2358
rect -1309 -2438 -10 -2422
rect -1309 -2502 -94 -2438
rect -30 -2502 -10 -2438
rect -1309 -2550 -10 -2502
rect 70 -1398 1369 -1350
rect 70 -1462 1285 -1398
rect 1349 -1462 1369 -1398
rect 70 -1478 1369 -1462
rect 70 -1542 1285 -1478
rect 1349 -1542 1369 -1478
rect 70 -1558 1369 -1542
rect 70 -1622 1285 -1558
rect 1349 -1622 1369 -1558
rect 70 -1638 1369 -1622
rect 70 -1702 1285 -1638
rect 1349 -1702 1369 -1638
rect 70 -1718 1369 -1702
rect 70 -1782 1285 -1718
rect 1349 -1782 1369 -1718
rect 70 -1798 1369 -1782
rect 70 -1862 1285 -1798
rect 1349 -1862 1369 -1798
rect 70 -1878 1369 -1862
rect 70 -1942 1285 -1878
rect 1349 -1942 1369 -1878
rect 70 -1958 1369 -1942
rect 70 -2022 1285 -1958
rect 1349 -2022 1369 -1958
rect 70 -2038 1369 -2022
rect 70 -2102 1285 -2038
rect 1349 -2102 1369 -2038
rect 70 -2118 1369 -2102
rect 70 -2182 1285 -2118
rect 1349 -2182 1369 -2118
rect 70 -2198 1369 -2182
rect 70 -2262 1285 -2198
rect 1349 -2262 1369 -2198
rect 70 -2278 1369 -2262
rect 70 -2342 1285 -2278
rect 1349 -2342 1369 -2278
rect 70 -2358 1369 -2342
rect 70 -2422 1285 -2358
rect 1349 -2422 1369 -2358
rect 70 -2438 1369 -2422
rect 70 -2502 1285 -2438
rect 1349 -2502 1369 -2438
rect 70 -2550 1369 -2502
rect 1449 -1398 2748 -1350
rect 1449 -1462 2664 -1398
rect 2728 -1462 2748 -1398
rect 1449 -1478 2748 -1462
rect 1449 -1542 2664 -1478
rect 2728 -1542 2748 -1478
rect 1449 -1558 2748 -1542
rect 1449 -1622 2664 -1558
rect 2728 -1622 2748 -1558
rect 1449 -1638 2748 -1622
rect 1449 -1702 2664 -1638
rect 2728 -1702 2748 -1638
rect 1449 -1718 2748 -1702
rect 1449 -1782 2664 -1718
rect 2728 -1782 2748 -1718
rect 1449 -1798 2748 -1782
rect 1449 -1862 2664 -1798
rect 2728 -1862 2748 -1798
rect 1449 -1878 2748 -1862
rect 1449 -1942 2664 -1878
rect 2728 -1942 2748 -1878
rect 1449 -1958 2748 -1942
rect 1449 -2022 2664 -1958
rect 2728 -2022 2748 -1958
rect 1449 -2038 2748 -2022
rect 1449 -2102 2664 -2038
rect 2728 -2102 2748 -2038
rect 1449 -2118 2748 -2102
rect 1449 -2182 2664 -2118
rect 2728 -2182 2748 -2118
rect 1449 -2198 2748 -2182
rect 1449 -2262 2664 -2198
rect 2728 -2262 2748 -2198
rect 1449 -2278 2748 -2262
rect 1449 -2342 2664 -2278
rect 2728 -2342 2748 -2278
rect 1449 -2358 2748 -2342
rect 1449 -2422 2664 -2358
rect 2728 -2422 2748 -2358
rect 1449 -2438 2748 -2422
rect 1449 -2502 2664 -2438
rect 2728 -2502 2748 -2438
rect 1449 -2550 2748 -2502
<< via3 >>
rect -1473 2438 -1409 2502
rect -1473 2358 -1409 2422
rect -1473 2278 -1409 2342
rect -1473 2198 -1409 2262
rect -1473 2118 -1409 2182
rect -1473 2038 -1409 2102
rect -1473 1958 -1409 2022
rect -1473 1878 -1409 1942
rect -1473 1798 -1409 1862
rect -1473 1718 -1409 1782
rect -1473 1638 -1409 1702
rect -1473 1558 -1409 1622
rect -1473 1478 -1409 1542
rect -1473 1398 -1409 1462
rect -94 2438 -30 2502
rect -94 2358 -30 2422
rect -94 2278 -30 2342
rect -94 2198 -30 2262
rect -94 2118 -30 2182
rect -94 2038 -30 2102
rect -94 1958 -30 2022
rect -94 1878 -30 1942
rect -94 1798 -30 1862
rect -94 1718 -30 1782
rect -94 1638 -30 1702
rect -94 1558 -30 1622
rect -94 1478 -30 1542
rect -94 1398 -30 1462
rect 1285 2438 1349 2502
rect 1285 2358 1349 2422
rect 1285 2278 1349 2342
rect 1285 2198 1349 2262
rect 1285 2118 1349 2182
rect 1285 2038 1349 2102
rect 1285 1958 1349 2022
rect 1285 1878 1349 1942
rect 1285 1798 1349 1862
rect 1285 1718 1349 1782
rect 1285 1638 1349 1702
rect 1285 1558 1349 1622
rect 1285 1478 1349 1542
rect 1285 1398 1349 1462
rect 2664 2438 2728 2502
rect 2664 2358 2728 2422
rect 2664 2278 2728 2342
rect 2664 2198 2728 2262
rect 2664 2118 2728 2182
rect 2664 2038 2728 2102
rect 2664 1958 2728 2022
rect 2664 1878 2728 1942
rect 2664 1798 2728 1862
rect 2664 1718 2728 1782
rect 2664 1638 2728 1702
rect 2664 1558 2728 1622
rect 2664 1478 2728 1542
rect 2664 1398 2728 1462
rect -1473 1138 -1409 1202
rect -1473 1058 -1409 1122
rect -1473 978 -1409 1042
rect -1473 898 -1409 962
rect -1473 818 -1409 882
rect -1473 738 -1409 802
rect -1473 658 -1409 722
rect -1473 578 -1409 642
rect -1473 498 -1409 562
rect -1473 418 -1409 482
rect -1473 338 -1409 402
rect -1473 258 -1409 322
rect -1473 178 -1409 242
rect -1473 98 -1409 162
rect -94 1138 -30 1202
rect -94 1058 -30 1122
rect -94 978 -30 1042
rect -94 898 -30 962
rect -94 818 -30 882
rect -94 738 -30 802
rect -94 658 -30 722
rect -94 578 -30 642
rect -94 498 -30 562
rect -94 418 -30 482
rect -94 338 -30 402
rect -94 258 -30 322
rect -94 178 -30 242
rect -94 98 -30 162
rect 1285 1138 1349 1202
rect 1285 1058 1349 1122
rect 1285 978 1349 1042
rect 1285 898 1349 962
rect 1285 818 1349 882
rect 1285 738 1349 802
rect 1285 658 1349 722
rect 1285 578 1349 642
rect 1285 498 1349 562
rect 1285 418 1349 482
rect 1285 338 1349 402
rect 1285 258 1349 322
rect 1285 178 1349 242
rect 1285 98 1349 162
rect 2664 1138 2728 1202
rect 2664 1058 2728 1122
rect 2664 978 2728 1042
rect 2664 898 2728 962
rect 2664 818 2728 882
rect 2664 738 2728 802
rect 2664 658 2728 722
rect 2664 578 2728 642
rect 2664 498 2728 562
rect 2664 418 2728 482
rect 2664 338 2728 402
rect 2664 258 2728 322
rect 2664 178 2728 242
rect 2664 98 2728 162
rect -1473 -162 -1409 -98
rect -1473 -242 -1409 -178
rect -1473 -322 -1409 -258
rect -1473 -402 -1409 -338
rect -1473 -482 -1409 -418
rect -1473 -562 -1409 -498
rect -1473 -642 -1409 -578
rect -1473 -722 -1409 -658
rect -1473 -802 -1409 -738
rect -1473 -882 -1409 -818
rect -1473 -962 -1409 -898
rect -1473 -1042 -1409 -978
rect -1473 -1122 -1409 -1058
rect -1473 -1202 -1409 -1138
rect -94 -162 -30 -98
rect -94 -242 -30 -178
rect -94 -322 -30 -258
rect -94 -402 -30 -338
rect -94 -482 -30 -418
rect -94 -562 -30 -498
rect -94 -642 -30 -578
rect -94 -722 -30 -658
rect -94 -802 -30 -738
rect -94 -882 -30 -818
rect -94 -962 -30 -898
rect -94 -1042 -30 -978
rect -94 -1122 -30 -1058
rect -94 -1202 -30 -1138
rect 1285 -162 1349 -98
rect 1285 -242 1349 -178
rect 1285 -322 1349 -258
rect 1285 -402 1349 -338
rect 1285 -482 1349 -418
rect 1285 -562 1349 -498
rect 1285 -642 1349 -578
rect 1285 -722 1349 -658
rect 1285 -802 1349 -738
rect 1285 -882 1349 -818
rect 1285 -962 1349 -898
rect 1285 -1042 1349 -978
rect 1285 -1122 1349 -1058
rect 1285 -1202 1349 -1138
rect 2664 -162 2728 -98
rect 2664 -242 2728 -178
rect 2664 -322 2728 -258
rect 2664 -402 2728 -338
rect 2664 -482 2728 -418
rect 2664 -562 2728 -498
rect 2664 -642 2728 -578
rect 2664 -722 2728 -658
rect 2664 -802 2728 -738
rect 2664 -882 2728 -818
rect 2664 -962 2728 -898
rect 2664 -1042 2728 -978
rect 2664 -1122 2728 -1058
rect 2664 -1202 2728 -1138
rect -1473 -1462 -1409 -1398
rect -1473 -1542 -1409 -1478
rect -1473 -1622 -1409 -1558
rect -1473 -1702 -1409 -1638
rect -1473 -1782 -1409 -1718
rect -1473 -1862 -1409 -1798
rect -1473 -1942 -1409 -1878
rect -1473 -2022 -1409 -1958
rect -1473 -2102 -1409 -2038
rect -1473 -2182 -1409 -2118
rect -1473 -2262 -1409 -2198
rect -1473 -2342 -1409 -2278
rect -1473 -2422 -1409 -2358
rect -1473 -2502 -1409 -2438
rect -94 -1462 -30 -1398
rect -94 -1542 -30 -1478
rect -94 -1622 -30 -1558
rect -94 -1702 -30 -1638
rect -94 -1782 -30 -1718
rect -94 -1862 -30 -1798
rect -94 -1942 -30 -1878
rect -94 -2022 -30 -1958
rect -94 -2102 -30 -2038
rect -94 -2182 -30 -2118
rect -94 -2262 -30 -2198
rect -94 -2342 -30 -2278
rect -94 -2422 -30 -2358
rect -94 -2502 -30 -2438
rect 1285 -1462 1349 -1398
rect 1285 -1542 1349 -1478
rect 1285 -1622 1349 -1558
rect 1285 -1702 1349 -1638
rect 1285 -1782 1349 -1718
rect 1285 -1862 1349 -1798
rect 1285 -1942 1349 -1878
rect 1285 -2022 1349 -1958
rect 1285 -2102 1349 -2038
rect 1285 -2182 1349 -2118
rect 1285 -2262 1349 -2198
rect 1285 -2342 1349 -2278
rect 1285 -2422 1349 -2358
rect 1285 -2502 1349 -2438
rect 2664 -1462 2728 -1398
rect 2664 -1542 2728 -1478
rect 2664 -1622 2728 -1558
rect 2664 -1702 2728 -1638
rect 2664 -1782 2728 -1718
rect 2664 -1862 2728 -1798
rect 2664 -1942 2728 -1878
rect 2664 -2022 2728 -1958
rect 2664 -2102 2728 -2038
rect 2664 -2182 2728 -2118
rect 2664 -2262 2728 -2198
rect 2664 -2342 2728 -2278
rect 2664 -2422 2728 -2358
rect 2664 -2502 2728 -2438
<< mimcap >>
rect -2588 2382 -1588 2450
rect -2588 1518 -2520 2382
rect -1656 1518 -1588 2382
rect -2588 1450 -1588 1518
rect -1209 2382 -209 2450
rect -1209 1518 -1141 2382
rect -277 1518 -209 2382
rect -1209 1450 -209 1518
rect 170 2382 1170 2450
rect 170 1518 238 2382
rect 1102 1518 1170 2382
rect 170 1450 1170 1518
rect 1549 2382 2549 2450
rect 1549 1518 1617 2382
rect 2481 1518 2549 2382
rect 1549 1450 2549 1518
rect -2588 1082 -1588 1150
rect -2588 218 -2520 1082
rect -1656 218 -1588 1082
rect -2588 150 -1588 218
rect -1209 1082 -209 1150
rect -1209 218 -1141 1082
rect -277 218 -209 1082
rect -1209 150 -209 218
rect 170 1082 1170 1150
rect 170 218 238 1082
rect 1102 218 1170 1082
rect 170 150 1170 218
rect 1549 1082 2549 1150
rect 1549 218 1617 1082
rect 2481 218 2549 1082
rect 1549 150 2549 218
rect -2588 -218 -1588 -150
rect -2588 -1082 -2520 -218
rect -1656 -1082 -1588 -218
rect -2588 -1150 -1588 -1082
rect -1209 -218 -209 -150
rect -1209 -1082 -1141 -218
rect -277 -1082 -209 -218
rect -1209 -1150 -209 -1082
rect 170 -218 1170 -150
rect 170 -1082 238 -218
rect 1102 -1082 1170 -218
rect 170 -1150 1170 -1082
rect 1549 -218 2549 -150
rect 1549 -1082 1617 -218
rect 2481 -1082 2549 -218
rect 1549 -1150 2549 -1082
rect -2588 -1518 -1588 -1450
rect -2588 -2382 -2520 -1518
rect -1656 -2382 -1588 -1518
rect -2588 -2450 -1588 -2382
rect -1209 -1518 -209 -1450
rect -1209 -2382 -1141 -1518
rect -277 -2382 -209 -1518
rect -1209 -2450 -209 -2382
rect 170 -1518 1170 -1450
rect 170 -2382 238 -1518
rect 1102 -2382 1170 -1518
rect 170 -2450 1170 -2382
rect 1549 -1518 2549 -1450
rect 1549 -2382 1617 -1518
rect 2481 -2382 2549 -1518
rect 1549 -2450 2549 -2382
<< mimcapcontact >>
rect -2520 1518 -1656 2382
rect -1141 1518 -277 2382
rect 238 1518 1102 2382
rect 1617 1518 2481 2382
rect -2520 218 -1656 1082
rect -1141 218 -277 1082
rect 238 218 1102 1082
rect 1617 218 2481 1082
rect -2520 -1082 -1656 -218
rect -1141 -1082 -277 -218
rect 238 -1082 1102 -218
rect 1617 -1082 2481 -218
rect -2520 -2382 -1656 -1518
rect -1141 -2382 -277 -1518
rect 238 -2382 1102 -1518
rect 1617 -2382 2481 -1518
<< metal4 >>
rect -2549 2382 -1627 2600
rect -2549 1518 -2520 2382
rect -1656 1518 -1627 2382
rect -2549 1082 -1627 1518
rect -2549 218 -2520 1082
rect -1656 218 -1627 1082
rect -2549 -218 -1627 218
rect -2549 -1082 -2520 -218
rect -1656 -1082 -1627 -218
rect -2549 -1518 -1627 -1082
rect -2549 -2382 -2520 -1518
rect -1656 -2382 -1627 -1518
rect -2549 -2939 -1627 -2382
rect -1520 2538 -1416 2600
rect -1520 2502 -1393 2538
rect -1520 2438 -1473 2502
rect -1409 2438 -1393 2502
rect -1520 2422 -1393 2438
rect -1520 2358 -1473 2422
rect -1409 2358 -1393 2422
rect -1520 2342 -1393 2358
rect -1520 2278 -1473 2342
rect -1409 2278 -1393 2342
rect -1520 2262 -1393 2278
rect -1520 2198 -1473 2262
rect -1409 2198 -1393 2262
rect -1520 2182 -1393 2198
rect -1520 2118 -1473 2182
rect -1409 2118 -1393 2182
rect -1520 2102 -1393 2118
rect -1520 2038 -1473 2102
rect -1409 2038 -1393 2102
rect -1520 2022 -1393 2038
rect -1520 1958 -1473 2022
rect -1409 1958 -1393 2022
rect -1520 1942 -1393 1958
rect -1520 1878 -1473 1942
rect -1409 1878 -1393 1942
rect -1520 1862 -1393 1878
rect -1520 1798 -1473 1862
rect -1409 1798 -1393 1862
rect -1520 1782 -1393 1798
rect -1520 1718 -1473 1782
rect -1409 1718 -1393 1782
rect -1520 1702 -1393 1718
rect -1520 1638 -1473 1702
rect -1409 1638 -1393 1702
rect -1520 1622 -1393 1638
rect -1520 1558 -1473 1622
rect -1409 1558 -1393 1622
rect -1520 1542 -1393 1558
rect -1520 1478 -1473 1542
rect -1409 1478 -1393 1542
rect -1520 1462 -1393 1478
rect -1520 1398 -1473 1462
rect -1409 1398 -1393 1462
rect -1520 1362 -1393 1398
rect -1170 2382 -248 2600
rect -1170 1518 -1141 2382
rect -277 1518 -248 2382
rect -1520 1238 -1416 1362
rect -1520 1202 -1393 1238
rect -1520 1138 -1473 1202
rect -1409 1138 -1393 1202
rect -1520 1122 -1393 1138
rect -1520 1058 -1473 1122
rect -1409 1058 -1393 1122
rect -1520 1042 -1393 1058
rect -1520 978 -1473 1042
rect -1409 978 -1393 1042
rect -1520 962 -1393 978
rect -1520 898 -1473 962
rect -1409 898 -1393 962
rect -1520 882 -1393 898
rect -1520 818 -1473 882
rect -1409 818 -1393 882
rect -1520 802 -1393 818
rect -1520 738 -1473 802
rect -1409 738 -1393 802
rect -1520 722 -1393 738
rect -1520 658 -1473 722
rect -1409 658 -1393 722
rect -1520 642 -1393 658
rect -1520 578 -1473 642
rect -1409 578 -1393 642
rect -1520 562 -1393 578
rect -1520 498 -1473 562
rect -1409 498 -1393 562
rect -1520 482 -1393 498
rect -1520 418 -1473 482
rect -1409 418 -1393 482
rect -1520 402 -1393 418
rect -1520 338 -1473 402
rect -1409 338 -1393 402
rect -1520 322 -1393 338
rect -1520 258 -1473 322
rect -1409 258 -1393 322
rect -1520 242 -1393 258
rect -1520 178 -1473 242
rect -1409 178 -1393 242
rect -1520 162 -1393 178
rect -1520 98 -1473 162
rect -1409 98 -1393 162
rect -1520 62 -1393 98
rect -1170 1082 -248 1518
rect -1170 218 -1141 1082
rect -277 218 -248 1082
rect -1520 -62 -1416 62
rect -1520 -98 -1393 -62
rect -1520 -162 -1473 -98
rect -1409 -162 -1393 -98
rect -1520 -178 -1393 -162
rect -1520 -242 -1473 -178
rect -1409 -242 -1393 -178
rect -1520 -258 -1393 -242
rect -1520 -322 -1473 -258
rect -1409 -322 -1393 -258
rect -1520 -338 -1393 -322
rect -1520 -402 -1473 -338
rect -1409 -402 -1393 -338
rect -1520 -418 -1393 -402
rect -1520 -482 -1473 -418
rect -1409 -482 -1393 -418
rect -1520 -498 -1393 -482
rect -1520 -562 -1473 -498
rect -1409 -562 -1393 -498
rect -1520 -578 -1393 -562
rect -1520 -642 -1473 -578
rect -1409 -642 -1393 -578
rect -1520 -658 -1393 -642
rect -1520 -722 -1473 -658
rect -1409 -722 -1393 -658
rect -1520 -738 -1393 -722
rect -1520 -802 -1473 -738
rect -1409 -802 -1393 -738
rect -1520 -818 -1393 -802
rect -1520 -882 -1473 -818
rect -1409 -882 -1393 -818
rect -1520 -898 -1393 -882
rect -1520 -962 -1473 -898
rect -1409 -962 -1393 -898
rect -1520 -978 -1393 -962
rect -1520 -1042 -1473 -978
rect -1409 -1042 -1393 -978
rect -1520 -1058 -1393 -1042
rect -1520 -1122 -1473 -1058
rect -1409 -1122 -1393 -1058
rect -1520 -1138 -1393 -1122
rect -1520 -1202 -1473 -1138
rect -1409 -1202 -1393 -1138
rect -1520 -1238 -1393 -1202
rect -1170 -218 -248 218
rect -1170 -1082 -1141 -218
rect -277 -1082 -248 -218
rect -1520 -1362 -1416 -1238
rect -1520 -1398 -1393 -1362
rect -1520 -1462 -1473 -1398
rect -1409 -1462 -1393 -1398
rect -1520 -1478 -1393 -1462
rect -1520 -1542 -1473 -1478
rect -1409 -1542 -1393 -1478
rect -1520 -1558 -1393 -1542
rect -1520 -1622 -1473 -1558
rect -1409 -1622 -1393 -1558
rect -1520 -1638 -1393 -1622
rect -1520 -1702 -1473 -1638
rect -1409 -1702 -1393 -1638
rect -1520 -1718 -1393 -1702
rect -1520 -1782 -1473 -1718
rect -1409 -1782 -1393 -1718
rect -1520 -1798 -1393 -1782
rect -1520 -1862 -1473 -1798
rect -1409 -1862 -1393 -1798
rect -1520 -1878 -1393 -1862
rect -1520 -1942 -1473 -1878
rect -1409 -1942 -1393 -1878
rect -1520 -1958 -1393 -1942
rect -1520 -2022 -1473 -1958
rect -1409 -2022 -1393 -1958
rect -1520 -2038 -1393 -2022
rect -1520 -2102 -1473 -2038
rect -1409 -2102 -1393 -2038
rect -1520 -2118 -1393 -2102
rect -1520 -2182 -1473 -2118
rect -1409 -2182 -1393 -2118
rect -1520 -2198 -1393 -2182
rect -1520 -2262 -1473 -2198
rect -1409 -2262 -1393 -2198
rect -1520 -2278 -1393 -2262
rect -1520 -2342 -1473 -2278
rect -1409 -2342 -1393 -2278
rect -1520 -2358 -1393 -2342
rect -1520 -2422 -1473 -2358
rect -1409 -2422 -1393 -2358
rect -1520 -2438 -1393 -2422
rect -1520 -2502 -1473 -2438
rect -1409 -2502 -1393 -2438
rect -1520 -2538 -1393 -2502
rect -1170 -1518 -248 -1082
rect -1170 -2382 -1141 -1518
rect -277 -2382 -248 -1518
rect -1520 -2600 -1416 -2538
rect -1170 -2936 -248 -2382
rect -141 2538 -37 2600
rect -141 2502 -14 2538
rect -141 2438 -94 2502
rect -30 2438 -14 2502
rect -141 2422 -14 2438
rect -141 2358 -94 2422
rect -30 2358 -14 2422
rect -141 2342 -14 2358
rect -141 2278 -94 2342
rect -30 2278 -14 2342
rect -141 2262 -14 2278
rect -141 2198 -94 2262
rect -30 2198 -14 2262
rect -141 2182 -14 2198
rect -141 2118 -94 2182
rect -30 2118 -14 2182
rect -141 2102 -14 2118
rect -141 2038 -94 2102
rect -30 2038 -14 2102
rect -141 2022 -14 2038
rect -141 1958 -94 2022
rect -30 1958 -14 2022
rect -141 1942 -14 1958
rect -141 1878 -94 1942
rect -30 1878 -14 1942
rect -141 1862 -14 1878
rect -141 1798 -94 1862
rect -30 1798 -14 1862
rect -141 1782 -14 1798
rect -141 1718 -94 1782
rect -30 1718 -14 1782
rect -141 1702 -14 1718
rect -141 1638 -94 1702
rect -30 1638 -14 1702
rect -141 1622 -14 1638
rect -141 1558 -94 1622
rect -30 1558 -14 1622
rect -141 1542 -14 1558
rect -141 1478 -94 1542
rect -30 1478 -14 1542
rect -141 1462 -14 1478
rect -141 1398 -94 1462
rect -30 1398 -14 1462
rect -141 1362 -14 1398
rect 209 2382 1131 2600
rect 209 1518 238 2382
rect 1102 1518 1131 2382
rect -141 1238 -37 1362
rect -141 1202 -14 1238
rect -141 1138 -94 1202
rect -30 1138 -14 1202
rect -141 1122 -14 1138
rect -141 1058 -94 1122
rect -30 1058 -14 1122
rect -141 1042 -14 1058
rect -141 978 -94 1042
rect -30 978 -14 1042
rect -141 962 -14 978
rect -141 898 -94 962
rect -30 898 -14 962
rect -141 882 -14 898
rect -141 818 -94 882
rect -30 818 -14 882
rect -141 802 -14 818
rect -141 738 -94 802
rect -30 738 -14 802
rect -141 722 -14 738
rect -141 658 -94 722
rect -30 658 -14 722
rect -141 642 -14 658
rect -141 578 -94 642
rect -30 578 -14 642
rect -141 562 -14 578
rect -141 498 -94 562
rect -30 498 -14 562
rect -141 482 -14 498
rect -141 418 -94 482
rect -30 418 -14 482
rect -141 402 -14 418
rect -141 338 -94 402
rect -30 338 -14 402
rect -141 322 -14 338
rect -141 258 -94 322
rect -30 258 -14 322
rect -141 242 -14 258
rect -141 178 -94 242
rect -30 178 -14 242
rect -141 162 -14 178
rect -141 98 -94 162
rect -30 98 -14 162
rect -141 62 -14 98
rect 209 1082 1131 1518
rect 209 218 238 1082
rect 1102 218 1131 1082
rect -141 -62 -37 62
rect -141 -98 -14 -62
rect -141 -162 -94 -98
rect -30 -162 -14 -98
rect -141 -178 -14 -162
rect -141 -242 -94 -178
rect -30 -242 -14 -178
rect -141 -258 -14 -242
rect -141 -322 -94 -258
rect -30 -322 -14 -258
rect -141 -338 -14 -322
rect -141 -402 -94 -338
rect -30 -402 -14 -338
rect -141 -418 -14 -402
rect -141 -482 -94 -418
rect -30 -482 -14 -418
rect -141 -498 -14 -482
rect -141 -562 -94 -498
rect -30 -562 -14 -498
rect -141 -578 -14 -562
rect -141 -642 -94 -578
rect -30 -642 -14 -578
rect -141 -658 -14 -642
rect -141 -722 -94 -658
rect -30 -722 -14 -658
rect -141 -738 -14 -722
rect -141 -802 -94 -738
rect -30 -802 -14 -738
rect -141 -818 -14 -802
rect -141 -882 -94 -818
rect -30 -882 -14 -818
rect -141 -898 -14 -882
rect -141 -962 -94 -898
rect -30 -962 -14 -898
rect -141 -978 -14 -962
rect -141 -1042 -94 -978
rect -30 -1042 -14 -978
rect -141 -1058 -14 -1042
rect -141 -1122 -94 -1058
rect -30 -1122 -14 -1058
rect -141 -1138 -14 -1122
rect -141 -1202 -94 -1138
rect -30 -1202 -14 -1138
rect -141 -1238 -14 -1202
rect 209 -218 1131 218
rect 209 -1082 238 -218
rect 1102 -1082 1131 -218
rect -141 -1362 -37 -1238
rect -141 -1398 -14 -1362
rect -141 -1462 -94 -1398
rect -30 -1462 -14 -1398
rect -141 -1478 -14 -1462
rect -141 -1542 -94 -1478
rect -30 -1542 -14 -1478
rect -141 -1558 -14 -1542
rect -141 -1622 -94 -1558
rect -30 -1622 -14 -1558
rect -141 -1638 -14 -1622
rect -141 -1702 -94 -1638
rect -30 -1702 -14 -1638
rect -141 -1718 -14 -1702
rect -141 -1782 -94 -1718
rect -30 -1782 -14 -1718
rect -141 -1798 -14 -1782
rect -141 -1862 -94 -1798
rect -30 -1862 -14 -1798
rect -141 -1878 -14 -1862
rect -141 -1942 -94 -1878
rect -30 -1942 -14 -1878
rect -141 -1958 -14 -1942
rect -141 -2022 -94 -1958
rect -30 -2022 -14 -1958
rect -141 -2038 -14 -2022
rect -141 -2102 -94 -2038
rect -30 -2102 -14 -2038
rect -141 -2118 -14 -2102
rect -141 -2182 -94 -2118
rect -30 -2182 -14 -2118
rect -141 -2198 -14 -2182
rect -141 -2262 -94 -2198
rect -30 -2262 -14 -2198
rect -141 -2278 -14 -2262
rect -141 -2342 -94 -2278
rect -30 -2342 -14 -2278
rect -141 -2358 -14 -2342
rect -141 -2422 -94 -2358
rect -30 -2422 -14 -2358
rect -141 -2438 -14 -2422
rect -141 -2502 -94 -2438
rect -30 -2502 -14 -2438
rect -141 -2538 -14 -2502
rect 209 -1518 1131 -1082
rect 209 -2382 238 -1518
rect 1102 -2382 1131 -1518
rect -141 -2600 -37 -2538
rect 209 -2917 1131 -2382
rect 1238 2538 1342 2600
rect 1238 2502 1365 2538
rect 1238 2438 1285 2502
rect 1349 2438 1365 2502
rect 1238 2422 1365 2438
rect 1238 2358 1285 2422
rect 1349 2358 1365 2422
rect 1238 2342 1365 2358
rect 1238 2278 1285 2342
rect 1349 2278 1365 2342
rect 1238 2262 1365 2278
rect 1238 2198 1285 2262
rect 1349 2198 1365 2262
rect 1238 2182 1365 2198
rect 1238 2118 1285 2182
rect 1349 2118 1365 2182
rect 1238 2102 1365 2118
rect 1238 2038 1285 2102
rect 1349 2038 1365 2102
rect 1238 2022 1365 2038
rect 1238 1958 1285 2022
rect 1349 1958 1365 2022
rect 1238 1942 1365 1958
rect 1238 1878 1285 1942
rect 1349 1878 1365 1942
rect 1238 1862 1365 1878
rect 1238 1798 1285 1862
rect 1349 1798 1365 1862
rect 1238 1782 1365 1798
rect 1238 1718 1285 1782
rect 1349 1718 1365 1782
rect 1238 1702 1365 1718
rect 1238 1638 1285 1702
rect 1349 1638 1365 1702
rect 1238 1622 1365 1638
rect 1238 1558 1285 1622
rect 1349 1558 1365 1622
rect 1238 1542 1365 1558
rect 1238 1478 1285 1542
rect 1349 1478 1365 1542
rect 1238 1462 1365 1478
rect 1238 1398 1285 1462
rect 1349 1398 1365 1462
rect 1238 1362 1365 1398
rect 1588 2382 2510 2600
rect 1588 1518 1617 2382
rect 2481 1518 2510 2382
rect 1238 1238 1342 1362
rect 1238 1202 1365 1238
rect 1238 1138 1285 1202
rect 1349 1138 1365 1202
rect 1238 1122 1365 1138
rect 1238 1058 1285 1122
rect 1349 1058 1365 1122
rect 1238 1042 1365 1058
rect 1238 978 1285 1042
rect 1349 978 1365 1042
rect 1238 962 1365 978
rect 1238 898 1285 962
rect 1349 898 1365 962
rect 1238 882 1365 898
rect 1238 818 1285 882
rect 1349 818 1365 882
rect 1238 802 1365 818
rect 1238 738 1285 802
rect 1349 738 1365 802
rect 1238 722 1365 738
rect 1238 658 1285 722
rect 1349 658 1365 722
rect 1238 642 1365 658
rect 1238 578 1285 642
rect 1349 578 1365 642
rect 1238 562 1365 578
rect 1238 498 1285 562
rect 1349 498 1365 562
rect 1238 482 1365 498
rect 1238 418 1285 482
rect 1349 418 1365 482
rect 1238 402 1365 418
rect 1238 338 1285 402
rect 1349 338 1365 402
rect 1238 322 1365 338
rect 1238 258 1285 322
rect 1349 258 1365 322
rect 1238 242 1365 258
rect 1238 178 1285 242
rect 1349 178 1365 242
rect 1238 162 1365 178
rect 1238 98 1285 162
rect 1349 98 1365 162
rect 1238 62 1365 98
rect 1588 1082 2510 1518
rect 1588 218 1617 1082
rect 2481 218 2510 1082
rect 1238 -62 1342 62
rect 1238 -98 1365 -62
rect 1238 -162 1285 -98
rect 1349 -162 1365 -98
rect 1238 -178 1365 -162
rect 1238 -242 1285 -178
rect 1349 -242 1365 -178
rect 1238 -258 1365 -242
rect 1238 -322 1285 -258
rect 1349 -322 1365 -258
rect 1238 -338 1365 -322
rect 1238 -402 1285 -338
rect 1349 -402 1365 -338
rect 1238 -418 1365 -402
rect 1238 -482 1285 -418
rect 1349 -482 1365 -418
rect 1238 -498 1365 -482
rect 1238 -562 1285 -498
rect 1349 -562 1365 -498
rect 1238 -578 1365 -562
rect 1238 -642 1285 -578
rect 1349 -642 1365 -578
rect 1238 -658 1365 -642
rect 1238 -722 1285 -658
rect 1349 -722 1365 -658
rect 1238 -738 1365 -722
rect 1238 -802 1285 -738
rect 1349 -802 1365 -738
rect 1238 -818 1365 -802
rect 1238 -882 1285 -818
rect 1349 -882 1365 -818
rect 1238 -898 1365 -882
rect 1238 -962 1285 -898
rect 1349 -962 1365 -898
rect 1238 -978 1365 -962
rect 1238 -1042 1285 -978
rect 1349 -1042 1365 -978
rect 1238 -1058 1365 -1042
rect 1238 -1122 1285 -1058
rect 1349 -1122 1365 -1058
rect 1238 -1138 1365 -1122
rect 1238 -1202 1285 -1138
rect 1349 -1202 1365 -1138
rect 1238 -1238 1365 -1202
rect 1588 -218 2510 218
rect 1588 -1082 1617 -218
rect 2481 -1082 2510 -218
rect 1238 -1362 1342 -1238
rect 1238 -1398 1365 -1362
rect 1238 -1462 1285 -1398
rect 1349 -1462 1365 -1398
rect 1238 -1478 1365 -1462
rect 1238 -1542 1285 -1478
rect 1349 -1542 1365 -1478
rect 1238 -1558 1365 -1542
rect 1238 -1622 1285 -1558
rect 1349 -1622 1365 -1558
rect 1238 -1638 1365 -1622
rect 1238 -1702 1285 -1638
rect 1349 -1702 1365 -1638
rect 1238 -1718 1365 -1702
rect 1238 -1782 1285 -1718
rect 1349 -1782 1365 -1718
rect 1238 -1798 1365 -1782
rect 1238 -1862 1285 -1798
rect 1349 -1862 1365 -1798
rect 1238 -1878 1365 -1862
rect 1238 -1942 1285 -1878
rect 1349 -1942 1365 -1878
rect 1238 -1958 1365 -1942
rect 1238 -2022 1285 -1958
rect 1349 -2022 1365 -1958
rect 1238 -2038 1365 -2022
rect 1238 -2102 1285 -2038
rect 1349 -2102 1365 -2038
rect 1238 -2118 1365 -2102
rect 1238 -2182 1285 -2118
rect 1349 -2182 1365 -2118
rect 1238 -2198 1365 -2182
rect 1238 -2262 1285 -2198
rect 1349 -2262 1365 -2198
rect 1238 -2278 1365 -2262
rect 1238 -2342 1285 -2278
rect 1349 -2342 1365 -2278
rect 1238 -2358 1365 -2342
rect 1238 -2422 1285 -2358
rect 1349 -2422 1365 -2358
rect 1238 -2438 1365 -2422
rect 1238 -2502 1285 -2438
rect 1349 -2502 1365 -2438
rect 1238 -2538 1365 -2502
rect 1588 -1518 2510 -1082
rect 1588 -2382 1617 -1518
rect 2481 -2382 2510 -1518
rect 1238 -2600 1342 -2538
rect 1588 -2945 2510 -2382
rect 2617 2538 2721 2600
rect 2617 2502 2744 2538
rect 2617 2438 2664 2502
rect 2728 2438 2744 2502
rect 2617 2422 2744 2438
rect 2617 2358 2664 2422
rect 2728 2358 2744 2422
rect 2617 2342 2744 2358
rect 2617 2278 2664 2342
rect 2728 2278 2744 2342
rect 2617 2262 2744 2278
rect 2617 2198 2664 2262
rect 2728 2198 2744 2262
rect 2617 2182 2744 2198
rect 2617 2118 2664 2182
rect 2728 2118 2744 2182
rect 2617 2102 2744 2118
rect 2617 2038 2664 2102
rect 2728 2038 2744 2102
rect 2617 2022 2744 2038
rect 2617 1958 2664 2022
rect 2728 1958 2744 2022
rect 2617 1942 2744 1958
rect 2617 1878 2664 1942
rect 2728 1878 2744 1942
rect 2617 1862 2744 1878
rect 2617 1798 2664 1862
rect 2728 1798 2744 1862
rect 2617 1782 2744 1798
rect 2617 1718 2664 1782
rect 2728 1718 2744 1782
rect 2617 1702 2744 1718
rect 2617 1638 2664 1702
rect 2728 1638 2744 1702
rect 2617 1622 2744 1638
rect 2617 1558 2664 1622
rect 2728 1558 2744 1622
rect 2617 1542 2744 1558
rect 2617 1478 2664 1542
rect 2728 1478 2744 1542
rect 2617 1462 2744 1478
rect 2617 1398 2664 1462
rect 2728 1398 2744 1462
rect 2617 1362 2744 1398
rect 2617 1238 2721 1362
rect 2617 1202 2744 1238
rect 2617 1138 2664 1202
rect 2728 1138 2744 1202
rect 2617 1122 2744 1138
rect 2617 1058 2664 1122
rect 2728 1058 2744 1122
rect 2617 1042 2744 1058
rect 2617 978 2664 1042
rect 2728 978 2744 1042
rect 2617 962 2744 978
rect 2617 898 2664 962
rect 2728 898 2744 962
rect 2617 882 2744 898
rect 2617 818 2664 882
rect 2728 818 2744 882
rect 2617 802 2744 818
rect 2617 738 2664 802
rect 2728 738 2744 802
rect 2617 722 2744 738
rect 2617 658 2664 722
rect 2728 658 2744 722
rect 2617 642 2744 658
rect 2617 578 2664 642
rect 2728 578 2744 642
rect 2617 562 2744 578
rect 2617 498 2664 562
rect 2728 498 2744 562
rect 2617 482 2744 498
rect 2617 418 2664 482
rect 2728 418 2744 482
rect 2617 402 2744 418
rect 2617 338 2664 402
rect 2728 338 2744 402
rect 2617 322 2744 338
rect 2617 258 2664 322
rect 2728 258 2744 322
rect 2617 242 2744 258
rect 2617 178 2664 242
rect 2728 178 2744 242
rect 2617 162 2744 178
rect 2617 98 2664 162
rect 2728 98 2744 162
rect 2617 62 2744 98
rect 2617 -62 2721 62
rect 2617 -98 2744 -62
rect 2617 -162 2664 -98
rect 2728 -162 2744 -98
rect 2617 -178 2744 -162
rect 2617 -242 2664 -178
rect 2728 -242 2744 -178
rect 2617 -258 2744 -242
rect 2617 -322 2664 -258
rect 2728 -322 2744 -258
rect 2617 -338 2744 -322
rect 2617 -402 2664 -338
rect 2728 -402 2744 -338
rect 2617 -418 2744 -402
rect 2617 -482 2664 -418
rect 2728 -482 2744 -418
rect 2617 -498 2744 -482
rect 2617 -562 2664 -498
rect 2728 -562 2744 -498
rect 2617 -578 2744 -562
rect 2617 -642 2664 -578
rect 2728 -642 2744 -578
rect 2617 -658 2744 -642
rect 2617 -722 2664 -658
rect 2728 -722 2744 -658
rect 2617 -738 2744 -722
rect 2617 -802 2664 -738
rect 2728 -802 2744 -738
rect 2617 -818 2744 -802
rect 2617 -882 2664 -818
rect 2728 -882 2744 -818
rect 2617 -898 2744 -882
rect 2617 -962 2664 -898
rect 2728 -962 2744 -898
rect 2617 -978 2744 -962
rect 2617 -1042 2664 -978
rect 2728 -1042 2744 -978
rect 2617 -1058 2744 -1042
rect 2617 -1122 2664 -1058
rect 2728 -1122 2744 -1058
rect 2617 -1138 2744 -1122
rect 2617 -1202 2664 -1138
rect 2728 -1202 2744 -1138
rect 2617 -1238 2744 -1202
rect 2617 -1362 2721 -1238
rect 2617 -1398 2744 -1362
rect 2617 -1462 2664 -1398
rect 2728 -1462 2744 -1398
rect 2617 -1478 2744 -1462
rect 2617 -1542 2664 -1478
rect 2728 -1542 2744 -1478
rect 2617 -1558 2744 -1542
rect 2617 -1622 2664 -1558
rect 2728 -1622 2744 -1558
rect 2617 -1638 2744 -1622
rect 2617 -1702 2664 -1638
rect 2728 -1702 2744 -1638
rect 2617 -1718 2744 -1702
rect 2617 -1782 2664 -1718
rect 2728 -1782 2744 -1718
rect 2617 -1798 2744 -1782
rect 2617 -1862 2664 -1798
rect 2728 -1862 2744 -1798
rect 2617 -1878 2744 -1862
rect 2617 -1942 2664 -1878
rect 2728 -1942 2744 -1878
rect 2617 -1958 2744 -1942
rect 2617 -2022 2664 -1958
rect 2728 -2022 2744 -1958
rect 2617 -2038 2744 -2022
rect 2617 -2102 2664 -2038
rect 2728 -2102 2744 -2038
rect 2617 -2118 2744 -2102
rect 2617 -2182 2664 -2118
rect 2728 -2182 2744 -2118
rect 2617 -2198 2744 -2182
rect 2617 -2262 2664 -2198
rect 2728 -2262 2744 -2198
rect 2617 -2278 2744 -2262
rect 2617 -2342 2664 -2278
rect 2728 -2342 2744 -2278
rect 2617 -2358 2744 -2342
rect 2617 -2422 2664 -2358
rect 2728 -2422 2744 -2358
rect 2617 -2438 2744 -2422
rect 2617 -2502 2664 -2438
rect 2728 -2502 2744 -2438
rect 2617 -2538 2744 -2502
rect 2617 -2600 2721 -2538
<< properties >>
string FIXED_BBOX 1329 1350 2529 2550
<< end >>
