magic
tech sky130A
timestamp 1664679546
<< nwell >>
rect -62 -61 62 61
<< pmos >>
rect -15 -30 15 30
<< pdiff >>
rect -44 24 -15 30
rect -44 -24 -38 24
rect -21 -24 -15 24
rect -44 -30 -15 -24
rect 15 24 44 30
rect 15 -24 21 24
rect 38 -24 44 24
rect 15 -30 44 -24
<< pdiffc >>
rect -38 -24 -21 24
rect 21 -24 38 24
<< poly >>
rect -15 30 15 43
rect -15 -43 15 -30
<< locali >>
rect -38 24 -21 32
rect -38 -32 -21 -24
rect 21 24 38 32
rect 21 -32 38 -24
<< viali >>
rect -38 -24 -21 24
rect 21 -24 38 24
<< metal1 >>
rect -41 24 -18 30
rect -41 -24 -38 24
rect -21 -24 -18 24
rect -41 -30 -18 -24
rect 18 24 41 30
rect 18 -24 21 24
rect 38 -24 41 24
rect 18 -30 41 -24
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.6 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
