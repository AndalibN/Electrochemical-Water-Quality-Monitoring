magic
tech sky130A
timestamp 1667954557
<< nmos >>
rect -15 -175 15 175
<< ndiff >>
rect -44 169 -15 175
rect -44 -169 -38 169
rect -21 -169 -15 169
rect -44 -175 -15 -169
rect 15 169 44 175
rect 15 -169 21 169
rect 38 -169 44 169
rect 15 -175 44 -169
<< ndiffc >>
rect -38 -169 -21 169
rect 21 -169 38 169
<< poly >>
rect -15 175 15 188
rect -15 -188 15 -175
<< locali >>
rect -38 169 -21 177
rect -38 -177 -21 -169
rect 21 169 38 177
rect 21 -177 38 -169
<< viali >>
rect -38 -169 -21 169
rect 21 -169 38 169
<< metal1 >>
rect -41 169 -18 175
rect -41 -169 -38 169
rect -21 -169 -18 169
rect -41 -175 -18 -169
rect 18 169 41 175
rect 18 -169 21 169
rect 38 -169 41 169
rect 18 -175 41 -169
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.5 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
