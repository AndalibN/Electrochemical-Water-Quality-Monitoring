magic
tech sky130A
magscale 1 2
timestamp 1666398315
<< nwell >>
rect 750 2052 1598 2236
rect 1550 1618 1574 1620
rect 1516 1586 1540 1590
<< psubdiff >>
rect 750 1040 1598 1054
rect 750 996 792 1040
rect 1548 996 1598 1040
rect 750 978 1598 996
<< nsubdiff >>
rect 786 2174 1562 2200
rect 786 2140 806 2174
rect 1542 2140 1562 2174
rect 786 2110 1562 2140
<< psubdiffcont >>
rect 792 996 1548 1040
<< nsubdiffcont >>
rect 806 2140 1542 2174
<< poly >>
rect 860 1344 928 1544
rect 1140 1344 1208 1544
rect 1420 1344 1488 1544
<< locali >>
rect 788 2174 1558 2182
rect 788 2140 806 2174
rect 1542 2140 1558 2174
rect 788 2130 1558 2140
rect 798 1964 832 2130
rect 1078 1960 1112 2130
rect 1358 1966 1392 2130
rect 978 1380 1012 1620
rect 1262 1380 1296 1620
rect 1550 1618 1574 1620
rect 1540 1590 1574 1618
rect 1516 1586 1574 1590
rect 1540 1380 1574 1586
rect 750 1346 942 1380
rect 978 1346 1226 1380
rect 1262 1346 1506 1380
rect 1540 1346 1598 1380
rect 978 1312 1012 1346
rect 1262 1312 1296 1346
rect 1540 1312 1574 1346
rect 954 1278 1012 1312
rect 1238 1308 1296 1312
rect 1238 1276 1260 1308
rect 1262 1278 1296 1308
rect 1518 1276 1574 1312
rect 796 1042 830 1130
rect 1080 1042 1114 1136
rect 1360 1042 1394 1132
rect 776 1040 1582 1042
rect 776 996 792 1040
rect 1548 996 1582 1040
<< metal1 >>
rect 978 1380 1012 1620
rect 1262 1380 1296 1620
rect 1550 1618 1574 1620
rect 1540 1590 1574 1618
rect 1516 1586 1574 1590
rect 1540 1380 1574 1586
rect 750 1346 942 1380
rect 978 1346 1226 1380
rect 1262 1346 1506 1380
rect 1540 1346 1598 1380
rect 978 1312 1012 1346
rect 1262 1312 1296 1346
rect 1540 1312 1574 1346
rect 954 1278 1012 1312
rect 1238 1308 1296 1312
rect 1238 1276 1260 1308
rect 1262 1278 1296 1308
rect 1518 1276 1574 1312
use sky130_fd_pr__pfet_01v8_G3UWY6  XM1
timestamp 1666397798
transform 1 0 894 0 1 1754
box -144 -264 144 298
use sky130_fd_pr__pfet_01v8_G3UWY6  XM2
timestamp 1666397798
transform 1 0 1174 0 1 1754
box -144 -264 144 298
use sky130_fd_pr__nfet_01v8_N5USK7  XM4
timestamp 1666397798
transform 1 0 892 0 1 1239
box -108 -157 108 157
use sky130_fd_pr__nfet_01v8_WSTS35  XM6
timestamp 1666397798
transform -1 0 1456 0 1 1239
box -108 -157 108 157
use sky130_fd_pr__nfet_01v8_N5USK7  sky130_fd_pr__nfet_01v8_N5USK7_0
timestamp 1666397798
transform 1 0 1176 0 1 1239
box -108 -157 108 157
use sky130_fd_pr__pfet_01v8_G3UWY6  sky130_fd_pr__pfet_01v8_G3UWY6_0
timestamp 1666397798
transform 1 0 1454 0 1 1754
box -144 -264 144 298
<< labels >>
rlabel metal1 1598 1362 1598 1362 3 OUT
port 1 e
rlabel metal1 750 1362 750 1362 7 IN
port 2 w
rlabel psubdiffcont 804 1018 804 1018 7 GND
port 3 w
rlabel nsubdiffcont 828 2158 828 2158 7 VDD
port 4 w
<< end >>
