magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -184 -1457 184 1395
<< nmos >>
rect -100 -1431 100 1369
<< ndiff >>
rect -158 1346 -100 1369
rect -158 1312 -146 1346
rect -112 1312 -100 1346
rect -158 1278 -100 1312
rect -158 1244 -146 1278
rect -112 1244 -100 1278
rect -158 1210 -100 1244
rect -158 1176 -146 1210
rect -112 1176 -100 1210
rect -158 1142 -100 1176
rect -158 1108 -146 1142
rect -112 1108 -100 1142
rect -158 1074 -100 1108
rect -158 1040 -146 1074
rect -112 1040 -100 1074
rect -158 1006 -100 1040
rect -158 972 -146 1006
rect -112 972 -100 1006
rect -158 938 -100 972
rect -158 904 -146 938
rect -112 904 -100 938
rect -158 870 -100 904
rect -158 836 -146 870
rect -112 836 -100 870
rect -158 802 -100 836
rect -158 768 -146 802
rect -112 768 -100 802
rect -158 734 -100 768
rect -158 700 -146 734
rect -112 700 -100 734
rect -158 666 -100 700
rect -158 632 -146 666
rect -112 632 -100 666
rect -158 598 -100 632
rect -158 564 -146 598
rect -112 564 -100 598
rect -158 530 -100 564
rect -158 496 -146 530
rect -112 496 -100 530
rect -158 462 -100 496
rect -158 428 -146 462
rect -112 428 -100 462
rect -158 394 -100 428
rect -158 360 -146 394
rect -112 360 -100 394
rect -158 326 -100 360
rect -158 292 -146 326
rect -112 292 -100 326
rect -158 258 -100 292
rect -158 224 -146 258
rect -112 224 -100 258
rect -158 190 -100 224
rect -158 156 -146 190
rect -112 156 -100 190
rect -158 122 -100 156
rect -158 88 -146 122
rect -112 88 -100 122
rect -158 54 -100 88
rect -158 20 -146 54
rect -112 20 -100 54
rect -158 -14 -100 20
rect -158 -48 -146 -14
rect -112 -48 -100 -14
rect -158 -82 -100 -48
rect -158 -116 -146 -82
rect -112 -116 -100 -82
rect -158 -150 -100 -116
rect -158 -184 -146 -150
rect -112 -184 -100 -150
rect -158 -218 -100 -184
rect -158 -252 -146 -218
rect -112 -252 -100 -218
rect -158 -286 -100 -252
rect -158 -320 -146 -286
rect -112 -320 -100 -286
rect -158 -354 -100 -320
rect -158 -388 -146 -354
rect -112 -388 -100 -354
rect -158 -422 -100 -388
rect -158 -456 -146 -422
rect -112 -456 -100 -422
rect -158 -490 -100 -456
rect -158 -524 -146 -490
rect -112 -524 -100 -490
rect -158 -558 -100 -524
rect -158 -592 -146 -558
rect -112 -592 -100 -558
rect -158 -626 -100 -592
rect -158 -660 -146 -626
rect -112 -660 -100 -626
rect -158 -694 -100 -660
rect -158 -728 -146 -694
rect -112 -728 -100 -694
rect -158 -762 -100 -728
rect -158 -796 -146 -762
rect -112 -796 -100 -762
rect -158 -830 -100 -796
rect -158 -864 -146 -830
rect -112 -864 -100 -830
rect -158 -898 -100 -864
rect -158 -932 -146 -898
rect -112 -932 -100 -898
rect -158 -966 -100 -932
rect -158 -1000 -146 -966
rect -112 -1000 -100 -966
rect -158 -1034 -100 -1000
rect -158 -1068 -146 -1034
rect -112 -1068 -100 -1034
rect -158 -1102 -100 -1068
rect -158 -1136 -146 -1102
rect -112 -1136 -100 -1102
rect -158 -1170 -100 -1136
rect -158 -1204 -146 -1170
rect -112 -1204 -100 -1170
rect -158 -1238 -100 -1204
rect -158 -1272 -146 -1238
rect -112 -1272 -100 -1238
rect -158 -1306 -100 -1272
rect -158 -1340 -146 -1306
rect -112 -1340 -100 -1306
rect -158 -1374 -100 -1340
rect -158 -1408 -146 -1374
rect -112 -1408 -100 -1374
rect -158 -1431 -100 -1408
rect 100 1346 158 1369
rect 100 1312 112 1346
rect 146 1312 158 1346
rect 100 1278 158 1312
rect 100 1244 112 1278
rect 146 1244 158 1278
rect 100 1210 158 1244
rect 100 1176 112 1210
rect 146 1176 158 1210
rect 100 1142 158 1176
rect 100 1108 112 1142
rect 146 1108 158 1142
rect 100 1074 158 1108
rect 100 1040 112 1074
rect 146 1040 158 1074
rect 100 1006 158 1040
rect 100 972 112 1006
rect 146 972 158 1006
rect 100 938 158 972
rect 100 904 112 938
rect 146 904 158 938
rect 100 870 158 904
rect 100 836 112 870
rect 146 836 158 870
rect 100 802 158 836
rect 100 768 112 802
rect 146 768 158 802
rect 100 734 158 768
rect 100 700 112 734
rect 146 700 158 734
rect 100 666 158 700
rect 100 632 112 666
rect 146 632 158 666
rect 100 598 158 632
rect 100 564 112 598
rect 146 564 158 598
rect 100 530 158 564
rect 100 496 112 530
rect 146 496 158 530
rect 100 462 158 496
rect 100 428 112 462
rect 146 428 158 462
rect 100 394 158 428
rect 100 360 112 394
rect 146 360 158 394
rect 100 326 158 360
rect 100 292 112 326
rect 146 292 158 326
rect 100 258 158 292
rect 100 224 112 258
rect 146 224 158 258
rect 100 190 158 224
rect 100 156 112 190
rect 146 156 158 190
rect 100 122 158 156
rect 100 88 112 122
rect 146 88 158 122
rect 100 54 158 88
rect 100 20 112 54
rect 146 20 158 54
rect 100 -14 158 20
rect 100 -48 112 -14
rect 146 -48 158 -14
rect 100 -82 158 -48
rect 100 -116 112 -82
rect 146 -116 158 -82
rect 100 -150 158 -116
rect 100 -184 112 -150
rect 146 -184 158 -150
rect 100 -218 158 -184
rect 100 -252 112 -218
rect 146 -252 158 -218
rect 100 -286 158 -252
rect 100 -320 112 -286
rect 146 -320 158 -286
rect 100 -354 158 -320
rect 100 -388 112 -354
rect 146 -388 158 -354
rect 100 -422 158 -388
rect 100 -456 112 -422
rect 146 -456 158 -422
rect 100 -490 158 -456
rect 100 -524 112 -490
rect 146 -524 158 -490
rect 100 -558 158 -524
rect 100 -592 112 -558
rect 146 -592 158 -558
rect 100 -626 158 -592
rect 100 -660 112 -626
rect 146 -660 158 -626
rect 100 -694 158 -660
rect 100 -728 112 -694
rect 146 -728 158 -694
rect 100 -762 158 -728
rect 100 -796 112 -762
rect 146 -796 158 -762
rect 100 -830 158 -796
rect 100 -864 112 -830
rect 146 -864 158 -830
rect 100 -898 158 -864
rect 100 -932 112 -898
rect 146 -932 158 -898
rect 100 -966 158 -932
rect 100 -1000 112 -966
rect 146 -1000 158 -966
rect 100 -1034 158 -1000
rect 100 -1068 112 -1034
rect 146 -1068 158 -1034
rect 100 -1102 158 -1068
rect 100 -1136 112 -1102
rect 146 -1136 158 -1102
rect 100 -1170 158 -1136
rect 100 -1204 112 -1170
rect 146 -1204 158 -1170
rect 100 -1238 158 -1204
rect 100 -1272 112 -1238
rect 146 -1272 158 -1238
rect 100 -1306 158 -1272
rect 100 -1340 112 -1306
rect 146 -1340 158 -1306
rect 100 -1374 158 -1340
rect 100 -1408 112 -1374
rect 146 -1408 158 -1374
rect 100 -1431 158 -1408
<< ndiffc >>
rect -146 1312 -112 1346
rect -146 1244 -112 1278
rect -146 1176 -112 1210
rect -146 1108 -112 1142
rect -146 1040 -112 1074
rect -146 972 -112 1006
rect -146 904 -112 938
rect -146 836 -112 870
rect -146 768 -112 802
rect -146 700 -112 734
rect -146 632 -112 666
rect -146 564 -112 598
rect -146 496 -112 530
rect -146 428 -112 462
rect -146 360 -112 394
rect -146 292 -112 326
rect -146 224 -112 258
rect -146 156 -112 190
rect -146 88 -112 122
rect -146 20 -112 54
rect -146 -48 -112 -14
rect -146 -116 -112 -82
rect -146 -184 -112 -150
rect -146 -252 -112 -218
rect -146 -320 -112 -286
rect -146 -388 -112 -354
rect -146 -456 -112 -422
rect -146 -524 -112 -490
rect -146 -592 -112 -558
rect -146 -660 -112 -626
rect -146 -728 -112 -694
rect -146 -796 -112 -762
rect -146 -864 -112 -830
rect -146 -932 -112 -898
rect -146 -1000 -112 -966
rect -146 -1068 -112 -1034
rect -146 -1136 -112 -1102
rect -146 -1204 -112 -1170
rect -146 -1272 -112 -1238
rect -146 -1340 -112 -1306
rect -146 -1408 -112 -1374
rect 112 1312 146 1346
rect 112 1244 146 1278
rect 112 1176 146 1210
rect 112 1108 146 1142
rect 112 1040 146 1074
rect 112 972 146 1006
rect 112 904 146 938
rect 112 836 146 870
rect 112 768 146 802
rect 112 700 146 734
rect 112 632 146 666
rect 112 564 146 598
rect 112 496 146 530
rect 112 428 146 462
rect 112 360 146 394
rect 112 292 146 326
rect 112 224 146 258
rect 112 156 146 190
rect 112 88 146 122
rect 112 20 146 54
rect 112 -48 146 -14
rect 112 -116 146 -82
rect 112 -184 146 -150
rect 112 -252 146 -218
rect 112 -320 146 -286
rect 112 -388 146 -354
rect 112 -456 146 -422
rect 112 -524 146 -490
rect 112 -592 146 -558
rect 112 -660 146 -626
rect 112 -728 146 -694
rect 112 -796 146 -762
rect 112 -864 146 -830
rect 112 -932 146 -898
rect 112 -1000 146 -966
rect 112 -1068 146 -1034
rect 112 -1136 146 -1102
rect 112 -1204 146 -1170
rect 112 -1272 146 -1238
rect 112 -1340 146 -1306
rect 112 -1408 146 -1374
<< poly >>
rect -100 1441 100 1457
rect -100 1407 -51 1441
rect -17 1407 17 1441
rect 51 1407 100 1441
rect -100 1369 100 1407
rect -100 -1457 100 -1431
<< polycont >>
rect -51 1407 -17 1441
rect 17 1407 51 1441
<< locali >>
rect -100 1407 -53 1441
rect -17 1407 17 1441
rect 53 1407 100 1441
rect -146 1354 -112 1373
rect -146 1282 -112 1312
rect -146 1210 -112 1244
rect -146 1142 -112 1176
rect -146 1074 -112 1104
rect -146 1006 -112 1032
rect -146 938 -112 960
rect -146 870 -112 888
rect -146 802 -112 816
rect -146 734 -112 744
rect -146 666 -112 672
rect -146 598 -112 600
rect -146 562 -112 564
rect -146 490 -112 496
rect -146 418 -112 428
rect -146 346 -112 360
rect -146 274 -112 292
rect -146 202 -112 224
rect -146 130 -112 156
rect -146 58 -112 88
rect -146 -14 -112 20
rect -146 -82 -112 -48
rect -146 -150 -112 -120
rect -146 -218 -112 -192
rect -146 -286 -112 -264
rect -146 -354 -112 -336
rect -146 -422 -112 -408
rect -146 -490 -112 -480
rect -146 -558 -112 -552
rect -146 -626 -112 -624
rect -146 -662 -112 -660
rect -146 -734 -112 -728
rect -146 -806 -112 -796
rect -146 -878 -112 -864
rect -146 -950 -112 -932
rect -146 -1022 -112 -1000
rect -146 -1094 -112 -1068
rect -146 -1166 -112 -1136
rect -146 -1238 -112 -1204
rect -146 -1306 -112 -1272
rect -146 -1374 -112 -1344
rect -146 -1435 -112 -1416
rect 112 1354 146 1373
rect 112 1282 146 1312
rect 112 1210 146 1244
rect 112 1142 146 1176
rect 112 1074 146 1104
rect 112 1006 146 1032
rect 112 938 146 960
rect 112 870 146 888
rect 112 802 146 816
rect 112 734 146 744
rect 112 666 146 672
rect 112 598 146 600
rect 112 562 146 564
rect 112 490 146 496
rect 112 418 146 428
rect 112 346 146 360
rect 112 274 146 292
rect 112 202 146 224
rect 112 130 146 156
rect 112 58 146 88
rect 112 -14 146 20
rect 112 -82 146 -48
rect 112 -150 146 -120
rect 112 -218 146 -192
rect 112 -286 146 -264
rect 112 -354 146 -336
rect 112 -422 146 -408
rect 112 -490 146 -480
rect 112 -558 146 -552
rect 112 -626 146 -624
rect 112 -662 146 -660
rect 112 -734 146 -728
rect 112 -806 146 -796
rect 112 -878 146 -864
rect 112 -950 146 -932
rect 112 -1022 146 -1000
rect 112 -1094 146 -1068
rect 112 -1166 146 -1136
rect 112 -1238 146 -1204
rect 112 -1306 146 -1272
rect 112 -1374 146 -1344
rect 112 -1435 146 -1416
<< viali >>
rect -53 1407 -51 1441
rect -51 1407 -19 1441
rect 19 1407 51 1441
rect 51 1407 53 1441
rect -146 1346 -112 1354
rect -146 1320 -112 1346
rect -146 1278 -112 1282
rect -146 1248 -112 1278
rect -146 1176 -112 1210
rect -146 1108 -112 1138
rect -146 1104 -112 1108
rect -146 1040 -112 1066
rect -146 1032 -112 1040
rect -146 972 -112 994
rect -146 960 -112 972
rect -146 904 -112 922
rect -146 888 -112 904
rect -146 836 -112 850
rect -146 816 -112 836
rect -146 768 -112 778
rect -146 744 -112 768
rect -146 700 -112 706
rect -146 672 -112 700
rect -146 632 -112 634
rect -146 600 -112 632
rect -146 530 -112 562
rect -146 528 -112 530
rect -146 462 -112 490
rect -146 456 -112 462
rect -146 394 -112 418
rect -146 384 -112 394
rect -146 326 -112 346
rect -146 312 -112 326
rect -146 258 -112 274
rect -146 240 -112 258
rect -146 190 -112 202
rect -146 168 -112 190
rect -146 122 -112 130
rect -146 96 -112 122
rect -146 54 -112 58
rect -146 24 -112 54
rect -146 -48 -112 -14
rect -146 -116 -112 -86
rect -146 -120 -112 -116
rect -146 -184 -112 -158
rect -146 -192 -112 -184
rect -146 -252 -112 -230
rect -146 -264 -112 -252
rect -146 -320 -112 -302
rect -146 -336 -112 -320
rect -146 -388 -112 -374
rect -146 -408 -112 -388
rect -146 -456 -112 -446
rect -146 -480 -112 -456
rect -146 -524 -112 -518
rect -146 -552 -112 -524
rect -146 -592 -112 -590
rect -146 -624 -112 -592
rect -146 -694 -112 -662
rect -146 -696 -112 -694
rect -146 -762 -112 -734
rect -146 -768 -112 -762
rect -146 -830 -112 -806
rect -146 -840 -112 -830
rect -146 -898 -112 -878
rect -146 -912 -112 -898
rect -146 -966 -112 -950
rect -146 -984 -112 -966
rect -146 -1034 -112 -1022
rect -146 -1056 -112 -1034
rect -146 -1102 -112 -1094
rect -146 -1128 -112 -1102
rect -146 -1170 -112 -1166
rect -146 -1200 -112 -1170
rect -146 -1272 -112 -1238
rect -146 -1340 -112 -1310
rect -146 -1344 -112 -1340
rect -146 -1408 -112 -1382
rect -146 -1416 -112 -1408
rect 112 1346 146 1354
rect 112 1320 146 1346
rect 112 1278 146 1282
rect 112 1248 146 1278
rect 112 1176 146 1210
rect 112 1108 146 1138
rect 112 1104 146 1108
rect 112 1040 146 1066
rect 112 1032 146 1040
rect 112 972 146 994
rect 112 960 146 972
rect 112 904 146 922
rect 112 888 146 904
rect 112 836 146 850
rect 112 816 146 836
rect 112 768 146 778
rect 112 744 146 768
rect 112 700 146 706
rect 112 672 146 700
rect 112 632 146 634
rect 112 600 146 632
rect 112 530 146 562
rect 112 528 146 530
rect 112 462 146 490
rect 112 456 146 462
rect 112 394 146 418
rect 112 384 146 394
rect 112 326 146 346
rect 112 312 146 326
rect 112 258 146 274
rect 112 240 146 258
rect 112 190 146 202
rect 112 168 146 190
rect 112 122 146 130
rect 112 96 146 122
rect 112 54 146 58
rect 112 24 146 54
rect 112 -48 146 -14
rect 112 -116 146 -86
rect 112 -120 146 -116
rect 112 -184 146 -158
rect 112 -192 146 -184
rect 112 -252 146 -230
rect 112 -264 146 -252
rect 112 -320 146 -302
rect 112 -336 146 -320
rect 112 -388 146 -374
rect 112 -408 146 -388
rect 112 -456 146 -446
rect 112 -480 146 -456
rect 112 -524 146 -518
rect 112 -552 146 -524
rect 112 -592 146 -590
rect 112 -624 146 -592
rect 112 -694 146 -662
rect 112 -696 146 -694
rect 112 -762 146 -734
rect 112 -768 146 -762
rect 112 -830 146 -806
rect 112 -840 146 -830
rect 112 -898 146 -878
rect 112 -912 146 -898
rect 112 -966 146 -950
rect 112 -984 146 -966
rect 112 -1034 146 -1022
rect 112 -1056 146 -1034
rect 112 -1102 146 -1094
rect 112 -1128 146 -1102
rect 112 -1170 146 -1166
rect 112 -1200 146 -1170
rect 112 -1272 146 -1238
rect 112 -1340 146 -1310
rect 112 -1344 146 -1340
rect 112 -1408 146 -1382
rect 112 -1416 146 -1408
<< metal1 >>
rect -96 1441 96 1447
rect -96 1407 -53 1441
rect -19 1407 19 1441
rect 53 1407 96 1441
rect -96 1401 96 1407
rect -152 1354 -106 1369
rect -152 1320 -146 1354
rect -112 1320 -106 1354
rect -152 1282 -106 1320
rect -152 1248 -146 1282
rect -112 1248 -106 1282
rect -152 1210 -106 1248
rect -152 1176 -146 1210
rect -112 1176 -106 1210
rect -152 1138 -106 1176
rect -152 1104 -146 1138
rect -112 1104 -106 1138
rect -152 1066 -106 1104
rect -152 1032 -146 1066
rect -112 1032 -106 1066
rect -152 994 -106 1032
rect -152 960 -146 994
rect -112 960 -106 994
rect -152 922 -106 960
rect -152 888 -146 922
rect -112 888 -106 922
rect -152 850 -106 888
rect -152 816 -146 850
rect -112 816 -106 850
rect -152 778 -106 816
rect -152 744 -146 778
rect -112 744 -106 778
rect -152 706 -106 744
rect -152 672 -146 706
rect -112 672 -106 706
rect -152 634 -106 672
rect -152 600 -146 634
rect -112 600 -106 634
rect -152 562 -106 600
rect -152 528 -146 562
rect -112 528 -106 562
rect -152 490 -106 528
rect -152 456 -146 490
rect -112 456 -106 490
rect -152 418 -106 456
rect -152 384 -146 418
rect -112 384 -106 418
rect -152 346 -106 384
rect -152 312 -146 346
rect -112 312 -106 346
rect -152 274 -106 312
rect -152 240 -146 274
rect -112 240 -106 274
rect -152 202 -106 240
rect -152 168 -146 202
rect -112 168 -106 202
rect -152 130 -106 168
rect -152 96 -146 130
rect -112 96 -106 130
rect -152 58 -106 96
rect -152 24 -146 58
rect -112 24 -106 58
rect -152 -14 -106 24
rect -152 -48 -146 -14
rect -112 -48 -106 -14
rect -152 -86 -106 -48
rect -152 -120 -146 -86
rect -112 -120 -106 -86
rect -152 -158 -106 -120
rect -152 -192 -146 -158
rect -112 -192 -106 -158
rect -152 -230 -106 -192
rect -152 -264 -146 -230
rect -112 -264 -106 -230
rect -152 -302 -106 -264
rect -152 -336 -146 -302
rect -112 -336 -106 -302
rect -152 -374 -106 -336
rect -152 -408 -146 -374
rect -112 -408 -106 -374
rect -152 -446 -106 -408
rect -152 -480 -146 -446
rect -112 -480 -106 -446
rect -152 -518 -106 -480
rect -152 -552 -146 -518
rect -112 -552 -106 -518
rect -152 -590 -106 -552
rect -152 -624 -146 -590
rect -112 -624 -106 -590
rect -152 -662 -106 -624
rect -152 -696 -146 -662
rect -112 -696 -106 -662
rect -152 -734 -106 -696
rect -152 -768 -146 -734
rect -112 -768 -106 -734
rect -152 -806 -106 -768
rect -152 -840 -146 -806
rect -112 -840 -106 -806
rect -152 -878 -106 -840
rect -152 -912 -146 -878
rect -112 -912 -106 -878
rect -152 -950 -106 -912
rect -152 -984 -146 -950
rect -112 -984 -106 -950
rect -152 -1022 -106 -984
rect -152 -1056 -146 -1022
rect -112 -1056 -106 -1022
rect -152 -1094 -106 -1056
rect -152 -1128 -146 -1094
rect -112 -1128 -106 -1094
rect -152 -1166 -106 -1128
rect -152 -1200 -146 -1166
rect -112 -1200 -106 -1166
rect -152 -1238 -106 -1200
rect -152 -1272 -146 -1238
rect -112 -1272 -106 -1238
rect -152 -1310 -106 -1272
rect -152 -1344 -146 -1310
rect -112 -1344 -106 -1310
rect -152 -1382 -106 -1344
rect -152 -1416 -146 -1382
rect -112 -1416 -106 -1382
rect -152 -1431 -106 -1416
rect 106 1354 152 1369
rect 106 1320 112 1354
rect 146 1320 152 1354
rect 106 1282 152 1320
rect 106 1248 112 1282
rect 146 1248 152 1282
rect 106 1210 152 1248
rect 106 1176 112 1210
rect 146 1176 152 1210
rect 106 1138 152 1176
rect 106 1104 112 1138
rect 146 1104 152 1138
rect 106 1066 152 1104
rect 106 1032 112 1066
rect 146 1032 152 1066
rect 106 994 152 1032
rect 106 960 112 994
rect 146 960 152 994
rect 106 922 152 960
rect 106 888 112 922
rect 146 888 152 922
rect 106 850 152 888
rect 106 816 112 850
rect 146 816 152 850
rect 106 778 152 816
rect 106 744 112 778
rect 146 744 152 778
rect 106 706 152 744
rect 106 672 112 706
rect 146 672 152 706
rect 106 634 152 672
rect 106 600 112 634
rect 146 600 152 634
rect 106 562 152 600
rect 106 528 112 562
rect 146 528 152 562
rect 106 490 152 528
rect 106 456 112 490
rect 146 456 152 490
rect 106 418 152 456
rect 106 384 112 418
rect 146 384 152 418
rect 106 346 152 384
rect 106 312 112 346
rect 146 312 152 346
rect 106 274 152 312
rect 106 240 112 274
rect 146 240 152 274
rect 106 202 152 240
rect 106 168 112 202
rect 146 168 152 202
rect 106 130 152 168
rect 106 96 112 130
rect 146 96 152 130
rect 106 58 152 96
rect 106 24 112 58
rect 146 24 152 58
rect 106 -14 152 24
rect 106 -48 112 -14
rect 146 -48 152 -14
rect 106 -86 152 -48
rect 106 -120 112 -86
rect 146 -120 152 -86
rect 106 -158 152 -120
rect 106 -192 112 -158
rect 146 -192 152 -158
rect 106 -230 152 -192
rect 106 -264 112 -230
rect 146 -264 152 -230
rect 106 -302 152 -264
rect 106 -336 112 -302
rect 146 -336 152 -302
rect 106 -374 152 -336
rect 106 -408 112 -374
rect 146 -408 152 -374
rect 106 -446 152 -408
rect 106 -480 112 -446
rect 146 -480 152 -446
rect 106 -518 152 -480
rect 106 -552 112 -518
rect 146 -552 152 -518
rect 106 -590 152 -552
rect 106 -624 112 -590
rect 146 -624 152 -590
rect 106 -662 152 -624
rect 106 -696 112 -662
rect 146 -696 152 -662
rect 106 -734 152 -696
rect 106 -768 112 -734
rect 146 -768 152 -734
rect 106 -806 152 -768
rect 106 -840 112 -806
rect 146 -840 152 -806
rect 106 -878 152 -840
rect 106 -912 112 -878
rect 146 -912 152 -878
rect 106 -950 152 -912
rect 106 -984 112 -950
rect 146 -984 152 -950
rect 106 -1022 152 -984
rect 106 -1056 112 -1022
rect 146 -1056 152 -1022
rect 106 -1094 152 -1056
rect 106 -1128 112 -1094
rect 146 -1128 152 -1094
rect 106 -1166 152 -1128
rect 106 -1200 112 -1166
rect 146 -1200 152 -1166
rect 106 -1238 152 -1200
rect 106 -1272 112 -1238
rect 146 -1272 152 -1238
rect 106 -1310 152 -1272
rect 106 -1344 112 -1310
rect 146 -1344 152 -1310
rect 106 -1382 152 -1344
rect 106 -1416 112 -1382
rect 146 -1416 152 -1382
rect 106 -1431 152 -1416
<< end >>
