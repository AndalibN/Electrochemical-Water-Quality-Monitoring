magic
tech sky130A
magscale 1 2
timestamp 1666707788
<< nwell >>
rect -396 -2219 396 2219
<< pmos >>
rect -200 -2000 200 2000
<< pdiff >>
rect -258 1988 -200 2000
rect -258 -1988 -246 1988
rect -212 -1988 -200 1988
rect -258 -2000 -200 -1988
rect 200 1988 258 2000
rect 200 -1988 212 1988
rect 246 -1988 258 1988
rect 200 -2000 258 -1988
<< pdiffc >>
rect -246 -1988 -212 1988
rect 212 -1988 246 1988
<< nsubdiff >>
rect -360 2149 -264 2183
rect 264 2149 360 2183
rect -360 2087 -326 2149
rect 326 2087 360 2149
rect -360 -2149 -326 -2087
rect 326 -2149 360 -2087
rect -360 -2183 -264 -2149
rect 264 -2183 360 -2149
<< nsubdiffcont >>
rect -264 2149 264 2183
rect -360 -2087 -326 2087
rect 326 -2087 360 2087
rect -264 -2183 264 -2149
<< poly >>
rect -200 2081 200 2097
rect -200 2047 -184 2081
rect 184 2047 200 2081
rect -200 2000 200 2047
rect -200 -2047 200 -2000
rect -200 -2081 -184 -2047
rect 184 -2081 200 -2047
rect -200 -2097 200 -2081
<< polycont >>
rect -184 2047 184 2081
rect -184 -2081 184 -2047
<< locali >>
rect -360 2149 -264 2183
rect 264 2149 360 2183
rect -360 2087 -326 2149
rect 326 2087 360 2149
rect -200 2047 -184 2081
rect 184 2047 200 2081
rect -246 1988 -212 2004
rect -246 -2004 -212 -1988
rect 212 1988 246 2004
rect 212 -2004 246 -1988
rect -200 -2081 -184 -2047
rect 184 -2081 200 -2047
rect -360 -2149 -326 -2087
rect 326 -2149 360 -2087
rect -360 -2183 -264 -2149
rect 264 -2183 360 -2149
<< viali >>
rect -184 2047 184 2081
rect -246 -1988 -212 1988
rect 212 -1988 246 1988
rect -184 -2081 184 -2047
<< metal1 >>
rect -196 2081 196 2087
rect -196 2047 -184 2081
rect 184 2047 196 2081
rect -196 2041 196 2047
rect -252 1988 -206 2000
rect -252 -1988 -246 1988
rect -212 -1988 -206 1988
rect -252 -2000 -206 -1988
rect 206 1988 252 2000
rect 206 -1988 212 1988
rect 246 -1988 252 1988
rect 206 -2000 252 -1988
rect -196 -2047 196 -2041
rect -196 -2081 -184 -2047
rect 184 -2081 196 -2047
rect -196 -2087 196 -2081
<< properties >>
string FIXED_BBOX -343 -2166 343 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
