magic
tech sky130A
magscale 1 2
timestamp 1668099713
<< metal1 >>
rect 3470 -9588 4018 -9574
rect 3470 -9662 4442 -9588
rect 3470 -10144 4018 -9662
rect 3470 -10512 3546 -10144
rect 3966 -10512 4018 -10144
rect 3470 -10558 4018 -10512
<< via1 >>
rect 3546 -10512 3966 -10144
<< metal2 >>
rect 3354 -10144 4130 -10056
rect 3354 -10512 3546 -10144
rect 3966 -10512 4130 -10144
rect 3354 -11474 4130 -10512
rect 3412 -11928 4092 -11474
rect 3412 -12370 3462 -11928
rect 4024 -12370 4092 -11928
rect 3412 -12412 4092 -12370
<< via2 >>
rect 3462 -12370 4024 -11928
<< metal3 >>
rect 3416 -11928 4084 -11876
rect 3416 -12370 3462 -11928
rect 4024 -12370 4084 -11928
rect 3416 -12804 4084 -12370
rect 2468 -12946 4084 -12804
rect 2468 -13494 2528 -12946
rect 2970 -13494 4084 -12946
rect 2468 -13602 4084 -13494
<< via3 >>
rect 2528 -13494 2970 -12946
<< metal4 >>
rect 63148 51650 69836 55118
rect -3652 -12006 -1110 -8826
rect 2030 -12888 3016 -12886
rect 1292 -12946 3016 -12888
rect 1292 -12974 2528 -12946
rect 1770 -13494 2528 -12974
rect 2970 -13494 3016 -12946
rect 1770 -13538 3016 -13494
rect 1292 -13604 3016 -13538
rect 1292 -13606 2278 -13604
<< via4 >>
rect 1292 -13538 1770 -12974
<< metal5 >>
rect -3566 -12974 1854 -12834
rect -3566 -13538 1292 -12974
rect 1770 -13538 1854 -12974
rect -3566 -13622 1854 -13538
use ind700p_1  ind700p_1_0
timestamp 1667951165
transform -1 0 -20110 0 -1 -11320
box -17300 -8000 14700 8000
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_0
timestamp 1667951165
transform 0 1 4684 1 0 -9625
box -37 -502 37 502
<< labels >>
rlabel metal4 -2554 -11370 -1110 -9578 1 A
port 1 n
<< end >>
