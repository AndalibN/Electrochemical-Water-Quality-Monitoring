magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< metal3 >>
rect -775 697 774 725
rect -775 -697 690 697
rect 754 -697 774 697
rect -775 -725 774 -697
<< via3 >>
rect 690 -697 754 697
<< mimcap >>
rect -675 585 575 625
rect -675 -585 -635 585
rect 535 -585 575 585
rect -675 -625 575 -585
<< mimcapcontact >>
rect -635 -585 535 585
<< metal4 >>
rect 674 697 770 713
rect -636 585 536 586
rect -636 -585 -635 585
rect 535 -585 536 585
rect -636 -586 536 -585
rect 674 -697 690 697
rect 754 -697 770 697
rect 674 -713 770 -697
<< properties >>
string FIXED_BBOX -775 -725 675 725
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6.25 l 6.25 val 82.875 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
