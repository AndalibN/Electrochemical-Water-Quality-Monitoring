magic
tech sky130A
timestamp 1668127436
<< metal4 >>
rect -5047 -18154 -3263 -16349
rect -9283 -32265 -7548 -32248
rect -9283 -33725 -9270 -32265
rect -7589 -33725 -7548 -32265
rect -9283 -35818 -7548 -33725
rect -9029 -36011 -7627 -35818
rect -5849 -39011 -2022 -38868
rect -5849 -39532 -5759 -39011
rect -4789 -39532 -2022 -39011
rect -5849 -39712 -2022 -39532
<< via4 >>
rect -9270 -33725 -7589 -32265
rect -5759 -39532 -4789 -39011
<< metal5 >>
rect -14641 16963 -4527 18800
rect -6559 13401 -4722 13449
rect -11997 -7891 -10160 13361
rect -6559 11594 -2464 13401
rect -11997 -10722 -10236 -7891
rect -11997 -11577 -10196 -10722
rect -6559 -10965 -4722 11594
rect -10605 -11620 -10196 -11577
rect -6560 -11051 -4722 -10965
rect -6560 -12756 -5245 -11051
rect -9338 -32265 -7501 -15153
rect -9338 -33725 -9270 -32265
rect -7589 -33725 -7501 -32265
rect -9338 -34086 -7501 -33725
rect -8670 -36812 -7689 -36577
rect -8670 -37144 -7681 -36812
rect -8224 -38920 -7681 -37144
rect -8224 -39011 -4741 -38920
rect -8224 -39532 -5759 -39011
rect -4789 -39532 -4741 -39011
rect -8224 -39631 -4741 -39532
rect -8119 -39638 -4741 -39631
rect -1506 -39887 -993 -39461
rect -1572 -41747 -935 -41010
<< mrdlcontact >>
rect -1572 -41010 -935 -39887
use ind2p69  ind2p69_0
timestamp 1667951165
transform -1 0 -37941 0 -1 5162
box -26600 -22500 2700 2500
use ind2p69  ind2p69_1
timestamp 1667951165
transform 1 0 20835 0 1 25200
box -26600 -22500 2700 2500
use ind2p69  ind2p69_2
timestamp 1667951165
transform 1 0 20923 0 1 -4557
box -26600 -22500 2700 2500
use ind2p69  ind2p69_3
timestamp 1667951165
transform -1 0 -35289 0 -1 -23359
box -26600 -22500 2700 2500
use ind700p_1  ind700p_1_0
timestamp 1667951165
transform 0 1 -2255 1 0 -31008
box -8650 -4000 7350 4000
use ind700p_1  ind700p_1_1
timestamp 1667951165
transform -1 0 -17253 0 -1 -35839
box -8650 -4000 7350 4000
<< labels >>
rlabel metal4 -5042 -18137 -4621 -16362 1 E
port 1 n
rlabel metal5 -1572 -41747 -941 -41388 1 F
port 2 n
<< properties >>
string LEFview true
string device primitive
<< end >>
