magic
tech sky130A
magscale 1 2
timestamp 1666402782
<< metal3 >>
rect -1850 572 1849 600
rect -1850 -572 1765 572
rect 1829 -572 1849 572
rect -1850 -600 1849 -572
<< via3 >>
rect 1765 -572 1829 572
<< mimcap >>
rect -1750 460 1650 500
rect -1750 -460 -1710 460
rect 1610 -460 1650 460
rect -1750 -500 1650 -460
<< mimcapcontact >>
rect -1710 -460 1610 460
<< metal4 >>
rect 1749 572 1845 588
rect -1711 460 1611 461
rect -1711 -460 -1710 460
rect 1610 -460 1611 460
rect -1711 -461 1611 -460
rect 1749 -572 1765 572
rect 1829 -572 1845 572
rect 1749 -588 1845 -572
<< properties >>
string FIXED_BBOX -1850 -600 1750 600
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17.0 l 5.0 val 178.36 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
