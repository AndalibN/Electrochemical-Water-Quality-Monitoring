magic
tech sky130A
magscale 1 2
timestamp 1667266911
<< nwell >>
rect -1123 -300 1123 300
<< pmos >>
rect -1029 -200 -29 200
rect 29 -200 1029 200
<< pdiff >>
rect -1087 188 -1029 200
rect -1087 -188 -1075 188
rect -1041 -188 -1029 188
rect -1087 -200 -1029 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 1029 188 1087 200
rect 1029 -188 1041 188
rect 1075 -188 1087 188
rect 1029 -200 1087 -188
<< pdiffc >>
rect -1075 -188 -1041 188
rect -17 -188 17 188
rect 1041 -188 1075 188
<< poly >>
rect -1029 281 -29 297
rect -1029 247 -1013 281
rect -45 247 -29 281
rect -1029 200 -29 247
rect 29 281 1029 297
rect 29 247 45 281
rect 1013 247 1029 281
rect 29 200 1029 247
rect -1029 -247 -29 -200
rect -1029 -281 -1013 -247
rect -45 -281 -29 -247
rect -1029 -297 -29 -281
rect 29 -247 1029 -200
rect 29 -281 45 -247
rect 1013 -281 1029 -247
rect 29 -297 1029 -281
<< polycont >>
rect -1013 247 -45 281
rect 45 247 1013 281
rect -1013 -281 -45 -247
rect 45 -281 1013 -247
<< locali >>
rect -1029 247 -1013 281
rect -45 247 -29 281
rect 29 247 45 281
rect 1013 247 1029 281
rect -1075 188 -1041 204
rect -1075 -204 -1041 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 1041 188 1075 204
rect 1041 -204 1075 -188
rect -1029 -281 -1013 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 1013 -281 1029 -247
<< viali >>
rect -1013 247 -45 281
rect 45 247 1013 281
rect -1075 -188 -1041 188
rect -17 -188 17 188
rect 1041 -188 1075 188
rect -1013 -281 -45 -247
rect 45 -281 1013 -247
<< metal1 >>
rect -1025 281 -33 287
rect -1025 247 -1013 281
rect -45 247 -33 281
rect -1025 241 -33 247
rect 33 281 1025 287
rect 33 247 45 281
rect 1013 247 1025 281
rect 33 241 1025 247
rect -1081 188 -1035 200
rect -1081 -188 -1075 188
rect -1041 -188 -1035 188
rect -1081 -200 -1035 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 1035 188 1081 200
rect 1035 -188 1041 188
rect 1075 -188 1081 188
rect 1035 -200 1081 -188
rect -1025 -247 -33 -241
rect -1025 -281 -1013 -247
rect -45 -281 -33 -247
rect -1025 -287 -33 -281
rect 33 -247 1025 -241
rect 33 -281 45 -247
rect 1013 -281 1025 -247
rect 33 -287 1025 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 5.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
