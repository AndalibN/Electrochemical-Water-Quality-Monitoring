magic
tech sky130A
timestamp 1667443905
<< nmos >>
rect -100 -1000 100 1000
<< ndiff >>
rect -129 994 -100 1000
rect -129 -994 -123 994
rect -106 -994 -100 994
rect -129 -1000 -100 -994
rect 100 994 129 1000
rect 100 -994 106 994
rect 123 -994 129 994
rect 100 -1000 129 -994
<< ndiffc >>
rect -123 -994 -106 994
rect 106 -994 123 994
<< poly >>
rect -100 1036 100 1044
rect -100 1019 -92 1036
rect 92 1019 100 1036
rect -100 1000 100 1019
rect -100 -1019 100 -1000
rect -100 -1036 -92 -1019
rect 92 -1036 100 -1019
rect -100 -1044 100 -1036
<< polycont >>
rect -92 1019 92 1036
rect -92 -1036 92 -1019
<< locali >>
rect -100 1019 -92 1036
rect 92 1019 100 1036
rect -123 994 -106 1002
rect -123 -1002 -106 -994
rect 106 994 123 1002
rect 106 -1002 123 -994
rect -100 -1036 -92 -1019
rect 92 -1036 100 -1019
<< viali >>
rect -92 1019 92 1036
rect -123 -994 -106 994
rect 106 -994 123 994
rect -92 -1036 92 -1019
<< metal1 >>
rect -98 1036 98 1039
rect -98 1019 -92 1036
rect 92 1019 98 1036
rect -98 1016 98 1019
rect -126 994 -103 1000
rect -126 -994 -123 994
rect -106 -994 -103 994
rect -126 -1000 -103 -994
rect 103 994 126 1000
rect 103 -994 106 994
rect 123 -994 126 994
rect 103 -1000 126 -994
rect -98 -1019 98 -1016
rect -98 -1036 -92 -1019
rect 92 -1036 98 -1019
rect -98 -1039 98 -1036
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
