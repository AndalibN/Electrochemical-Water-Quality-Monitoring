magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -3568 3332 -1849 3390
rect -3568 3268 -1933 3332
rect -1869 3268 -1849 3332
rect -3568 3252 -1849 3268
rect -3568 3188 -1933 3252
rect -1869 3188 -1849 3252
rect -3568 3172 -1849 3188
rect -3568 3108 -1933 3172
rect -1869 3108 -1849 3172
rect -3568 3092 -1849 3108
rect -3568 3028 -1933 3092
rect -1869 3028 -1849 3092
rect -3568 3012 -1849 3028
rect -3568 2948 -1933 3012
rect -1869 2948 -1849 3012
rect -3568 2932 -1849 2948
rect -3568 2868 -1933 2932
rect -1869 2868 -1849 2932
rect -3568 2852 -1849 2868
rect -3568 2788 -1933 2852
rect -1869 2788 -1849 2852
rect -3568 2772 -1849 2788
rect -3568 2708 -1933 2772
rect -1869 2708 -1849 2772
rect -3568 2692 -1849 2708
rect -3568 2628 -1933 2692
rect -1869 2628 -1849 2692
rect -3568 2612 -1849 2628
rect -3568 2548 -1933 2612
rect -1869 2548 -1849 2612
rect -3568 2532 -1849 2548
rect -3568 2468 -1933 2532
rect -1869 2468 -1849 2532
rect -3568 2452 -1849 2468
rect -3568 2388 -1933 2452
rect -1869 2388 -1849 2452
rect -3568 2372 -1849 2388
rect -3568 2308 -1933 2372
rect -1869 2308 -1849 2372
rect -3568 2292 -1849 2308
rect -3568 2228 -1933 2292
rect -1869 2228 -1849 2292
rect -3568 2212 -1849 2228
rect -3568 2148 -1933 2212
rect -1869 2148 -1849 2212
rect -3568 2132 -1849 2148
rect -3568 2068 -1933 2132
rect -1869 2068 -1849 2132
rect -3568 2052 -1849 2068
rect -3568 1988 -1933 2052
rect -1869 1988 -1849 2052
rect -3568 1972 -1849 1988
rect -3568 1908 -1933 1972
rect -1869 1908 -1849 1972
rect -3568 1892 -1849 1908
rect -3568 1828 -1933 1892
rect -1869 1828 -1849 1892
rect -3568 1770 -1849 1828
rect -1729 3332 -10 3390
rect -1729 3268 -94 3332
rect -30 3268 -10 3332
rect -1729 3252 -10 3268
rect -1729 3188 -94 3252
rect -30 3188 -10 3252
rect -1729 3172 -10 3188
rect -1729 3108 -94 3172
rect -30 3108 -10 3172
rect -1729 3092 -10 3108
rect -1729 3028 -94 3092
rect -30 3028 -10 3092
rect -1729 3012 -10 3028
rect -1729 2948 -94 3012
rect -30 2948 -10 3012
rect -1729 2932 -10 2948
rect -1729 2868 -94 2932
rect -30 2868 -10 2932
rect -1729 2852 -10 2868
rect -1729 2788 -94 2852
rect -30 2788 -10 2852
rect -1729 2772 -10 2788
rect -1729 2708 -94 2772
rect -30 2708 -10 2772
rect -1729 2692 -10 2708
rect -1729 2628 -94 2692
rect -30 2628 -10 2692
rect -1729 2612 -10 2628
rect -1729 2548 -94 2612
rect -30 2548 -10 2612
rect -1729 2532 -10 2548
rect -1729 2468 -94 2532
rect -30 2468 -10 2532
rect -1729 2452 -10 2468
rect -1729 2388 -94 2452
rect -30 2388 -10 2452
rect -1729 2372 -10 2388
rect -1729 2308 -94 2372
rect -30 2308 -10 2372
rect -1729 2292 -10 2308
rect -1729 2228 -94 2292
rect -30 2228 -10 2292
rect -1729 2212 -10 2228
rect -1729 2148 -94 2212
rect -30 2148 -10 2212
rect -1729 2132 -10 2148
rect -1729 2068 -94 2132
rect -30 2068 -10 2132
rect -1729 2052 -10 2068
rect -1729 1988 -94 2052
rect -30 1988 -10 2052
rect -1729 1972 -10 1988
rect -1729 1908 -94 1972
rect -30 1908 -10 1972
rect -1729 1892 -10 1908
rect -1729 1828 -94 1892
rect -30 1828 -10 1892
rect -1729 1770 -10 1828
rect 110 3332 1829 3390
rect 110 3268 1745 3332
rect 1809 3268 1829 3332
rect 110 3252 1829 3268
rect 110 3188 1745 3252
rect 1809 3188 1829 3252
rect 110 3172 1829 3188
rect 110 3108 1745 3172
rect 1809 3108 1829 3172
rect 110 3092 1829 3108
rect 110 3028 1745 3092
rect 1809 3028 1829 3092
rect 110 3012 1829 3028
rect 110 2948 1745 3012
rect 1809 2948 1829 3012
rect 110 2932 1829 2948
rect 110 2868 1745 2932
rect 1809 2868 1829 2932
rect 110 2852 1829 2868
rect 110 2788 1745 2852
rect 1809 2788 1829 2852
rect 110 2772 1829 2788
rect 110 2708 1745 2772
rect 1809 2708 1829 2772
rect 110 2692 1829 2708
rect 110 2628 1745 2692
rect 1809 2628 1829 2692
rect 110 2612 1829 2628
rect 110 2548 1745 2612
rect 1809 2548 1829 2612
rect 110 2532 1829 2548
rect 110 2468 1745 2532
rect 1809 2468 1829 2532
rect 110 2452 1829 2468
rect 110 2388 1745 2452
rect 1809 2388 1829 2452
rect 110 2372 1829 2388
rect 110 2308 1745 2372
rect 1809 2308 1829 2372
rect 110 2292 1829 2308
rect 110 2228 1745 2292
rect 1809 2228 1829 2292
rect 110 2212 1829 2228
rect 110 2148 1745 2212
rect 1809 2148 1829 2212
rect 110 2132 1829 2148
rect 110 2068 1745 2132
rect 1809 2068 1829 2132
rect 110 2052 1829 2068
rect 110 1988 1745 2052
rect 1809 1988 1829 2052
rect 110 1972 1829 1988
rect 110 1908 1745 1972
rect 1809 1908 1829 1972
rect 110 1892 1829 1908
rect 110 1828 1745 1892
rect 1809 1828 1829 1892
rect 110 1770 1829 1828
rect 1949 3332 3668 3390
rect 1949 3268 3584 3332
rect 3648 3268 3668 3332
rect 1949 3252 3668 3268
rect 1949 3188 3584 3252
rect 3648 3188 3668 3252
rect 1949 3172 3668 3188
rect 1949 3108 3584 3172
rect 3648 3108 3668 3172
rect 1949 3092 3668 3108
rect 1949 3028 3584 3092
rect 3648 3028 3668 3092
rect 1949 3012 3668 3028
rect 1949 2948 3584 3012
rect 3648 2948 3668 3012
rect 1949 2932 3668 2948
rect 1949 2868 3584 2932
rect 3648 2868 3668 2932
rect 1949 2852 3668 2868
rect 1949 2788 3584 2852
rect 3648 2788 3668 2852
rect 1949 2772 3668 2788
rect 1949 2708 3584 2772
rect 3648 2708 3668 2772
rect 1949 2692 3668 2708
rect 1949 2628 3584 2692
rect 3648 2628 3668 2692
rect 1949 2612 3668 2628
rect 1949 2548 3584 2612
rect 3648 2548 3668 2612
rect 1949 2532 3668 2548
rect 1949 2468 3584 2532
rect 3648 2468 3668 2532
rect 1949 2452 3668 2468
rect 1949 2388 3584 2452
rect 3648 2388 3668 2452
rect 1949 2372 3668 2388
rect 1949 2308 3584 2372
rect 3648 2308 3668 2372
rect 1949 2292 3668 2308
rect 1949 2228 3584 2292
rect 3648 2228 3668 2292
rect 1949 2212 3668 2228
rect 1949 2148 3584 2212
rect 3648 2148 3668 2212
rect 1949 2132 3668 2148
rect 1949 2068 3584 2132
rect 3648 2068 3668 2132
rect 1949 2052 3668 2068
rect 1949 1988 3584 2052
rect 3648 1988 3668 2052
rect 1949 1972 3668 1988
rect 1949 1908 3584 1972
rect 3648 1908 3668 1972
rect 1949 1892 3668 1908
rect 1949 1828 3584 1892
rect 3648 1828 3668 1892
rect 1949 1770 3668 1828
rect -3568 1612 -1849 1670
rect -3568 1548 -1933 1612
rect -1869 1548 -1849 1612
rect -3568 1532 -1849 1548
rect -3568 1468 -1933 1532
rect -1869 1468 -1849 1532
rect -3568 1452 -1849 1468
rect -3568 1388 -1933 1452
rect -1869 1388 -1849 1452
rect -3568 1372 -1849 1388
rect -3568 1308 -1933 1372
rect -1869 1308 -1849 1372
rect -3568 1292 -1849 1308
rect -3568 1228 -1933 1292
rect -1869 1228 -1849 1292
rect -3568 1212 -1849 1228
rect -3568 1148 -1933 1212
rect -1869 1148 -1849 1212
rect -3568 1132 -1849 1148
rect -3568 1068 -1933 1132
rect -1869 1068 -1849 1132
rect -3568 1052 -1849 1068
rect -3568 988 -1933 1052
rect -1869 988 -1849 1052
rect -3568 972 -1849 988
rect -3568 908 -1933 972
rect -1869 908 -1849 972
rect -3568 892 -1849 908
rect -3568 828 -1933 892
rect -1869 828 -1849 892
rect -3568 812 -1849 828
rect -3568 748 -1933 812
rect -1869 748 -1849 812
rect -3568 732 -1849 748
rect -3568 668 -1933 732
rect -1869 668 -1849 732
rect -3568 652 -1849 668
rect -3568 588 -1933 652
rect -1869 588 -1849 652
rect -3568 572 -1849 588
rect -3568 508 -1933 572
rect -1869 508 -1849 572
rect -3568 492 -1849 508
rect -3568 428 -1933 492
rect -1869 428 -1849 492
rect -3568 412 -1849 428
rect -3568 348 -1933 412
rect -1869 348 -1849 412
rect -3568 332 -1849 348
rect -3568 268 -1933 332
rect -1869 268 -1849 332
rect -3568 252 -1849 268
rect -3568 188 -1933 252
rect -1869 188 -1849 252
rect -3568 172 -1849 188
rect -3568 108 -1933 172
rect -1869 108 -1849 172
rect -3568 50 -1849 108
rect -1729 1612 -10 1670
rect -1729 1548 -94 1612
rect -30 1548 -10 1612
rect -1729 1532 -10 1548
rect -1729 1468 -94 1532
rect -30 1468 -10 1532
rect -1729 1452 -10 1468
rect -1729 1388 -94 1452
rect -30 1388 -10 1452
rect -1729 1372 -10 1388
rect -1729 1308 -94 1372
rect -30 1308 -10 1372
rect -1729 1292 -10 1308
rect -1729 1228 -94 1292
rect -30 1228 -10 1292
rect -1729 1212 -10 1228
rect -1729 1148 -94 1212
rect -30 1148 -10 1212
rect -1729 1132 -10 1148
rect -1729 1068 -94 1132
rect -30 1068 -10 1132
rect -1729 1052 -10 1068
rect -1729 988 -94 1052
rect -30 988 -10 1052
rect -1729 972 -10 988
rect -1729 908 -94 972
rect -30 908 -10 972
rect -1729 892 -10 908
rect -1729 828 -94 892
rect -30 828 -10 892
rect -1729 812 -10 828
rect -1729 748 -94 812
rect -30 748 -10 812
rect -1729 732 -10 748
rect -1729 668 -94 732
rect -30 668 -10 732
rect -1729 652 -10 668
rect -1729 588 -94 652
rect -30 588 -10 652
rect -1729 572 -10 588
rect -1729 508 -94 572
rect -30 508 -10 572
rect -1729 492 -10 508
rect -1729 428 -94 492
rect -30 428 -10 492
rect -1729 412 -10 428
rect -1729 348 -94 412
rect -30 348 -10 412
rect -1729 332 -10 348
rect -1729 268 -94 332
rect -30 268 -10 332
rect -1729 252 -10 268
rect -1729 188 -94 252
rect -30 188 -10 252
rect -1729 172 -10 188
rect -1729 108 -94 172
rect -30 108 -10 172
rect -1729 50 -10 108
rect 110 1612 1829 1670
rect 110 1548 1745 1612
rect 1809 1548 1829 1612
rect 110 1532 1829 1548
rect 110 1468 1745 1532
rect 1809 1468 1829 1532
rect 110 1452 1829 1468
rect 110 1388 1745 1452
rect 1809 1388 1829 1452
rect 110 1372 1829 1388
rect 110 1308 1745 1372
rect 1809 1308 1829 1372
rect 110 1292 1829 1308
rect 110 1228 1745 1292
rect 1809 1228 1829 1292
rect 110 1212 1829 1228
rect 110 1148 1745 1212
rect 1809 1148 1829 1212
rect 110 1132 1829 1148
rect 110 1068 1745 1132
rect 1809 1068 1829 1132
rect 110 1052 1829 1068
rect 110 988 1745 1052
rect 1809 988 1829 1052
rect 110 972 1829 988
rect 110 908 1745 972
rect 1809 908 1829 972
rect 110 892 1829 908
rect 110 828 1745 892
rect 1809 828 1829 892
rect 110 812 1829 828
rect 110 748 1745 812
rect 1809 748 1829 812
rect 110 732 1829 748
rect 110 668 1745 732
rect 1809 668 1829 732
rect 110 652 1829 668
rect 110 588 1745 652
rect 1809 588 1829 652
rect 110 572 1829 588
rect 110 508 1745 572
rect 1809 508 1829 572
rect 110 492 1829 508
rect 110 428 1745 492
rect 1809 428 1829 492
rect 110 412 1829 428
rect 110 348 1745 412
rect 1809 348 1829 412
rect 110 332 1829 348
rect 110 268 1745 332
rect 1809 268 1829 332
rect 110 252 1829 268
rect 110 188 1745 252
rect 1809 188 1829 252
rect 110 172 1829 188
rect 110 108 1745 172
rect 1809 108 1829 172
rect 110 50 1829 108
rect 1949 1612 3668 1670
rect 1949 1548 3584 1612
rect 3648 1548 3668 1612
rect 1949 1532 3668 1548
rect 1949 1468 3584 1532
rect 3648 1468 3668 1532
rect 1949 1452 3668 1468
rect 1949 1388 3584 1452
rect 3648 1388 3668 1452
rect 1949 1372 3668 1388
rect 1949 1308 3584 1372
rect 3648 1308 3668 1372
rect 1949 1292 3668 1308
rect 1949 1228 3584 1292
rect 3648 1228 3668 1292
rect 1949 1212 3668 1228
rect 1949 1148 3584 1212
rect 3648 1148 3668 1212
rect 1949 1132 3668 1148
rect 1949 1068 3584 1132
rect 3648 1068 3668 1132
rect 1949 1052 3668 1068
rect 1949 988 3584 1052
rect 3648 988 3668 1052
rect 1949 972 3668 988
rect 1949 908 3584 972
rect 3648 908 3668 972
rect 1949 892 3668 908
rect 1949 828 3584 892
rect 3648 828 3668 892
rect 1949 812 3668 828
rect 1949 748 3584 812
rect 3648 748 3668 812
rect 1949 732 3668 748
rect 1949 668 3584 732
rect 3648 668 3668 732
rect 1949 652 3668 668
rect 1949 588 3584 652
rect 3648 588 3668 652
rect 1949 572 3668 588
rect 1949 508 3584 572
rect 3648 508 3668 572
rect 1949 492 3668 508
rect 1949 428 3584 492
rect 3648 428 3668 492
rect 1949 412 3668 428
rect 1949 348 3584 412
rect 3648 348 3668 412
rect 1949 332 3668 348
rect 1949 268 3584 332
rect 3648 268 3668 332
rect 1949 252 3668 268
rect 1949 188 3584 252
rect 3648 188 3668 252
rect 1949 172 3668 188
rect 1949 108 3584 172
rect 3648 108 3668 172
rect 1949 50 3668 108
rect -3568 -108 -1849 -50
rect -3568 -172 -1933 -108
rect -1869 -172 -1849 -108
rect -3568 -188 -1849 -172
rect -3568 -252 -1933 -188
rect -1869 -252 -1849 -188
rect -3568 -268 -1849 -252
rect -3568 -332 -1933 -268
rect -1869 -332 -1849 -268
rect -3568 -348 -1849 -332
rect -3568 -412 -1933 -348
rect -1869 -412 -1849 -348
rect -3568 -428 -1849 -412
rect -3568 -492 -1933 -428
rect -1869 -492 -1849 -428
rect -3568 -508 -1849 -492
rect -3568 -572 -1933 -508
rect -1869 -572 -1849 -508
rect -3568 -588 -1849 -572
rect -3568 -652 -1933 -588
rect -1869 -652 -1849 -588
rect -3568 -668 -1849 -652
rect -3568 -732 -1933 -668
rect -1869 -732 -1849 -668
rect -3568 -748 -1849 -732
rect -3568 -812 -1933 -748
rect -1869 -812 -1849 -748
rect -3568 -828 -1849 -812
rect -3568 -892 -1933 -828
rect -1869 -892 -1849 -828
rect -3568 -908 -1849 -892
rect -3568 -972 -1933 -908
rect -1869 -972 -1849 -908
rect -3568 -988 -1849 -972
rect -3568 -1052 -1933 -988
rect -1869 -1052 -1849 -988
rect -3568 -1068 -1849 -1052
rect -3568 -1132 -1933 -1068
rect -1869 -1132 -1849 -1068
rect -3568 -1148 -1849 -1132
rect -3568 -1212 -1933 -1148
rect -1869 -1212 -1849 -1148
rect -3568 -1228 -1849 -1212
rect -3568 -1292 -1933 -1228
rect -1869 -1292 -1849 -1228
rect -3568 -1308 -1849 -1292
rect -3568 -1372 -1933 -1308
rect -1869 -1372 -1849 -1308
rect -3568 -1388 -1849 -1372
rect -3568 -1452 -1933 -1388
rect -1869 -1452 -1849 -1388
rect -3568 -1468 -1849 -1452
rect -3568 -1532 -1933 -1468
rect -1869 -1532 -1849 -1468
rect -3568 -1548 -1849 -1532
rect -3568 -1612 -1933 -1548
rect -1869 -1612 -1849 -1548
rect -3568 -1670 -1849 -1612
rect -1729 -108 -10 -50
rect -1729 -172 -94 -108
rect -30 -172 -10 -108
rect -1729 -188 -10 -172
rect -1729 -252 -94 -188
rect -30 -252 -10 -188
rect -1729 -268 -10 -252
rect -1729 -332 -94 -268
rect -30 -332 -10 -268
rect -1729 -348 -10 -332
rect -1729 -412 -94 -348
rect -30 -412 -10 -348
rect -1729 -428 -10 -412
rect -1729 -492 -94 -428
rect -30 -492 -10 -428
rect -1729 -508 -10 -492
rect -1729 -572 -94 -508
rect -30 -572 -10 -508
rect -1729 -588 -10 -572
rect -1729 -652 -94 -588
rect -30 -652 -10 -588
rect -1729 -668 -10 -652
rect -1729 -732 -94 -668
rect -30 -732 -10 -668
rect -1729 -748 -10 -732
rect -1729 -812 -94 -748
rect -30 -812 -10 -748
rect -1729 -828 -10 -812
rect -1729 -892 -94 -828
rect -30 -892 -10 -828
rect -1729 -908 -10 -892
rect -1729 -972 -94 -908
rect -30 -972 -10 -908
rect -1729 -988 -10 -972
rect -1729 -1052 -94 -988
rect -30 -1052 -10 -988
rect -1729 -1068 -10 -1052
rect -1729 -1132 -94 -1068
rect -30 -1132 -10 -1068
rect -1729 -1148 -10 -1132
rect -1729 -1212 -94 -1148
rect -30 -1212 -10 -1148
rect -1729 -1228 -10 -1212
rect -1729 -1292 -94 -1228
rect -30 -1292 -10 -1228
rect -1729 -1308 -10 -1292
rect -1729 -1372 -94 -1308
rect -30 -1372 -10 -1308
rect -1729 -1388 -10 -1372
rect -1729 -1452 -94 -1388
rect -30 -1452 -10 -1388
rect -1729 -1468 -10 -1452
rect -1729 -1532 -94 -1468
rect -30 -1532 -10 -1468
rect -1729 -1548 -10 -1532
rect -1729 -1612 -94 -1548
rect -30 -1612 -10 -1548
rect -1729 -1670 -10 -1612
rect 110 -108 1829 -50
rect 110 -172 1745 -108
rect 1809 -172 1829 -108
rect 110 -188 1829 -172
rect 110 -252 1745 -188
rect 1809 -252 1829 -188
rect 110 -268 1829 -252
rect 110 -332 1745 -268
rect 1809 -332 1829 -268
rect 110 -348 1829 -332
rect 110 -412 1745 -348
rect 1809 -412 1829 -348
rect 110 -428 1829 -412
rect 110 -492 1745 -428
rect 1809 -492 1829 -428
rect 110 -508 1829 -492
rect 110 -572 1745 -508
rect 1809 -572 1829 -508
rect 110 -588 1829 -572
rect 110 -652 1745 -588
rect 1809 -652 1829 -588
rect 110 -668 1829 -652
rect 110 -732 1745 -668
rect 1809 -732 1829 -668
rect 110 -748 1829 -732
rect 110 -812 1745 -748
rect 1809 -812 1829 -748
rect 110 -828 1829 -812
rect 110 -892 1745 -828
rect 1809 -892 1829 -828
rect 110 -908 1829 -892
rect 110 -972 1745 -908
rect 1809 -972 1829 -908
rect 110 -988 1829 -972
rect 110 -1052 1745 -988
rect 1809 -1052 1829 -988
rect 110 -1068 1829 -1052
rect 110 -1132 1745 -1068
rect 1809 -1132 1829 -1068
rect 110 -1148 1829 -1132
rect 110 -1212 1745 -1148
rect 1809 -1212 1829 -1148
rect 110 -1228 1829 -1212
rect 110 -1292 1745 -1228
rect 1809 -1292 1829 -1228
rect 110 -1308 1829 -1292
rect 110 -1372 1745 -1308
rect 1809 -1372 1829 -1308
rect 110 -1388 1829 -1372
rect 110 -1452 1745 -1388
rect 1809 -1452 1829 -1388
rect 110 -1468 1829 -1452
rect 110 -1532 1745 -1468
rect 1809 -1532 1829 -1468
rect 110 -1548 1829 -1532
rect 110 -1612 1745 -1548
rect 1809 -1612 1829 -1548
rect 110 -1670 1829 -1612
rect 1949 -108 3668 -50
rect 1949 -172 3584 -108
rect 3648 -172 3668 -108
rect 1949 -188 3668 -172
rect 1949 -252 3584 -188
rect 3648 -252 3668 -188
rect 1949 -268 3668 -252
rect 1949 -332 3584 -268
rect 3648 -332 3668 -268
rect 1949 -348 3668 -332
rect 1949 -412 3584 -348
rect 3648 -412 3668 -348
rect 1949 -428 3668 -412
rect 1949 -492 3584 -428
rect 3648 -492 3668 -428
rect 1949 -508 3668 -492
rect 1949 -572 3584 -508
rect 3648 -572 3668 -508
rect 1949 -588 3668 -572
rect 1949 -652 3584 -588
rect 3648 -652 3668 -588
rect 1949 -668 3668 -652
rect 1949 -732 3584 -668
rect 3648 -732 3668 -668
rect 1949 -748 3668 -732
rect 1949 -812 3584 -748
rect 3648 -812 3668 -748
rect 1949 -828 3668 -812
rect 1949 -892 3584 -828
rect 3648 -892 3668 -828
rect 1949 -908 3668 -892
rect 1949 -972 3584 -908
rect 3648 -972 3668 -908
rect 1949 -988 3668 -972
rect 1949 -1052 3584 -988
rect 3648 -1052 3668 -988
rect 1949 -1068 3668 -1052
rect 1949 -1132 3584 -1068
rect 3648 -1132 3668 -1068
rect 1949 -1148 3668 -1132
rect 1949 -1212 3584 -1148
rect 3648 -1212 3668 -1148
rect 1949 -1228 3668 -1212
rect 1949 -1292 3584 -1228
rect 3648 -1292 3668 -1228
rect 1949 -1308 3668 -1292
rect 1949 -1372 3584 -1308
rect 3648 -1372 3668 -1308
rect 1949 -1388 3668 -1372
rect 1949 -1452 3584 -1388
rect 3648 -1452 3668 -1388
rect 1949 -1468 3668 -1452
rect 1949 -1532 3584 -1468
rect 3648 -1532 3668 -1468
rect 1949 -1548 3668 -1532
rect 1949 -1612 3584 -1548
rect 3648 -1612 3668 -1548
rect 1949 -1670 3668 -1612
rect -3568 -1828 -1849 -1770
rect -3568 -1892 -1933 -1828
rect -1869 -1892 -1849 -1828
rect -3568 -1908 -1849 -1892
rect -3568 -1972 -1933 -1908
rect -1869 -1972 -1849 -1908
rect -3568 -1988 -1849 -1972
rect -3568 -2052 -1933 -1988
rect -1869 -2052 -1849 -1988
rect -3568 -2068 -1849 -2052
rect -3568 -2132 -1933 -2068
rect -1869 -2132 -1849 -2068
rect -3568 -2148 -1849 -2132
rect -3568 -2212 -1933 -2148
rect -1869 -2212 -1849 -2148
rect -3568 -2228 -1849 -2212
rect -3568 -2292 -1933 -2228
rect -1869 -2292 -1849 -2228
rect -3568 -2308 -1849 -2292
rect -3568 -2372 -1933 -2308
rect -1869 -2372 -1849 -2308
rect -3568 -2388 -1849 -2372
rect -3568 -2452 -1933 -2388
rect -1869 -2452 -1849 -2388
rect -3568 -2468 -1849 -2452
rect -3568 -2532 -1933 -2468
rect -1869 -2532 -1849 -2468
rect -3568 -2548 -1849 -2532
rect -3568 -2612 -1933 -2548
rect -1869 -2612 -1849 -2548
rect -3568 -2628 -1849 -2612
rect -3568 -2692 -1933 -2628
rect -1869 -2692 -1849 -2628
rect -3568 -2708 -1849 -2692
rect -3568 -2772 -1933 -2708
rect -1869 -2772 -1849 -2708
rect -3568 -2788 -1849 -2772
rect -3568 -2852 -1933 -2788
rect -1869 -2852 -1849 -2788
rect -3568 -2868 -1849 -2852
rect -3568 -2932 -1933 -2868
rect -1869 -2932 -1849 -2868
rect -3568 -2948 -1849 -2932
rect -3568 -3012 -1933 -2948
rect -1869 -3012 -1849 -2948
rect -3568 -3028 -1849 -3012
rect -3568 -3092 -1933 -3028
rect -1869 -3092 -1849 -3028
rect -3568 -3108 -1849 -3092
rect -3568 -3172 -1933 -3108
rect -1869 -3172 -1849 -3108
rect -3568 -3188 -1849 -3172
rect -3568 -3252 -1933 -3188
rect -1869 -3252 -1849 -3188
rect -3568 -3268 -1849 -3252
rect -3568 -3332 -1933 -3268
rect -1869 -3332 -1849 -3268
rect -3568 -3390 -1849 -3332
rect -1729 -1828 -10 -1770
rect -1729 -1892 -94 -1828
rect -30 -1892 -10 -1828
rect -1729 -1908 -10 -1892
rect -1729 -1972 -94 -1908
rect -30 -1972 -10 -1908
rect -1729 -1988 -10 -1972
rect -1729 -2052 -94 -1988
rect -30 -2052 -10 -1988
rect -1729 -2068 -10 -2052
rect -1729 -2132 -94 -2068
rect -30 -2132 -10 -2068
rect -1729 -2148 -10 -2132
rect -1729 -2212 -94 -2148
rect -30 -2212 -10 -2148
rect -1729 -2228 -10 -2212
rect -1729 -2292 -94 -2228
rect -30 -2292 -10 -2228
rect -1729 -2308 -10 -2292
rect -1729 -2372 -94 -2308
rect -30 -2372 -10 -2308
rect -1729 -2388 -10 -2372
rect -1729 -2452 -94 -2388
rect -30 -2452 -10 -2388
rect -1729 -2468 -10 -2452
rect -1729 -2532 -94 -2468
rect -30 -2532 -10 -2468
rect -1729 -2548 -10 -2532
rect -1729 -2612 -94 -2548
rect -30 -2612 -10 -2548
rect -1729 -2628 -10 -2612
rect -1729 -2692 -94 -2628
rect -30 -2692 -10 -2628
rect -1729 -2708 -10 -2692
rect -1729 -2772 -94 -2708
rect -30 -2772 -10 -2708
rect -1729 -2788 -10 -2772
rect -1729 -2852 -94 -2788
rect -30 -2852 -10 -2788
rect -1729 -2868 -10 -2852
rect -1729 -2932 -94 -2868
rect -30 -2932 -10 -2868
rect -1729 -2948 -10 -2932
rect -1729 -3012 -94 -2948
rect -30 -3012 -10 -2948
rect -1729 -3028 -10 -3012
rect -1729 -3092 -94 -3028
rect -30 -3092 -10 -3028
rect -1729 -3108 -10 -3092
rect -1729 -3172 -94 -3108
rect -30 -3172 -10 -3108
rect -1729 -3188 -10 -3172
rect -1729 -3252 -94 -3188
rect -30 -3252 -10 -3188
rect -1729 -3268 -10 -3252
rect -1729 -3332 -94 -3268
rect -30 -3332 -10 -3268
rect -1729 -3390 -10 -3332
rect 110 -1828 1829 -1770
rect 110 -1892 1745 -1828
rect 1809 -1892 1829 -1828
rect 110 -1908 1829 -1892
rect 110 -1972 1745 -1908
rect 1809 -1972 1829 -1908
rect 110 -1988 1829 -1972
rect 110 -2052 1745 -1988
rect 1809 -2052 1829 -1988
rect 110 -2068 1829 -2052
rect 110 -2132 1745 -2068
rect 1809 -2132 1829 -2068
rect 110 -2148 1829 -2132
rect 110 -2212 1745 -2148
rect 1809 -2212 1829 -2148
rect 110 -2228 1829 -2212
rect 110 -2292 1745 -2228
rect 1809 -2292 1829 -2228
rect 110 -2308 1829 -2292
rect 110 -2372 1745 -2308
rect 1809 -2372 1829 -2308
rect 110 -2388 1829 -2372
rect 110 -2452 1745 -2388
rect 1809 -2452 1829 -2388
rect 110 -2468 1829 -2452
rect 110 -2532 1745 -2468
rect 1809 -2532 1829 -2468
rect 110 -2548 1829 -2532
rect 110 -2612 1745 -2548
rect 1809 -2612 1829 -2548
rect 110 -2628 1829 -2612
rect 110 -2692 1745 -2628
rect 1809 -2692 1829 -2628
rect 110 -2708 1829 -2692
rect 110 -2772 1745 -2708
rect 1809 -2772 1829 -2708
rect 110 -2788 1829 -2772
rect 110 -2852 1745 -2788
rect 1809 -2852 1829 -2788
rect 110 -2868 1829 -2852
rect 110 -2932 1745 -2868
rect 1809 -2932 1829 -2868
rect 110 -2948 1829 -2932
rect 110 -3012 1745 -2948
rect 1809 -3012 1829 -2948
rect 110 -3028 1829 -3012
rect 110 -3092 1745 -3028
rect 1809 -3092 1829 -3028
rect 110 -3108 1829 -3092
rect 110 -3172 1745 -3108
rect 1809 -3172 1829 -3108
rect 110 -3188 1829 -3172
rect 110 -3252 1745 -3188
rect 1809 -3252 1829 -3188
rect 110 -3268 1829 -3252
rect 110 -3332 1745 -3268
rect 1809 -3332 1829 -3268
rect 110 -3390 1829 -3332
rect 1949 -1828 3668 -1770
rect 1949 -1892 3584 -1828
rect 3648 -1892 3668 -1828
rect 1949 -1908 3668 -1892
rect 1949 -1972 3584 -1908
rect 3648 -1972 3668 -1908
rect 1949 -1988 3668 -1972
rect 1949 -2052 3584 -1988
rect 3648 -2052 3668 -1988
rect 1949 -2068 3668 -2052
rect 1949 -2132 3584 -2068
rect 3648 -2132 3668 -2068
rect 1949 -2148 3668 -2132
rect 1949 -2212 3584 -2148
rect 3648 -2212 3668 -2148
rect 1949 -2228 3668 -2212
rect 1949 -2292 3584 -2228
rect 3648 -2292 3668 -2228
rect 1949 -2308 3668 -2292
rect 1949 -2372 3584 -2308
rect 3648 -2372 3668 -2308
rect 1949 -2388 3668 -2372
rect 1949 -2452 3584 -2388
rect 3648 -2452 3668 -2388
rect 1949 -2468 3668 -2452
rect 1949 -2532 3584 -2468
rect 3648 -2532 3668 -2468
rect 1949 -2548 3668 -2532
rect 1949 -2612 3584 -2548
rect 3648 -2612 3668 -2548
rect 1949 -2628 3668 -2612
rect 1949 -2692 3584 -2628
rect 3648 -2692 3668 -2628
rect 1949 -2708 3668 -2692
rect 1949 -2772 3584 -2708
rect 3648 -2772 3668 -2708
rect 1949 -2788 3668 -2772
rect 1949 -2852 3584 -2788
rect 3648 -2852 3668 -2788
rect 1949 -2868 3668 -2852
rect 1949 -2932 3584 -2868
rect 3648 -2932 3668 -2868
rect 1949 -2948 3668 -2932
rect 1949 -3012 3584 -2948
rect 3648 -3012 3668 -2948
rect 1949 -3028 3668 -3012
rect 1949 -3092 3584 -3028
rect 3648 -3092 3668 -3028
rect 1949 -3108 3668 -3092
rect 1949 -3172 3584 -3108
rect 3648 -3172 3668 -3108
rect 1949 -3188 3668 -3172
rect 1949 -3252 3584 -3188
rect 3648 -3252 3668 -3188
rect 1949 -3268 3668 -3252
rect 1949 -3332 3584 -3268
rect 3648 -3332 3668 -3268
rect 1949 -3390 3668 -3332
<< via3 >>
rect -1933 3268 -1869 3332
rect -1933 3188 -1869 3252
rect -1933 3108 -1869 3172
rect -1933 3028 -1869 3092
rect -1933 2948 -1869 3012
rect -1933 2868 -1869 2932
rect -1933 2788 -1869 2852
rect -1933 2708 -1869 2772
rect -1933 2628 -1869 2692
rect -1933 2548 -1869 2612
rect -1933 2468 -1869 2532
rect -1933 2388 -1869 2452
rect -1933 2308 -1869 2372
rect -1933 2228 -1869 2292
rect -1933 2148 -1869 2212
rect -1933 2068 -1869 2132
rect -1933 1988 -1869 2052
rect -1933 1908 -1869 1972
rect -1933 1828 -1869 1892
rect -94 3268 -30 3332
rect -94 3188 -30 3252
rect -94 3108 -30 3172
rect -94 3028 -30 3092
rect -94 2948 -30 3012
rect -94 2868 -30 2932
rect -94 2788 -30 2852
rect -94 2708 -30 2772
rect -94 2628 -30 2692
rect -94 2548 -30 2612
rect -94 2468 -30 2532
rect -94 2388 -30 2452
rect -94 2308 -30 2372
rect -94 2228 -30 2292
rect -94 2148 -30 2212
rect -94 2068 -30 2132
rect -94 1988 -30 2052
rect -94 1908 -30 1972
rect -94 1828 -30 1892
rect 1745 3268 1809 3332
rect 1745 3188 1809 3252
rect 1745 3108 1809 3172
rect 1745 3028 1809 3092
rect 1745 2948 1809 3012
rect 1745 2868 1809 2932
rect 1745 2788 1809 2852
rect 1745 2708 1809 2772
rect 1745 2628 1809 2692
rect 1745 2548 1809 2612
rect 1745 2468 1809 2532
rect 1745 2388 1809 2452
rect 1745 2308 1809 2372
rect 1745 2228 1809 2292
rect 1745 2148 1809 2212
rect 1745 2068 1809 2132
rect 1745 1988 1809 2052
rect 1745 1908 1809 1972
rect 1745 1828 1809 1892
rect 3584 3268 3648 3332
rect 3584 3188 3648 3252
rect 3584 3108 3648 3172
rect 3584 3028 3648 3092
rect 3584 2948 3648 3012
rect 3584 2868 3648 2932
rect 3584 2788 3648 2852
rect 3584 2708 3648 2772
rect 3584 2628 3648 2692
rect 3584 2548 3648 2612
rect 3584 2468 3648 2532
rect 3584 2388 3648 2452
rect 3584 2308 3648 2372
rect 3584 2228 3648 2292
rect 3584 2148 3648 2212
rect 3584 2068 3648 2132
rect 3584 1988 3648 2052
rect 3584 1908 3648 1972
rect 3584 1828 3648 1892
rect -1933 1548 -1869 1612
rect -1933 1468 -1869 1532
rect -1933 1388 -1869 1452
rect -1933 1308 -1869 1372
rect -1933 1228 -1869 1292
rect -1933 1148 -1869 1212
rect -1933 1068 -1869 1132
rect -1933 988 -1869 1052
rect -1933 908 -1869 972
rect -1933 828 -1869 892
rect -1933 748 -1869 812
rect -1933 668 -1869 732
rect -1933 588 -1869 652
rect -1933 508 -1869 572
rect -1933 428 -1869 492
rect -1933 348 -1869 412
rect -1933 268 -1869 332
rect -1933 188 -1869 252
rect -1933 108 -1869 172
rect -94 1548 -30 1612
rect -94 1468 -30 1532
rect -94 1388 -30 1452
rect -94 1308 -30 1372
rect -94 1228 -30 1292
rect -94 1148 -30 1212
rect -94 1068 -30 1132
rect -94 988 -30 1052
rect -94 908 -30 972
rect -94 828 -30 892
rect -94 748 -30 812
rect -94 668 -30 732
rect -94 588 -30 652
rect -94 508 -30 572
rect -94 428 -30 492
rect -94 348 -30 412
rect -94 268 -30 332
rect -94 188 -30 252
rect -94 108 -30 172
rect 1745 1548 1809 1612
rect 1745 1468 1809 1532
rect 1745 1388 1809 1452
rect 1745 1308 1809 1372
rect 1745 1228 1809 1292
rect 1745 1148 1809 1212
rect 1745 1068 1809 1132
rect 1745 988 1809 1052
rect 1745 908 1809 972
rect 1745 828 1809 892
rect 1745 748 1809 812
rect 1745 668 1809 732
rect 1745 588 1809 652
rect 1745 508 1809 572
rect 1745 428 1809 492
rect 1745 348 1809 412
rect 1745 268 1809 332
rect 1745 188 1809 252
rect 1745 108 1809 172
rect 3584 1548 3648 1612
rect 3584 1468 3648 1532
rect 3584 1388 3648 1452
rect 3584 1308 3648 1372
rect 3584 1228 3648 1292
rect 3584 1148 3648 1212
rect 3584 1068 3648 1132
rect 3584 988 3648 1052
rect 3584 908 3648 972
rect 3584 828 3648 892
rect 3584 748 3648 812
rect 3584 668 3648 732
rect 3584 588 3648 652
rect 3584 508 3648 572
rect 3584 428 3648 492
rect 3584 348 3648 412
rect 3584 268 3648 332
rect 3584 188 3648 252
rect 3584 108 3648 172
rect -1933 -172 -1869 -108
rect -1933 -252 -1869 -188
rect -1933 -332 -1869 -268
rect -1933 -412 -1869 -348
rect -1933 -492 -1869 -428
rect -1933 -572 -1869 -508
rect -1933 -652 -1869 -588
rect -1933 -732 -1869 -668
rect -1933 -812 -1869 -748
rect -1933 -892 -1869 -828
rect -1933 -972 -1869 -908
rect -1933 -1052 -1869 -988
rect -1933 -1132 -1869 -1068
rect -1933 -1212 -1869 -1148
rect -1933 -1292 -1869 -1228
rect -1933 -1372 -1869 -1308
rect -1933 -1452 -1869 -1388
rect -1933 -1532 -1869 -1468
rect -1933 -1612 -1869 -1548
rect -94 -172 -30 -108
rect -94 -252 -30 -188
rect -94 -332 -30 -268
rect -94 -412 -30 -348
rect -94 -492 -30 -428
rect -94 -572 -30 -508
rect -94 -652 -30 -588
rect -94 -732 -30 -668
rect -94 -812 -30 -748
rect -94 -892 -30 -828
rect -94 -972 -30 -908
rect -94 -1052 -30 -988
rect -94 -1132 -30 -1068
rect -94 -1212 -30 -1148
rect -94 -1292 -30 -1228
rect -94 -1372 -30 -1308
rect -94 -1452 -30 -1388
rect -94 -1532 -30 -1468
rect -94 -1612 -30 -1548
rect 1745 -172 1809 -108
rect 1745 -252 1809 -188
rect 1745 -332 1809 -268
rect 1745 -412 1809 -348
rect 1745 -492 1809 -428
rect 1745 -572 1809 -508
rect 1745 -652 1809 -588
rect 1745 -732 1809 -668
rect 1745 -812 1809 -748
rect 1745 -892 1809 -828
rect 1745 -972 1809 -908
rect 1745 -1052 1809 -988
rect 1745 -1132 1809 -1068
rect 1745 -1212 1809 -1148
rect 1745 -1292 1809 -1228
rect 1745 -1372 1809 -1308
rect 1745 -1452 1809 -1388
rect 1745 -1532 1809 -1468
rect 1745 -1612 1809 -1548
rect 3584 -172 3648 -108
rect 3584 -252 3648 -188
rect 3584 -332 3648 -268
rect 3584 -412 3648 -348
rect 3584 -492 3648 -428
rect 3584 -572 3648 -508
rect 3584 -652 3648 -588
rect 3584 -732 3648 -668
rect 3584 -812 3648 -748
rect 3584 -892 3648 -828
rect 3584 -972 3648 -908
rect 3584 -1052 3648 -988
rect 3584 -1132 3648 -1068
rect 3584 -1212 3648 -1148
rect 3584 -1292 3648 -1228
rect 3584 -1372 3648 -1308
rect 3584 -1452 3648 -1388
rect 3584 -1532 3648 -1468
rect 3584 -1612 3648 -1548
rect -1933 -1892 -1869 -1828
rect -1933 -1972 -1869 -1908
rect -1933 -2052 -1869 -1988
rect -1933 -2132 -1869 -2068
rect -1933 -2212 -1869 -2148
rect -1933 -2292 -1869 -2228
rect -1933 -2372 -1869 -2308
rect -1933 -2452 -1869 -2388
rect -1933 -2532 -1869 -2468
rect -1933 -2612 -1869 -2548
rect -1933 -2692 -1869 -2628
rect -1933 -2772 -1869 -2708
rect -1933 -2852 -1869 -2788
rect -1933 -2932 -1869 -2868
rect -1933 -3012 -1869 -2948
rect -1933 -3092 -1869 -3028
rect -1933 -3172 -1869 -3108
rect -1933 -3252 -1869 -3188
rect -1933 -3332 -1869 -3268
rect -94 -1892 -30 -1828
rect -94 -1972 -30 -1908
rect -94 -2052 -30 -1988
rect -94 -2132 -30 -2068
rect -94 -2212 -30 -2148
rect -94 -2292 -30 -2228
rect -94 -2372 -30 -2308
rect -94 -2452 -30 -2388
rect -94 -2532 -30 -2468
rect -94 -2612 -30 -2548
rect -94 -2692 -30 -2628
rect -94 -2772 -30 -2708
rect -94 -2852 -30 -2788
rect -94 -2932 -30 -2868
rect -94 -3012 -30 -2948
rect -94 -3092 -30 -3028
rect -94 -3172 -30 -3108
rect -94 -3252 -30 -3188
rect -94 -3332 -30 -3268
rect 1745 -1892 1809 -1828
rect 1745 -1972 1809 -1908
rect 1745 -2052 1809 -1988
rect 1745 -2132 1809 -2068
rect 1745 -2212 1809 -2148
rect 1745 -2292 1809 -2228
rect 1745 -2372 1809 -2308
rect 1745 -2452 1809 -2388
rect 1745 -2532 1809 -2468
rect 1745 -2612 1809 -2548
rect 1745 -2692 1809 -2628
rect 1745 -2772 1809 -2708
rect 1745 -2852 1809 -2788
rect 1745 -2932 1809 -2868
rect 1745 -3012 1809 -2948
rect 1745 -3092 1809 -3028
rect 1745 -3172 1809 -3108
rect 1745 -3252 1809 -3188
rect 1745 -3332 1809 -3268
rect 3584 -1892 3648 -1828
rect 3584 -1972 3648 -1908
rect 3584 -2052 3648 -1988
rect 3584 -2132 3648 -2068
rect 3584 -2212 3648 -2148
rect 3584 -2292 3648 -2228
rect 3584 -2372 3648 -2308
rect 3584 -2452 3648 -2388
rect 3584 -2532 3648 -2468
rect 3584 -2612 3648 -2548
rect 3584 -2692 3648 -2628
rect 3584 -2772 3648 -2708
rect 3584 -2852 3648 -2788
rect 3584 -2932 3648 -2868
rect 3584 -3012 3648 -2948
rect 3584 -3092 3648 -3028
rect 3584 -3172 3648 -3108
rect 3584 -3252 3648 -3188
rect 3584 -3332 3648 -3268
<< mimcap >>
rect -3468 3212 -2048 3290
rect -3468 1948 -3390 3212
rect -2126 1948 -2048 3212
rect -3468 1870 -2048 1948
rect -1629 3212 -209 3290
rect -1629 1948 -1551 3212
rect -287 1948 -209 3212
rect -1629 1870 -209 1948
rect 210 3212 1630 3290
rect 210 1948 288 3212
rect 1552 1948 1630 3212
rect 210 1870 1630 1948
rect 2049 3212 3469 3290
rect 2049 1948 2127 3212
rect 3391 1948 3469 3212
rect 2049 1870 3469 1948
rect -3468 1492 -2048 1570
rect -3468 228 -3390 1492
rect -2126 228 -2048 1492
rect -3468 150 -2048 228
rect -1629 1492 -209 1570
rect -1629 228 -1551 1492
rect -287 228 -209 1492
rect -1629 150 -209 228
rect 210 1492 1630 1570
rect 210 228 288 1492
rect 1552 228 1630 1492
rect 210 150 1630 228
rect 2049 1492 3469 1570
rect 2049 228 2127 1492
rect 3391 228 3469 1492
rect 2049 150 3469 228
rect -3468 -228 -2048 -150
rect -3468 -1492 -3390 -228
rect -2126 -1492 -2048 -228
rect -3468 -1570 -2048 -1492
rect -1629 -228 -209 -150
rect -1629 -1492 -1551 -228
rect -287 -1492 -209 -228
rect -1629 -1570 -209 -1492
rect 210 -228 1630 -150
rect 210 -1492 288 -228
rect 1552 -1492 1630 -228
rect 210 -1570 1630 -1492
rect 2049 -228 3469 -150
rect 2049 -1492 2127 -228
rect 3391 -1492 3469 -228
rect 2049 -1570 3469 -1492
rect -3468 -1948 -2048 -1870
rect -3468 -3212 -3390 -1948
rect -2126 -3212 -2048 -1948
rect -3468 -3290 -2048 -3212
rect -1629 -1948 -209 -1870
rect -1629 -3212 -1551 -1948
rect -287 -3212 -209 -1948
rect -1629 -3290 -209 -3212
rect 210 -1948 1630 -1870
rect 210 -3212 288 -1948
rect 1552 -3212 1630 -1948
rect 210 -3290 1630 -3212
rect 2049 -1948 3469 -1870
rect 2049 -3212 2127 -1948
rect 3391 -3212 3469 -1948
rect 2049 -3290 3469 -3212
<< mimcapcontact >>
rect -3390 1948 -2126 3212
rect -1551 1948 -287 3212
rect 288 1948 1552 3212
rect 2127 1948 3391 3212
rect -3390 228 -2126 1492
rect -1551 228 -287 1492
rect 288 228 1552 1492
rect 2127 228 3391 1492
rect -3390 -1492 -2126 -228
rect -1551 -1492 -287 -228
rect 288 -1492 1552 -228
rect 2127 -1492 3391 -228
rect -3390 -3212 -2126 -1948
rect -1551 -3212 -287 -1948
rect 288 -3212 1552 -1948
rect 2127 -3212 3391 -1948
<< metal4 >>
rect -3429 3212 -2087 3440
rect -3429 1948 -3390 3212
rect -2126 1948 -2087 3212
rect -3429 1492 -2087 1948
rect -3429 228 -3390 1492
rect -2126 228 -2087 1492
rect -3429 -228 -2087 228
rect -3429 -1492 -3390 -228
rect -2126 -1492 -2087 -228
rect -3429 -1948 -2087 -1492
rect -3429 -3212 -3390 -1948
rect -2126 -3212 -2087 -1948
rect -3429 -3740 -2087 -3212
rect -1980 3332 -1853 3729
rect -1980 3268 -1933 3332
rect -1869 3268 -1853 3332
rect -1980 3252 -1853 3268
rect -1980 3188 -1933 3252
rect -1869 3188 -1853 3252
rect -1980 3172 -1853 3188
rect -1980 3108 -1933 3172
rect -1869 3108 -1853 3172
rect -1980 3092 -1853 3108
rect -1980 3028 -1933 3092
rect -1869 3028 -1853 3092
rect -1980 3012 -1853 3028
rect -1980 2948 -1933 3012
rect -1869 2948 -1853 3012
rect -1980 2932 -1853 2948
rect -1980 2868 -1933 2932
rect -1869 2868 -1853 2932
rect -1980 2852 -1853 2868
rect -1980 2788 -1933 2852
rect -1869 2788 -1853 2852
rect -1980 2772 -1853 2788
rect -1980 2708 -1933 2772
rect -1869 2708 -1853 2772
rect -1980 2692 -1853 2708
rect -1980 2628 -1933 2692
rect -1869 2628 -1853 2692
rect -1980 2612 -1853 2628
rect -1980 2548 -1933 2612
rect -1869 2548 -1853 2612
rect -1980 2532 -1853 2548
rect -1980 2468 -1933 2532
rect -1869 2468 -1853 2532
rect -1980 2452 -1853 2468
rect -1980 2388 -1933 2452
rect -1869 2388 -1853 2452
rect -1980 2372 -1853 2388
rect -1980 2308 -1933 2372
rect -1869 2308 -1853 2372
rect -1980 2292 -1853 2308
rect -1980 2228 -1933 2292
rect -1869 2228 -1853 2292
rect -1980 2212 -1853 2228
rect -1980 2148 -1933 2212
rect -1869 2148 -1853 2212
rect -1980 2132 -1853 2148
rect -1980 2068 -1933 2132
rect -1869 2068 -1853 2132
rect -1980 2052 -1853 2068
rect -1980 1988 -1933 2052
rect -1869 1988 -1853 2052
rect -1980 1972 -1853 1988
rect -1980 1908 -1933 1972
rect -1869 1908 -1853 1972
rect -1980 1892 -1853 1908
rect -1980 1828 -1933 1892
rect -1869 1828 -1853 1892
rect -1980 1612 -1853 1828
rect -1980 1548 -1933 1612
rect -1869 1548 -1853 1612
rect -1980 1532 -1853 1548
rect -1980 1468 -1933 1532
rect -1869 1468 -1853 1532
rect -1980 1452 -1853 1468
rect -1980 1388 -1933 1452
rect -1869 1388 -1853 1452
rect -1980 1372 -1853 1388
rect -1980 1308 -1933 1372
rect -1869 1308 -1853 1372
rect -1980 1292 -1853 1308
rect -1980 1228 -1933 1292
rect -1869 1228 -1853 1292
rect -1980 1212 -1853 1228
rect -1980 1148 -1933 1212
rect -1869 1148 -1853 1212
rect -1980 1132 -1853 1148
rect -1980 1068 -1933 1132
rect -1869 1068 -1853 1132
rect -1980 1052 -1853 1068
rect -1980 988 -1933 1052
rect -1869 988 -1853 1052
rect -1980 972 -1853 988
rect -1980 908 -1933 972
rect -1869 908 -1853 972
rect -1980 892 -1853 908
rect -1980 828 -1933 892
rect -1869 828 -1853 892
rect -1980 812 -1853 828
rect -1980 748 -1933 812
rect -1869 748 -1853 812
rect -1980 732 -1853 748
rect -1980 668 -1933 732
rect -1869 668 -1853 732
rect -1980 652 -1853 668
rect -1980 588 -1933 652
rect -1869 588 -1853 652
rect -1980 572 -1853 588
rect -1980 508 -1933 572
rect -1869 508 -1853 572
rect -1980 492 -1853 508
rect -1980 428 -1933 492
rect -1869 428 -1853 492
rect -1980 412 -1853 428
rect -1980 348 -1933 412
rect -1869 348 -1853 412
rect -1980 332 -1853 348
rect -1980 268 -1933 332
rect -1869 268 -1853 332
rect -1980 252 -1853 268
rect -1980 188 -1933 252
rect -1869 188 -1853 252
rect -1980 172 -1853 188
rect -1980 108 -1933 172
rect -1869 108 -1853 172
rect -1980 -108 -1853 108
rect -1980 -172 -1933 -108
rect -1869 -172 -1853 -108
rect -1980 -188 -1853 -172
rect -1980 -252 -1933 -188
rect -1869 -252 -1853 -188
rect -1980 -268 -1853 -252
rect -1980 -332 -1933 -268
rect -1869 -332 -1853 -268
rect -1980 -348 -1853 -332
rect -1980 -412 -1933 -348
rect -1869 -412 -1853 -348
rect -1980 -428 -1853 -412
rect -1980 -492 -1933 -428
rect -1869 -492 -1853 -428
rect -1980 -508 -1853 -492
rect -1980 -572 -1933 -508
rect -1869 -572 -1853 -508
rect -1980 -588 -1853 -572
rect -1980 -652 -1933 -588
rect -1869 -652 -1853 -588
rect -1980 -668 -1853 -652
rect -1980 -732 -1933 -668
rect -1869 -732 -1853 -668
rect -1980 -748 -1853 -732
rect -1980 -812 -1933 -748
rect -1869 -812 -1853 -748
rect -1980 -828 -1853 -812
rect -1980 -892 -1933 -828
rect -1869 -892 -1853 -828
rect -1980 -908 -1853 -892
rect -1980 -972 -1933 -908
rect -1869 -972 -1853 -908
rect -1980 -988 -1853 -972
rect -1980 -1052 -1933 -988
rect -1869 -1052 -1853 -988
rect -1980 -1068 -1853 -1052
rect -1980 -1132 -1933 -1068
rect -1869 -1132 -1853 -1068
rect -1980 -1148 -1853 -1132
rect -1980 -1212 -1933 -1148
rect -1869 -1212 -1853 -1148
rect -1980 -1228 -1853 -1212
rect -1980 -1292 -1933 -1228
rect -1869 -1292 -1853 -1228
rect -1980 -1308 -1853 -1292
rect -1980 -1372 -1933 -1308
rect -1869 -1372 -1853 -1308
rect -1980 -1388 -1853 -1372
rect -1980 -1452 -1933 -1388
rect -1869 -1452 -1853 -1388
rect -1980 -1468 -1853 -1452
rect -1980 -1532 -1933 -1468
rect -1869 -1532 -1853 -1468
rect -1980 -1548 -1853 -1532
rect -1980 -1612 -1933 -1548
rect -1869 -1612 -1853 -1548
rect -1980 -1828 -1853 -1612
rect -1980 -1892 -1933 -1828
rect -1869 -1892 -1853 -1828
rect -1980 -1908 -1853 -1892
rect -1980 -1972 -1933 -1908
rect -1869 -1972 -1853 -1908
rect -1980 -1988 -1853 -1972
rect -1980 -2052 -1933 -1988
rect -1869 -2052 -1853 -1988
rect -1980 -2068 -1853 -2052
rect -1980 -2132 -1933 -2068
rect -1869 -2132 -1853 -2068
rect -1980 -2148 -1853 -2132
rect -1980 -2212 -1933 -2148
rect -1869 -2212 -1853 -2148
rect -1980 -2228 -1853 -2212
rect -1980 -2292 -1933 -2228
rect -1869 -2292 -1853 -2228
rect -1980 -2308 -1853 -2292
rect -1980 -2372 -1933 -2308
rect -1869 -2372 -1853 -2308
rect -1980 -2388 -1853 -2372
rect -1980 -2452 -1933 -2388
rect -1869 -2452 -1853 -2388
rect -1980 -2468 -1853 -2452
rect -1980 -2532 -1933 -2468
rect -1869 -2532 -1853 -2468
rect -1980 -2548 -1853 -2532
rect -1980 -2612 -1933 -2548
rect -1869 -2612 -1853 -2548
rect -1980 -2628 -1853 -2612
rect -1980 -2692 -1933 -2628
rect -1869 -2692 -1853 -2628
rect -1980 -2708 -1853 -2692
rect -1980 -2772 -1933 -2708
rect -1869 -2772 -1853 -2708
rect -1980 -2788 -1853 -2772
rect -1980 -2852 -1933 -2788
rect -1869 -2852 -1853 -2788
rect -1980 -2868 -1853 -2852
rect -1980 -2932 -1933 -2868
rect -1869 -2932 -1853 -2868
rect -1980 -2948 -1853 -2932
rect -1980 -3012 -1933 -2948
rect -1869 -3012 -1853 -2948
rect -1980 -3028 -1853 -3012
rect -1980 -3092 -1933 -3028
rect -1869 -3092 -1853 -3028
rect -1980 -3108 -1853 -3092
rect -1980 -3172 -1933 -3108
rect -1869 -3172 -1853 -3108
rect -1980 -3188 -1853 -3172
rect -1980 -3252 -1933 -3188
rect -1869 -3252 -1853 -3188
rect -1980 -3268 -1853 -3252
rect -1980 -3332 -1933 -3268
rect -1869 -3332 -1853 -3268
rect -1980 -3378 -1853 -3332
rect -1590 3212 -248 3440
rect -1590 1948 -1551 3212
rect -287 1948 -248 3212
rect -1590 1492 -248 1948
rect -1590 228 -1551 1492
rect -287 228 -248 1492
rect -1590 -228 -248 228
rect -1590 -1492 -1551 -228
rect -287 -1492 -248 -228
rect -1590 -1948 -248 -1492
rect -1590 -3212 -1551 -1948
rect -287 -3212 -248 -1948
rect -1590 -3697 -248 -3212
rect -141 3332 -14 3693
rect -141 3268 -94 3332
rect -30 3268 -14 3332
rect -141 3252 -14 3268
rect -141 3188 -94 3252
rect -30 3188 -14 3252
rect -141 3172 -14 3188
rect -141 3108 -94 3172
rect -30 3108 -14 3172
rect -141 3092 -14 3108
rect -141 3028 -94 3092
rect -30 3028 -14 3092
rect -141 3012 -14 3028
rect -141 2948 -94 3012
rect -30 2948 -14 3012
rect -141 2932 -14 2948
rect -141 2868 -94 2932
rect -30 2868 -14 2932
rect -141 2852 -14 2868
rect -141 2788 -94 2852
rect -30 2788 -14 2852
rect -141 2772 -14 2788
rect -141 2708 -94 2772
rect -30 2708 -14 2772
rect -141 2692 -14 2708
rect -141 2628 -94 2692
rect -30 2628 -14 2692
rect -141 2612 -14 2628
rect -141 2548 -94 2612
rect -30 2548 -14 2612
rect -141 2532 -14 2548
rect -141 2468 -94 2532
rect -30 2468 -14 2532
rect -141 2452 -14 2468
rect -141 2388 -94 2452
rect -30 2388 -14 2452
rect -141 2372 -14 2388
rect -141 2308 -94 2372
rect -30 2308 -14 2372
rect -141 2292 -14 2308
rect -141 2228 -94 2292
rect -30 2228 -14 2292
rect -141 2212 -14 2228
rect -141 2148 -94 2212
rect -30 2148 -14 2212
rect -141 2132 -14 2148
rect -141 2068 -94 2132
rect -30 2068 -14 2132
rect -141 2052 -14 2068
rect -141 1988 -94 2052
rect -30 1988 -14 2052
rect -141 1972 -14 1988
rect -141 1908 -94 1972
rect -30 1908 -14 1972
rect -141 1892 -14 1908
rect -141 1828 -94 1892
rect -30 1828 -14 1892
rect -141 1612 -14 1828
rect -141 1548 -94 1612
rect -30 1548 -14 1612
rect -141 1532 -14 1548
rect -141 1468 -94 1532
rect -30 1468 -14 1532
rect -141 1452 -14 1468
rect -141 1388 -94 1452
rect -30 1388 -14 1452
rect -141 1372 -14 1388
rect -141 1308 -94 1372
rect -30 1308 -14 1372
rect -141 1292 -14 1308
rect -141 1228 -94 1292
rect -30 1228 -14 1292
rect -141 1212 -14 1228
rect -141 1148 -94 1212
rect -30 1148 -14 1212
rect -141 1132 -14 1148
rect -141 1068 -94 1132
rect -30 1068 -14 1132
rect -141 1052 -14 1068
rect -141 988 -94 1052
rect -30 988 -14 1052
rect -141 972 -14 988
rect -141 908 -94 972
rect -30 908 -14 972
rect -141 892 -14 908
rect -141 828 -94 892
rect -30 828 -14 892
rect -141 812 -14 828
rect -141 748 -94 812
rect -30 748 -14 812
rect -141 732 -14 748
rect -141 668 -94 732
rect -30 668 -14 732
rect -141 652 -14 668
rect -141 588 -94 652
rect -30 588 -14 652
rect -141 572 -14 588
rect -141 508 -94 572
rect -30 508 -14 572
rect -141 492 -14 508
rect -141 428 -94 492
rect -30 428 -14 492
rect -141 412 -14 428
rect -141 348 -94 412
rect -30 348 -14 412
rect -141 332 -14 348
rect -141 268 -94 332
rect -30 268 -14 332
rect -141 252 -14 268
rect -141 188 -94 252
rect -30 188 -14 252
rect -141 172 -14 188
rect -141 108 -94 172
rect -30 108 -14 172
rect -141 -108 -14 108
rect -141 -172 -94 -108
rect -30 -172 -14 -108
rect -141 -188 -14 -172
rect -141 -252 -94 -188
rect -30 -252 -14 -188
rect -141 -268 -14 -252
rect -141 -332 -94 -268
rect -30 -332 -14 -268
rect -141 -348 -14 -332
rect -141 -412 -94 -348
rect -30 -412 -14 -348
rect -141 -428 -14 -412
rect -141 -492 -94 -428
rect -30 -492 -14 -428
rect -141 -508 -14 -492
rect -141 -572 -94 -508
rect -30 -572 -14 -508
rect -141 -588 -14 -572
rect -141 -652 -94 -588
rect -30 -652 -14 -588
rect -141 -668 -14 -652
rect -141 -732 -94 -668
rect -30 -732 -14 -668
rect -141 -748 -14 -732
rect -141 -812 -94 -748
rect -30 -812 -14 -748
rect -141 -828 -14 -812
rect -141 -892 -94 -828
rect -30 -892 -14 -828
rect -141 -908 -14 -892
rect -141 -972 -94 -908
rect -30 -972 -14 -908
rect -141 -988 -14 -972
rect -141 -1052 -94 -988
rect -30 -1052 -14 -988
rect -141 -1068 -14 -1052
rect -141 -1132 -94 -1068
rect -30 -1132 -14 -1068
rect -141 -1148 -14 -1132
rect -141 -1212 -94 -1148
rect -30 -1212 -14 -1148
rect -141 -1228 -14 -1212
rect -141 -1292 -94 -1228
rect -30 -1292 -14 -1228
rect -141 -1308 -14 -1292
rect -141 -1372 -94 -1308
rect -30 -1372 -14 -1308
rect -141 -1388 -14 -1372
rect -141 -1452 -94 -1388
rect -30 -1452 -14 -1388
rect -141 -1468 -14 -1452
rect -141 -1532 -94 -1468
rect -30 -1532 -14 -1468
rect -141 -1548 -14 -1532
rect -141 -1612 -94 -1548
rect -30 -1612 -14 -1548
rect -141 -1828 -14 -1612
rect -141 -1892 -94 -1828
rect -30 -1892 -14 -1828
rect -141 -1908 -14 -1892
rect -141 -1972 -94 -1908
rect -30 -1972 -14 -1908
rect -141 -1988 -14 -1972
rect -141 -2052 -94 -1988
rect -30 -2052 -14 -1988
rect -141 -2068 -14 -2052
rect -141 -2132 -94 -2068
rect -30 -2132 -14 -2068
rect -141 -2148 -14 -2132
rect -141 -2212 -94 -2148
rect -30 -2212 -14 -2148
rect -141 -2228 -14 -2212
rect -141 -2292 -94 -2228
rect -30 -2292 -14 -2228
rect -141 -2308 -14 -2292
rect -141 -2372 -94 -2308
rect -30 -2372 -14 -2308
rect -141 -2388 -14 -2372
rect -141 -2452 -94 -2388
rect -30 -2452 -14 -2388
rect -141 -2468 -14 -2452
rect -141 -2532 -94 -2468
rect -30 -2532 -14 -2468
rect -141 -2548 -14 -2532
rect -141 -2612 -94 -2548
rect -30 -2612 -14 -2548
rect -141 -2628 -14 -2612
rect -141 -2692 -94 -2628
rect -30 -2692 -14 -2628
rect -141 -2708 -14 -2692
rect -141 -2772 -94 -2708
rect -30 -2772 -14 -2708
rect -141 -2788 -14 -2772
rect -141 -2852 -94 -2788
rect -30 -2852 -14 -2788
rect -141 -2868 -14 -2852
rect -141 -2932 -94 -2868
rect -30 -2932 -14 -2868
rect -141 -2948 -14 -2932
rect -141 -3012 -94 -2948
rect -30 -3012 -14 -2948
rect -141 -3028 -14 -3012
rect -141 -3092 -94 -3028
rect -30 -3092 -14 -3028
rect -141 -3108 -14 -3092
rect -141 -3172 -94 -3108
rect -30 -3172 -14 -3108
rect -141 -3188 -14 -3172
rect -141 -3252 -94 -3188
rect -30 -3252 -14 -3188
rect -141 -3268 -14 -3252
rect -141 -3332 -94 -3268
rect -30 -3332 -14 -3268
rect -141 -3378 -14 -3332
rect 249 3212 1591 3440
rect 249 1948 288 3212
rect 1552 1948 1591 3212
rect 249 1492 1591 1948
rect 249 228 288 1492
rect 1552 228 1591 1492
rect 249 -228 1591 228
rect 249 -1492 288 -228
rect 1552 -1492 1591 -228
rect 249 -1948 1591 -1492
rect 249 -3212 288 -1948
rect 1552 -3212 1591 -1948
rect 249 -3730 1591 -3212
rect 1698 3332 1825 3705
rect 1698 3268 1745 3332
rect 1809 3268 1825 3332
rect 1698 3252 1825 3268
rect 1698 3188 1745 3252
rect 1809 3188 1825 3252
rect 1698 3172 1825 3188
rect 1698 3108 1745 3172
rect 1809 3108 1825 3172
rect 1698 3092 1825 3108
rect 1698 3028 1745 3092
rect 1809 3028 1825 3092
rect 1698 3012 1825 3028
rect 1698 2948 1745 3012
rect 1809 2948 1825 3012
rect 1698 2932 1825 2948
rect 1698 2868 1745 2932
rect 1809 2868 1825 2932
rect 1698 2852 1825 2868
rect 1698 2788 1745 2852
rect 1809 2788 1825 2852
rect 1698 2772 1825 2788
rect 1698 2708 1745 2772
rect 1809 2708 1825 2772
rect 1698 2692 1825 2708
rect 1698 2628 1745 2692
rect 1809 2628 1825 2692
rect 1698 2612 1825 2628
rect 1698 2548 1745 2612
rect 1809 2548 1825 2612
rect 1698 2532 1825 2548
rect 1698 2468 1745 2532
rect 1809 2468 1825 2532
rect 1698 2452 1825 2468
rect 1698 2388 1745 2452
rect 1809 2388 1825 2452
rect 1698 2372 1825 2388
rect 1698 2308 1745 2372
rect 1809 2308 1825 2372
rect 1698 2292 1825 2308
rect 1698 2228 1745 2292
rect 1809 2228 1825 2292
rect 1698 2212 1825 2228
rect 1698 2148 1745 2212
rect 1809 2148 1825 2212
rect 1698 2132 1825 2148
rect 1698 2068 1745 2132
rect 1809 2068 1825 2132
rect 1698 2052 1825 2068
rect 1698 1988 1745 2052
rect 1809 1988 1825 2052
rect 1698 1972 1825 1988
rect 1698 1908 1745 1972
rect 1809 1908 1825 1972
rect 1698 1892 1825 1908
rect 1698 1828 1745 1892
rect 1809 1828 1825 1892
rect 1698 1612 1825 1828
rect 1698 1548 1745 1612
rect 1809 1548 1825 1612
rect 1698 1532 1825 1548
rect 1698 1468 1745 1532
rect 1809 1468 1825 1532
rect 1698 1452 1825 1468
rect 1698 1388 1745 1452
rect 1809 1388 1825 1452
rect 1698 1372 1825 1388
rect 1698 1308 1745 1372
rect 1809 1308 1825 1372
rect 1698 1292 1825 1308
rect 1698 1228 1745 1292
rect 1809 1228 1825 1292
rect 1698 1212 1825 1228
rect 1698 1148 1745 1212
rect 1809 1148 1825 1212
rect 1698 1132 1825 1148
rect 1698 1068 1745 1132
rect 1809 1068 1825 1132
rect 1698 1052 1825 1068
rect 1698 988 1745 1052
rect 1809 988 1825 1052
rect 1698 972 1825 988
rect 1698 908 1745 972
rect 1809 908 1825 972
rect 1698 892 1825 908
rect 1698 828 1745 892
rect 1809 828 1825 892
rect 1698 812 1825 828
rect 1698 748 1745 812
rect 1809 748 1825 812
rect 1698 732 1825 748
rect 1698 668 1745 732
rect 1809 668 1825 732
rect 1698 652 1825 668
rect 1698 588 1745 652
rect 1809 588 1825 652
rect 1698 572 1825 588
rect 1698 508 1745 572
rect 1809 508 1825 572
rect 1698 492 1825 508
rect 1698 428 1745 492
rect 1809 428 1825 492
rect 1698 412 1825 428
rect 1698 348 1745 412
rect 1809 348 1825 412
rect 1698 332 1825 348
rect 1698 268 1745 332
rect 1809 268 1825 332
rect 1698 252 1825 268
rect 1698 188 1745 252
rect 1809 188 1825 252
rect 1698 172 1825 188
rect 1698 108 1745 172
rect 1809 108 1825 172
rect 1698 -108 1825 108
rect 1698 -172 1745 -108
rect 1809 -172 1825 -108
rect 1698 -188 1825 -172
rect 1698 -252 1745 -188
rect 1809 -252 1825 -188
rect 1698 -268 1825 -252
rect 1698 -332 1745 -268
rect 1809 -332 1825 -268
rect 1698 -348 1825 -332
rect 1698 -412 1745 -348
rect 1809 -412 1825 -348
rect 1698 -428 1825 -412
rect 1698 -492 1745 -428
rect 1809 -492 1825 -428
rect 1698 -508 1825 -492
rect 1698 -572 1745 -508
rect 1809 -572 1825 -508
rect 1698 -588 1825 -572
rect 1698 -652 1745 -588
rect 1809 -652 1825 -588
rect 1698 -668 1825 -652
rect 1698 -732 1745 -668
rect 1809 -732 1825 -668
rect 1698 -748 1825 -732
rect 1698 -812 1745 -748
rect 1809 -812 1825 -748
rect 1698 -828 1825 -812
rect 1698 -892 1745 -828
rect 1809 -892 1825 -828
rect 1698 -908 1825 -892
rect 1698 -972 1745 -908
rect 1809 -972 1825 -908
rect 1698 -988 1825 -972
rect 1698 -1052 1745 -988
rect 1809 -1052 1825 -988
rect 1698 -1068 1825 -1052
rect 1698 -1132 1745 -1068
rect 1809 -1132 1825 -1068
rect 1698 -1148 1825 -1132
rect 1698 -1212 1745 -1148
rect 1809 -1212 1825 -1148
rect 1698 -1228 1825 -1212
rect 1698 -1292 1745 -1228
rect 1809 -1292 1825 -1228
rect 1698 -1308 1825 -1292
rect 1698 -1372 1745 -1308
rect 1809 -1372 1825 -1308
rect 1698 -1388 1825 -1372
rect 1698 -1452 1745 -1388
rect 1809 -1452 1825 -1388
rect 1698 -1468 1825 -1452
rect 1698 -1532 1745 -1468
rect 1809 -1532 1825 -1468
rect 1698 -1548 1825 -1532
rect 1698 -1612 1745 -1548
rect 1809 -1612 1825 -1548
rect 1698 -1828 1825 -1612
rect 1698 -1892 1745 -1828
rect 1809 -1892 1825 -1828
rect 1698 -1908 1825 -1892
rect 1698 -1972 1745 -1908
rect 1809 -1972 1825 -1908
rect 1698 -1988 1825 -1972
rect 1698 -2052 1745 -1988
rect 1809 -2052 1825 -1988
rect 1698 -2068 1825 -2052
rect 1698 -2132 1745 -2068
rect 1809 -2132 1825 -2068
rect 1698 -2148 1825 -2132
rect 1698 -2212 1745 -2148
rect 1809 -2212 1825 -2148
rect 1698 -2228 1825 -2212
rect 1698 -2292 1745 -2228
rect 1809 -2292 1825 -2228
rect 1698 -2308 1825 -2292
rect 1698 -2372 1745 -2308
rect 1809 -2372 1825 -2308
rect 1698 -2388 1825 -2372
rect 1698 -2452 1745 -2388
rect 1809 -2452 1825 -2388
rect 1698 -2468 1825 -2452
rect 1698 -2532 1745 -2468
rect 1809 -2532 1825 -2468
rect 1698 -2548 1825 -2532
rect 1698 -2612 1745 -2548
rect 1809 -2612 1825 -2548
rect 1698 -2628 1825 -2612
rect 1698 -2692 1745 -2628
rect 1809 -2692 1825 -2628
rect 1698 -2708 1825 -2692
rect 1698 -2772 1745 -2708
rect 1809 -2772 1825 -2708
rect 1698 -2788 1825 -2772
rect 1698 -2852 1745 -2788
rect 1809 -2852 1825 -2788
rect 1698 -2868 1825 -2852
rect 1698 -2932 1745 -2868
rect 1809 -2932 1825 -2868
rect 1698 -2948 1825 -2932
rect 1698 -3012 1745 -2948
rect 1809 -3012 1825 -2948
rect 1698 -3028 1825 -3012
rect 1698 -3092 1745 -3028
rect 1809 -3092 1825 -3028
rect 1698 -3108 1825 -3092
rect 1698 -3172 1745 -3108
rect 1809 -3172 1825 -3108
rect 1698 -3188 1825 -3172
rect 1698 -3252 1745 -3188
rect 1809 -3252 1825 -3188
rect 1698 -3268 1825 -3252
rect 1698 -3332 1745 -3268
rect 1809 -3332 1825 -3268
rect 1698 -3378 1825 -3332
rect 2088 3212 3430 3440
rect 2088 1948 2127 3212
rect 3391 1948 3430 3212
rect 2088 1492 3430 1948
rect 2088 228 2127 1492
rect 3391 228 3430 1492
rect 2088 -228 3430 228
rect 2088 -1492 2127 -228
rect 3391 -1492 3430 -228
rect 2088 -1948 3430 -1492
rect 2088 -3212 2127 -1948
rect 3391 -3212 3430 -1948
rect 2088 -3814 3430 -3212
rect 3537 3332 3664 3729
rect 3537 3268 3584 3332
rect 3648 3268 3664 3332
rect 3537 3252 3664 3268
rect 3537 3188 3584 3252
rect 3648 3188 3664 3252
rect 3537 3172 3664 3188
rect 3537 3108 3584 3172
rect 3648 3108 3664 3172
rect 3537 3092 3664 3108
rect 3537 3028 3584 3092
rect 3648 3028 3664 3092
rect 3537 3012 3664 3028
rect 3537 2948 3584 3012
rect 3648 2948 3664 3012
rect 3537 2932 3664 2948
rect 3537 2868 3584 2932
rect 3648 2868 3664 2932
rect 3537 2852 3664 2868
rect 3537 2788 3584 2852
rect 3648 2788 3664 2852
rect 3537 2772 3664 2788
rect 3537 2708 3584 2772
rect 3648 2708 3664 2772
rect 3537 2692 3664 2708
rect 3537 2628 3584 2692
rect 3648 2628 3664 2692
rect 3537 2612 3664 2628
rect 3537 2548 3584 2612
rect 3648 2548 3664 2612
rect 3537 2532 3664 2548
rect 3537 2468 3584 2532
rect 3648 2468 3664 2532
rect 3537 2452 3664 2468
rect 3537 2388 3584 2452
rect 3648 2388 3664 2452
rect 3537 2372 3664 2388
rect 3537 2308 3584 2372
rect 3648 2308 3664 2372
rect 3537 2292 3664 2308
rect 3537 2228 3584 2292
rect 3648 2228 3664 2292
rect 3537 2212 3664 2228
rect 3537 2148 3584 2212
rect 3648 2148 3664 2212
rect 3537 2132 3664 2148
rect 3537 2068 3584 2132
rect 3648 2068 3664 2132
rect 3537 2052 3664 2068
rect 3537 1988 3584 2052
rect 3648 1988 3664 2052
rect 3537 1972 3664 1988
rect 3537 1908 3584 1972
rect 3648 1908 3664 1972
rect 3537 1892 3664 1908
rect 3537 1828 3584 1892
rect 3648 1828 3664 1892
rect 3537 1612 3664 1828
rect 3537 1548 3584 1612
rect 3648 1548 3664 1612
rect 3537 1532 3664 1548
rect 3537 1468 3584 1532
rect 3648 1468 3664 1532
rect 3537 1452 3664 1468
rect 3537 1388 3584 1452
rect 3648 1388 3664 1452
rect 3537 1372 3664 1388
rect 3537 1308 3584 1372
rect 3648 1308 3664 1372
rect 3537 1292 3664 1308
rect 3537 1228 3584 1292
rect 3648 1228 3664 1292
rect 3537 1212 3664 1228
rect 3537 1148 3584 1212
rect 3648 1148 3664 1212
rect 3537 1132 3664 1148
rect 3537 1068 3584 1132
rect 3648 1068 3664 1132
rect 3537 1052 3664 1068
rect 3537 988 3584 1052
rect 3648 988 3664 1052
rect 3537 972 3664 988
rect 3537 908 3584 972
rect 3648 908 3664 972
rect 3537 892 3664 908
rect 3537 828 3584 892
rect 3648 828 3664 892
rect 3537 812 3664 828
rect 3537 748 3584 812
rect 3648 748 3664 812
rect 3537 732 3664 748
rect 3537 668 3584 732
rect 3648 668 3664 732
rect 3537 652 3664 668
rect 3537 588 3584 652
rect 3648 588 3664 652
rect 3537 572 3664 588
rect 3537 508 3584 572
rect 3648 508 3664 572
rect 3537 492 3664 508
rect 3537 428 3584 492
rect 3648 428 3664 492
rect 3537 412 3664 428
rect 3537 348 3584 412
rect 3648 348 3664 412
rect 3537 332 3664 348
rect 3537 268 3584 332
rect 3648 268 3664 332
rect 3537 252 3664 268
rect 3537 188 3584 252
rect 3648 188 3664 252
rect 3537 172 3664 188
rect 3537 108 3584 172
rect 3648 108 3664 172
rect 3537 -108 3664 108
rect 3537 -172 3584 -108
rect 3648 -172 3664 -108
rect 3537 -188 3664 -172
rect 3537 -252 3584 -188
rect 3648 -252 3664 -188
rect 3537 -268 3664 -252
rect 3537 -332 3584 -268
rect 3648 -332 3664 -268
rect 3537 -348 3664 -332
rect 3537 -412 3584 -348
rect 3648 -412 3664 -348
rect 3537 -428 3664 -412
rect 3537 -492 3584 -428
rect 3648 -492 3664 -428
rect 3537 -508 3664 -492
rect 3537 -572 3584 -508
rect 3648 -572 3664 -508
rect 3537 -588 3664 -572
rect 3537 -652 3584 -588
rect 3648 -652 3664 -588
rect 3537 -668 3664 -652
rect 3537 -732 3584 -668
rect 3648 -732 3664 -668
rect 3537 -748 3664 -732
rect 3537 -812 3584 -748
rect 3648 -812 3664 -748
rect 3537 -828 3664 -812
rect 3537 -892 3584 -828
rect 3648 -892 3664 -828
rect 3537 -908 3664 -892
rect 3537 -972 3584 -908
rect 3648 -972 3664 -908
rect 3537 -988 3664 -972
rect 3537 -1052 3584 -988
rect 3648 -1052 3664 -988
rect 3537 -1068 3664 -1052
rect 3537 -1132 3584 -1068
rect 3648 -1132 3664 -1068
rect 3537 -1148 3664 -1132
rect 3537 -1212 3584 -1148
rect 3648 -1212 3664 -1148
rect 3537 -1228 3664 -1212
rect 3537 -1292 3584 -1228
rect 3648 -1292 3664 -1228
rect 3537 -1308 3664 -1292
rect 3537 -1372 3584 -1308
rect 3648 -1372 3664 -1308
rect 3537 -1388 3664 -1372
rect 3537 -1452 3584 -1388
rect 3648 -1452 3664 -1388
rect 3537 -1468 3664 -1452
rect 3537 -1532 3584 -1468
rect 3648 -1532 3664 -1468
rect 3537 -1548 3664 -1532
rect 3537 -1612 3584 -1548
rect 3648 -1612 3664 -1548
rect 3537 -1828 3664 -1612
rect 3537 -1892 3584 -1828
rect 3648 -1892 3664 -1828
rect 3537 -1908 3664 -1892
rect 3537 -1972 3584 -1908
rect 3648 -1972 3664 -1908
rect 3537 -1988 3664 -1972
rect 3537 -2052 3584 -1988
rect 3648 -2052 3664 -1988
rect 3537 -2068 3664 -2052
rect 3537 -2132 3584 -2068
rect 3648 -2132 3664 -2068
rect 3537 -2148 3664 -2132
rect 3537 -2212 3584 -2148
rect 3648 -2212 3664 -2148
rect 3537 -2228 3664 -2212
rect 3537 -2292 3584 -2228
rect 3648 -2292 3664 -2228
rect 3537 -2308 3664 -2292
rect 3537 -2372 3584 -2308
rect 3648 -2372 3664 -2308
rect 3537 -2388 3664 -2372
rect 3537 -2452 3584 -2388
rect 3648 -2452 3664 -2388
rect 3537 -2468 3664 -2452
rect 3537 -2532 3584 -2468
rect 3648 -2532 3664 -2468
rect 3537 -2548 3664 -2532
rect 3537 -2612 3584 -2548
rect 3648 -2612 3664 -2548
rect 3537 -2628 3664 -2612
rect 3537 -2692 3584 -2628
rect 3648 -2692 3664 -2628
rect 3537 -2708 3664 -2692
rect 3537 -2772 3584 -2708
rect 3648 -2772 3664 -2708
rect 3537 -2788 3664 -2772
rect 3537 -2852 3584 -2788
rect 3648 -2852 3664 -2788
rect 3537 -2868 3664 -2852
rect 3537 -2932 3584 -2868
rect 3648 -2932 3664 -2868
rect 3537 -2948 3664 -2932
rect 3537 -3012 3584 -2948
rect 3648 -3012 3664 -2948
rect 3537 -3028 3664 -3012
rect 3537 -3092 3584 -3028
rect 3648 -3092 3664 -3028
rect 3537 -3108 3664 -3092
rect 3537 -3172 3584 -3108
rect 3648 -3172 3664 -3108
rect 3537 -3188 3664 -3172
rect 3537 -3252 3584 -3188
rect 3648 -3252 3664 -3188
rect 3537 -3268 3664 -3252
rect 3537 -3332 3584 -3268
rect 3648 -3332 3664 -3268
rect 3537 -3378 3664 -3332
<< properties >>
string FIXED_BBOX 1749 1770 3369 3390
<< end >>
