magic
tech sky130A
timestamp 1666407406
<< nmos >>
rect -15 -285 15 285
<< ndiff >>
rect -44 279 -15 285
rect -44 -279 -38 279
rect -21 -279 -15 279
rect -44 -285 -15 -279
rect 15 279 44 285
rect 15 -279 21 279
rect 38 -279 44 279
rect 15 -285 44 -279
<< ndiffc >>
rect -38 -279 -21 279
rect 21 -279 38 279
<< poly >>
rect -15 285 15 298
rect -15 -298 15 -285
<< locali >>
rect -38 279 -21 287
rect -38 -287 -21 -279
rect 21 279 38 287
rect 21 -287 38 -279
<< viali >>
rect -38 -279 -21 279
rect 21 -279 38 279
<< metal1 >>
rect -41 279 -18 285
rect -41 -279 -38 279
rect -21 -279 -18 279
rect -41 -285 -18 -279
rect 18 279 41 285
rect 18 -279 21 279
rect 38 -279 41 279
rect 18 -285 41 -279
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.7 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
