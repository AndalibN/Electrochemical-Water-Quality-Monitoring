magic
tech sky130A
magscale 1 2
timestamp 1667328903
use sky130_fd_pr__res_xhigh_po_0p35_QTYTGM  sky130_fd_pr__res_xhigh_po_0p35_QTYTGM_0
timestamp 1667328903
transform 0 -1 1432 1 0 673
box -1134 -1432 673 1432
<< labels >>
rlabel space 1298 -334 1298 -334 7 gnd
rlabel space 216 34 216 34 7 top
<< end >>
