magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -294 -2514 294 2548
<< pmos >>
rect -200 -2414 200 2486
<< pdiff >>
rect -258 2467 -200 2486
rect -258 2433 -246 2467
rect -212 2433 -200 2467
rect -258 2399 -200 2433
rect -258 2365 -246 2399
rect -212 2365 -200 2399
rect -258 2331 -200 2365
rect -258 2297 -246 2331
rect -212 2297 -200 2331
rect -258 2263 -200 2297
rect -258 2229 -246 2263
rect -212 2229 -200 2263
rect -258 2195 -200 2229
rect -258 2161 -246 2195
rect -212 2161 -200 2195
rect -258 2127 -200 2161
rect -258 2093 -246 2127
rect -212 2093 -200 2127
rect -258 2059 -200 2093
rect -258 2025 -246 2059
rect -212 2025 -200 2059
rect -258 1991 -200 2025
rect -258 1957 -246 1991
rect -212 1957 -200 1991
rect -258 1923 -200 1957
rect -258 1889 -246 1923
rect -212 1889 -200 1923
rect -258 1855 -200 1889
rect -258 1821 -246 1855
rect -212 1821 -200 1855
rect -258 1787 -200 1821
rect -258 1753 -246 1787
rect -212 1753 -200 1787
rect -258 1719 -200 1753
rect -258 1685 -246 1719
rect -212 1685 -200 1719
rect -258 1651 -200 1685
rect -258 1617 -246 1651
rect -212 1617 -200 1651
rect -258 1583 -200 1617
rect -258 1549 -246 1583
rect -212 1549 -200 1583
rect -258 1515 -200 1549
rect -258 1481 -246 1515
rect -212 1481 -200 1515
rect -258 1447 -200 1481
rect -258 1413 -246 1447
rect -212 1413 -200 1447
rect -258 1379 -200 1413
rect -258 1345 -246 1379
rect -212 1345 -200 1379
rect -258 1311 -200 1345
rect -258 1277 -246 1311
rect -212 1277 -200 1311
rect -258 1243 -200 1277
rect -258 1209 -246 1243
rect -212 1209 -200 1243
rect -258 1175 -200 1209
rect -258 1141 -246 1175
rect -212 1141 -200 1175
rect -258 1107 -200 1141
rect -258 1073 -246 1107
rect -212 1073 -200 1107
rect -258 1039 -200 1073
rect -258 1005 -246 1039
rect -212 1005 -200 1039
rect -258 971 -200 1005
rect -258 937 -246 971
rect -212 937 -200 971
rect -258 903 -200 937
rect -258 869 -246 903
rect -212 869 -200 903
rect -258 835 -200 869
rect -258 801 -246 835
rect -212 801 -200 835
rect -258 767 -200 801
rect -258 733 -246 767
rect -212 733 -200 767
rect -258 699 -200 733
rect -258 665 -246 699
rect -212 665 -200 699
rect -258 631 -200 665
rect -258 597 -246 631
rect -212 597 -200 631
rect -258 563 -200 597
rect -258 529 -246 563
rect -212 529 -200 563
rect -258 495 -200 529
rect -258 461 -246 495
rect -212 461 -200 495
rect -258 427 -200 461
rect -258 393 -246 427
rect -212 393 -200 427
rect -258 359 -200 393
rect -258 325 -246 359
rect -212 325 -200 359
rect -258 291 -200 325
rect -258 257 -246 291
rect -212 257 -200 291
rect -258 223 -200 257
rect -258 189 -246 223
rect -212 189 -200 223
rect -258 155 -200 189
rect -258 121 -246 155
rect -212 121 -200 155
rect -258 87 -200 121
rect -258 53 -246 87
rect -212 53 -200 87
rect -258 19 -200 53
rect -258 -15 -246 19
rect -212 -15 -200 19
rect -258 -49 -200 -15
rect -258 -83 -246 -49
rect -212 -83 -200 -49
rect -258 -117 -200 -83
rect -258 -151 -246 -117
rect -212 -151 -200 -117
rect -258 -185 -200 -151
rect -258 -219 -246 -185
rect -212 -219 -200 -185
rect -258 -253 -200 -219
rect -258 -287 -246 -253
rect -212 -287 -200 -253
rect -258 -321 -200 -287
rect -258 -355 -246 -321
rect -212 -355 -200 -321
rect -258 -389 -200 -355
rect -258 -423 -246 -389
rect -212 -423 -200 -389
rect -258 -457 -200 -423
rect -258 -491 -246 -457
rect -212 -491 -200 -457
rect -258 -525 -200 -491
rect -258 -559 -246 -525
rect -212 -559 -200 -525
rect -258 -593 -200 -559
rect -258 -627 -246 -593
rect -212 -627 -200 -593
rect -258 -661 -200 -627
rect -258 -695 -246 -661
rect -212 -695 -200 -661
rect -258 -729 -200 -695
rect -258 -763 -246 -729
rect -212 -763 -200 -729
rect -258 -797 -200 -763
rect -258 -831 -246 -797
rect -212 -831 -200 -797
rect -258 -865 -200 -831
rect -258 -899 -246 -865
rect -212 -899 -200 -865
rect -258 -933 -200 -899
rect -258 -967 -246 -933
rect -212 -967 -200 -933
rect -258 -1001 -200 -967
rect -258 -1035 -246 -1001
rect -212 -1035 -200 -1001
rect -258 -1069 -200 -1035
rect -258 -1103 -246 -1069
rect -212 -1103 -200 -1069
rect -258 -1137 -200 -1103
rect -258 -1171 -246 -1137
rect -212 -1171 -200 -1137
rect -258 -1205 -200 -1171
rect -258 -1239 -246 -1205
rect -212 -1239 -200 -1205
rect -258 -1273 -200 -1239
rect -258 -1307 -246 -1273
rect -212 -1307 -200 -1273
rect -258 -1341 -200 -1307
rect -258 -1375 -246 -1341
rect -212 -1375 -200 -1341
rect -258 -1409 -200 -1375
rect -258 -1443 -246 -1409
rect -212 -1443 -200 -1409
rect -258 -1477 -200 -1443
rect -258 -1511 -246 -1477
rect -212 -1511 -200 -1477
rect -258 -1545 -200 -1511
rect -258 -1579 -246 -1545
rect -212 -1579 -200 -1545
rect -258 -1613 -200 -1579
rect -258 -1647 -246 -1613
rect -212 -1647 -200 -1613
rect -258 -1681 -200 -1647
rect -258 -1715 -246 -1681
rect -212 -1715 -200 -1681
rect -258 -1749 -200 -1715
rect -258 -1783 -246 -1749
rect -212 -1783 -200 -1749
rect -258 -1817 -200 -1783
rect -258 -1851 -246 -1817
rect -212 -1851 -200 -1817
rect -258 -1885 -200 -1851
rect -258 -1919 -246 -1885
rect -212 -1919 -200 -1885
rect -258 -1953 -200 -1919
rect -258 -1987 -246 -1953
rect -212 -1987 -200 -1953
rect -258 -2021 -200 -1987
rect -258 -2055 -246 -2021
rect -212 -2055 -200 -2021
rect -258 -2089 -200 -2055
rect -258 -2123 -246 -2089
rect -212 -2123 -200 -2089
rect -258 -2157 -200 -2123
rect -258 -2191 -246 -2157
rect -212 -2191 -200 -2157
rect -258 -2225 -200 -2191
rect -258 -2259 -246 -2225
rect -212 -2259 -200 -2225
rect -258 -2293 -200 -2259
rect -258 -2327 -246 -2293
rect -212 -2327 -200 -2293
rect -258 -2361 -200 -2327
rect -258 -2395 -246 -2361
rect -212 -2395 -200 -2361
rect -258 -2414 -200 -2395
rect 200 2467 258 2486
rect 200 2433 212 2467
rect 246 2433 258 2467
rect 200 2399 258 2433
rect 200 2365 212 2399
rect 246 2365 258 2399
rect 200 2331 258 2365
rect 200 2297 212 2331
rect 246 2297 258 2331
rect 200 2263 258 2297
rect 200 2229 212 2263
rect 246 2229 258 2263
rect 200 2195 258 2229
rect 200 2161 212 2195
rect 246 2161 258 2195
rect 200 2127 258 2161
rect 200 2093 212 2127
rect 246 2093 258 2127
rect 200 2059 258 2093
rect 200 2025 212 2059
rect 246 2025 258 2059
rect 200 1991 258 2025
rect 200 1957 212 1991
rect 246 1957 258 1991
rect 200 1923 258 1957
rect 200 1889 212 1923
rect 246 1889 258 1923
rect 200 1855 258 1889
rect 200 1821 212 1855
rect 246 1821 258 1855
rect 200 1787 258 1821
rect 200 1753 212 1787
rect 246 1753 258 1787
rect 200 1719 258 1753
rect 200 1685 212 1719
rect 246 1685 258 1719
rect 200 1651 258 1685
rect 200 1617 212 1651
rect 246 1617 258 1651
rect 200 1583 258 1617
rect 200 1549 212 1583
rect 246 1549 258 1583
rect 200 1515 258 1549
rect 200 1481 212 1515
rect 246 1481 258 1515
rect 200 1447 258 1481
rect 200 1413 212 1447
rect 246 1413 258 1447
rect 200 1379 258 1413
rect 200 1345 212 1379
rect 246 1345 258 1379
rect 200 1311 258 1345
rect 200 1277 212 1311
rect 246 1277 258 1311
rect 200 1243 258 1277
rect 200 1209 212 1243
rect 246 1209 258 1243
rect 200 1175 258 1209
rect 200 1141 212 1175
rect 246 1141 258 1175
rect 200 1107 258 1141
rect 200 1073 212 1107
rect 246 1073 258 1107
rect 200 1039 258 1073
rect 200 1005 212 1039
rect 246 1005 258 1039
rect 200 971 258 1005
rect 200 937 212 971
rect 246 937 258 971
rect 200 903 258 937
rect 200 869 212 903
rect 246 869 258 903
rect 200 835 258 869
rect 200 801 212 835
rect 246 801 258 835
rect 200 767 258 801
rect 200 733 212 767
rect 246 733 258 767
rect 200 699 258 733
rect 200 665 212 699
rect 246 665 258 699
rect 200 631 258 665
rect 200 597 212 631
rect 246 597 258 631
rect 200 563 258 597
rect 200 529 212 563
rect 246 529 258 563
rect 200 495 258 529
rect 200 461 212 495
rect 246 461 258 495
rect 200 427 258 461
rect 200 393 212 427
rect 246 393 258 427
rect 200 359 258 393
rect 200 325 212 359
rect 246 325 258 359
rect 200 291 258 325
rect 200 257 212 291
rect 246 257 258 291
rect 200 223 258 257
rect 200 189 212 223
rect 246 189 258 223
rect 200 155 258 189
rect 200 121 212 155
rect 246 121 258 155
rect 200 87 258 121
rect 200 53 212 87
rect 246 53 258 87
rect 200 19 258 53
rect 200 -15 212 19
rect 246 -15 258 19
rect 200 -49 258 -15
rect 200 -83 212 -49
rect 246 -83 258 -49
rect 200 -117 258 -83
rect 200 -151 212 -117
rect 246 -151 258 -117
rect 200 -185 258 -151
rect 200 -219 212 -185
rect 246 -219 258 -185
rect 200 -253 258 -219
rect 200 -287 212 -253
rect 246 -287 258 -253
rect 200 -321 258 -287
rect 200 -355 212 -321
rect 246 -355 258 -321
rect 200 -389 258 -355
rect 200 -423 212 -389
rect 246 -423 258 -389
rect 200 -457 258 -423
rect 200 -491 212 -457
rect 246 -491 258 -457
rect 200 -525 258 -491
rect 200 -559 212 -525
rect 246 -559 258 -525
rect 200 -593 258 -559
rect 200 -627 212 -593
rect 246 -627 258 -593
rect 200 -661 258 -627
rect 200 -695 212 -661
rect 246 -695 258 -661
rect 200 -729 258 -695
rect 200 -763 212 -729
rect 246 -763 258 -729
rect 200 -797 258 -763
rect 200 -831 212 -797
rect 246 -831 258 -797
rect 200 -865 258 -831
rect 200 -899 212 -865
rect 246 -899 258 -865
rect 200 -933 258 -899
rect 200 -967 212 -933
rect 246 -967 258 -933
rect 200 -1001 258 -967
rect 200 -1035 212 -1001
rect 246 -1035 258 -1001
rect 200 -1069 258 -1035
rect 200 -1103 212 -1069
rect 246 -1103 258 -1069
rect 200 -1137 258 -1103
rect 200 -1171 212 -1137
rect 246 -1171 258 -1137
rect 200 -1205 258 -1171
rect 200 -1239 212 -1205
rect 246 -1239 258 -1205
rect 200 -1273 258 -1239
rect 200 -1307 212 -1273
rect 246 -1307 258 -1273
rect 200 -1341 258 -1307
rect 200 -1375 212 -1341
rect 246 -1375 258 -1341
rect 200 -1409 258 -1375
rect 200 -1443 212 -1409
rect 246 -1443 258 -1409
rect 200 -1477 258 -1443
rect 200 -1511 212 -1477
rect 246 -1511 258 -1477
rect 200 -1545 258 -1511
rect 200 -1579 212 -1545
rect 246 -1579 258 -1545
rect 200 -1613 258 -1579
rect 200 -1647 212 -1613
rect 246 -1647 258 -1613
rect 200 -1681 258 -1647
rect 200 -1715 212 -1681
rect 246 -1715 258 -1681
rect 200 -1749 258 -1715
rect 200 -1783 212 -1749
rect 246 -1783 258 -1749
rect 200 -1817 258 -1783
rect 200 -1851 212 -1817
rect 246 -1851 258 -1817
rect 200 -1885 258 -1851
rect 200 -1919 212 -1885
rect 246 -1919 258 -1885
rect 200 -1953 258 -1919
rect 200 -1987 212 -1953
rect 246 -1987 258 -1953
rect 200 -2021 258 -1987
rect 200 -2055 212 -2021
rect 246 -2055 258 -2021
rect 200 -2089 258 -2055
rect 200 -2123 212 -2089
rect 246 -2123 258 -2089
rect 200 -2157 258 -2123
rect 200 -2191 212 -2157
rect 246 -2191 258 -2157
rect 200 -2225 258 -2191
rect 200 -2259 212 -2225
rect 246 -2259 258 -2225
rect 200 -2293 258 -2259
rect 200 -2327 212 -2293
rect 246 -2327 258 -2293
rect 200 -2361 258 -2327
rect 200 -2395 212 -2361
rect 246 -2395 258 -2361
rect 200 -2414 258 -2395
<< pdiffc >>
rect -246 2433 -212 2467
rect -246 2365 -212 2399
rect -246 2297 -212 2331
rect -246 2229 -212 2263
rect -246 2161 -212 2195
rect -246 2093 -212 2127
rect -246 2025 -212 2059
rect -246 1957 -212 1991
rect -246 1889 -212 1923
rect -246 1821 -212 1855
rect -246 1753 -212 1787
rect -246 1685 -212 1719
rect -246 1617 -212 1651
rect -246 1549 -212 1583
rect -246 1481 -212 1515
rect -246 1413 -212 1447
rect -246 1345 -212 1379
rect -246 1277 -212 1311
rect -246 1209 -212 1243
rect -246 1141 -212 1175
rect -246 1073 -212 1107
rect -246 1005 -212 1039
rect -246 937 -212 971
rect -246 869 -212 903
rect -246 801 -212 835
rect -246 733 -212 767
rect -246 665 -212 699
rect -246 597 -212 631
rect -246 529 -212 563
rect -246 461 -212 495
rect -246 393 -212 427
rect -246 325 -212 359
rect -246 257 -212 291
rect -246 189 -212 223
rect -246 121 -212 155
rect -246 53 -212 87
rect -246 -15 -212 19
rect -246 -83 -212 -49
rect -246 -151 -212 -117
rect -246 -219 -212 -185
rect -246 -287 -212 -253
rect -246 -355 -212 -321
rect -246 -423 -212 -389
rect -246 -491 -212 -457
rect -246 -559 -212 -525
rect -246 -627 -212 -593
rect -246 -695 -212 -661
rect -246 -763 -212 -729
rect -246 -831 -212 -797
rect -246 -899 -212 -865
rect -246 -967 -212 -933
rect -246 -1035 -212 -1001
rect -246 -1103 -212 -1069
rect -246 -1171 -212 -1137
rect -246 -1239 -212 -1205
rect -246 -1307 -212 -1273
rect -246 -1375 -212 -1341
rect -246 -1443 -212 -1409
rect -246 -1511 -212 -1477
rect -246 -1579 -212 -1545
rect -246 -1647 -212 -1613
rect -246 -1715 -212 -1681
rect -246 -1783 -212 -1749
rect -246 -1851 -212 -1817
rect -246 -1919 -212 -1885
rect -246 -1987 -212 -1953
rect -246 -2055 -212 -2021
rect -246 -2123 -212 -2089
rect -246 -2191 -212 -2157
rect -246 -2259 -212 -2225
rect -246 -2327 -212 -2293
rect -246 -2395 -212 -2361
rect 212 2433 246 2467
rect 212 2365 246 2399
rect 212 2297 246 2331
rect 212 2229 246 2263
rect 212 2161 246 2195
rect 212 2093 246 2127
rect 212 2025 246 2059
rect 212 1957 246 1991
rect 212 1889 246 1923
rect 212 1821 246 1855
rect 212 1753 246 1787
rect 212 1685 246 1719
rect 212 1617 246 1651
rect 212 1549 246 1583
rect 212 1481 246 1515
rect 212 1413 246 1447
rect 212 1345 246 1379
rect 212 1277 246 1311
rect 212 1209 246 1243
rect 212 1141 246 1175
rect 212 1073 246 1107
rect 212 1005 246 1039
rect 212 937 246 971
rect 212 869 246 903
rect 212 801 246 835
rect 212 733 246 767
rect 212 665 246 699
rect 212 597 246 631
rect 212 529 246 563
rect 212 461 246 495
rect 212 393 246 427
rect 212 325 246 359
rect 212 257 246 291
rect 212 189 246 223
rect 212 121 246 155
rect 212 53 246 87
rect 212 -15 246 19
rect 212 -83 246 -49
rect 212 -151 246 -117
rect 212 -219 246 -185
rect 212 -287 246 -253
rect 212 -355 246 -321
rect 212 -423 246 -389
rect 212 -491 246 -457
rect 212 -559 246 -525
rect 212 -627 246 -593
rect 212 -695 246 -661
rect 212 -763 246 -729
rect 212 -831 246 -797
rect 212 -899 246 -865
rect 212 -967 246 -933
rect 212 -1035 246 -1001
rect 212 -1103 246 -1069
rect 212 -1171 246 -1137
rect 212 -1239 246 -1205
rect 212 -1307 246 -1273
rect 212 -1375 246 -1341
rect 212 -1443 246 -1409
rect 212 -1511 246 -1477
rect 212 -1579 246 -1545
rect 212 -1647 246 -1613
rect 212 -1715 246 -1681
rect 212 -1783 246 -1749
rect 212 -1851 246 -1817
rect 212 -1919 246 -1885
rect 212 -1987 246 -1953
rect 212 -2055 246 -2021
rect 212 -2123 246 -2089
rect 212 -2191 246 -2157
rect 212 -2259 246 -2225
rect 212 -2327 246 -2293
rect 212 -2395 246 -2361
<< poly >>
rect -200 2486 200 2512
rect -200 -2461 200 -2414
rect -200 -2495 -153 -2461
rect -119 -2495 -85 -2461
rect -51 -2495 -17 -2461
rect 17 -2495 51 -2461
rect 85 -2495 119 -2461
rect 153 -2495 200 -2461
rect -200 -2511 200 -2495
<< polycont >>
rect -153 -2495 -119 -2461
rect -85 -2495 -51 -2461
rect -17 -2495 17 -2461
rect 51 -2495 85 -2461
rect 119 -2495 153 -2461
<< locali >>
rect -246 2467 -212 2490
rect -246 2399 -212 2431
rect -246 2331 -212 2359
rect -246 2263 -212 2287
rect -246 2195 -212 2215
rect -246 2127 -212 2143
rect -246 2059 -212 2071
rect -246 1991 -212 1999
rect -246 1923 -212 1927
rect -246 1817 -212 1821
rect -246 1745 -212 1753
rect -246 1673 -212 1685
rect -246 1601 -212 1617
rect -246 1529 -212 1549
rect -246 1457 -212 1481
rect -246 1385 -212 1413
rect -246 1313 -212 1345
rect -246 1243 -212 1277
rect -246 1175 -212 1207
rect -246 1107 -212 1135
rect -246 1039 -212 1063
rect -246 971 -212 991
rect -246 903 -212 919
rect -246 835 -212 847
rect -246 767 -212 775
rect -246 699 -212 703
rect -246 593 -212 597
rect -246 521 -212 529
rect -246 449 -212 461
rect -246 377 -212 393
rect -246 305 -212 325
rect -246 233 -212 257
rect -246 161 -212 189
rect -246 89 -212 121
rect -246 19 -212 53
rect -246 -49 -212 -17
rect -246 -117 -212 -89
rect -246 -185 -212 -161
rect -246 -253 -212 -233
rect -246 -321 -212 -305
rect -246 -389 -212 -377
rect -246 -457 -212 -449
rect -246 -525 -212 -521
rect -246 -631 -212 -627
rect -246 -703 -212 -695
rect -246 -775 -212 -763
rect -246 -847 -212 -831
rect -246 -919 -212 -899
rect -246 -991 -212 -967
rect -246 -1063 -212 -1035
rect -246 -1135 -212 -1103
rect -246 -1205 -212 -1171
rect -246 -1273 -212 -1241
rect -246 -1341 -212 -1313
rect -246 -1409 -212 -1385
rect -246 -1477 -212 -1457
rect -246 -1545 -212 -1529
rect -246 -1613 -212 -1601
rect -246 -1681 -212 -1673
rect -246 -1749 -212 -1745
rect -246 -1855 -212 -1851
rect -246 -1927 -212 -1919
rect -246 -1999 -212 -1987
rect -246 -2071 -212 -2055
rect -246 -2143 -212 -2123
rect -246 -2215 -212 -2191
rect -246 -2287 -212 -2259
rect -246 -2359 -212 -2327
rect -246 -2418 -212 -2395
rect 212 2467 246 2490
rect 212 2399 246 2431
rect 212 2331 246 2359
rect 212 2263 246 2287
rect 212 2195 246 2215
rect 212 2127 246 2143
rect 212 2059 246 2071
rect 212 1991 246 1999
rect 212 1923 246 1927
rect 212 1817 246 1821
rect 212 1745 246 1753
rect 212 1673 246 1685
rect 212 1601 246 1617
rect 212 1529 246 1549
rect 212 1457 246 1481
rect 212 1385 246 1413
rect 212 1313 246 1345
rect 212 1243 246 1277
rect 212 1175 246 1207
rect 212 1107 246 1135
rect 212 1039 246 1063
rect 212 971 246 991
rect 212 903 246 919
rect 212 835 246 847
rect 212 767 246 775
rect 212 699 246 703
rect 212 593 246 597
rect 212 521 246 529
rect 212 449 246 461
rect 212 377 246 393
rect 212 305 246 325
rect 212 233 246 257
rect 212 161 246 189
rect 212 89 246 121
rect 212 19 246 53
rect 212 -49 246 -17
rect 212 -117 246 -89
rect 212 -185 246 -161
rect 212 -253 246 -233
rect 212 -321 246 -305
rect 212 -389 246 -377
rect 212 -457 246 -449
rect 212 -525 246 -521
rect 212 -631 246 -627
rect 212 -703 246 -695
rect 212 -775 246 -763
rect 212 -847 246 -831
rect 212 -919 246 -899
rect 212 -991 246 -967
rect 212 -1063 246 -1035
rect 212 -1135 246 -1103
rect 212 -1205 246 -1171
rect 212 -1273 246 -1241
rect 212 -1341 246 -1313
rect 212 -1409 246 -1385
rect 212 -1477 246 -1457
rect 212 -1545 246 -1529
rect 212 -1613 246 -1601
rect 212 -1681 246 -1673
rect 212 -1749 246 -1745
rect 212 -1855 246 -1851
rect 212 -1927 246 -1919
rect 212 -1999 246 -1987
rect 212 -2071 246 -2055
rect 212 -2143 246 -2123
rect 212 -2215 246 -2191
rect 212 -2287 246 -2259
rect 212 -2359 246 -2327
rect 212 -2418 246 -2395
rect -200 -2495 -161 -2461
rect -119 -2495 -89 -2461
rect -51 -2495 -17 -2461
rect 17 -2495 51 -2461
rect 89 -2495 119 -2461
rect 161 -2495 200 -2461
<< viali >>
rect -246 2433 -212 2465
rect -246 2431 -212 2433
rect -246 2365 -212 2393
rect -246 2359 -212 2365
rect -246 2297 -212 2321
rect -246 2287 -212 2297
rect -246 2229 -212 2249
rect -246 2215 -212 2229
rect -246 2161 -212 2177
rect -246 2143 -212 2161
rect -246 2093 -212 2105
rect -246 2071 -212 2093
rect -246 2025 -212 2033
rect -246 1999 -212 2025
rect -246 1957 -212 1961
rect -246 1927 -212 1957
rect -246 1855 -212 1889
rect -246 1787 -212 1817
rect -246 1783 -212 1787
rect -246 1719 -212 1745
rect -246 1711 -212 1719
rect -246 1651 -212 1673
rect -246 1639 -212 1651
rect -246 1583 -212 1601
rect -246 1567 -212 1583
rect -246 1515 -212 1529
rect -246 1495 -212 1515
rect -246 1447 -212 1457
rect -246 1423 -212 1447
rect -246 1379 -212 1385
rect -246 1351 -212 1379
rect -246 1311 -212 1313
rect -246 1279 -212 1311
rect -246 1209 -212 1241
rect -246 1207 -212 1209
rect -246 1141 -212 1169
rect -246 1135 -212 1141
rect -246 1073 -212 1097
rect -246 1063 -212 1073
rect -246 1005 -212 1025
rect -246 991 -212 1005
rect -246 937 -212 953
rect -246 919 -212 937
rect -246 869 -212 881
rect -246 847 -212 869
rect -246 801 -212 809
rect -246 775 -212 801
rect -246 733 -212 737
rect -246 703 -212 733
rect -246 631 -212 665
rect -246 563 -212 593
rect -246 559 -212 563
rect -246 495 -212 521
rect -246 487 -212 495
rect -246 427 -212 449
rect -246 415 -212 427
rect -246 359 -212 377
rect -246 343 -212 359
rect -246 291 -212 305
rect -246 271 -212 291
rect -246 223 -212 233
rect -246 199 -212 223
rect -246 155 -212 161
rect -246 127 -212 155
rect -246 87 -212 89
rect -246 55 -212 87
rect -246 -15 -212 17
rect -246 -17 -212 -15
rect -246 -83 -212 -55
rect -246 -89 -212 -83
rect -246 -151 -212 -127
rect -246 -161 -212 -151
rect -246 -219 -212 -199
rect -246 -233 -212 -219
rect -246 -287 -212 -271
rect -246 -305 -212 -287
rect -246 -355 -212 -343
rect -246 -377 -212 -355
rect -246 -423 -212 -415
rect -246 -449 -212 -423
rect -246 -491 -212 -487
rect -246 -521 -212 -491
rect -246 -593 -212 -559
rect -246 -661 -212 -631
rect -246 -665 -212 -661
rect -246 -729 -212 -703
rect -246 -737 -212 -729
rect -246 -797 -212 -775
rect -246 -809 -212 -797
rect -246 -865 -212 -847
rect -246 -881 -212 -865
rect -246 -933 -212 -919
rect -246 -953 -212 -933
rect -246 -1001 -212 -991
rect -246 -1025 -212 -1001
rect -246 -1069 -212 -1063
rect -246 -1097 -212 -1069
rect -246 -1137 -212 -1135
rect -246 -1169 -212 -1137
rect -246 -1239 -212 -1207
rect -246 -1241 -212 -1239
rect -246 -1307 -212 -1279
rect -246 -1313 -212 -1307
rect -246 -1375 -212 -1351
rect -246 -1385 -212 -1375
rect -246 -1443 -212 -1423
rect -246 -1457 -212 -1443
rect -246 -1511 -212 -1495
rect -246 -1529 -212 -1511
rect -246 -1579 -212 -1567
rect -246 -1601 -212 -1579
rect -246 -1647 -212 -1639
rect -246 -1673 -212 -1647
rect -246 -1715 -212 -1711
rect -246 -1745 -212 -1715
rect -246 -1817 -212 -1783
rect -246 -1885 -212 -1855
rect -246 -1889 -212 -1885
rect -246 -1953 -212 -1927
rect -246 -1961 -212 -1953
rect -246 -2021 -212 -1999
rect -246 -2033 -212 -2021
rect -246 -2089 -212 -2071
rect -246 -2105 -212 -2089
rect -246 -2157 -212 -2143
rect -246 -2177 -212 -2157
rect -246 -2225 -212 -2215
rect -246 -2249 -212 -2225
rect -246 -2293 -212 -2287
rect -246 -2321 -212 -2293
rect -246 -2361 -212 -2359
rect -246 -2393 -212 -2361
rect 212 2433 246 2465
rect 212 2431 246 2433
rect 212 2365 246 2393
rect 212 2359 246 2365
rect 212 2297 246 2321
rect 212 2287 246 2297
rect 212 2229 246 2249
rect 212 2215 246 2229
rect 212 2161 246 2177
rect 212 2143 246 2161
rect 212 2093 246 2105
rect 212 2071 246 2093
rect 212 2025 246 2033
rect 212 1999 246 2025
rect 212 1957 246 1961
rect 212 1927 246 1957
rect 212 1855 246 1889
rect 212 1787 246 1817
rect 212 1783 246 1787
rect 212 1719 246 1745
rect 212 1711 246 1719
rect 212 1651 246 1673
rect 212 1639 246 1651
rect 212 1583 246 1601
rect 212 1567 246 1583
rect 212 1515 246 1529
rect 212 1495 246 1515
rect 212 1447 246 1457
rect 212 1423 246 1447
rect 212 1379 246 1385
rect 212 1351 246 1379
rect 212 1311 246 1313
rect 212 1279 246 1311
rect 212 1209 246 1241
rect 212 1207 246 1209
rect 212 1141 246 1169
rect 212 1135 246 1141
rect 212 1073 246 1097
rect 212 1063 246 1073
rect 212 1005 246 1025
rect 212 991 246 1005
rect 212 937 246 953
rect 212 919 246 937
rect 212 869 246 881
rect 212 847 246 869
rect 212 801 246 809
rect 212 775 246 801
rect 212 733 246 737
rect 212 703 246 733
rect 212 631 246 665
rect 212 563 246 593
rect 212 559 246 563
rect 212 495 246 521
rect 212 487 246 495
rect 212 427 246 449
rect 212 415 246 427
rect 212 359 246 377
rect 212 343 246 359
rect 212 291 246 305
rect 212 271 246 291
rect 212 223 246 233
rect 212 199 246 223
rect 212 155 246 161
rect 212 127 246 155
rect 212 87 246 89
rect 212 55 246 87
rect 212 -15 246 17
rect 212 -17 246 -15
rect 212 -83 246 -55
rect 212 -89 246 -83
rect 212 -151 246 -127
rect 212 -161 246 -151
rect 212 -219 246 -199
rect 212 -233 246 -219
rect 212 -287 246 -271
rect 212 -305 246 -287
rect 212 -355 246 -343
rect 212 -377 246 -355
rect 212 -423 246 -415
rect 212 -449 246 -423
rect 212 -491 246 -487
rect 212 -521 246 -491
rect 212 -593 246 -559
rect 212 -661 246 -631
rect 212 -665 246 -661
rect 212 -729 246 -703
rect 212 -737 246 -729
rect 212 -797 246 -775
rect 212 -809 246 -797
rect 212 -865 246 -847
rect 212 -881 246 -865
rect 212 -933 246 -919
rect 212 -953 246 -933
rect 212 -1001 246 -991
rect 212 -1025 246 -1001
rect 212 -1069 246 -1063
rect 212 -1097 246 -1069
rect 212 -1137 246 -1135
rect 212 -1169 246 -1137
rect 212 -1239 246 -1207
rect 212 -1241 246 -1239
rect 212 -1307 246 -1279
rect 212 -1313 246 -1307
rect 212 -1375 246 -1351
rect 212 -1385 246 -1375
rect 212 -1443 246 -1423
rect 212 -1457 246 -1443
rect 212 -1511 246 -1495
rect 212 -1529 246 -1511
rect 212 -1579 246 -1567
rect 212 -1601 246 -1579
rect 212 -1647 246 -1639
rect 212 -1673 246 -1647
rect 212 -1715 246 -1711
rect 212 -1745 246 -1715
rect 212 -1817 246 -1783
rect 212 -1885 246 -1855
rect 212 -1889 246 -1885
rect 212 -1953 246 -1927
rect 212 -1961 246 -1953
rect 212 -2021 246 -1999
rect 212 -2033 246 -2021
rect 212 -2089 246 -2071
rect 212 -2105 246 -2089
rect 212 -2157 246 -2143
rect 212 -2177 246 -2157
rect 212 -2225 246 -2215
rect 212 -2249 246 -2225
rect 212 -2293 246 -2287
rect 212 -2321 246 -2293
rect 212 -2361 246 -2359
rect 212 -2393 246 -2361
rect -161 -2495 -153 -2461
rect -153 -2495 -127 -2461
rect -89 -2495 -85 -2461
rect -85 -2495 -55 -2461
rect -17 -2495 17 -2461
rect 55 -2495 85 -2461
rect 85 -2495 89 -2461
rect 127 -2495 153 -2461
rect 153 -2495 161 -2461
<< metal1 >>
rect -252 2465 -206 2486
rect -252 2431 -246 2465
rect -212 2431 -206 2465
rect -252 2393 -206 2431
rect -252 2359 -246 2393
rect -212 2359 -206 2393
rect -252 2321 -206 2359
rect -252 2287 -246 2321
rect -212 2287 -206 2321
rect -252 2249 -206 2287
rect -252 2215 -246 2249
rect -212 2215 -206 2249
rect -252 2177 -206 2215
rect -252 2143 -246 2177
rect -212 2143 -206 2177
rect -252 2105 -206 2143
rect -252 2071 -246 2105
rect -212 2071 -206 2105
rect -252 2033 -206 2071
rect -252 1999 -246 2033
rect -212 1999 -206 2033
rect -252 1961 -206 1999
rect -252 1927 -246 1961
rect -212 1927 -206 1961
rect -252 1889 -206 1927
rect -252 1855 -246 1889
rect -212 1855 -206 1889
rect -252 1817 -206 1855
rect -252 1783 -246 1817
rect -212 1783 -206 1817
rect -252 1745 -206 1783
rect -252 1711 -246 1745
rect -212 1711 -206 1745
rect -252 1673 -206 1711
rect -252 1639 -246 1673
rect -212 1639 -206 1673
rect -252 1601 -206 1639
rect -252 1567 -246 1601
rect -212 1567 -206 1601
rect -252 1529 -206 1567
rect -252 1495 -246 1529
rect -212 1495 -206 1529
rect -252 1457 -206 1495
rect -252 1423 -246 1457
rect -212 1423 -206 1457
rect -252 1385 -206 1423
rect -252 1351 -246 1385
rect -212 1351 -206 1385
rect -252 1313 -206 1351
rect -252 1279 -246 1313
rect -212 1279 -206 1313
rect -252 1241 -206 1279
rect -252 1207 -246 1241
rect -212 1207 -206 1241
rect -252 1169 -206 1207
rect -252 1135 -246 1169
rect -212 1135 -206 1169
rect -252 1097 -206 1135
rect -252 1063 -246 1097
rect -212 1063 -206 1097
rect -252 1025 -206 1063
rect -252 991 -246 1025
rect -212 991 -206 1025
rect -252 953 -206 991
rect -252 919 -246 953
rect -212 919 -206 953
rect -252 881 -206 919
rect -252 847 -246 881
rect -212 847 -206 881
rect -252 809 -206 847
rect -252 775 -246 809
rect -212 775 -206 809
rect -252 737 -206 775
rect -252 703 -246 737
rect -212 703 -206 737
rect -252 665 -206 703
rect -252 631 -246 665
rect -212 631 -206 665
rect -252 593 -206 631
rect -252 559 -246 593
rect -212 559 -206 593
rect -252 521 -206 559
rect -252 487 -246 521
rect -212 487 -206 521
rect -252 449 -206 487
rect -252 415 -246 449
rect -212 415 -206 449
rect -252 377 -206 415
rect -252 343 -246 377
rect -212 343 -206 377
rect -252 305 -206 343
rect -252 271 -246 305
rect -212 271 -206 305
rect -252 233 -206 271
rect -252 199 -246 233
rect -212 199 -206 233
rect -252 161 -206 199
rect -252 127 -246 161
rect -212 127 -206 161
rect -252 89 -206 127
rect -252 55 -246 89
rect -212 55 -206 89
rect -252 17 -206 55
rect -252 -17 -246 17
rect -212 -17 -206 17
rect -252 -55 -206 -17
rect -252 -89 -246 -55
rect -212 -89 -206 -55
rect -252 -127 -206 -89
rect -252 -161 -246 -127
rect -212 -161 -206 -127
rect -252 -199 -206 -161
rect -252 -233 -246 -199
rect -212 -233 -206 -199
rect -252 -271 -206 -233
rect -252 -305 -246 -271
rect -212 -305 -206 -271
rect -252 -343 -206 -305
rect -252 -377 -246 -343
rect -212 -377 -206 -343
rect -252 -415 -206 -377
rect -252 -449 -246 -415
rect -212 -449 -206 -415
rect -252 -487 -206 -449
rect -252 -521 -246 -487
rect -212 -521 -206 -487
rect -252 -559 -206 -521
rect -252 -593 -246 -559
rect -212 -593 -206 -559
rect -252 -631 -206 -593
rect -252 -665 -246 -631
rect -212 -665 -206 -631
rect -252 -703 -206 -665
rect -252 -737 -246 -703
rect -212 -737 -206 -703
rect -252 -775 -206 -737
rect -252 -809 -246 -775
rect -212 -809 -206 -775
rect -252 -847 -206 -809
rect -252 -881 -246 -847
rect -212 -881 -206 -847
rect -252 -919 -206 -881
rect -252 -953 -246 -919
rect -212 -953 -206 -919
rect -252 -991 -206 -953
rect -252 -1025 -246 -991
rect -212 -1025 -206 -991
rect -252 -1063 -206 -1025
rect -252 -1097 -246 -1063
rect -212 -1097 -206 -1063
rect -252 -1135 -206 -1097
rect -252 -1169 -246 -1135
rect -212 -1169 -206 -1135
rect -252 -1207 -206 -1169
rect -252 -1241 -246 -1207
rect -212 -1241 -206 -1207
rect -252 -1279 -206 -1241
rect -252 -1313 -246 -1279
rect -212 -1313 -206 -1279
rect -252 -1351 -206 -1313
rect -252 -1385 -246 -1351
rect -212 -1385 -206 -1351
rect -252 -1423 -206 -1385
rect -252 -1457 -246 -1423
rect -212 -1457 -206 -1423
rect -252 -1495 -206 -1457
rect -252 -1529 -246 -1495
rect -212 -1529 -206 -1495
rect -252 -1567 -206 -1529
rect -252 -1601 -246 -1567
rect -212 -1601 -206 -1567
rect -252 -1639 -206 -1601
rect -252 -1673 -246 -1639
rect -212 -1673 -206 -1639
rect -252 -1711 -206 -1673
rect -252 -1745 -246 -1711
rect -212 -1745 -206 -1711
rect -252 -1783 -206 -1745
rect -252 -1817 -246 -1783
rect -212 -1817 -206 -1783
rect -252 -1855 -206 -1817
rect -252 -1889 -246 -1855
rect -212 -1889 -206 -1855
rect -252 -1927 -206 -1889
rect -252 -1961 -246 -1927
rect -212 -1961 -206 -1927
rect -252 -1999 -206 -1961
rect -252 -2033 -246 -1999
rect -212 -2033 -206 -1999
rect -252 -2071 -206 -2033
rect -252 -2105 -246 -2071
rect -212 -2105 -206 -2071
rect -252 -2143 -206 -2105
rect -252 -2177 -246 -2143
rect -212 -2177 -206 -2143
rect -252 -2215 -206 -2177
rect -252 -2249 -246 -2215
rect -212 -2249 -206 -2215
rect -252 -2287 -206 -2249
rect -252 -2321 -246 -2287
rect -212 -2321 -206 -2287
rect -252 -2359 -206 -2321
rect -252 -2393 -246 -2359
rect -212 -2393 -206 -2359
rect -252 -2414 -206 -2393
rect 206 2465 252 2486
rect 206 2431 212 2465
rect 246 2431 252 2465
rect 206 2393 252 2431
rect 206 2359 212 2393
rect 246 2359 252 2393
rect 206 2321 252 2359
rect 206 2287 212 2321
rect 246 2287 252 2321
rect 206 2249 252 2287
rect 206 2215 212 2249
rect 246 2215 252 2249
rect 206 2177 252 2215
rect 206 2143 212 2177
rect 246 2143 252 2177
rect 206 2105 252 2143
rect 206 2071 212 2105
rect 246 2071 252 2105
rect 206 2033 252 2071
rect 206 1999 212 2033
rect 246 1999 252 2033
rect 206 1961 252 1999
rect 206 1927 212 1961
rect 246 1927 252 1961
rect 206 1889 252 1927
rect 206 1855 212 1889
rect 246 1855 252 1889
rect 206 1817 252 1855
rect 206 1783 212 1817
rect 246 1783 252 1817
rect 206 1745 252 1783
rect 206 1711 212 1745
rect 246 1711 252 1745
rect 206 1673 252 1711
rect 206 1639 212 1673
rect 246 1639 252 1673
rect 206 1601 252 1639
rect 206 1567 212 1601
rect 246 1567 252 1601
rect 206 1529 252 1567
rect 206 1495 212 1529
rect 246 1495 252 1529
rect 206 1457 252 1495
rect 206 1423 212 1457
rect 246 1423 252 1457
rect 206 1385 252 1423
rect 206 1351 212 1385
rect 246 1351 252 1385
rect 206 1313 252 1351
rect 206 1279 212 1313
rect 246 1279 252 1313
rect 206 1241 252 1279
rect 206 1207 212 1241
rect 246 1207 252 1241
rect 206 1169 252 1207
rect 206 1135 212 1169
rect 246 1135 252 1169
rect 206 1097 252 1135
rect 206 1063 212 1097
rect 246 1063 252 1097
rect 206 1025 252 1063
rect 206 991 212 1025
rect 246 991 252 1025
rect 206 953 252 991
rect 206 919 212 953
rect 246 919 252 953
rect 206 881 252 919
rect 206 847 212 881
rect 246 847 252 881
rect 206 809 252 847
rect 206 775 212 809
rect 246 775 252 809
rect 206 737 252 775
rect 206 703 212 737
rect 246 703 252 737
rect 206 665 252 703
rect 206 631 212 665
rect 246 631 252 665
rect 206 593 252 631
rect 206 559 212 593
rect 246 559 252 593
rect 206 521 252 559
rect 206 487 212 521
rect 246 487 252 521
rect 206 449 252 487
rect 206 415 212 449
rect 246 415 252 449
rect 206 377 252 415
rect 206 343 212 377
rect 246 343 252 377
rect 206 305 252 343
rect 206 271 212 305
rect 246 271 252 305
rect 206 233 252 271
rect 206 199 212 233
rect 246 199 252 233
rect 206 161 252 199
rect 206 127 212 161
rect 246 127 252 161
rect 206 89 252 127
rect 206 55 212 89
rect 246 55 252 89
rect 206 17 252 55
rect 206 -17 212 17
rect 246 -17 252 17
rect 206 -55 252 -17
rect 206 -89 212 -55
rect 246 -89 252 -55
rect 206 -127 252 -89
rect 206 -161 212 -127
rect 246 -161 252 -127
rect 206 -199 252 -161
rect 206 -233 212 -199
rect 246 -233 252 -199
rect 206 -271 252 -233
rect 206 -305 212 -271
rect 246 -305 252 -271
rect 206 -343 252 -305
rect 206 -377 212 -343
rect 246 -377 252 -343
rect 206 -415 252 -377
rect 206 -449 212 -415
rect 246 -449 252 -415
rect 206 -487 252 -449
rect 206 -521 212 -487
rect 246 -521 252 -487
rect 206 -559 252 -521
rect 206 -593 212 -559
rect 246 -593 252 -559
rect 206 -631 252 -593
rect 206 -665 212 -631
rect 246 -665 252 -631
rect 206 -703 252 -665
rect 206 -737 212 -703
rect 246 -737 252 -703
rect 206 -775 252 -737
rect 206 -809 212 -775
rect 246 -809 252 -775
rect 206 -847 252 -809
rect 206 -881 212 -847
rect 246 -881 252 -847
rect 206 -919 252 -881
rect 206 -953 212 -919
rect 246 -953 252 -919
rect 206 -991 252 -953
rect 206 -1025 212 -991
rect 246 -1025 252 -991
rect 206 -1063 252 -1025
rect 206 -1097 212 -1063
rect 246 -1097 252 -1063
rect 206 -1135 252 -1097
rect 206 -1169 212 -1135
rect 246 -1169 252 -1135
rect 206 -1207 252 -1169
rect 206 -1241 212 -1207
rect 246 -1241 252 -1207
rect 206 -1279 252 -1241
rect 206 -1313 212 -1279
rect 246 -1313 252 -1279
rect 206 -1351 252 -1313
rect 206 -1385 212 -1351
rect 246 -1385 252 -1351
rect 206 -1423 252 -1385
rect 206 -1457 212 -1423
rect 246 -1457 252 -1423
rect 206 -1495 252 -1457
rect 206 -1529 212 -1495
rect 246 -1529 252 -1495
rect 206 -1567 252 -1529
rect 206 -1601 212 -1567
rect 246 -1601 252 -1567
rect 206 -1639 252 -1601
rect 206 -1673 212 -1639
rect 246 -1673 252 -1639
rect 206 -1711 252 -1673
rect 206 -1745 212 -1711
rect 246 -1745 252 -1711
rect 206 -1783 252 -1745
rect 206 -1817 212 -1783
rect 246 -1817 252 -1783
rect 206 -1855 252 -1817
rect 206 -1889 212 -1855
rect 246 -1889 252 -1855
rect 206 -1927 252 -1889
rect 206 -1961 212 -1927
rect 246 -1961 252 -1927
rect 206 -1999 252 -1961
rect 206 -2033 212 -1999
rect 246 -2033 252 -1999
rect 206 -2071 252 -2033
rect 206 -2105 212 -2071
rect 246 -2105 252 -2071
rect 206 -2143 252 -2105
rect 206 -2177 212 -2143
rect 246 -2177 252 -2143
rect 206 -2215 252 -2177
rect 206 -2249 212 -2215
rect 246 -2249 252 -2215
rect 206 -2287 252 -2249
rect 206 -2321 212 -2287
rect 246 -2321 252 -2287
rect 206 -2359 252 -2321
rect 206 -2393 212 -2359
rect 246 -2393 252 -2359
rect 206 -2414 252 -2393
rect -196 -2461 196 -2455
rect -196 -2495 -161 -2461
rect -127 -2495 -89 -2461
rect -55 -2495 -17 -2461
rect 17 -2495 55 -2461
rect 89 -2495 127 -2461
rect 161 -2495 196 -2461
rect -196 -2501 196 -2495
<< end >>
