magic
tech sky130A
magscale 1 2
timestamp 1664683715
<< error_p >>
rect -29 -71 29 -65
rect -29 -105 -17 -71
rect -29 -111 29 -105
<< nwell >>
rect -124 -124 124 158
<< pmos >>
rect -30 -24 30 96
<< pdiff >>
rect -88 84 -30 96
rect -88 -12 -76 84
rect -42 -12 -30 84
rect -88 -24 -30 -12
rect 30 84 88 96
rect 30 -12 42 84
rect 76 -12 88 84
rect 30 -24 88 -12
<< pdiffc >>
rect -76 -12 -42 84
rect 42 -12 76 84
<< poly >>
rect -30 96 30 122
rect -30 -55 30 -24
rect -33 -71 33 -55
rect -33 -105 -17 -71
rect 17 -105 33 -71
rect -33 -121 33 -105
<< polycont >>
rect -17 -105 17 -71
<< locali >>
rect -76 84 -42 100
rect -76 -28 -42 -12
rect 42 84 76 100
rect 42 -28 76 -12
rect -33 -105 -17 -71
rect 17 -105 33 -71
<< viali >>
rect -76 -12 -42 84
rect 42 -12 76 84
rect -17 -105 17 -71
<< metal1 >>
rect -82 84 -36 96
rect -82 -12 -76 84
rect -42 -12 -36 84
rect -82 -24 -36 -12
rect 36 84 82 96
rect 36 -12 42 84
rect 76 -12 82 84
rect 36 -24 82 -12
rect -29 -71 29 -65
rect -29 -105 -17 -71
rect 17 -105 29 -71
rect -29 -111 29 -105
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.6 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
