magic
tech sky130A
magscale 1 2
timestamp 1668324311
<< nwell >>
rect -2498 1724 1462 2367
rect -2498 -716 1465 1724
<< psubdiff >>
rect -2704 -3040 -2680 -2614
rect 2114 -3040 2138 -2614
<< nsubdiff >>
rect -2383 2156 1387 2229
rect -2383 2155 -985 2156
rect -2383 2154 -1423 2155
rect -1347 2154 -985 2155
rect -909 2154 1387 2156
rect -2383 1995 -2253 2154
rect 1292 1995 1387 2154
rect -2383 1895 1387 1995
<< psubdiffcont >>
rect -2680 -3040 2114 -2614
<< nsubdiffcont >>
rect -1423 2154 -1347 2155
rect -985 2154 -909 2156
rect -2253 1995 1292 2154
<< poly >>
rect -2634 1870 -2562 1888
rect -2634 1834 -2616 1870
rect -2582 1846 -2562 1870
rect -2582 1834 -982 1846
rect -2634 1816 -982 1834
rect -2628 1772 -2556 1773
rect -2628 1755 -1304 1772
rect -2628 1719 -2610 1755
rect -2576 1742 -1304 1755
rect -2576 1719 -2556 1742
rect -2628 1701 -2556 1719
rect -1348 1640 -1304 1742
rect -1012 1549 -982 1816
rect -733 1742 -653 1746
rect -733 1729 712 1742
rect -733 1693 -713 1729
rect -671 1693 712 1729
rect -733 1685 712 1693
rect -733 1676 -653 1685
rect -250 1615 -170 1628
rect -250 1611 482 1615
rect -250 1608 -230 1611
rect -535 1575 -230 1608
rect -188 1575 482 1611
rect -535 1566 482 1575
rect -535 1506 -475 1566
rect -417 1506 -357 1566
rect -250 1558 -170 1566
rect 422 1436 482 1566
rect 652 1457 712 1685
rect -653 -508 -593 -460
rect -299 -508 -239 -460
rect 40 -508 364 -507
rect -653 -548 364 -508
rect 899 -597 1083 -550
rect -289 -1053 1169 -1023
rect -289 -1147 -250 -1053
rect 499 -1159 557 -1053
rect 1113 -1156 1169 -1053
rect -1358 -1863 -1065 -1807
rect -534 -1874 -472 -1813
rect 115 -1874 175 -1809
rect -534 -1922 175 -1874
rect 116 -1935 175 -1922
rect 883 -1935 926 -1820
rect 116 -1979 926 -1935
<< polycont >>
rect -2616 1834 -2582 1870
rect -2610 1719 -2576 1755
rect -713 1693 -671 1729
rect -230 1575 -188 1611
<< locali >>
rect -2310 2156 1335 2190
rect -2310 2155 -985 2156
rect -2310 2154 -1423 2155
rect -1347 2154 -985 2155
rect -909 2154 1335 2156
rect -2310 1995 -2253 2154
rect 1292 1995 1335 2154
rect -2310 1948 1335 1995
rect -2634 1870 -2562 1888
rect -2634 1834 -2616 1870
rect -2582 1834 -2562 1870
rect -2634 1816 -2562 1834
rect -2628 1755 -2556 1773
rect -2628 1719 -2610 1755
rect -2576 1719 -2556 1755
rect -2628 1701 -2556 1719
rect -733 1729 -653 1746
rect -733 1693 -713 1729
rect -671 1693 -653 1729
rect -733 1676 -653 1693
rect -250 1611 -170 1628
rect -2186 1531 -1944 1585
rect -250 1575 -230 1611
rect -188 1575 -170 1611
rect -250 1558 -170 1575
rect -2002 -818 -1944 1531
rect -1342 -566 -1308 -483
rect 258 -566 292 1419
rect -1342 -600 292 -566
rect 258 -708 292 -600
rect 818 -514 888 44
rect 1092 -513 1163 29
rect 818 -610 864 -514
rect 812 -625 864 -610
rect 812 -626 872 -625
rect 812 -660 824 -626
rect 858 -660 872 -626
rect 812 -668 872 -660
rect 812 -673 864 -668
rect 915 -708 949 -557
rect 1117 -614 1163 -513
rect 1116 -628 1170 -614
rect 1116 -662 1124 -628
rect 1158 -662 1170 -628
rect 1116 -674 1170 -662
rect 258 -742 949 -708
rect -2003 -822 -1944 -818
rect -2003 -867 -1998 -822
rect -1949 -836 -1944 -822
rect -1949 -867 44 -836
rect -2003 -870 44 -867
rect -2003 -872 -1944 -870
rect 9 -988 44 -870
rect 9 -1018 427 -988
rect 10 -1022 427 -1018
rect 10 -1146 44 -1022
rect 393 -1153 427 -1022
rect -1171 -1894 -1137 -1197
rect -935 -1755 -901 -1165
rect -960 -1789 -901 -1755
rect -699 -1750 -665 -1181
rect 794 -1184 836 -742
rect 934 -823 992 -809
rect 934 -857 946 -823
rect 980 -857 992 -823
rect 934 -870 992 -857
rect 1117 -813 1163 -674
rect 1323 -813 1394 -801
rect 1117 -822 1394 -813
rect 1117 -859 1336 -822
rect 1372 -859 1394 -822
rect -699 -1789 -640 -1750
rect -227 -1771 -193 -1195
rect 794 -1467 863 -1184
rect 940 -1329 986 -870
rect 1323 -873 1394 -859
rect 1331 -914 1378 -873
rect 1332 -1130 1378 -914
rect 1332 -1264 1414 -1130
rect -960 -1894 -926 -1789
rect -674 -1894 -640 -1789
rect -1171 -1928 -640 -1894
rect -2696 -3040 -2680 -2614
rect 2114 -3040 2130 -2614
<< viali >>
rect -1712 2065 -1667 2107
rect -1525 2094 -1480 2136
rect -1408 2101 -1363 2143
rect -970 2102 -925 2144
rect -468 2088 -423 2130
rect 123 2089 168 2131
rect 478 2091 523 2133
rect 598 2089 643 2131
rect 959 2089 1004 2131
rect 1224 2086 1269 2128
rect -2616 1834 -2582 1870
rect -2610 1719 -2576 1755
rect -713 1693 -671 1729
rect -230 1575 -188 1611
rect 824 -660 858 -626
rect 1124 -662 1158 -628
rect -1998 -867 -1949 -822
rect -296 -1149 -244 -1097
rect 946 -857 980 -823
rect 1336 -859 1372 -822
rect -2397 -2835 -2352 -2793
rect -1866 -2834 -1821 -2792
rect -2524 -2880 -2479 -2838
rect -1424 -2840 -1379 -2798
rect -1058 -2840 -1013 -2798
rect -239 -2835 -194 -2793
rect 577 -2838 622 -2796
rect 1200 -2831 1245 -2789
rect 1608 -2826 1653 -2784
rect 1877 -2822 1922 -2780
<< metal1 >>
rect -1539 2136 -1465 2145
rect -1726 2107 -1652 2116
rect -1726 2065 -1712 2107
rect -1667 2065 -1652 2107
rect -1539 2094 -1525 2136
rect -1480 2094 -1465 2136
rect -1539 2082 -1465 2094
rect -1422 2143 -1348 2152
rect -1422 2101 -1408 2143
rect -1363 2101 -1348 2143
rect -1422 2089 -1348 2101
rect -984 2144 -910 2153
rect -984 2102 -970 2144
rect -925 2102 -910 2144
rect -984 2090 -910 2102
rect -482 2130 -408 2139
rect -1726 2050 -1652 2065
rect -2634 1879 -2562 1888
rect -2634 1827 -2622 1879
rect -2570 1827 -2562 1879
rect -2634 1816 -2562 1827
rect -2628 1764 -2556 1773
rect -2628 1712 -2616 1764
rect -2564 1712 -2556 1764
rect -2628 1701 -2556 1712
rect -5586 1610 -5458 1618
rect -5586 1580 -5576 1610
rect -5638 1530 -5576 1580
rect -5586 1510 -5576 1530
rect -5464 1580 -5458 1610
rect -3928 1610 -3800 1618
rect -3928 1580 -3918 1610
rect -5464 1530 -3918 1580
rect -5464 1510 -5458 1530
rect -5586 1502 -5458 1510
rect -4711 1276 -4648 1530
rect -3928 1510 -3918 1530
rect -3806 1595 -3800 1610
rect -3806 1580 -3790 1595
rect -2190 1583 -2127 1584
rect -2309 1580 -2242 1581
rect -3806 1528 -2242 1580
rect -3806 1517 -3790 1528
rect -3806 1510 -3800 1517
rect -3928 1502 -3800 1510
rect -3059 1295 -2988 1528
rect -2190 1526 -2126 1583
rect -2189 1525 -2126 1526
rect -1702 1322 -1668 2050
rect -1517 1707 -1483 2082
rect -1530 1700 -1467 1707
rect -1530 1648 -1524 1700
rect -1472 1648 -1467 1700
rect -1530 1640 -1467 1648
rect -1401 1345 -1367 2089
rect -962 1493 -928 2090
rect -482 2088 -468 2130
rect -423 2088 -408 2130
rect -482 2076 -408 2088
rect 109 2131 183 2140
rect 109 2089 123 2131
rect 168 2089 183 2131
rect 109 2077 183 2089
rect 464 2133 538 2142
rect 464 2091 478 2133
rect 523 2091 538 2133
rect 464 2079 538 2091
rect 584 2131 658 2140
rect 584 2089 598 2131
rect 643 2089 658 2131
rect -733 1729 -653 1746
rect -733 1693 -713 1729
rect -671 1693 -653 1729
rect -733 1676 -653 1693
rect -699 1561 -665 1676
rect -888 1527 -665 1561
rect -962 1465 -913 1493
rect -947 1331 -913 1465
rect -4976 478 -4879 781
rect -3318 541 -3212 844
rect -4976 371 -4878 478
rect -5384 243 -5326 251
rect -4972 247 -4878 371
rect -5384 191 -5378 243
rect -5326 226 -5311 243
rect -5326 198 -5309 226
rect -5326 191 -5311 198
rect -5384 183 -5311 191
rect -4972 195 -4958 247
rect -4906 195 -4878 247
rect -5384 182 -5326 183
rect -5378 -2848 -5326 182
rect -4972 171 -4878 195
rect -5268 66 -5140 74
rect -5268 36 -5258 66
rect -5282 -14 -5258 36
rect -5268 -34 -5258 -14
rect -5146 36 -5140 66
rect -4714 40 -4645 456
rect -3314 261 -3220 541
rect -3314 209 -3292 261
rect -3240 209 -3220 261
rect -3314 182 -3220 209
rect -3610 66 -3482 74
rect -4716 36 -4644 40
rect -3610 36 -3600 66
rect -5146 -14 -4644 36
rect -3624 -14 -3600 36
rect -5146 -34 -5140 -14
rect -5268 -42 -5140 -34
rect -4982 -876 -4925 -14
rect -4714 -21 -4645 -14
rect -3610 -34 -3600 -14
rect -3488 36 -3482 66
rect -3059 68 -2988 430
rect -3059 36 -2986 68
rect -3488 -14 -2986 36
rect -3488 -34 -3482 -14
rect -3610 -42 -3482 -34
rect -3216 -724 -3145 -14
rect -2369 -41 -2323 -40
rect -2369 -198 -2320 -41
rect -3218 -730 -3145 -724
rect -3218 -782 -3212 -730
rect -3160 -782 -3145 -730
rect -3218 -788 -3145 -782
rect -3215 -791 -3145 -788
rect -2368 -390 -2320 -198
rect -4986 -883 -4915 -876
rect -4988 -889 -4915 -883
rect -4988 -941 -4982 -889
rect -4930 -941 -4915 -889
rect -4988 -947 -4915 -941
rect -4985 -950 -4915 -947
rect -4982 -957 -4925 -950
rect -2368 -1248 -2333 -390
rect -2236 -484 -2202 -264
rect -2237 -491 -2174 -484
rect -2237 -544 -2232 -491
rect -2180 -544 -2174 -491
rect -2237 -550 -2174 -544
rect -2118 -1187 -2083 -130
rect -1866 -395 -1787 0
rect -1866 -491 -1802 -395
rect -1290 -406 -1236 -94
rect -1774 -483 -1711 -427
rect -1866 -544 -1859 -491
rect -1807 -544 -1802 -491
rect -1866 -550 -1802 -544
rect -1772 -601 -1716 -483
rect -1358 -496 -1292 -434
rect -1264 -524 -1236 -406
rect -1065 -474 -1031 612
rect -829 -474 -795 -145
rect -1065 -507 -783 -474
rect -1283 -550 -1236 -524
rect -1775 -611 -1711 -601
rect -1775 -664 -1768 -611
rect -1716 -664 -1711 -611
rect -1775 -670 -1711 -664
rect -2010 -810 -1938 -809
rect -2012 -813 -1938 -810
rect -2012 -870 -2003 -813
rect -1945 -870 -1938 -813
rect -2012 -879 -1938 -870
rect -2257 -1233 -1694 -1187
rect -2519 -1302 -2285 -1248
rect -2519 -1303 -2400 -1302
rect -2519 -1631 -2473 -1303
rect -2257 -1328 -2225 -1233
rect -2272 -1512 -2225 -1328
rect -2389 -2774 -2361 -1519
rect -1401 -1526 -1367 -1203
rect -1861 -1864 -1822 -1526
rect -1679 -1678 -1643 -1677
rect -1679 -1856 -1632 -1678
rect -1861 -2773 -1833 -1864
rect -1668 -1868 -1632 -1856
rect -1664 -1961 -1632 -1868
rect -1414 -1789 -1367 -1526
rect -1665 -1970 -1596 -1961
rect -1665 -2022 -1654 -1970
rect -1602 -2022 -1596 -1970
rect -1665 -2029 -1596 -2022
rect -2413 -2793 -2334 -2774
rect -2540 -2838 -2462 -2819
rect -2540 -2848 -2524 -2838
rect -5378 -2876 -2524 -2848
rect -2540 -2880 -2524 -2876
rect -2479 -2880 -2462 -2838
rect -2413 -2835 -2397 -2793
rect -2352 -2835 -2334 -2793
rect -2413 -2855 -2334 -2835
rect -1882 -2792 -1803 -2773
rect -1414 -2779 -1386 -1789
rect -1283 -1817 -1249 -550
rect -817 -731 -783 -507
rect -699 -635 -665 1527
rect -463 -428 -429 2076
rect -242 1611 -176 1623
rect -242 1575 -230 1611
rect -188 1575 -176 1611
rect -242 1563 -176 1575
rect -227 955 -193 1563
rect -228 -428 -193 955
rect -699 -669 -547 -635
rect -834 -737 -770 -731
rect -834 -789 -828 -737
rect -776 -789 -770 -737
rect -834 -795 -770 -789
rect -1053 -1482 -1019 -1197
rect -1358 -1857 -1249 -1817
rect -1358 -1863 -1292 -1857
rect -1054 -2186 -1019 -1482
rect -817 -1773 -783 -795
rect -581 -1773 -547 -669
rect -228 -939 -194 -428
rect -109 -492 -75 497
rect 129 -439 163 2077
rect 494 -477 528 2079
rect 584 2077 658 2089
rect 945 2131 1019 2140
rect 1242 2137 1276 2141
rect 945 2089 959 2131
rect 1004 2089 1019 2131
rect 945 2077 1019 2089
rect 1210 2128 1284 2137
rect 1210 2086 1224 2128
rect 1269 2086 1284 2128
rect 606 -477 637 2077
rect 974 1405 1008 2077
rect 1210 2074 1284 2086
rect 1242 1551 1276 2074
rect 1229 1544 1292 1551
rect 1229 1492 1235 1544
rect 1287 1492 1292 1544
rect 1229 1484 1292 1492
rect 4339 -3 4488 12
rect 4339 -103 4356 -3
rect 4468 -103 4488 -3
rect 4339 -120 4488 -103
rect 4318 -266 4470 -248
rect 4318 -278 4341 -266
rect 4141 -279 4341 -278
rect -109 -538 113 -492
rect 69 -868 104 -538
rect 69 -904 353 -868
rect -228 -972 221 -939
rect -423 -996 -359 -990
rect -423 -1048 -417 -996
rect -365 -1048 -359 -996
rect -423 -1054 -359 -1048
rect 187 -1044 221 -972
rect -404 -1100 -370 -1054
rect 187 -1076 234 -1044
rect -308 -1094 -231 -1082
rect -421 -1155 -353 -1100
rect -308 -1149 -296 -1094
rect -244 -1111 -231 -1094
rect -244 -1145 -77 -1111
rect -244 -1149 -231 -1145
rect -308 -1156 -231 -1149
rect -6 -1154 59 -1100
rect 203 -1104 234 -1076
rect 114 -1152 234 -1104
rect -308 -1157 -232 -1156
rect 203 -1180 234 -1152
rect 187 -1223 234 -1180
rect 325 -1187 353 -904
rect 723 -974 769 -304
rect 1914 -347 4341 -279
rect 899 -597 965 -543
rect 1018 -597 1084 -543
rect 812 -625 872 -610
rect 1116 -625 1170 -614
rect 812 -626 1170 -625
rect 812 -660 824 -626
rect 858 -628 1170 -626
rect 858 -660 1124 -628
rect 812 -662 1124 -660
rect 1158 -662 1170 -628
rect 812 -668 1170 -662
rect 812 -673 872 -668
rect 1116 -674 1170 -668
rect 1179 -772 1811 -744
rect 934 -821 992 -809
rect 1179 -821 1209 -772
rect 934 -823 1209 -821
rect 934 -857 946 -823
rect 980 -857 1209 -823
rect 1323 -807 1394 -801
rect 934 -870 992 -857
rect 1323 -859 1336 -807
rect 1388 -859 1394 -807
rect 1323 -873 1394 -859
rect 1771 -938 1811 -772
rect 1914 -797 1968 -347
rect 4318 -367 4341 -347
rect 4447 -367 4470 -266
rect 4318 -391 4470 -367
rect 1911 -803 1975 -797
rect 1911 -855 1917 -803
rect 1969 -855 1975 -803
rect 1911 -861 1975 -855
rect 1771 -974 2421 -938
rect 723 -1016 1602 -974
rect 1421 -1050 1490 -1044
rect 1550 -1048 1602 -1016
rect 381 -1161 443 -1104
rect 499 -1161 561 -1104
rect 1112 -1158 1174 -1101
rect 1421 -1102 1430 -1050
rect 1482 -1102 1490 -1050
rect 1421 -1106 1490 -1102
rect 1540 -1104 1860 -1048
rect 1738 -1134 1768 -1104
rect 325 -1215 368 -1187
rect -469 -1725 -422 -1489
rect -469 -1782 -402 -1725
rect -892 -1865 -709 -1815
rect -818 -2038 -784 -1865
rect -538 -1870 -472 -1813
rect -831 -2045 -768 -2038
rect -831 -2097 -825 -2045
rect -773 -2097 -768 -2045
rect -831 -2105 -768 -2097
rect -1054 -2779 -1020 -2186
rect -442 -2389 -402 -1782
rect -452 -2395 -388 -2389
rect -452 -2447 -446 -2395
rect -394 -2447 -388 -2395
rect -452 -2453 -388 -2447
rect -227 -2774 -193 -1527
rect -52 -1750 -15 -1489
rect -52 -1964 -14 -1750
rect 187 -1771 221 -1223
rect 334 -1309 368 -1215
rect 570 -1791 620 -1400
rect 1738 -1418 1786 -1134
rect 1182 -1788 1236 -1513
rect 377 -1822 439 -1821
rect 377 -1878 443 -1822
rect 496 -1876 558 -1819
rect -60 -1971 5 -1964
rect -60 -2023 -54 -1971
rect -2 -2023 5 -1971
rect -60 -2030 5 -2023
rect -1882 -2834 -1866 -2792
rect -1821 -2834 -1803 -2792
rect -1882 -2854 -1803 -2834
rect -1440 -2798 -1361 -2779
rect -1440 -2840 -1424 -2798
rect -1379 -2840 -1361 -2798
rect -1440 -2860 -1361 -2840
rect -1074 -2798 -995 -2779
rect -1074 -2840 -1058 -2798
rect -1013 -2840 -995 -2798
rect -1074 -2860 -995 -2840
rect -255 -2793 -176 -2774
rect 586 -2777 620 -1791
rect 874 -1872 936 -1818
rect 992 -1872 1054 -1818
rect 1110 -1870 1172 -1816
rect 994 -2010 1052 -1872
rect 990 -2016 1054 -2010
rect 990 -2068 996 -2016
rect 1048 -2068 1054 -2016
rect 990 -2074 1054 -2068
rect 1202 -2770 1236 -1788
rect 1622 -2765 1656 -1511
rect 1876 -2761 1910 -1511
rect 2381 -2529 2421 -974
rect 3389 -2455 3665 -2427
rect 3389 -2529 3420 -2455
rect 2381 -2585 3420 -2529
rect 3389 -2656 3420 -2585
rect 3630 -2656 3665 -2455
rect 3389 -2682 3665 -2656
rect -255 -2835 -239 -2793
rect -194 -2835 -176 -2793
rect -255 -2855 -176 -2835
rect 561 -2796 640 -2777
rect 561 -2838 577 -2796
rect 622 -2838 640 -2796
rect 561 -2858 640 -2838
rect 1184 -2789 1263 -2770
rect 1184 -2831 1200 -2789
rect 1245 -2831 1263 -2789
rect 1184 -2851 1263 -2831
rect 1592 -2784 1671 -2765
rect 1592 -2826 1608 -2784
rect 1653 -2826 1671 -2784
rect 1592 -2846 1671 -2826
rect 1861 -2780 1940 -2761
rect 1861 -2822 1877 -2780
rect 1922 -2822 1940 -2780
rect 1861 -2842 1940 -2822
rect -2540 -2899 -2462 -2880
<< via1 >>
rect -2622 1870 -2570 1879
rect -2622 1834 -2616 1870
rect -2616 1834 -2582 1870
rect -2582 1834 -2570 1870
rect -2622 1827 -2570 1834
rect -2616 1755 -2564 1764
rect -2616 1719 -2610 1755
rect -2610 1719 -2576 1755
rect -2576 1719 -2564 1755
rect -2616 1712 -2564 1719
rect -5576 1510 -5464 1610
rect -3918 1510 -3806 1610
rect -1524 1648 -1472 1700
rect -5378 191 -5326 243
rect -4958 195 -4906 247
rect -5258 -34 -5146 66
rect -3292 209 -3240 261
rect -3600 -34 -3488 66
rect -3212 -782 -3160 -730
rect -4982 -941 -4930 -889
rect -2232 -544 -2180 -491
rect -1859 -544 -1807 -491
rect -1768 -664 -1716 -611
rect -2003 -822 -1945 -813
rect -2003 -867 -1998 -822
rect -1998 -867 -1949 -822
rect -1949 -867 -1945 -822
rect -2003 -870 -1945 -867
rect -1654 -2022 -1602 -1970
rect -828 -789 -776 -737
rect 1235 1492 1287 1544
rect 4356 -103 4468 -3
rect -417 -1048 -365 -996
rect -296 -1097 -244 -1094
rect -296 -1146 -244 -1097
rect 1336 -822 1388 -807
rect 1336 -859 1372 -822
rect 1372 -859 1388 -822
rect 4341 -367 4447 -266
rect 1917 -855 1969 -803
rect 1430 -1102 1482 -1050
rect -825 -2097 -773 -2045
rect -446 -2447 -394 -2395
rect -54 -2023 -2 -1971
rect 996 -2068 1048 -2016
rect 3420 -2656 3630 -2455
<< metal2 >>
rect 3307 2269 3482 2282
rect 3307 2238 3327 2269
rect 1620 2175 3327 2238
rect -7106 1875 -6904 2003
rect -2634 1879 -2562 1888
rect -7106 1874 -5382 1875
rect -2634 1874 -2622 1879
rect -7106 1827 -2622 1874
rect -2570 1827 -2562 1879
rect -7106 1825 -2562 1827
rect -6929 1823 -2562 1825
rect -5699 1822 -2562 1823
rect -2634 1816 -2562 1822
rect -2628 1764 -2556 1773
rect -7113 1760 -6911 1762
rect -7113 1758 -5391 1760
rect -2628 1758 -2616 1764
rect -7113 1712 -2616 1758
rect -2564 1712 -2556 1764
rect -7113 1708 -2556 1712
rect -7113 1584 -6911 1708
rect -5706 1706 -2556 1708
rect -2628 1701 -2556 1706
rect -1537 1702 -1460 1715
rect -1537 1646 -1526 1702
rect -1470 1646 -1460 1702
rect -1537 1630 -1460 1646
rect -5592 1614 -5448 1626
rect -5592 1506 -5582 1614
rect -5460 1506 -5448 1614
rect -5592 1496 -5448 1506
rect -3934 1614 -3790 1626
rect -3934 1506 -3924 1614
rect -3802 1506 -3790 1614
rect -3934 1496 -3790 1506
rect 1222 1546 1299 1559
rect 1222 1490 1233 1546
rect 1289 1490 1299 1546
rect 1222 1474 1299 1490
rect -3302 261 -3230 284
rect -5384 243 -5309 255
rect -5384 191 -5378 243
rect -5326 232 -5309 243
rect -4964 247 -4900 253
rect -4964 232 -4958 247
rect -5326 202 -4958 232
rect -5326 191 -5309 202
rect -5384 182 -5309 191
rect -4964 195 -4958 202
rect -4906 232 -4900 247
rect -3302 232 -3292 261
rect -4906 209 -3292 232
rect -3240 209 -3230 261
rect -4906 202 -3230 209
rect -4906 195 -4900 202
rect -3302 197 -3230 202
rect -4964 189 -4900 195
rect -5274 70 -5130 82
rect -5274 -38 -5264 70
rect -5142 -38 -5130 70
rect -5274 -48 -5130 -38
rect -3616 70 -3472 82
rect -3616 -38 -3606 70
rect -3484 -38 -3472 70
rect -3616 -48 -3472 -38
rect -7102 -125 -6900 -67
rect -7102 -167 -5503 -125
rect -7102 -245 -6900 -167
rect -7112 -536 -6910 -449
rect -7112 -567 -5711 -536
rect -7112 -627 -6910 -567
rect -5758 -821 -5711 -567
rect -5565 -619 -5503 -167
rect -2237 -491 -2174 -484
rect -2237 -544 -2232 -491
rect -2180 -508 -2174 -491
rect -1866 -491 -1802 -481
rect -1866 -508 -1859 -491
rect -2180 -544 -1859 -508
rect -1807 -544 -1802 -491
rect -2237 -550 -1802 -544
rect -1775 -611 -1711 -601
rect -5565 -620 -2200 -619
rect -1775 -620 -1768 -611
rect -5565 -660 -1768 -620
rect -5397 -661 -1768 -660
rect -1775 -664 -1768 -661
rect -1716 -664 -1711 -611
rect -1775 -670 -1711 -664
rect 1620 -692 1659 2175
rect 3307 2143 3327 2175
rect 3463 2234 3482 2269
rect 5065 2234 5267 2292
rect 3463 2171 5267 2234
rect 3463 2143 3482 2171
rect 3307 2129 3482 2143
rect 5065 2114 5267 2171
rect 4339 1 4485 12
rect 4339 -23 4352 1
rect 993 -722 1659 -692
rect 2297 -78 4352 -23
rect -3218 -730 -3154 -724
rect -3218 -782 -3212 -730
rect -3160 -745 -3154 -730
rect -834 -737 -770 -731
rect -834 -745 -828 -737
rect -3160 -778 -828 -745
rect -3160 -782 -3154 -778
rect -3218 -788 -3154 -782
rect -834 -789 -828 -778
rect -776 -748 -770 -737
rect 993 -748 1027 -722
rect -776 -778 1027 -748
rect -776 -789 -770 -778
rect -834 -795 -770 -789
rect -2012 -813 -1939 -806
rect -5758 -822 -3975 -821
rect -5758 -823 -2435 -822
rect -2012 -823 -2003 -813
rect -5758 -852 -2003 -823
rect -5546 -853 -2003 -852
rect -5396 -854 -2003 -853
rect -2012 -870 -2003 -854
rect -1945 -870 -1939 -813
rect -2012 -875 -1939 -870
rect 1323 -807 1394 -801
rect 1323 -859 1336 -807
rect 1388 -815 1394 -807
rect 1911 -803 1975 -797
rect 1911 -815 1917 -803
rect 1388 -845 1917 -815
rect 1388 -859 1394 -845
rect 1323 -873 1394 -859
rect 1911 -855 1917 -845
rect 1969 -855 1975 -803
rect 1911 -861 1975 -855
rect -4988 -889 -4924 -883
rect -4988 -941 -4982 -889
rect -4930 -904 -4924 -889
rect 1332 -904 1378 -873
rect -4930 -934 1378 -904
rect 1422 -883 1496 -874
rect -4930 -941 -4924 -934
rect -4988 -947 -4924 -941
rect 1422 -939 1430 -883
rect 1486 -939 1496 -883
rect 1422 -943 1496 -939
rect 1422 -944 1494 -943
rect -7114 -1002 -6912 -986
rect -423 -996 -359 -990
rect -7114 -1003 -849 -1002
rect -423 -1003 -417 -996
rect -7114 -1032 -417 -1003
rect -7114 -1164 -6912 -1032
rect -5264 -1033 -417 -1032
rect -423 -1048 -417 -1033
rect -365 -1048 -359 -996
rect -423 -1054 -359 -1048
rect 1421 -1050 1494 -944
rect -308 -1094 -232 -1082
rect -5584 -1111 -728 -1110
rect -308 -1111 -296 -1094
rect -5584 -1144 -296 -1111
rect -7117 -1590 -6915 -1521
rect -5584 -1590 -5529 -1144
rect -5244 -1145 -296 -1144
rect -308 -1146 -296 -1145
rect -244 -1146 -232 -1094
rect 1421 -1102 1430 -1050
rect 1482 -1102 1494 -1050
rect 1421 -1105 1494 -1102
rect 1421 -1106 1490 -1105
rect -308 -1160 -232 -1146
rect -7117 -1637 -5529 -1590
rect -7117 -1699 -6915 -1637
rect -1665 -1968 -1596 -1961
rect -60 -1968 5 -1964
rect -1665 -1970 5 -1968
rect -1665 -2022 -1654 -1970
rect -1602 -1971 5 -1970
rect -1602 -2002 -54 -1971
rect -1602 -2022 -1596 -2002
rect -61 -2006 -54 -2002
rect -1665 -2029 -1596 -2022
rect -60 -2023 -54 -2006
rect -2 -2023 5 -1971
rect -60 -2030 5 -2023
rect 990 -2016 1054 -2010
rect 990 -2026 996 -2016
rect -838 -2043 -761 -2030
rect -7117 -2150 -6915 -2078
rect -838 -2099 -827 -2043
rect -771 -2099 -761 -2043
rect 989 -2056 996 -2026
rect 990 -2068 996 -2056
rect 1048 -2068 1054 -2016
rect 990 -2074 1054 -2068
rect -838 -2115 -761 -2099
rect -7117 -2151 612 -2150
rect 999 -2151 1045 -2074
rect -7117 -2197 1044 -2151
rect -7117 -2256 -6915 -2197
rect -5246 -2198 1044 -2197
rect -452 -2395 -388 -2389
rect -452 -2447 -446 -2395
rect -394 -2412 -388 -2395
rect 2297 -2412 2331 -78
rect 4339 -107 4352 -78
rect 4474 -107 4485 1
rect 4339 -118 4485 -107
rect 4340 -119 4484 -118
rect 4318 -266 4470 -248
rect 4318 -367 4341 -266
rect 4447 -282 4470 -266
rect 4925 -282 5127 -215
rect 4447 -345 5127 -282
rect 4447 -367 4470 -345
rect 4318 -391 4470 -367
rect 4925 -393 5127 -345
rect -394 -2446 2331 -2412
rect -394 -2447 -388 -2446
rect -452 -2453 -388 -2447
rect 3389 -2455 3665 -2427
rect 3389 -2656 3420 -2455
rect 3630 -2656 3665 -2455
rect 3389 -2682 3665 -2656
<< via2 >>
rect -1526 1700 -1470 1702
rect -1526 1648 -1524 1700
rect -1524 1648 -1472 1700
rect -1472 1648 -1470 1700
rect -1526 1646 -1470 1648
rect -5582 1610 -5460 1614
rect -5582 1510 -5576 1610
rect -5576 1510 -5464 1610
rect -5464 1510 -5460 1610
rect -5582 1506 -5460 1510
rect -3924 1610 -3802 1614
rect -3924 1510 -3918 1610
rect -3918 1510 -3806 1610
rect -3806 1510 -3802 1610
rect -3924 1506 -3802 1510
rect 1233 1544 1289 1546
rect 1233 1492 1235 1544
rect 1235 1492 1287 1544
rect 1287 1492 1289 1544
rect 1233 1490 1289 1492
rect -5264 66 -5142 70
rect -5264 -34 -5258 66
rect -5258 -34 -5146 66
rect -5146 -34 -5142 66
rect -5264 -38 -5142 -34
rect -3606 66 -3484 70
rect -3606 -34 -3600 66
rect -3600 -34 -3488 66
rect -3488 -34 -3484 66
rect -3606 -38 -3484 -34
rect 3327 2143 3463 2269
rect 4352 -3 4474 1
rect 1430 -939 1486 -883
rect -827 -2045 -771 -2043
rect -827 -2097 -825 -2045
rect -825 -2097 -773 -2045
rect -773 -2097 -771 -2045
rect -827 -2099 -771 -2097
rect 4352 -103 4356 -3
rect 4356 -103 4468 -3
rect 4468 -103 4474 -3
rect 4352 -107 4474 -103
rect 4341 -367 4447 -266
rect 3420 -2656 3630 -2455
<< metal3 >>
rect 3307 2269 3482 2282
rect 3307 2143 3327 2269
rect 3463 2143 3482 2269
rect 3307 2129 3482 2143
rect -1537 1702 -1460 1715
rect -1537 1646 -1526 1702
rect -1470 1646 -1460 1702
rect -1537 1630 -1460 1646
rect -5592 1618 -5450 1624
rect -5592 1502 -5586 1618
rect -5458 1502 -5450 1618
rect -5592 1496 -5450 1502
rect -3934 1618 -3792 1624
rect -3934 1502 -3928 1618
rect -3800 1502 -3792 1618
rect -3934 1496 -3792 1502
rect -5274 74 -5132 80
rect -5274 -42 -5268 74
rect -5140 -42 -5132 74
rect -5274 -48 -5132 -42
rect -3616 74 -3474 80
rect -3616 -42 -3610 74
rect -3482 -42 -3474 74
rect -3616 -48 -3474 -42
rect -1534 -2031 -1462 1630
rect 1222 1546 1299 1559
rect 1222 1490 1233 1546
rect 1289 1490 1299 1546
rect 1222 1474 1299 1490
rect 1230 -831 1293 1474
rect 4342 5 4484 11
rect 4342 -111 4350 5
rect 4478 -111 4484 5
rect 4342 -117 4484 -111
rect 4318 -266 4470 -248
rect 4318 -367 4341 -266
rect 4447 -367 4470 -266
rect 4318 -391 4470 -367
rect 1230 -883 1496 -831
rect 1230 -894 1430 -883
rect 1422 -939 1430 -894
rect 1486 -939 1496 -883
rect 1422 -944 1496 -939
rect -838 -2031 -761 -2030
rect -1534 -2043 -761 -2031
rect -1534 -2099 -827 -2043
rect -771 -2099 -761 -2043
rect -1534 -2112 -761 -2099
rect -838 -2115 -761 -2112
rect 3389 -2455 3665 -2427
rect 3389 -2656 3420 -2455
rect 3630 -2656 3665 -2455
rect 3389 -2682 3665 -2656
<< via3 >>
rect 3327 2143 3463 2269
rect -5586 1614 -5458 1618
rect -5586 1506 -5582 1614
rect -5582 1506 -5460 1614
rect -5460 1506 -5458 1614
rect -5586 1502 -5458 1506
rect -3928 1614 -3800 1618
rect -3928 1506 -3924 1614
rect -3924 1506 -3802 1614
rect -3802 1506 -3800 1614
rect -3928 1502 -3800 1506
rect -5268 70 -5140 74
rect -5268 -38 -5264 70
rect -5264 -38 -5142 70
rect -5142 -38 -5140 70
rect -5268 -42 -5140 -38
rect -3610 70 -3482 74
rect -3610 -38 -3606 70
rect -3606 -38 -3484 70
rect -3484 -38 -3482 70
rect -3610 -42 -3482 -38
rect 4350 1 4478 5
rect 4350 -107 4352 1
rect 4352 -107 4474 1
rect 4474 -107 4478 1
rect 4350 -111 4478 -107
rect 4341 -367 4447 -266
rect 3420 -2656 3630 -2455
<< metal4 >>
rect 3307 2269 3482 2282
rect 3307 2143 3327 2269
rect 3463 2143 3482 2269
rect 3307 2129 3482 2143
rect -5594 1618 -5448 1626
rect -5594 1502 -5586 1618
rect -5458 1502 -5448 1618
rect -5594 1496 -5448 1502
rect -3936 1618 -3790 1626
rect -3936 1502 -3928 1618
rect -3800 1502 -3790 1618
rect -3936 1496 -3790 1502
rect -5539 1259 -5476 1496
rect -5540 844 -5476 1259
rect -3880 981 -3817 1496
rect -3878 932 -3817 981
rect 3338 946 3443 2129
rect -5234 82 -5174 456
rect -3576 82 -3516 626
rect 4359 83 4465 1075
rect -5276 74 -5130 82
rect -5276 -42 -5268 74
rect -5140 -42 -5130 74
rect -5276 -48 -5130 -42
rect -3618 74 -3472 82
rect -3618 -42 -3610 74
rect -3482 -42 -3472 74
rect 4360 11 4466 83
rect -3618 -48 -3472 -42
rect 4340 5 4486 11
rect -5218 -60 -5158 -48
rect -3560 -60 -3500 -48
rect 4340 -111 4350 5
rect 4478 -111 4486 5
rect 4340 -119 4486 -111
rect 4318 -266 4470 -248
rect 4318 -367 4341 -266
rect 4447 -367 4470 -266
rect 4318 -391 4470 -367
rect 4350 -690 4435 -391
rect 3470 -2427 3582 -1531
rect 4354 -2073 4430 -690
rect 3389 -2455 3665 -2427
rect 3389 -2656 3420 -2455
rect 3630 -2656 3665 -2455
rect 3389 -2682 3665 -2656
use res20_046K  res20_046K_0
timestamp 1668144350
transform 1 0 -4718 0 1 145
box -274 0 74 1528
use res20_046K  res20_046K_1
timestamp 1668144350
transform 1 0 -3060 0 1 39
box -274 0 74 1528
use sky130_fd_pr__cap_mim_m3_1_2TJQJA  sky130_fd_pr__cap_mim_m3_1_2TJQJA_0
timestamp 1668227070
transform 1 0 -5510 0 1 715
box -356 -306 355 306
use sky130_fd_pr__cap_mim_m3_1_2TJQJA  sky130_fd_pr__cap_mim_m3_1_2TJQJA_1
timestamp 1668227070
transform 1 0 -3849 0 1 818
box -356 -306 355 306
use sky130_fd_pr__cap_mim_m3_1_UJT6R3  sky130_fd_pr__cap_mim_m3_1_UJT6R3_0
timestamp 1668228500
transform 1 0 3614 0 1 1014
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_UJT6R3  sky130_fd_pr__cap_mim_m3_1_UJT6R3_1
timestamp 1668228500
transform 1 0 3595 0 1 -1301
box -850 -800 849 800
use sky130_fd_pr__nfet_01v8_4LH4MW  sky130_fd_pr__nfet_01v8_4LH4MW_0
timestamp 1668300629
transform 1 0 -1036 0 1 -1486
box -147 -326 147 369
use sky130_fd_pr__nfet_01v8_DDE7UB  sky130_fd_pr__nfet_01v8_DDE7UB_0
timestamp 1668224055
transform 1 0 -1750 0 1 -1537
box -118 -357 118 357
use sky130_fd_pr__nfet_01v8_PW4FSF  sky130_fd_pr__nfet_01v8_PW4FSF_0
timestamp 1668225783
transform 1 0 411 0 1 -1489
box -88 -388 88 388
use sky130_fd_pr__nfet_01v8_PW4FSF  sky130_fd_pr__nfet_01v8_PW4FSF_1
timestamp 1668225783
transform 1 0 529 0 1 -1489
box -88 -388 88 388
use sky130_fd_pr__nfet_01v8_PW4FSF  sky130_fd_pr__nfet_01v8_PW4FSF_2
timestamp 1668225783
transform 1 0 1140 0 1 -1486
box -88 -388 88 388
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_0
timestamp 1668226193
transform 1 0 -1325 0 1 -1520
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_1
timestamp 1668226193
transform 1 0 -505 0 1 -1516
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_2
timestamp 1668226193
transform 1 0 904 0 1 -1517
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_PWLUNE  sky130_fd_pr__nfet_01v8_PWLUNE_3
timestamp 1668226193
transform 1 0 1022 0 1 -1517
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_QSQEJU  sky130_fd_pr__nfet_01v8_QSQEJU_0
timestamp 1668225108
transform 1 0 -121 0 1 -1454
box -118 -357 118 357
use sky130_fd_pr__nfet_01v8_QSSMMX  sky130_fd_pr__nfet_01v8_QSSMMX_0
timestamp 1668223655
transform 1 0 -2434 0 1 -1601
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_VXZ4X9  sky130_fd_pr__nfet_01v8_VXZ4X9_0
timestamp 1668226574
transform 1 0 1458 0 1 -1703
box -88 -657 88 657
use sky130_fd_pr__nfet_01v8_VXZ4X9  sky130_fd_pr__nfet_01v8_VXZ4X9_1
timestamp 1668226574
transform 1 0 1576 0 1 -1703
box -88 -657 88 657
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_0
timestamp 1668294244
transform 1 0 -2316 0 1 -1601
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_1
timestamp 1668294244
transform 1 0 145 0 1 -1454
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_2
timestamp 1668294244
transform 1 0 -387 0 1 -1454
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_3
timestamp 1668294244
transform 1 0 27 0 1 -1454
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_4
timestamp 1668294244
transform 1 0 1818 0 1 -1401
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_VXZEP9  sky130_fd_pr__nfet_01v8_VXZEP9_5
timestamp 1668294244
transform 1 0 -269 0 1 -1454
box -88 -357 88 357
use sky130_fd_pr__nfet_01v8_ZG8UN4  sky130_fd_pr__nfet_01v8_ZG8UN4_0
timestamp 1668299617
transform 1 0 -800 0 1 -1517
box -147 -357 147 398
use sky130_fd_pr__pfet_01v8_3AH94A  sky130_fd_pr__pfet_01v8_3AH94A_0
timestamp 1668221973
transform 1 0 -1744 0 1 525
box -124 -1024 124 1058
use sky130_fd_pr__pfet_01v8_BGAJ3C  sky130_fd_pr__pfet_01v8_BGAJ3C_0
timestamp 1668223390
transform 1 0 -2160 0 1 567
box -124 -1058 124 1024
use sky130_fd_pr__pfet_01v8_BGN7SB  sky130_fd_pr__pfet_01v8_BGN7SB_0
timestamp 1668299723
transform 1 0 -930 0 1 556
box -183 -1058 183 1024
use sky130_fd_pr__pfet_01v8_DLEZW3  sky130_fd_pr__pfet_01v8_DLEZW3_0
timestamp 1668221782
transform 1 0 -2278 0 1 567
box -124 -1058 124 1024
use sky130_fd_pr__pfet_01v8_FHN7S9  sky130_fd_pr__pfet_01v8_FHN7S9_0
timestamp 1668299617
transform 1 0 990 0 1 424
box -183 -1024 183 1058
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_0
timestamp 1668223090
transform 1 0 -623 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_1
timestamp 1668223090
transform 1 0 -505 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_2
timestamp 1668223090
transform 1 0 -387 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_3
timestamp 1668223090
transform 1 0 -269 0 1 520
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_4
timestamp 1668223090
transform 1 0 334 0 1 478
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_5
timestamp 1668223090
transform 1 0 452 0 1 478
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_JBAJ3C  sky130_fd_pr__pfet_01v8_JBAJ3C_6
timestamp 1668223090
transform 1 0 682 0 1 472
box -124 -1022 124 1022
use sky130_fd_pr__pfet_01v8_XLJZXD  sky130_fd_pr__pfet_01v8_XLJZXD_0
timestamp 1668221782
transform 1 0 -1325 0 1 579
box -124 -1084 124 1118
use sky130_fd_pr__pfet_01v8_ZF98YR  sky130_fd_pr__pfet_01v8_ZF98YR_0
timestamp 1668222928
transform 1 0 27 0 1 -7
box -184 -544 184 578
<< labels >>
rlabel nsubdiffcont -2216 2018 1290 2144 7 VDD
port 1 w
rlabel psubdiffcont -2612 -2948 2008 -2688 7 GND
port 2 w
rlabel metal2 -7093 -1680 -6944 -1550 1 Vbiasn
port 4 n
rlabel metal2 -7075 -218 -6925 -88 1 Vbp
port 5 n
rlabel metal2 -7090 -2230 -6948 -2100 1 Vin
port 6 n
rlabel metal2 -7085 -1145 -6943 -1015 1 Vip
port 7 n
rlabel metal2 -7086 -599 -6932 -465 1 Vcm
port 3 n
rlabel metal2 5089 2133 5240 2275 3 Vop
port 8 e
rlabel metal2 4948 -367 5103 -236 3 Von
port 9 e
rlabel metal2 -7080 1844 -6935 1987 7 Vabn
port 10 w
rlabel metal2 -7086 1611 -6936 1738 7 Vabp
port 11 w
<< end >>
