magic
tech sky130A
magscale 1 2
timestamp 1666707788
<< nwell >>
rect -296 -959 296 959
<< pmos >>
rect -100 -740 100 740
<< pdiff >>
rect -158 728 -100 740
rect -158 -728 -146 728
rect -112 -728 -100 728
rect -158 -740 -100 -728
rect 100 728 158 740
rect 100 -728 112 728
rect 146 -728 158 728
rect 100 -740 158 -728
<< pdiffc >>
rect -146 -728 -112 728
rect 112 -728 146 728
<< nsubdiff >>
rect -260 889 -164 923
rect 164 889 260 923
rect -260 827 -226 889
rect 226 827 260 889
rect -260 -889 -226 -827
rect 226 -889 260 -827
rect -260 -923 -164 -889
rect 164 -923 260 -889
<< nsubdiffcont >>
rect -164 889 164 923
rect -260 -827 -226 827
rect 226 -827 260 827
rect -164 -923 164 -889
<< poly >>
rect -100 821 100 837
rect -100 787 -84 821
rect 84 787 100 821
rect -100 740 100 787
rect -100 -787 100 -740
rect -100 -821 -84 -787
rect 84 -821 100 -787
rect -100 -837 100 -821
<< polycont >>
rect -84 787 84 821
rect -84 -821 84 -787
<< locali >>
rect -260 889 -164 923
rect 164 889 260 923
rect -260 827 -226 889
rect 226 827 260 889
rect -100 787 -84 821
rect 84 787 100 821
rect -146 728 -112 744
rect -146 -744 -112 -728
rect 112 728 146 744
rect 112 -744 146 -728
rect -100 -821 -84 -787
rect 84 -821 100 -787
rect -260 -889 -226 -827
rect 226 -889 260 -827
rect -260 -923 -164 -889
rect 164 -923 260 -889
<< viali >>
rect -84 787 84 821
rect -146 -728 -112 728
rect 112 -728 146 728
rect -84 -821 84 -787
<< metal1 >>
rect -96 821 96 827
rect -96 787 -84 821
rect 84 787 96 821
rect -96 781 96 787
rect -152 728 -106 740
rect -152 -728 -146 728
rect -112 -728 -106 728
rect -152 -740 -106 -728
rect 106 728 152 740
rect 106 -728 112 728
rect 146 -728 152 728
rect 106 -740 152 -728
rect -96 -787 96 -781
rect -96 -821 -84 -787
rect 84 -821 96 -787
rect -96 -827 96 -821
<< properties >>
string FIXED_BBOX -243 -906 243 906
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7.4 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
