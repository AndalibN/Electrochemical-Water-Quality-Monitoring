magic
tech sky130A
magscale 1 2
timestamp 1666402782
<< error_p >>
rect -29 822 29 828
rect -29 788 -17 822
rect -29 782 29 788
rect -29 -788 29 -782
rect -29 -822 -17 -788
rect -29 -828 29 -822
<< pwell >>
rect -226 -960 226 960
<< nmos >>
rect -30 -750 30 750
<< ndiff >>
rect -88 738 -30 750
rect -88 -738 -76 738
rect -42 -738 -30 738
rect -88 -750 -30 -738
rect 30 738 88 750
rect 30 -738 42 738
rect 76 -738 88 738
rect 30 -750 88 -738
<< ndiffc >>
rect -76 -738 -42 738
rect 42 -738 76 738
<< psubdiff >>
rect -190 890 -94 924
rect 94 890 190 924
rect -190 828 -156 890
rect 156 828 190 890
rect -190 -890 -156 -828
rect 156 -890 190 -828
rect -190 -924 -94 -890
rect 94 -924 190 -890
<< psubdiffcont >>
rect -94 890 94 924
rect -190 -828 -156 828
rect 156 -828 190 828
rect -94 -924 94 -890
<< poly >>
rect -33 822 33 838
rect -33 788 -17 822
rect 17 788 33 822
rect -33 772 33 788
rect -30 750 30 772
rect -30 -772 30 -750
rect -33 -788 33 -772
rect -33 -822 -17 -788
rect 17 -822 33 -788
rect -33 -838 33 -822
<< polycont >>
rect -17 788 17 822
rect -17 -822 17 -788
<< locali >>
rect -190 890 -94 924
rect 94 890 190 924
rect -190 828 -156 890
rect 156 828 190 890
rect -33 788 -17 822
rect 17 788 33 822
rect -76 738 -42 754
rect -76 -754 -42 -738
rect 42 738 76 754
rect 42 -754 76 -738
rect -33 -822 -17 -788
rect 17 -822 33 -788
rect -190 -890 -156 -828
rect 156 -890 190 -828
rect -190 -924 -94 -890
rect 94 -924 190 -890
<< viali >>
rect -17 788 17 822
rect -76 -738 -42 738
rect 42 -738 76 738
rect -17 -822 17 -788
<< metal1 >>
rect -29 822 29 828
rect -29 788 -17 822
rect 17 788 29 822
rect -29 782 29 788
rect -82 738 -36 750
rect -82 -738 -76 738
rect -42 -738 -36 738
rect -82 -750 -36 -738
rect 36 738 82 750
rect 36 -738 42 738
rect 76 -738 82 738
rect 36 -750 82 -738
rect -29 -788 29 -782
rect -29 -822 -17 -788
rect 17 -822 29 -788
rect -29 -828 29 -822
<< properties >>
string FIXED_BBOX -173 -907 173 907
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 7.5 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
