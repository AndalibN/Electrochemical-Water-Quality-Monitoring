magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 -811 29 -805
rect -29 -845 -17 -811
rect -29 -851 29 -845
<< nwell >>
rect -109 -864 109 898
<< pmos >>
rect -15 -764 15 836
<< pdiff >>
rect -73 801 -15 836
rect -73 767 -61 801
rect -27 767 -15 801
rect -73 733 -15 767
rect -73 699 -61 733
rect -27 699 -15 733
rect -73 665 -15 699
rect -73 631 -61 665
rect -27 631 -15 665
rect -73 597 -15 631
rect -73 563 -61 597
rect -27 563 -15 597
rect -73 529 -15 563
rect -73 495 -61 529
rect -27 495 -15 529
rect -73 461 -15 495
rect -73 427 -61 461
rect -27 427 -15 461
rect -73 393 -15 427
rect -73 359 -61 393
rect -27 359 -15 393
rect -73 325 -15 359
rect -73 291 -61 325
rect -27 291 -15 325
rect -73 257 -15 291
rect -73 223 -61 257
rect -27 223 -15 257
rect -73 189 -15 223
rect -73 155 -61 189
rect -27 155 -15 189
rect -73 121 -15 155
rect -73 87 -61 121
rect -27 87 -15 121
rect -73 53 -15 87
rect -73 19 -61 53
rect -27 19 -15 53
rect -73 -15 -15 19
rect -73 -49 -61 -15
rect -27 -49 -15 -15
rect -73 -83 -15 -49
rect -73 -117 -61 -83
rect -27 -117 -15 -83
rect -73 -151 -15 -117
rect -73 -185 -61 -151
rect -27 -185 -15 -151
rect -73 -219 -15 -185
rect -73 -253 -61 -219
rect -27 -253 -15 -219
rect -73 -287 -15 -253
rect -73 -321 -61 -287
rect -27 -321 -15 -287
rect -73 -355 -15 -321
rect -73 -389 -61 -355
rect -27 -389 -15 -355
rect -73 -423 -15 -389
rect -73 -457 -61 -423
rect -27 -457 -15 -423
rect -73 -491 -15 -457
rect -73 -525 -61 -491
rect -27 -525 -15 -491
rect -73 -559 -15 -525
rect -73 -593 -61 -559
rect -27 -593 -15 -559
rect -73 -627 -15 -593
rect -73 -661 -61 -627
rect -27 -661 -15 -627
rect -73 -695 -15 -661
rect -73 -729 -61 -695
rect -27 -729 -15 -695
rect -73 -764 -15 -729
rect 15 801 73 836
rect 15 767 27 801
rect 61 767 73 801
rect 15 733 73 767
rect 15 699 27 733
rect 61 699 73 733
rect 15 665 73 699
rect 15 631 27 665
rect 61 631 73 665
rect 15 597 73 631
rect 15 563 27 597
rect 61 563 73 597
rect 15 529 73 563
rect 15 495 27 529
rect 61 495 73 529
rect 15 461 73 495
rect 15 427 27 461
rect 61 427 73 461
rect 15 393 73 427
rect 15 359 27 393
rect 61 359 73 393
rect 15 325 73 359
rect 15 291 27 325
rect 61 291 73 325
rect 15 257 73 291
rect 15 223 27 257
rect 61 223 73 257
rect 15 189 73 223
rect 15 155 27 189
rect 61 155 73 189
rect 15 121 73 155
rect 15 87 27 121
rect 61 87 73 121
rect 15 53 73 87
rect 15 19 27 53
rect 61 19 73 53
rect 15 -15 73 19
rect 15 -49 27 -15
rect 61 -49 73 -15
rect 15 -83 73 -49
rect 15 -117 27 -83
rect 61 -117 73 -83
rect 15 -151 73 -117
rect 15 -185 27 -151
rect 61 -185 73 -151
rect 15 -219 73 -185
rect 15 -253 27 -219
rect 61 -253 73 -219
rect 15 -287 73 -253
rect 15 -321 27 -287
rect 61 -321 73 -287
rect 15 -355 73 -321
rect 15 -389 27 -355
rect 61 -389 73 -355
rect 15 -423 73 -389
rect 15 -457 27 -423
rect 61 -457 73 -423
rect 15 -491 73 -457
rect 15 -525 27 -491
rect 61 -525 73 -491
rect 15 -559 73 -525
rect 15 -593 27 -559
rect 61 -593 73 -559
rect 15 -627 73 -593
rect 15 -661 27 -627
rect 61 -661 73 -627
rect 15 -695 73 -661
rect 15 -729 27 -695
rect 61 -729 73 -695
rect 15 -764 73 -729
<< pdiffc >>
rect -61 767 -27 801
rect -61 699 -27 733
rect -61 631 -27 665
rect -61 563 -27 597
rect -61 495 -27 529
rect -61 427 -27 461
rect -61 359 -27 393
rect -61 291 -27 325
rect -61 223 -27 257
rect -61 155 -27 189
rect -61 87 -27 121
rect -61 19 -27 53
rect -61 -49 -27 -15
rect -61 -117 -27 -83
rect -61 -185 -27 -151
rect -61 -253 -27 -219
rect -61 -321 -27 -287
rect -61 -389 -27 -355
rect -61 -457 -27 -423
rect -61 -525 -27 -491
rect -61 -593 -27 -559
rect -61 -661 -27 -627
rect -61 -729 -27 -695
rect 27 767 61 801
rect 27 699 61 733
rect 27 631 61 665
rect 27 563 61 597
rect 27 495 61 529
rect 27 427 61 461
rect 27 359 61 393
rect 27 291 61 325
rect 27 223 61 257
rect 27 155 61 189
rect 27 87 61 121
rect 27 19 61 53
rect 27 -49 61 -15
rect 27 -117 61 -83
rect 27 -185 61 -151
rect 27 -253 61 -219
rect 27 -321 61 -287
rect 27 -389 61 -355
rect 27 -457 61 -423
rect 27 -525 61 -491
rect 27 -593 61 -559
rect 27 -661 61 -627
rect 27 -729 61 -695
<< poly >>
rect -15 836 15 862
rect -15 -795 15 -764
rect -33 -811 33 -795
rect -33 -845 -17 -811
rect 17 -845 33 -811
rect -33 -861 33 -845
<< polycont >>
rect -17 -845 17 -811
<< locali >>
rect -61 809 -27 840
rect -61 737 -27 767
rect -61 665 -27 699
rect -61 597 -27 631
rect -61 529 -27 559
rect -61 461 -27 487
rect -61 393 -27 415
rect -61 325 -27 343
rect -61 257 -27 271
rect -61 189 -27 199
rect -61 121 -27 127
rect -61 53 -27 55
rect -61 17 -27 19
rect -61 -55 -27 -49
rect -61 -127 -27 -117
rect -61 -199 -27 -185
rect -61 -271 -27 -253
rect -61 -343 -27 -321
rect -61 -415 -27 -389
rect -61 -487 -27 -457
rect -61 -559 -27 -525
rect -61 -627 -27 -593
rect -61 -695 -27 -665
rect -61 -768 -27 -737
rect 27 809 61 840
rect 27 737 61 767
rect 27 665 61 699
rect 27 597 61 631
rect 27 529 61 559
rect 27 461 61 487
rect 27 393 61 415
rect 27 325 61 343
rect 27 257 61 271
rect 27 189 61 199
rect 27 121 61 127
rect 27 53 61 55
rect 27 17 61 19
rect 27 -55 61 -49
rect 27 -127 61 -117
rect 27 -199 61 -185
rect 27 -271 61 -253
rect 27 -343 61 -321
rect 27 -415 61 -389
rect 27 -487 61 -457
rect 27 -559 61 -525
rect 27 -627 61 -593
rect 27 -695 61 -665
rect 27 -768 61 -737
rect -33 -845 -17 -811
rect 17 -845 33 -811
<< viali >>
rect -61 801 -27 809
rect -61 775 -27 801
rect -61 733 -27 737
rect -61 703 -27 733
rect -61 631 -27 665
rect -61 563 -27 593
rect -61 559 -27 563
rect -61 495 -27 521
rect -61 487 -27 495
rect -61 427 -27 449
rect -61 415 -27 427
rect -61 359 -27 377
rect -61 343 -27 359
rect -61 291 -27 305
rect -61 271 -27 291
rect -61 223 -27 233
rect -61 199 -27 223
rect -61 155 -27 161
rect -61 127 -27 155
rect -61 87 -27 89
rect -61 55 -27 87
rect -61 -15 -27 17
rect -61 -17 -27 -15
rect -61 -83 -27 -55
rect -61 -89 -27 -83
rect -61 -151 -27 -127
rect -61 -161 -27 -151
rect -61 -219 -27 -199
rect -61 -233 -27 -219
rect -61 -287 -27 -271
rect -61 -305 -27 -287
rect -61 -355 -27 -343
rect -61 -377 -27 -355
rect -61 -423 -27 -415
rect -61 -449 -27 -423
rect -61 -491 -27 -487
rect -61 -521 -27 -491
rect -61 -593 -27 -559
rect -61 -661 -27 -631
rect -61 -665 -27 -661
rect -61 -729 -27 -703
rect -61 -737 -27 -729
rect 27 801 61 809
rect 27 775 61 801
rect 27 733 61 737
rect 27 703 61 733
rect 27 631 61 665
rect 27 563 61 593
rect 27 559 61 563
rect 27 495 61 521
rect 27 487 61 495
rect 27 427 61 449
rect 27 415 61 427
rect 27 359 61 377
rect 27 343 61 359
rect 27 291 61 305
rect 27 271 61 291
rect 27 223 61 233
rect 27 199 61 223
rect 27 155 61 161
rect 27 127 61 155
rect 27 87 61 89
rect 27 55 61 87
rect 27 -15 61 17
rect 27 -17 61 -15
rect 27 -83 61 -55
rect 27 -89 61 -83
rect 27 -151 61 -127
rect 27 -161 61 -151
rect 27 -219 61 -199
rect 27 -233 61 -219
rect 27 -287 61 -271
rect 27 -305 61 -287
rect 27 -355 61 -343
rect 27 -377 61 -355
rect 27 -423 61 -415
rect 27 -449 61 -423
rect 27 -491 61 -487
rect 27 -521 61 -491
rect 27 -593 61 -559
rect 27 -661 61 -631
rect 27 -665 61 -661
rect 27 -729 61 -703
rect 27 -737 61 -729
rect -17 -845 17 -811
<< metal1 >>
rect -67 809 -21 836
rect -67 775 -61 809
rect -27 775 -21 809
rect -67 737 -21 775
rect -67 703 -61 737
rect -27 703 -21 737
rect -67 665 -21 703
rect -67 631 -61 665
rect -27 631 -21 665
rect -67 593 -21 631
rect -67 559 -61 593
rect -27 559 -21 593
rect -67 521 -21 559
rect -67 487 -61 521
rect -27 487 -21 521
rect -67 449 -21 487
rect -67 415 -61 449
rect -27 415 -21 449
rect -67 377 -21 415
rect -67 343 -61 377
rect -27 343 -21 377
rect -67 305 -21 343
rect -67 271 -61 305
rect -27 271 -21 305
rect -67 233 -21 271
rect -67 199 -61 233
rect -27 199 -21 233
rect -67 161 -21 199
rect -67 127 -61 161
rect -27 127 -21 161
rect -67 89 -21 127
rect -67 55 -61 89
rect -27 55 -21 89
rect -67 17 -21 55
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -55 -21 -17
rect -67 -89 -61 -55
rect -27 -89 -21 -55
rect -67 -127 -21 -89
rect -67 -161 -61 -127
rect -27 -161 -21 -127
rect -67 -199 -21 -161
rect -67 -233 -61 -199
rect -27 -233 -21 -199
rect -67 -271 -21 -233
rect -67 -305 -61 -271
rect -27 -305 -21 -271
rect -67 -343 -21 -305
rect -67 -377 -61 -343
rect -27 -377 -21 -343
rect -67 -415 -21 -377
rect -67 -449 -61 -415
rect -27 -449 -21 -415
rect -67 -487 -21 -449
rect -67 -521 -61 -487
rect -27 -521 -21 -487
rect -67 -559 -21 -521
rect -67 -593 -61 -559
rect -27 -593 -21 -559
rect -67 -631 -21 -593
rect -67 -665 -61 -631
rect -27 -665 -21 -631
rect -67 -703 -21 -665
rect -67 -737 -61 -703
rect -27 -737 -21 -703
rect -67 -764 -21 -737
rect 21 809 67 836
rect 21 775 27 809
rect 61 775 67 809
rect 21 737 67 775
rect 21 703 27 737
rect 61 703 67 737
rect 21 665 67 703
rect 21 631 27 665
rect 61 631 67 665
rect 21 593 67 631
rect 21 559 27 593
rect 61 559 67 593
rect 21 521 67 559
rect 21 487 27 521
rect 61 487 67 521
rect 21 449 67 487
rect 21 415 27 449
rect 61 415 67 449
rect 21 377 67 415
rect 21 343 27 377
rect 61 343 67 377
rect 21 305 67 343
rect 21 271 27 305
rect 61 271 67 305
rect 21 233 67 271
rect 21 199 27 233
rect 61 199 67 233
rect 21 161 67 199
rect 21 127 27 161
rect 61 127 67 161
rect 21 89 67 127
rect 21 55 27 89
rect 61 55 67 89
rect 21 17 67 55
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -55 67 -17
rect 21 -89 27 -55
rect 61 -89 67 -55
rect 21 -127 67 -89
rect 21 -161 27 -127
rect 61 -161 67 -127
rect 21 -199 67 -161
rect 21 -233 27 -199
rect 61 -233 67 -199
rect 21 -271 67 -233
rect 21 -305 27 -271
rect 61 -305 67 -271
rect 21 -343 67 -305
rect 21 -377 27 -343
rect 61 -377 67 -343
rect 21 -415 67 -377
rect 21 -449 27 -415
rect 61 -449 67 -415
rect 21 -487 67 -449
rect 21 -521 27 -487
rect 61 -521 67 -487
rect 21 -559 67 -521
rect 21 -593 27 -559
rect 61 -593 67 -559
rect 21 -631 67 -593
rect 21 -665 27 -631
rect 61 -665 67 -631
rect 21 -703 67 -665
rect 21 -737 27 -703
rect 61 -737 67 -703
rect 21 -764 67 -737
rect -29 -811 29 -805
rect -29 -845 -17 -811
rect 17 -845 29 -811
rect -29 -851 29 -845
<< end >>
