magic
tech sky130A
timestamp 1668374365
<< nmos >>
rect -1639 -4000 -1609 4000
rect -1523 -4000 -1493 4000
rect -1407 -4000 -1377 4000
rect -1291 -4000 -1261 4000
rect -1175 -4000 -1145 4000
rect -1059 -4000 -1029 4000
rect -943 -4000 -913 4000
rect -827 -4000 -797 4000
rect -711 -4000 -681 4000
rect -595 -4000 -565 4000
rect -479 -4000 -449 4000
rect -363 -4000 -333 4000
rect -247 -4000 -217 4000
rect -131 -4000 -101 4000
rect -15 -4000 15 4000
rect 101 -4000 131 4000
rect 217 -4000 247 4000
rect 333 -4000 363 4000
rect 449 -4000 479 4000
rect 565 -4000 595 4000
rect 681 -4000 711 4000
rect 797 -4000 827 4000
rect 913 -4000 943 4000
rect 1029 -4000 1059 4000
rect 1145 -4000 1175 4000
rect 1261 -4000 1291 4000
rect 1377 -4000 1407 4000
rect 1493 -4000 1523 4000
rect 1609 -4000 1639 4000
<< ndiff >>
rect -1668 3994 -1639 4000
rect -1668 -3994 -1662 3994
rect -1645 -3994 -1639 3994
rect -1668 -4000 -1639 -3994
rect -1609 3994 -1580 4000
rect -1609 -3994 -1603 3994
rect -1586 -3994 -1580 3994
rect -1609 -4000 -1580 -3994
rect -1552 3994 -1523 4000
rect -1552 -3994 -1546 3994
rect -1529 -3994 -1523 3994
rect -1552 -4000 -1523 -3994
rect -1493 3994 -1464 4000
rect -1493 -3994 -1487 3994
rect -1470 -3994 -1464 3994
rect -1493 -4000 -1464 -3994
rect -1436 3994 -1407 4000
rect -1436 -3994 -1430 3994
rect -1413 -3994 -1407 3994
rect -1436 -4000 -1407 -3994
rect -1377 3994 -1348 4000
rect -1377 -3994 -1371 3994
rect -1354 -3994 -1348 3994
rect -1377 -4000 -1348 -3994
rect -1320 3994 -1291 4000
rect -1320 -3994 -1314 3994
rect -1297 -3994 -1291 3994
rect -1320 -4000 -1291 -3994
rect -1261 3994 -1232 4000
rect -1261 -3994 -1255 3994
rect -1238 -3994 -1232 3994
rect -1261 -4000 -1232 -3994
rect -1204 3994 -1175 4000
rect -1204 -3994 -1198 3994
rect -1181 -3994 -1175 3994
rect -1204 -4000 -1175 -3994
rect -1145 3994 -1116 4000
rect -1145 -3994 -1139 3994
rect -1122 -3994 -1116 3994
rect -1145 -4000 -1116 -3994
rect -1088 3994 -1059 4000
rect -1088 -3994 -1082 3994
rect -1065 -3994 -1059 3994
rect -1088 -4000 -1059 -3994
rect -1029 3994 -1000 4000
rect -1029 -3994 -1023 3994
rect -1006 -3994 -1000 3994
rect -1029 -4000 -1000 -3994
rect -972 3994 -943 4000
rect -972 -3994 -966 3994
rect -949 -3994 -943 3994
rect -972 -4000 -943 -3994
rect -913 3994 -884 4000
rect -913 -3994 -907 3994
rect -890 -3994 -884 3994
rect -913 -4000 -884 -3994
rect -856 3994 -827 4000
rect -856 -3994 -850 3994
rect -833 -3994 -827 3994
rect -856 -4000 -827 -3994
rect -797 3994 -768 4000
rect -797 -3994 -791 3994
rect -774 -3994 -768 3994
rect -797 -4000 -768 -3994
rect -740 3994 -711 4000
rect -740 -3994 -734 3994
rect -717 -3994 -711 3994
rect -740 -4000 -711 -3994
rect -681 3994 -652 4000
rect -681 -3994 -675 3994
rect -658 -3994 -652 3994
rect -681 -4000 -652 -3994
rect -624 3994 -595 4000
rect -624 -3994 -618 3994
rect -601 -3994 -595 3994
rect -624 -4000 -595 -3994
rect -565 3994 -536 4000
rect -565 -3994 -559 3994
rect -542 -3994 -536 3994
rect -565 -4000 -536 -3994
rect -508 3994 -479 4000
rect -508 -3994 -502 3994
rect -485 -3994 -479 3994
rect -508 -4000 -479 -3994
rect -449 3994 -420 4000
rect -449 -3994 -443 3994
rect -426 -3994 -420 3994
rect -449 -4000 -420 -3994
rect -392 3994 -363 4000
rect -392 -3994 -386 3994
rect -369 -3994 -363 3994
rect -392 -4000 -363 -3994
rect -333 3994 -304 4000
rect -333 -3994 -327 3994
rect -310 -3994 -304 3994
rect -333 -4000 -304 -3994
rect -276 3994 -247 4000
rect -276 -3994 -270 3994
rect -253 -3994 -247 3994
rect -276 -4000 -247 -3994
rect -217 3994 -188 4000
rect -217 -3994 -211 3994
rect -194 -3994 -188 3994
rect -217 -4000 -188 -3994
rect -160 3994 -131 4000
rect -160 -3994 -154 3994
rect -137 -3994 -131 3994
rect -160 -4000 -131 -3994
rect -101 3994 -72 4000
rect -101 -3994 -95 3994
rect -78 -3994 -72 3994
rect -101 -4000 -72 -3994
rect -44 3994 -15 4000
rect -44 -3994 -38 3994
rect -21 -3994 -15 3994
rect -44 -4000 -15 -3994
rect 15 3994 44 4000
rect 15 -3994 21 3994
rect 38 -3994 44 3994
rect 15 -4000 44 -3994
rect 72 3994 101 4000
rect 72 -3994 78 3994
rect 95 -3994 101 3994
rect 72 -4000 101 -3994
rect 131 3994 160 4000
rect 131 -3994 137 3994
rect 154 -3994 160 3994
rect 131 -4000 160 -3994
rect 188 3994 217 4000
rect 188 -3994 194 3994
rect 211 -3994 217 3994
rect 188 -4000 217 -3994
rect 247 3994 276 4000
rect 247 -3994 253 3994
rect 270 -3994 276 3994
rect 247 -4000 276 -3994
rect 304 3994 333 4000
rect 304 -3994 310 3994
rect 327 -3994 333 3994
rect 304 -4000 333 -3994
rect 363 3994 392 4000
rect 363 -3994 369 3994
rect 386 -3994 392 3994
rect 363 -4000 392 -3994
rect 420 3994 449 4000
rect 420 -3994 426 3994
rect 443 -3994 449 3994
rect 420 -4000 449 -3994
rect 479 3994 508 4000
rect 479 -3994 485 3994
rect 502 -3994 508 3994
rect 479 -4000 508 -3994
rect 536 3994 565 4000
rect 536 -3994 542 3994
rect 559 -3994 565 3994
rect 536 -4000 565 -3994
rect 595 3994 624 4000
rect 595 -3994 601 3994
rect 618 -3994 624 3994
rect 595 -4000 624 -3994
rect 652 3994 681 4000
rect 652 -3994 658 3994
rect 675 -3994 681 3994
rect 652 -4000 681 -3994
rect 711 3994 740 4000
rect 711 -3994 717 3994
rect 734 -3994 740 3994
rect 711 -4000 740 -3994
rect 768 3994 797 4000
rect 768 -3994 774 3994
rect 791 -3994 797 3994
rect 768 -4000 797 -3994
rect 827 3994 856 4000
rect 827 -3994 833 3994
rect 850 -3994 856 3994
rect 827 -4000 856 -3994
rect 884 3994 913 4000
rect 884 -3994 890 3994
rect 907 -3994 913 3994
rect 884 -4000 913 -3994
rect 943 3994 972 4000
rect 943 -3994 949 3994
rect 966 -3994 972 3994
rect 943 -4000 972 -3994
rect 1000 3994 1029 4000
rect 1000 -3994 1006 3994
rect 1023 -3994 1029 3994
rect 1000 -4000 1029 -3994
rect 1059 3994 1088 4000
rect 1059 -3994 1065 3994
rect 1082 -3994 1088 3994
rect 1059 -4000 1088 -3994
rect 1116 3994 1145 4000
rect 1116 -3994 1122 3994
rect 1139 -3994 1145 3994
rect 1116 -4000 1145 -3994
rect 1175 3994 1204 4000
rect 1175 -3994 1181 3994
rect 1198 -3994 1204 3994
rect 1175 -4000 1204 -3994
rect 1232 3994 1261 4000
rect 1232 -3994 1238 3994
rect 1255 -3994 1261 3994
rect 1232 -4000 1261 -3994
rect 1291 3994 1320 4000
rect 1291 -3994 1297 3994
rect 1314 -3994 1320 3994
rect 1291 -4000 1320 -3994
rect 1348 3994 1377 4000
rect 1348 -3994 1354 3994
rect 1371 -3994 1377 3994
rect 1348 -4000 1377 -3994
rect 1407 3994 1436 4000
rect 1407 -3994 1413 3994
rect 1430 -3994 1436 3994
rect 1407 -4000 1436 -3994
rect 1464 3994 1493 4000
rect 1464 -3994 1470 3994
rect 1487 -3994 1493 3994
rect 1464 -4000 1493 -3994
rect 1523 3994 1552 4000
rect 1523 -3994 1529 3994
rect 1546 -3994 1552 3994
rect 1523 -4000 1552 -3994
rect 1580 3994 1609 4000
rect 1580 -3994 1586 3994
rect 1603 -3994 1609 3994
rect 1580 -4000 1609 -3994
rect 1639 3994 1668 4000
rect 1639 -3994 1645 3994
rect 1662 -3994 1668 3994
rect 1639 -4000 1668 -3994
<< ndiffc >>
rect -1662 -3994 -1645 3994
rect -1603 -3994 -1586 3994
rect -1546 -3994 -1529 3994
rect -1487 -3994 -1470 3994
rect -1430 -3994 -1413 3994
rect -1371 -3994 -1354 3994
rect -1314 -3994 -1297 3994
rect -1255 -3994 -1238 3994
rect -1198 -3994 -1181 3994
rect -1139 -3994 -1122 3994
rect -1082 -3994 -1065 3994
rect -1023 -3994 -1006 3994
rect -966 -3994 -949 3994
rect -907 -3994 -890 3994
rect -850 -3994 -833 3994
rect -791 -3994 -774 3994
rect -734 -3994 -717 3994
rect -675 -3994 -658 3994
rect -618 -3994 -601 3994
rect -559 -3994 -542 3994
rect -502 -3994 -485 3994
rect -443 -3994 -426 3994
rect -386 -3994 -369 3994
rect -327 -3994 -310 3994
rect -270 -3994 -253 3994
rect -211 -3994 -194 3994
rect -154 -3994 -137 3994
rect -95 -3994 -78 3994
rect -38 -3994 -21 3994
rect 21 -3994 38 3994
rect 78 -3994 95 3994
rect 137 -3994 154 3994
rect 194 -3994 211 3994
rect 253 -3994 270 3994
rect 310 -3994 327 3994
rect 369 -3994 386 3994
rect 426 -3994 443 3994
rect 485 -3994 502 3994
rect 542 -3994 559 3994
rect 601 -3994 618 3994
rect 658 -3994 675 3994
rect 717 -3994 734 3994
rect 774 -3994 791 3994
rect 833 -3994 850 3994
rect 890 -3994 907 3994
rect 949 -3994 966 3994
rect 1006 -3994 1023 3994
rect 1065 -3994 1082 3994
rect 1122 -3994 1139 3994
rect 1181 -3994 1198 3994
rect 1238 -3994 1255 3994
rect 1297 -3994 1314 3994
rect 1354 -3994 1371 3994
rect 1413 -3994 1430 3994
rect 1470 -3994 1487 3994
rect 1529 -3994 1546 3994
rect 1586 -3994 1603 3994
rect 1645 -3994 1662 3994
<< poly >>
rect -1639 4000 -1609 4013
rect -1523 4000 -1493 4013
rect -1407 4000 -1377 4013
rect -1291 4000 -1261 4013
rect -1175 4000 -1145 4013
rect -1059 4000 -1029 4013
rect -943 4000 -913 4013
rect -827 4000 -797 4013
rect -711 4000 -681 4013
rect -595 4000 -565 4013
rect -479 4000 -449 4013
rect -363 4000 -333 4013
rect -247 4000 -217 4013
rect -131 4000 -101 4013
rect -15 4000 15 4013
rect 101 4000 131 4013
rect 217 4000 247 4013
rect 333 4000 363 4013
rect 449 4000 479 4013
rect 565 4000 595 4013
rect 681 4000 711 4013
rect 797 4000 827 4013
rect 913 4000 943 4013
rect 1029 4000 1059 4013
rect 1145 4000 1175 4013
rect 1261 4000 1291 4013
rect 1377 4000 1407 4013
rect 1493 4000 1523 4013
rect 1609 4000 1639 4013
rect -1639 -4013 -1609 -4000
rect -1523 -4013 -1493 -4000
rect -1407 -4013 -1377 -4000
rect -1291 -4013 -1261 -4000
rect -1175 -4013 -1145 -4000
rect -1059 -4013 -1029 -4000
rect -943 -4013 -913 -4000
rect -827 -4013 -797 -4000
rect -711 -4013 -681 -4000
rect -595 -4013 -565 -4000
rect -479 -4013 -449 -4000
rect -363 -4013 -333 -4000
rect -247 -4013 -217 -4000
rect -131 -4013 -101 -4000
rect -15 -4013 15 -4000
rect 101 -4013 131 -4000
rect 217 -4013 247 -4000
rect 333 -4013 363 -4000
rect 449 -4013 479 -4000
rect 565 -4013 595 -4000
rect 681 -4013 711 -4000
rect 797 -4013 827 -4000
rect 913 -4013 943 -4000
rect 1029 -4013 1059 -4000
rect 1145 -4013 1175 -4000
rect 1261 -4013 1291 -4000
rect 1377 -4013 1407 -4000
rect 1493 -4013 1523 -4000
rect 1609 -4013 1639 -4000
<< locali >>
rect -1662 3994 -1645 4002
rect -1662 -4002 -1645 -3994
rect -1603 3994 -1586 4002
rect -1603 -4002 -1586 -3994
rect -1546 3994 -1529 4002
rect -1546 -4002 -1529 -3994
rect -1487 3994 -1470 4002
rect -1487 -4002 -1470 -3994
rect -1430 3994 -1413 4002
rect -1430 -4002 -1413 -3994
rect -1371 3994 -1354 4002
rect -1371 -4002 -1354 -3994
rect -1314 3994 -1297 4002
rect -1314 -4002 -1297 -3994
rect -1255 3994 -1238 4002
rect -1255 -4002 -1238 -3994
rect -1198 3994 -1181 4002
rect -1198 -4002 -1181 -3994
rect -1139 3994 -1122 4002
rect -1139 -4002 -1122 -3994
rect -1082 3994 -1065 4002
rect -1082 -4002 -1065 -3994
rect -1023 3994 -1006 4002
rect -1023 -4002 -1006 -3994
rect -966 3994 -949 4002
rect -966 -4002 -949 -3994
rect -907 3994 -890 4002
rect -907 -4002 -890 -3994
rect -850 3994 -833 4002
rect -850 -4002 -833 -3994
rect -791 3994 -774 4002
rect -791 -4002 -774 -3994
rect -734 3994 -717 4002
rect -734 -4002 -717 -3994
rect -675 3994 -658 4002
rect -675 -4002 -658 -3994
rect -618 3994 -601 4002
rect -618 -4002 -601 -3994
rect -559 3994 -542 4002
rect -559 -4002 -542 -3994
rect -502 3994 -485 4002
rect -502 -4002 -485 -3994
rect -443 3994 -426 4002
rect -443 -4002 -426 -3994
rect -386 3994 -369 4002
rect -386 -4002 -369 -3994
rect -327 3994 -310 4002
rect -327 -4002 -310 -3994
rect -270 3994 -253 4002
rect -270 -4002 -253 -3994
rect -211 3994 -194 4002
rect -211 -4002 -194 -3994
rect -154 3994 -137 4002
rect -154 -4002 -137 -3994
rect -95 3994 -78 4002
rect -95 -4002 -78 -3994
rect -38 3994 -21 4002
rect -38 -4002 -21 -3994
rect 21 3994 38 4002
rect 21 -4002 38 -3994
rect 78 3994 95 4002
rect 78 -4002 95 -3994
rect 137 3994 154 4002
rect 137 -4002 154 -3994
rect 194 3994 211 4002
rect 194 -4002 211 -3994
rect 253 3994 270 4002
rect 253 -4002 270 -3994
rect 310 3994 327 4002
rect 310 -4002 327 -3994
rect 369 3994 386 4002
rect 369 -4002 386 -3994
rect 426 3994 443 4002
rect 426 -4002 443 -3994
rect 485 3994 502 4002
rect 485 -4002 502 -3994
rect 542 3994 559 4002
rect 542 -4002 559 -3994
rect 601 3994 618 4002
rect 601 -4002 618 -3994
rect 658 3994 675 4002
rect 658 -4002 675 -3994
rect 717 3994 734 4002
rect 717 -4002 734 -3994
rect 774 3994 791 4002
rect 774 -4002 791 -3994
rect 833 3994 850 4002
rect 833 -4002 850 -3994
rect 890 3994 907 4002
rect 890 -4002 907 -3994
rect 949 3994 966 4002
rect 949 -4002 966 -3994
rect 1006 3994 1023 4002
rect 1006 -4002 1023 -3994
rect 1065 3994 1082 4002
rect 1065 -4002 1082 -3994
rect 1122 3994 1139 4002
rect 1122 -4002 1139 -3994
rect 1181 3994 1198 4002
rect 1181 -4002 1198 -3994
rect 1238 3994 1255 4002
rect 1238 -4002 1255 -3994
rect 1297 3994 1314 4002
rect 1297 -4002 1314 -3994
rect 1354 3994 1371 4002
rect 1354 -4002 1371 -3994
rect 1413 3994 1430 4002
rect 1413 -4002 1430 -3994
rect 1470 3994 1487 4002
rect 1470 -4002 1487 -3994
rect 1529 3994 1546 4002
rect 1529 -4002 1546 -3994
rect 1586 3994 1603 4002
rect 1586 -4002 1603 -3994
rect 1645 3994 1662 4002
rect 1645 -4002 1662 -3994
<< viali >>
rect -1662 -3994 -1645 3994
rect -1603 -3994 -1586 3994
rect -1546 -3994 -1529 3994
rect -1487 -3994 -1470 3994
rect -1430 -3994 -1413 3994
rect -1371 -3994 -1354 3994
rect -1314 -3994 -1297 3994
rect -1255 -3994 -1238 3994
rect -1198 -3994 -1181 3994
rect -1139 -3994 -1122 3994
rect -1082 -3994 -1065 3994
rect -1023 -3994 -1006 3994
rect -966 -3994 -949 3994
rect -907 -3994 -890 3994
rect -850 -3994 -833 3994
rect -791 -3994 -774 3994
rect -734 -3994 -717 3994
rect -675 -3994 -658 3994
rect -618 -3994 -601 3994
rect -559 -3994 -542 3994
rect -502 -3994 -485 3994
rect -443 -3994 -426 3994
rect -386 -3994 -369 3994
rect -327 -3994 -310 3994
rect -270 -3994 -253 3994
rect -211 -3994 -194 3994
rect -154 -3994 -137 3994
rect -95 -3994 -78 3994
rect -38 -3994 -21 3994
rect 21 -3994 38 3994
rect 78 -3994 95 3994
rect 137 -3994 154 3994
rect 194 -3994 211 3994
rect 253 -3994 270 3994
rect 310 -3994 327 3994
rect 369 -3994 386 3994
rect 426 -3994 443 3994
rect 485 -3994 502 3994
rect 542 -3994 559 3994
rect 601 -3994 618 3994
rect 658 -3994 675 3994
rect 717 -3994 734 3994
rect 774 -3994 791 3994
rect 833 -3994 850 3994
rect 890 -3994 907 3994
rect 949 -3994 966 3994
rect 1006 -3994 1023 3994
rect 1065 -3994 1082 3994
rect 1122 -3994 1139 3994
rect 1181 -3994 1198 3994
rect 1238 -3994 1255 3994
rect 1297 -3994 1314 3994
rect 1354 -3994 1371 3994
rect 1413 -3994 1430 3994
rect 1470 -3994 1487 3994
rect 1529 -3994 1546 3994
rect 1586 -3994 1603 3994
rect 1645 -3994 1662 3994
<< metal1 >>
rect -1665 3994 -1642 4000
rect -1665 -3994 -1662 3994
rect -1645 -3994 -1642 3994
rect -1665 -4000 -1642 -3994
rect -1606 3994 -1583 4000
rect -1606 -3994 -1603 3994
rect -1586 -3994 -1583 3994
rect -1606 -4000 -1583 -3994
rect -1549 3994 -1526 4000
rect -1549 -3994 -1546 3994
rect -1529 -3994 -1526 3994
rect -1549 -4000 -1526 -3994
rect -1490 3994 -1467 4000
rect -1490 -3994 -1487 3994
rect -1470 -3994 -1467 3994
rect -1490 -4000 -1467 -3994
rect -1433 3994 -1410 4000
rect -1433 -3994 -1430 3994
rect -1413 -3994 -1410 3994
rect -1433 -4000 -1410 -3994
rect -1374 3994 -1351 4000
rect -1374 -3994 -1371 3994
rect -1354 -3994 -1351 3994
rect -1374 -4000 -1351 -3994
rect -1317 3994 -1294 4000
rect -1317 -3994 -1314 3994
rect -1297 -3994 -1294 3994
rect -1317 -4000 -1294 -3994
rect -1258 3994 -1235 4000
rect -1258 -3994 -1255 3994
rect -1238 -3994 -1235 3994
rect -1258 -4000 -1235 -3994
rect -1201 3994 -1178 4000
rect -1201 -3994 -1198 3994
rect -1181 -3994 -1178 3994
rect -1201 -4000 -1178 -3994
rect -1142 3994 -1119 4000
rect -1142 -3994 -1139 3994
rect -1122 -3994 -1119 3994
rect -1142 -4000 -1119 -3994
rect -1085 3994 -1062 4000
rect -1085 -3994 -1082 3994
rect -1065 -3994 -1062 3994
rect -1085 -4000 -1062 -3994
rect -1026 3994 -1003 4000
rect -1026 -3994 -1023 3994
rect -1006 -3994 -1003 3994
rect -1026 -4000 -1003 -3994
rect -969 3994 -946 4000
rect -969 -3994 -966 3994
rect -949 -3994 -946 3994
rect -969 -4000 -946 -3994
rect -910 3994 -887 4000
rect -910 -3994 -907 3994
rect -890 -3994 -887 3994
rect -910 -4000 -887 -3994
rect -853 3994 -830 4000
rect -853 -3994 -850 3994
rect -833 -3994 -830 3994
rect -853 -4000 -830 -3994
rect -794 3994 -771 4000
rect -794 -3994 -791 3994
rect -774 -3994 -771 3994
rect -794 -4000 -771 -3994
rect -737 3994 -714 4000
rect -737 -3994 -734 3994
rect -717 -3994 -714 3994
rect -737 -4000 -714 -3994
rect -678 3994 -655 4000
rect -678 -3994 -675 3994
rect -658 -3994 -655 3994
rect -678 -4000 -655 -3994
rect -621 3994 -598 4000
rect -621 -3994 -618 3994
rect -601 -3994 -598 3994
rect -621 -4000 -598 -3994
rect -562 3994 -539 4000
rect -562 -3994 -559 3994
rect -542 -3994 -539 3994
rect -562 -4000 -539 -3994
rect -505 3994 -482 4000
rect -505 -3994 -502 3994
rect -485 -3994 -482 3994
rect -505 -4000 -482 -3994
rect -446 3994 -423 4000
rect -446 -3994 -443 3994
rect -426 -3994 -423 3994
rect -446 -4000 -423 -3994
rect -389 3994 -366 4000
rect -389 -3994 -386 3994
rect -369 -3994 -366 3994
rect -389 -4000 -366 -3994
rect -330 3994 -307 4000
rect -330 -3994 -327 3994
rect -310 -3994 -307 3994
rect -330 -4000 -307 -3994
rect -273 3994 -250 4000
rect -273 -3994 -270 3994
rect -253 -3994 -250 3994
rect -273 -4000 -250 -3994
rect -214 3994 -191 4000
rect -214 -3994 -211 3994
rect -194 -3994 -191 3994
rect -214 -4000 -191 -3994
rect -157 3994 -134 4000
rect -157 -3994 -154 3994
rect -137 -3994 -134 3994
rect -157 -4000 -134 -3994
rect -98 3994 -75 4000
rect -98 -3994 -95 3994
rect -78 -3994 -75 3994
rect -98 -4000 -75 -3994
rect -41 3994 -18 4000
rect -41 -3994 -38 3994
rect -21 -3994 -18 3994
rect -41 -4000 -18 -3994
rect 18 3994 41 4000
rect 18 -3994 21 3994
rect 38 -3994 41 3994
rect 18 -4000 41 -3994
rect 75 3994 98 4000
rect 75 -3994 78 3994
rect 95 -3994 98 3994
rect 75 -4000 98 -3994
rect 134 3994 157 4000
rect 134 -3994 137 3994
rect 154 -3994 157 3994
rect 134 -4000 157 -3994
rect 191 3994 214 4000
rect 191 -3994 194 3994
rect 211 -3994 214 3994
rect 191 -4000 214 -3994
rect 250 3994 273 4000
rect 250 -3994 253 3994
rect 270 -3994 273 3994
rect 250 -4000 273 -3994
rect 307 3994 330 4000
rect 307 -3994 310 3994
rect 327 -3994 330 3994
rect 307 -4000 330 -3994
rect 366 3994 389 4000
rect 366 -3994 369 3994
rect 386 -3994 389 3994
rect 366 -4000 389 -3994
rect 423 3994 446 4000
rect 423 -3994 426 3994
rect 443 -3994 446 3994
rect 423 -4000 446 -3994
rect 482 3994 505 4000
rect 482 -3994 485 3994
rect 502 -3994 505 3994
rect 482 -4000 505 -3994
rect 539 3994 562 4000
rect 539 -3994 542 3994
rect 559 -3994 562 3994
rect 539 -4000 562 -3994
rect 598 3994 621 4000
rect 598 -3994 601 3994
rect 618 -3994 621 3994
rect 598 -4000 621 -3994
rect 655 3994 678 4000
rect 655 -3994 658 3994
rect 675 -3994 678 3994
rect 655 -4000 678 -3994
rect 714 3994 737 4000
rect 714 -3994 717 3994
rect 734 -3994 737 3994
rect 714 -4000 737 -3994
rect 771 3994 794 4000
rect 771 -3994 774 3994
rect 791 -3994 794 3994
rect 771 -4000 794 -3994
rect 830 3994 853 4000
rect 830 -3994 833 3994
rect 850 -3994 853 3994
rect 830 -4000 853 -3994
rect 887 3994 910 4000
rect 887 -3994 890 3994
rect 907 -3994 910 3994
rect 887 -4000 910 -3994
rect 946 3994 969 4000
rect 946 -3994 949 3994
rect 966 -3994 969 3994
rect 946 -4000 969 -3994
rect 1003 3994 1026 4000
rect 1003 -3994 1006 3994
rect 1023 -3994 1026 3994
rect 1003 -4000 1026 -3994
rect 1062 3994 1085 4000
rect 1062 -3994 1065 3994
rect 1082 -3994 1085 3994
rect 1062 -4000 1085 -3994
rect 1119 3994 1142 4000
rect 1119 -3994 1122 3994
rect 1139 -3994 1142 3994
rect 1119 -4000 1142 -3994
rect 1178 3994 1201 4000
rect 1178 -3994 1181 3994
rect 1198 -3994 1201 3994
rect 1178 -4000 1201 -3994
rect 1235 3994 1258 4000
rect 1235 -3994 1238 3994
rect 1255 -3994 1258 3994
rect 1235 -4000 1258 -3994
rect 1294 3994 1317 4000
rect 1294 -3994 1297 3994
rect 1314 -3994 1317 3994
rect 1294 -4000 1317 -3994
rect 1351 3994 1374 4000
rect 1351 -3994 1354 3994
rect 1371 -3994 1374 3994
rect 1351 -4000 1374 -3994
rect 1410 3994 1433 4000
rect 1410 -3994 1413 3994
rect 1430 -3994 1433 3994
rect 1410 -4000 1433 -3994
rect 1467 3994 1490 4000
rect 1467 -3994 1470 3994
rect 1487 -3994 1490 3994
rect 1467 -4000 1490 -3994
rect 1526 3994 1549 4000
rect 1526 -3994 1529 3994
rect 1546 -3994 1549 3994
rect 1526 -4000 1549 -3994
rect 1583 3994 1606 4000
rect 1583 -3994 1586 3994
rect 1603 -3994 1606 3994
rect 1583 -4000 1606 -3994
rect 1642 3994 1665 4000
rect 1642 -3994 1645 3994
rect 1662 -3994 1665 3994
rect 1642 -4000 1665 -3994
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 80 l 0.3 m 1 nf 29 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
