magic
tech sky130A
magscale 1 2
timestamp 1667395660
<< xpolycontact >>
rect -35 940 35 1372
rect -35 -1372 35 -940
<< xpolyres >>
rect -35 -940 35 940
<< viali >>
rect -19 957 19 1354
rect -19 -1354 19 -957
<< metal1 >>
rect -25 1354 25 1366
rect -25 957 -19 1354
rect 19 957 25 1354
rect -25 945 25 957
rect -25 -957 25 -945
rect -25 -1354 -19 -957
rect 19 -1354 25 -957
rect -25 -1366 25 -1354
<< res0p35 >>
rect -37 -942 37 942
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 9.4 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 54.789k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
