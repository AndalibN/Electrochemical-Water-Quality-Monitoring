magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -114 -376 114 376
<< nmos >>
rect -30 -350 30 350
<< ndiff >>
rect -88 323 -30 350
rect -88 289 -76 323
rect -42 289 -30 323
rect -88 255 -30 289
rect -88 221 -76 255
rect -42 221 -30 255
rect -88 187 -30 221
rect -88 153 -76 187
rect -42 153 -30 187
rect -88 119 -30 153
rect -88 85 -76 119
rect -42 85 -30 119
rect -88 51 -30 85
rect -88 17 -76 51
rect -42 17 -30 51
rect -88 -17 -30 17
rect -88 -51 -76 -17
rect -42 -51 -30 -17
rect -88 -85 -30 -51
rect -88 -119 -76 -85
rect -42 -119 -30 -85
rect -88 -153 -30 -119
rect -88 -187 -76 -153
rect -42 -187 -30 -153
rect -88 -221 -30 -187
rect -88 -255 -76 -221
rect -42 -255 -30 -221
rect -88 -289 -30 -255
rect -88 -323 -76 -289
rect -42 -323 -30 -289
rect -88 -350 -30 -323
rect 30 323 88 350
rect 30 289 42 323
rect 76 289 88 323
rect 30 255 88 289
rect 30 221 42 255
rect 76 221 88 255
rect 30 187 88 221
rect 30 153 42 187
rect 76 153 88 187
rect 30 119 88 153
rect 30 85 42 119
rect 76 85 88 119
rect 30 51 88 85
rect 30 17 42 51
rect 76 17 88 51
rect 30 -17 88 17
rect 30 -51 42 -17
rect 76 -51 88 -17
rect 30 -85 88 -51
rect 30 -119 42 -85
rect 76 -119 88 -85
rect 30 -153 88 -119
rect 30 -187 42 -153
rect 76 -187 88 -153
rect 30 -221 88 -187
rect 30 -255 42 -221
rect 76 -255 88 -221
rect 30 -289 88 -255
rect 30 -323 42 -289
rect 76 -323 88 -289
rect 30 -350 88 -323
<< ndiffc >>
rect -76 289 -42 323
rect -76 221 -42 255
rect -76 153 -42 187
rect -76 85 -42 119
rect -76 17 -42 51
rect -76 -51 -42 -17
rect -76 -119 -42 -85
rect -76 -187 -42 -153
rect -76 -255 -42 -221
rect -76 -323 -42 -289
rect 42 289 76 323
rect 42 221 76 255
rect 42 153 76 187
rect 42 85 76 119
rect 42 17 76 51
rect 42 -51 76 -17
rect 42 -119 76 -85
rect 42 -187 76 -153
rect 42 -255 76 -221
rect 42 -323 76 -289
<< poly >>
rect -30 350 30 376
rect -30 -376 30 -350
<< locali >>
rect -76 323 -42 354
rect -76 255 -42 271
rect -76 187 -42 199
rect -76 119 -42 127
rect -76 51 -42 55
rect -76 -55 -42 -51
rect -76 -127 -42 -119
rect -76 -199 -42 -187
rect -76 -271 -42 -255
rect -76 -354 -42 -323
rect 42 323 76 354
rect 42 255 76 271
rect 42 187 76 199
rect 42 119 76 127
rect 42 51 76 55
rect 42 -55 76 -51
rect 42 -127 76 -119
rect 42 -199 76 -187
rect 42 -271 76 -255
rect 42 -354 76 -323
<< viali >>
rect -76 289 -42 305
rect -76 271 -42 289
rect -76 221 -42 233
rect -76 199 -42 221
rect -76 153 -42 161
rect -76 127 -42 153
rect -76 85 -42 89
rect -76 55 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -55
rect -76 -89 -42 -85
rect -76 -153 -42 -127
rect -76 -161 -42 -153
rect -76 -221 -42 -199
rect -76 -233 -42 -221
rect -76 -289 -42 -271
rect -76 -305 -42 -289
rect 42 289 76 305
rect 42 271 76 289
rect 42 221 76 233
rect 42 199 76 221
rect 42 153 76 161
rect 42 127 76 153
rect 42 85 76 89
rect 42 55 76 85
rect 42 -17 76 17
rect 42 -85 76 -55
rect 42 -89 76 -85
rect 42 -153 76 -127
rect 42 -161 76 -153
rect 42 -221 76 -199
rect 42 -233 76 -221
rect 42 -289 76 -271
rect 42 -305 76 -289
<< metal1 >>
rect -82 305 -36 350
rect -82 271 -76 305
rect -42 271 -36 305
rect -82 233 -36 271
rect -82 199 -76 233
rect -42 199 -36 233
rect -82 161 -36 199
rect -82 127 -76 161
rect -42 127 -36 161
rect -82 89 -36 127
rect -82 55 -76 89
rect -42 55 -36 89
rect -82 17 -36 55
rect -82 -17 -76 17
rect -42 -17 -36 17
rect -82 -55 -36 -17
rect -82 -89 -76 -55
rect -42 -89 -36 -55
rect -82 -127 -36 -89
rect -82 -161 -76 -127
rect -42 -161 -36 -127
rect -82 -199 -36 -161
rect -82 -233 -76 -199
rect -42 -233 -36 -199
rect -82 -271 -36 -233
rect -82 -305 -76 -271
rect -42 -305 -36 -271
rect -82 -350 -36 -305
rect 36 305 82 350
rect 36 271 42 305
rect 76 271 82 305
rect 36 233 82 271
rect 36 199 42 233
rect 76 199 82 233
rect 36 161 82 199
rect 36 127 42 161
rect 76 127 82 161
rect 36 89 82 127
rect 36 55 42 89
rect 76 55 82 89
rect 36 17 82 55
rect 36 -17 42 17
rect 76 -17 82 17
rect 36 -55 82 -17
rect 36 -89 42 -55
rect 76 -89 82 -55
rect 36 -127 82 -89
rect 36 -161 42 -127
rect 76 -161 82 -127
rect 36 -199 82 -161
rect 36 -233 42 -199
rect 76 -233 82 -199
rect 36 -271 82 -233
rect 36 -305 42 -271
rect 76 -305 82 -271
rect 36 -350 82 -305
<< end >>
