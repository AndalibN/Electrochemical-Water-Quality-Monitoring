magic
tech sky130A
magscale 1 2
timestamp 1666404262
<< error_s >>
rect 1047 1423 1105 1429
rect 1293 1423 1351 1429
rect 1541 1423 1599 1429
rect 1047 1389 1059 1423
rect 1293 1389 1305 1423
rect 1541 1389 1553 1423
rect 1047 1383 1105 1389
rect 1293 1383 1351 1389
rect 1541 1383 1599 1389
rect 938 442 952 610
rect 1047 495 1105 501
rect 1293 495 1351 501
rect 1541 495 1599 501
rect 1047 461 1059 495
rect 1293 461 1305 495
rect 1541 461 1553 495
rect 1047 455 1105 461
rect 1293 455 1351 461
rect 1541 455 1599 461
rect 1106 294 1216 442
rect 1049 288 1216 294
rect 1049 284 1061 288
rect 1106 284 1216 288
rect 1048 240 1216 284
rect 1293 288 1351 294
rect 1511 288 1569 294
rect 1293 254 1305 288
rect 1511 254 1523 288
rect 1293 248 1351 254
rect 1511 248 1569 254
rect 1452 -184 1464 216
rect 1049 -222 1107 -216
rect 1293 -222 1351 -216
rect 1511 -222 1569 -216
rect 1049 -256 1061 -222
rect 1293 -256 1305 -222
rect 1511 -256 1523 -222
rect 1049 -262 1107 -256
rect 1293 -262 1351 -256
rect 1511 -262 1569 -256
<< nwell >>
rect 1046 452 1350 520
rect 1048 240 1106 452
<< poly >>
rect 1046 452 1350 520
rect 1048 302 1106 452
rect 1046 240 1352 302
use sky130_fd_pr__nfet_01v8_BYFWKT  XM2
timestamp 1666401230
transform 1 0 1540 0 1 16
box -88 -288 88 288
use sky130_fd_pr__pfet_01v8_6QH7WZ  XM3
timestamp 1666401230
transform 1 0 1570 0 1 942
box -124 -500 124 500
use sky130_fd_pr__pfet_01v8_6QH7WZ  XM4
timestamp 1666401230
transform 1 0 1322 0 1 942
box -124 -500 124 500
use sky130_fd_pr__nfet_01v8_BYFWKT  XM6
timestamp 1666401230
transform 1 0 1322 0 1 16
box -88 -288 88 288
use sky130_fd_pr__nfet_01v8_BYFWKT  sky130_fd_pr__nfet_01v8_BYFWKT_0
timestamp 1666401230
transform 1 0 1078 0 1 16
box -88 -288 88 288
use sky130_fd_pr__pfet_01v8_6QH7WZ  sky130_fd_pr__pfet_01v8_6QH7WZ_0
timestamp 1666401230
transform 1 0 1076 0 1 942
box -124 -500 124 500
<< end >>
