magic
timestamp 1668723770
<< checkpaint >>
rect 0 0 4985 2786
use sqr_ind_0p502n sqr_ind_0p502n_1
timestamp 1668723770
transform 1 0 -1415449 0 1 347524
box 1415449 -347524 1420434 -344739
<< end >>
