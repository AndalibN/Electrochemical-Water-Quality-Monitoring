magic
tech sky130A
magscale 1 2
timestamp 1666910672
<< nwell >>
rect -660 1420 550 1770
rect -660 810 550 1160
rect -660 200 550 550
rect -650 -410 560 -60
rect -650 -1020 560 -670
<< pmos >>
rect -473 1470 -433 1670
rect -375 1470 -335 1670
rect -277 1470 -237 1670
rect -179 1470 -139 1670
rect -81 1470 -41 1670
rect 17 1470 57 1670
rect 115 1470 155 1670
rect 213 1470 253 1670
rect 311 1470 351 1670
rect 409 1470 449 1670
rect -473 860 -433 1060
rect -375 860 -335 1060
rect -277 860 -237 1060
rect -179 860 -139 1060
rect -81 860 -41 1060
rect 17 860 57 1060
rect 115 860 155 1060
rect 213 860 253 1060
rect 311 860 351 1060
rect 409 860 449 1060
rect -473 250 -433 450
rect -375 250 -335 450
rect -277 250 -237 450
rect -179 250 -139 450
rect -81 250 -41 450
rect 17 250 57 450
rect 115 250 155 450
rect 213 250 253 450
rect 311 250 351 450
rect 409 250 449 450
rect -463 -360 -423 -160
rect -365 -360 -325 -160
rect -267 -360 -227 -160
rect -169 -360 -129 -160
rect -71 -360 -31 -160
rect 27 -360 67 -160
rect 125 -360 165 -160
rect 223 -360 263 -160
rect 321 -360 361 -160
rect 419 -360 459 -160
rect -463 -970 -423 -770
rect -365 -970 -325 -770
rect -267 -970 -227 -770
rect -169 -970 -129 -770
rect -71 -970 -31 -770
rect 27 -970 67 -770
rect 125 -970 165 -770
rect 223 -970 263 -770
rect 321 -970 361 -770
rect 419 -970 459 -770
<< pdiff >>
rect -531 1658 -473 1670
rect -531 1482 -519 1658
rect -485 1482 -473 1658
rect -531 1470 -473 1482
rect -433 1658 -375 1670
rect -433 1482 -421 1658
rect -387 1482 -375 1658
rect -433 1470 -375 1482
rect -335 1658 -277 1670
rect -335 1482 -323 1658
rect -289 1482 -277 1658
rect -335 1470 -277 1482
rect -237 1658 -179 1670
rect -237 1482 -225 1658
rect -191 1482 -179 1658
rect -237 1470 -179 1482
rect -139 1658 -81 1670
rect -139 1482 -127 1658
rect -93 1482 -81 1658
rect -139 1470 -81 1482
rect -41 1658 17 1670
rect -41 1482 -29 1658
rect 5 1482 17 1658
rect -41 1470 17 1482
rect 57 1658 115 1670
rect 57 1482 69 1658
rect 103 1482 115 1658
rect 57 1470 115 1482
rect 155 1658 213 1670
rect 155 1482 167 1658
rect 201 1482 213 1658
rect 155 1470 213 1482
rect 253 1658 311 1670
rect 253 1482 265 1658
rect 299 1482 311 1658
rect 253 1470 311 1482
rect 351 1658 409 1670
rect 351 1482 363 1658
rect 397 1482 409 1658
rect 351 1470 409 1482
rect 449 1658 507 1670
rect 449 1482 461 1658
rect 495 1482 507 1658
rect 449 1470 507 1482
rect -531 1048 -473 1060
rect -531 872 -519 1048
rect -485 872 -473 1048
rect -531 860 -473 872
rect -433 1048 -375 1060
rect -433 872 -421 1048
rect -387 872 -375 1048
rect -433 860 -375 872
rect -335 1048 -277 1060
rect -335 872 -323 1048
rect -289 872 -277 1048
rect -335 860 -277 872
rect -237 1048 -179 1060
rect -237 872 -225 1048
rect -191 872 -179 1048
rect -237 860 -179 872
rect -139 1048 -81 1060
rect -139 872 -127 1048
rect -93 872 -81 1048
rect -139 860 -81 872
rect -41 1048 17 1060
rect -41 872 -29 1048
rect 5 872 17 1048
rect -41 860 17 872
rect 57 1048 115 1060
rect 57 872 69 1048
rect 103 872 115 1048
rect 57 860 115 872
rect 155 1048 213 1060
rect 155 872 167 1048
rect 201 872 213 1048
rect 155 860 213 872
rect 253 1048 311 1060
rect 253 872 265 1048
rect 299 872 311 1048
rect 253 860 311 872
rect 351 1048 409 1060
rect 351 872 363 1048
rect 397 872 409 1048
rect 351 860 409 872
rect 449 1048 507 1060
rect 449 872 461 1048
rect 495 872 507 1048
rect 449 860 507 872
rect -531 438 -473 450
rect -531 262 -519 438
rect -485 262 -473 438
rect -531 250 -473 262
rect -433 438 -375 450
rect -433 262 -421 438
rect -387 262 -375 438
rect -433 250 -375 262
rect -335 438 -277 450
rect -335 262 -323 438
rect -289 262 -277 438
rect -335 250 -277 262
rect -237 438 -179 450
rect -237 262 -225 438
rect -191 262 -179 438
rect -237 250 -179 262
rect -139 438 -81 450
rect -139 262 -127 438
rect -93 262 -81 438
rect -139 250 -81 262
rect -41 438 17 450
rect -41 262 -29 438
rect 5 262 17 438
rect -41 250 17 262
rect 57 438 115 450
rect 57 262 69 438
rect 103 262 115 438
rect 57 250 115 262
rect 155 438 213 450
rect 155 262 167 438
rect 201 262 213 438
rect 155 250 213 262
rect 253 438 311 450
rect 253 262 265 438
rect 299 262 311 438
rect 253 250 311 262
rect 351 438 409 450
rect 351 262 363 438
rect 397 262 409 438
rect 351 250 409 262
rect 449 438 507 450
rect 449 262 461 438
rect 495 262 507 438
rect 449 250 507 262
rect -521 -172 -463 -160
rect -521 -348 -509 -172
rect -475 -348 -463 -172
rect -521 -360 -463 -348
rect -423 -172 -365 -160
rect -423 -348 -411 -172
rect -377 -348 -365 -172
rect -423 -360 -365 -348
rect -325 -172 -267 -160
rect -325 -348 -313 -172
rect -279 -348 -267 -172
rect -325 -360 -267 -348
rect -227 -172 -169 -160
rect -227 -348 -215 -172
rect -181 -348 -169 -172
rect -227 -360 -169 -348
rect -129 -172 -71 -160
rect -129 -348 -117 -172
rect -83 -348 -71 -172
rect -129 -360 -71 -348
rect -31 -172 27 -160
rect -31 -348 -19 -172
rect 15 -348 27 -172
rect -31 -360 27 -348
rect 67 -172 125 -160
rect 67 -348 79 -172
rect 113 -348 125 -172
rect 67 -360 125 -348
rect 165 -172 223 -160
rect 165 -348 177 -172
rect 211 -348 223 -172
rect 165 -360 223 -348
rect 263 -172 321 -160
rect 263 -348 275 -172
rect 309 -348 321 -172
rect 263 -360 321 -348
rect 361 -172 419 -160
rect 361 -348 373 -172
rect 407 -348 419 -172
rect 361 -360 419 -348
rect 459 -172 517 -160
rect 459 -348 471 -172
rect 505 -348 517 -172
rect 459 -360 517 -348
rect -521 -782 -463 -770
rect -521 -958 -509 -782
rect -475 -958 -463 -782
rect -521 -970 -463 -958
rect -423 -782 -365 -770
rect -423 -958 -411 -782
rect -377 -958 -365 -782
rect -423 -970 -365 -958
rect -325 -782 -267 -770
rect -325 -958 -313 -782
rect -279 -958 -267 -782
rect -325 -970 -267 -958
rect -227 -782 -169 -770
rect -227 -958 -215 -782
rect -181 -958 -169 -782
rect -227 -970 -169 -958
rect -129 -782 -71 -770
rect -129 -958 -117 -782
rect -83 -958 -71 -782
rect -129 -970 -71 -958
rect -31 -782 27 -770
rect -31 -958 -19 -782
rect 15 -958 27 -782
rect -31 -970 27 -958
rect 67 -782 125 -770
rect 67 -958 79 -782
rect 113 -958 125 -782
rect 67 -970 125 -958
rect 165 -782 223 -770
rect 165 -958 177 -782
rect 211 -958 223 -782
rect 165 -970 223 -958
rect 263 -782 321 -770
rect 263 -958 275 -782
rect 309 -958 321 -782
rect 263 -970 321 -958
rect 361 -782 419 -770
rect 361 -958 373 -782
rect 407 -958 419 -782
rect 361 -970 419 -958
rect 459 -782 517 -770
rect 459 -958 471 -782
rect 505 -958 517 -782
rect 459 -970 517 -958
<< pdiffc >>
rect -519 1482 -485 1658
rect -421 1482 -387 1658
rect -323 1482 -289 1658
rect -225 1482 -191 1658
rect -127 1482 -93 1658
rect -29 1482 5 1658
rect 69 1482 103 1658
rect 167 1482 201 1658
rect 265 1482 299 1658
rect 363 1482 397 1658
rect 461 1482 495 1658
rect -519 872 -485 1048
rect -421 872 -387 1048
rect -323 872 -289 1048
rect -225 872 -191 1048
rect -127 872 -93 1048
rect -29 872 5 1048
rect 69 872 103 1048
rect 167 872 201 1048
rect 265 872 299 1048
rect 363 872 397 1048
rect 461 872 495 1048
rect -519 262 -485 438
rect -421 262 -387 438
rect -323 262 -289 438
rect -225 262 -191 438
rect -127 262 -93 438
rect -29 262 5 438
rect 69 262 103 438
rect 167 262 201 438
rect 265 262 299 438
rect 363 262 397 438
rect 461 262 495 438
rect -509 -348 -475 -172
rect -411 -348 -377 -172
rect -313 -348 -279 -172
rect -215 -348 -181 -172
rect -117 -348 -83 -172
rect -19 -348 15 -172
rect 79 -348 113 -172
rect 177 -348 211 -172
rect 275 -348 309 -172
rect 373 -348 407 -172
rect 471 -348 505 -172
rect -509 -958 -475 -782
rect -411 -958 -377 -782
rect -313 -958 -279 -782
rect -215 -958 -181 -782
rect -117 -958 -83 -782
rect -19 -958 15 -782
rect 79 -958 113 -782
rect 177 -958 211 -782
rect 275 -958 309 -782
rect 373 -958 407 -782
rect 471 -958 505 -782
<< poly >>
rect -640 1730 -550 1750
rect -640 1715 450 1730
rect -640 1475 -615 1715
rect -580 1690 450 1715
rect -580 1475 -550 1690
rect -473 1670 -433 1690
rect -375 1670 -335 1690
rect -277 1670 -237 1690
rect -179 1670 -139 1690
rect -81 1670 -41 1690
rect 17 1670 57 1690
rect 115 1670 155 1690
rect 213 1670 253 1690
rect 311 1670 351 1690
rect 409 1670 449 1690
rect -640 1440 -550 1475
rect -473 1442 -433 1470
rect -375 1444 -335 1470
rect -277 1442 -237 1470
rect -179 1444 -139 1470
rect -81 1442 -41 1470
rect 17 1444 57 1470
rect 115 1442 155 1470
rect 213 1444 253 1470
rect 311 1442 351 1470
rect 409 1444 449 1470
rect -640 1120 -550 1140
rect -640 1105 450 1120
rect -640 865 -615 1105
rect -580 1080 450 1105
rect -580 865 -550 1080
rect -473 1060 -433 1080
rect -375 1060 -335 1080
rect -277 1060 -237 1080
rect -179 1060 -139 1080
rect -81 1060 -41 1080
rect 17 1060 57 1080
rect 115 1060 155 1080
rect 213 1060 253 1080
rect 311 1060 351 1080
rect 409 1060 449 1080
rect -640 830 -550 865
rect -473 832 -433 860
rect -375 834 -335 860
rect -277 832 -237 860
rect -179 834 -139 860
rect -81 832 -41 860
rect 17 834 57 860
rect 115 832 155 860
rect 213 834 253 860
rect 311 832 351 860
rect 409 834 449 860
rect -640 510 -550 530
rect -640 495 450 510
rect -640 255 -615 495
rect -580 470 450 495
rect -580 255 -550 470
rect -473 450 -433 470
rect -375 450 -335 470
rect -277 450 -237 470
rect -179 450 -139 470
rect -81 450 -41 470
rect 17 450 57 470
rect 115 450 155 470
rect 213 450 253 470
rect 311 450 351 470
rect 409 450 449 470
rect -640 220 -550 255
rect -473 222 -433 250
rect -375 224 -335 250
rect -277 222 -237 250
rect -179 224 -139 250
rect -81 222 -41 250
rect 17 224 57 250
rect 115 222 155 250
rect 213 224 253 250
rect 311 222 351 250
rect 409 224 449 250
rect -630 -100 -540 -80
rect -630 -115 460 -100
rect -630 -355 -605 -115
rect -570 -140 460 -115
rect -570 -355 -540 -140
rect -463 -160 -423 -140
rect -365 -160 -325 -140
rect -267 -160 -227 -140
rect -169 -160 -129 -140
rect -71 -160 -31 -140
rect 27 -160 67 -140
rect 125 -160 165 -140
rect 223 -160 263 -140
rect 321 -160 361 -140
rect 419 -160 459 -140
rect -630 -390 -540 -355
rect -463 -388 -423 -360
rect -365 -386 -325 -360
rect -267 -388 -227 -360
rect -169 -386 -129 -360
rect -71 -388 -31 -360
rect 27 -386 67 -360
rect 125 -388 165 -360
rect 223 -386 263 -360
rect 321 -388 361 -360
rect 419 -386 459 -360
rect -630 -710 -540 -690
rect -630 -725 460 -710
rect -630 -965 -605 -725
rect -570 -750 460 -725
rect -570 -965 -540 -750
rect -463 -770 -423 -750
rect -365 -770 -325 -750
rect -267 -770 -227 -750
rect -169 -770 -129 -750
rect -71 -770 -31 -750
rect 27 -770 67 -750
rect 125 -770 165 -750
rect 223 -770 263 -750
rect 321 -770 361 -750
rect 419 -770 459 -750
rect -630 -1000 -540 -965
rect -463 -998 -423 -970
rect -365 -996 -325 -970
rect -267 -998 -227 -970
rect -169 -996 -129 -970
rect -71 -998 -31 -970
rect 27 -996 67 -970
rect 125 -998 165 -970
rect 223 -996 263 -970
rect 321 -998 361 -970
rect 419 -996 459 -970
<< polycont >>
rect -615 1475 -580 1715
rect -615 865 -580 1105
rect -615 255 -580 495
rect -605 -355 -570 -115
rect -605 -965 -570 -725
<< locali >>
rect -630 1715 -560 1740
rect -630 1475 -615 1715
rect -580 1475 -560 1715
rect -630 1450 -560 1475
rect -519 1658 -485 1674
rect -519 1466 -485 1482
rect -421 1658 -387 1674
rect -421 1466 -387 1482
rect -323 1658 -289 1674
rect -323 1466 -289 1482
rect -225 1658 -191 1674
rect -225 1466 -191 1482
rect -127 1658 -93 1674
rect -127 1466 -93 1482
rect -29 1658 5 1674
rect -29 1466 5 1482
rect 69 1658 103 1674
rect 69 1466 103 1482
rect 167 1658 201 1674
rect 167 1466 201 1482
rect 265 1658 299 1674
rect 265 1466 299 1482
rect 363 1658 397 1674
rect 363 1466 397 1482
rect 461 1658 495 1674
rect 461 1466 495 1482
rect -630 1105 -560 1130
rect -630 865 -615 1105
rect -580 865 -560 1105
rect -630 840 -560 865
rect -519 1048 -485 1064
rect -519 856 -485 872
rect -421 1048 -387 1064
rect -421 856 -387 872
rect -323 1048 -289 1064
rect -323 856 -289 872
rect -225 1048 -191 1064
rect -225 856 -191 872
rect -127 1048 -93 1064
rect -127 856 -93 872
rect -29 1048 5 1064
rect -29 856 5 872
rect 69 1048 103 1064
rect 69 856 103 872
rect 167 1048 201 1064
rect 167 856 201 872
rect 265 1048 299 1064
rect 265 856 299 872
rect 363 1048 397 1064
rect 363 856 397 872
rect 461 1048 495 1064
rect 461 856 495 872
rect -630 495 -560 520
rect -630 255 -615 495
rect -580 255 -560 495
rect -630 230 -560 255
rect -519 438 -485 454
rect -519 246 -485 262
rect -421 438 -387 454
rect -421 246 -387 262
rect -323 438 -289 454
rect -323 246 -289 262
rect -225 438 -191 454
rect -225 246 -191 262
rect -127 438 -93 454
rect -127 246 -93 262
rect -29 438 5 454
rect -29 246 5 262
rect 69 438 103 454
rect 69 246 103 262
rect 167 438 201 454
rect 167 246 201 262
rect 265 438 299 454
rect 265 246 299 262
rect 363 438 397 454
rect 363 246 397 262
rect 461 438 495 454
rect 461 246 495 262
rect -620 -115 -550 -90
rect -620 -355 -605 -115
rect -570 -355 -550 -115
rect -620 -380 -550 -355
rect -509 -172 -475 -156
rect -509 -364 -475 -348
rect -411 -172 -377 -156
rect -411 -364 -377 -348
rect -313 -172 -279 -156
rect -313 -364 -279 -348
rect -215 -172 -181 -156
rect -215 -364 -181 -348
rect -117 -172 -83 -156
rect -117 -364 -83 -348
rect -19 -172 15 -156
rect -19 -364 15 -348
rect 79 -172 113 -156
rect 79 -364 113 -348
rect 177 -172 211 -156
rect 177 -364 211 -348
rect 275 -172 309 -156
rect 275 -364 309 -348
rect 373 -172 407 -156
rect 373 -364 407 -348
rect 471 -172 505 -156
rect 471 -364 505 -348
rect -620 -725 -550 -700
rect -620 -965 -605 -725
rect -570 -965 -550 -725
rect -620 -990 -550 -965
rect -509 -782 -475 -766
rect -509 -974 -475 -958
rect -411 -782 -377 -766
rect -411 -974 -377 -958
rect -313 -782 -279 -766
rect -313 -974 -279 -958
rect -215 -782 -181 -766
rect -215 -974 -181 -958
rect -117 -782 -83 -766
rect -117 -974 -83 -958
rect -19 -782 15 -766
rect -19 -974 15 -958
rect 79 -782 113 -766
rect 79 -974 113 -958
rect 177 -782 211 -766
rect 177 -974 211 -958
rect 275 -782 309 -766
rect 275 -974 309 -958
rect 373 -782 407 -766
rect 373 -974 407 -958
rect 471 -782 505 -766
rect 471 -974 505 -958
<< viali >>
rect -615 1475 -580 1715
rect -519 1482 -485 1658
rect -421 1482 -387 1658
rect -323 1482 -289 1658
rect -225 1482 -191 1658
rect -127 1482 -93 1658
rect -29 1482 5 1658
rect 69 1482 103 1658
rect 167 1482 201 1658
rect 265 1482 299 1658
rect 363 1482 397 1658
rect 461 1482 495 1658
rect -615 865 -580 1105
rect -519 872 -485 1048
rect -421 872 -387 1048
rect -323 872 -289 1048
rect -225 872 -191 1048
rect -127 872 -93 1048
rect -29 872 5 1048
rect 69 872 103 1048
rect 167 872 201 1048
rect 265 872 299 1048
rect 363 872 397 1048
rect 461 872 495 1048
rect -615 255 -580 495
rect -519 262 -485 438
rect -421 262 -387 438
rect -323 262 -289 438
rect -225 262 -191 438
rect -127 262 -93 438
rect -29 262 5 438
rect 69 262 103 438
rect 167 262 201 438
rect 265 262 299 438
rect 363 262 397 438
rect 461 262 495 438
rect -605 -355 -570 -115
rect -509 -348 -475 -172
rect -411 -348 -377 -172
rect -313 -348 -279 -172
rect -215 -348 -181 -172
rect -117 -348 -83 -172
rect -19 -348 15 -172
rect 79 -348 113 -172
rect 177 -348 211 -172
rect 275 -348 309 -172
rect 373 -348 407 -172
rect 471 -348 505 -172
rect -605 -965 -570 -725
rect -509 -958 -475 -782
rect -411 -958 -377 -782
rect -313 -958 -279 -782
rect -215 -958 -181 -782
rect -117 -958 -83 -782
rect -19 -958 15 -782
rect 79 -958 113 -782
rect 177 -958 211 -782
rect 275 -958 309 -782
rect 373 -958 407 -782
rect 471 -958 505 -782
<< metal1 >>
rect -625 1715 -565 1730
rect -625 1475 -615 1715
rect -580 1475 -565 1715
rect -625 1460 -565 1475
rect -525 1658 -479 1670
rect -525 1482 -519 1658
rect -485 1482 -479 1658
rect -525 1470 -479 1482
rect -427 1658 -381 1670
rect -427 1482 -421 1658
rect -387 1482 -381 1658
rect -427 1470 -381 1482
rect -329 1658 -283 1670
rect -329 1482 -323 1658
rect -289 1482 -283 1658
rect -329 1470 -283 1482
rect -231 1658 -185 1670
rect -231 1482 -225 1658
rect -191 1482 -185 1658
rect -231 1470 -185 1482
rect -133 1658 -87 1670
rect -133 1482 -127 1658
rect -93 1482 -87 1658
rect -133 1470 -87 1482
rect -35 1658 11 1670
rect -35 1482 -29 1658
rect 5 1482 11 1658
rect -35 1470 11 1482
rect 63 1658 109 1670
rect 63 1482 69 1658
rect 103 1482 109 1658
rect 63 1470 109 1482
rect 161 1658 207 1670
rect 161 1482 167 1658
rect 201 1482 207 1658
rect 161 1470 207 1482
rect 259 1658 305 1670
rect 259 1482 265 1658
rect 299 1482 305 1658
rect 259 1470 305 1482
rect 357 1658 403 1670
rect 357 1482 363 1658
rect 397 1482 403 1658
rect 357 1470 403 1482
rect 455 1658 501 1670
rect 455 1482 461 1658
rect 495 1482 501 1658
rect 455 1470 501 1482
rect -625 1105 -565 1120
rect -625 865 -615 1105
rect -580 865 -565 1105
rect -625 850 -565 865
rect -525 1048 -479 1060
rect -525 872 -519 1048
rect -485 872 -479 1048
rect -525 860 -479 872
rect -427 1048 -381 1060
rect -427 872 -421 1048
rect -387 872 -381 1048
rect -427 860 -381 872
rect -329 1048 -283 1060
rect -329 872 -323 1048
rect -289 872 -283 1048
rect -329 860 -283 872
rect -231 1048 -185 1060
rect -231 872 -225 1048
rect -191 872 -185 1048
rect -231 860 -185 872
rect -133 1048 -87 1060
rect -133 872 -127 1048
rect -93 872 -87 1048
rect -133 860 -87 872
rect -35 1048 11 1060
rect -35 872 -29 1048
rect 5 872 11 1048
rect -35 860 11 872
rect 63 1048 109 1060
rect 63 872 69 1048
rect 103 872 109 1048
rect 63 860 109 872
rect 161 1048 207 1060
rect 161 872 167 1048
rect 201 872 207 1048
rect 161 860 207 872
rect 259 1048 305 1060
rect 259 872 265 1048
rect 299 872 305 1048
rect 259 860 305 872
rect 357 1048 403 1060
rect 357 872 363 1048
rect 397 872 403 1048
rect 357 860 403 872
rect 455 1048 501 1060
rect 455 872 461 1048
rect 495 872 501 1048
rect 455 860 501 872
rect -625 495 -565 510
rect -625 255 -615 495
rect -580 255 -565 495
rect -625 240 -565 255
rect -525 438 -479 450
rect -525 262 -519 438
rect -485 262 -479 438
rect -525 250 -479 262
rect -427 438 -381 450
rect -427 262 -421 438
rect -387 262 -381 438
rect -427 250 -381 262
rect -329 438 -283 450
rect -329 262 -323 438
rect -289 262 -283 438
rect -329 250 -283 262
rect -231 438 -185 450
rect -231 262 -225 438
rect -191 262 -185 438
rect -231 250 -185 262
rect -133 438 -87 450
rect -133 262 -127 438
rect -93 262 -87 438
rect -133 250 -87 262
rect -35 438 11 450
rect -35 262 -29 438
rect 5 262 11 438
rect -35 250 11 262
rect 63 438 109 450
rect 63 262 69 438
rect 103 262 109 438
rect 63 250 109 262
rect 161 438 207 450
rect 161 262 167 438
rect 201 262 207 438
rect 161 250 207 262
rect 259 438 305 450
rect 259 262 265 438
rect 299 262 305 438
rect 259 250 305 262
rect 357 438 403 450
rect 357 262 363 438
rect 397 262 403 438
rect 357 250 403 262
rect 455 438 501 450
rect 455 262 461 438
rect 495 262 501 438
rect 455 250 501 262
rect -615 -115 -555 -100
rect -615 -355 -605 -115
rect -570 -355 -555 -115
rect -615 -370 -555 -355
rect -515 -172 -469 -160
rect -515 -348 -509 -172
rect -475 -348 -469 -172
rect -515 -360 -469 -348
rect -417 -172 -371 -160
rect -417 -348 -411 -172
rect -377 -348 -371 -172
rect -417 -360 -371 -348
rect -319 -172 -273 -160
rect -319 -348 -313 -172
rect -279 -348 -273 -172
rect -319 -360 -273 -348
rect -221 -172 -175 -160
rect -221 -348 -215 -172
rect -181 -348 -175 -172
rect -221 -360 -175 -348
rect -123 -172 -77 -160
rect -123 -348 -117 -172
rect -83 -348 -77 -172
rect -123 -360 -77 -348
rect -25 -172 21 -160
rect -25 -348 -19 -172
rect 15 -348 21 -172
rect -25 -360 21 -348
rect 73 -172 119 -160
rect 73 -348 79 -172
rect 113 -348 119 -172
rect 73 -360 119 -348
rect 171 -172 217 -160
rect 171 -348 177 -172
rect 211 -348 217 -172
rect 171 -360 217 -348
rect 269 -172 315 -160
rect 269 -348 275 -172
rect 309 -348 315 -172
rect 269 -360 315 -348
rect 367 -172 413 -160
rect 367 -348 373 -172
rect 407 -348 413 -172
rect 367 -360 413 -348
rect 465 -172 511 -160
rect 465 -348 471 -172
rect 505 -348 511 -172
rect 465 -360 511 -348
rect -615 -725 -555 -710
rect -615 -965 -605 -725
rect -570 -965 -555 -725
rect -615 -980 -555 -965
rect -515 -782 -469 -770
rect -515 -958 -509 -782
rect -475 -958 -469 -782
rect -515 -970 -469 -958
rect -417 -782 -371 -770
rect -417 -958 -411 -782
rect -377 -958 -371 -782
rect -417 -970 -371 -958
rect -319 -782 -273 -770
rect -319 -958 -313 -782
rect -279 -958 -273 -782
rect -319 -970 -273 -958
rect -221 -782 -175 -770
rect -221 -958 -215 -782
rect -181 -958 -175 -782
rect -221 -970 -175 -958
rect -123 -782 -77 -770
rect -123 -958 -117 -782
rect -83 -958 -77 -782
rect -123 -970 -77 -958
rect -25 -782 21 -770
rect -25 -958 -19 -782
rect 15 -958 21 -782
rect -25 -970 21 -958
rect 73 -782 119 -770
rect 73 -958 79 -782
rect 113 -958 119 -782
rect 73 -970 119 -958
rect 171 -782 217 -770
rect 171 -958 177 -782
rect 211 -958 217 -782
rect 171 -970 217 -958
rect 269 -782 315 -770
rect 269 -958 275 -782
rect 309 -958 315 -782
rect 269 -970 315 -958
rect 367 -782 413 -770
rect 367 -958 373 -782
rect 407 -958 413 -782
rect 367 -970 413 -958
rect 465 -782 511 -770
rect 465 -958 471 -782
rect 505 -958 511 -782
rect 465 -970 511 -958
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.2 m 5 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
