magic
tech sky130A
magscale 1 2
timestamp 1667053331
<< nwell >>
rect -194 -754 194 788
<< pmos >>
rect -100 -654 100 726
<< pdiff >>
rect -158 714 -100 726
rect -158 -642 -146 714
rect -112 -642 -100 714
rect -158 -654 -100 -642
rect 100 714 158 726
rect 100 -642 112 714
rect 146 -642 158 714
rect 100 -654 158 -642
<< pdiffc >>
rect -146 -642 -112 714
rect 112 -642 146 714
<< poly >>
rect -100 726 100 752
rect -100 -701 100 -654
rect -100 -735 -84 -701
rect 84 -735 100 -701
rect -100 -751 100 -735
<< polycont >>
rect -84 -735 84 -701
<< locali >>
rect -146 714 -112 730
rect -146 -658 -112 -642
rect 112 714 146 730
rect 112 -658 146 -642
rect -100 -735 -84 -701
rect 84 -735 100 -701
<< viali >>
rect -146 -642 -112 714
rect 112 -642 146 714
rect -84 -735 84 -701
<< metal1 >>
rect -152 714 -106 726
rect -152 -642 -146 714
rect -112 -642 -106 714
rect -152 -654 -106 -642
rect 106 714 152 726
rect 106 -642 112 714
rect 146 -642 152 714
rect 106 -654 152 -642
rect -96 -701 96 -695
rect -96 -735 -84 -701
rect 84 -735 96 -701
rect -96 -741 96 -735
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.9 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
