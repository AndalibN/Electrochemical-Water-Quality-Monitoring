magic
tech sky130A
magscale 1 2
timestamp 1667444078
<< nmos >>
rect -429 -2769 -29 2831
rect 29 -2769 429 2831
<< ndiff >>
rect -487 2819 -429 2831
rect -487 -2757 -475 2819
rect -441 -2757 -429 2819
rect -487 -2769 -429 -2757
rect -29 2819 29 2831
rect -29 -2757 -17 2819
rect 17 -2757 29 2819
rect -29 -2769 29 -2757
rect 429 2819 487 2831
rect 429 -2757 441 2819
rect 475 -2757 487 2819
rect 429 -2769 487 -2757
<< ndiffc >>
rect -475 -2757 -441 2819
rect -17 -2757 17 2819
rect 441 -2757 475 2819
<< poly >>
rect -429 2831 -29 2857
rect 29 2831 429 2857
rect -429 -2807 -29 -2769
rect -429 -2841 -413 -2807
rect -45 -2841 -29 -2807
rect -429 -2857 -29 -2841
rect 29 -2807 429 -2769
rect 29 -2841 45 -2807
rect 413 -2841 429 -2807
rect 29 -2857 429 -2841
<< polycont >>
rect -413 -2841 -45 -2807
rect 45 -2841 413 -2807
<< locali >>
rect -475 2819 -441 2835
rect -475 -2773 -441 -2757
rect -17 2819 17 2835
rect -17 -2773 17 -2757
rect 441 2819 475 2835
rect 441 -2773 475 -2757
rect -429 -2841 -413 -2807
rect -45 -2841 -29 -2807
rect 29 -2841 45 -2807
rect 413 -2841 429 -2807
<< viali >>
rect -475 -2757 -441 2819
rect -17 -2757 17 2819
rect 441 -2757 475 2819
rect -413 -2841 -45 -2807
rect 45 -2841 413 -2807
<< metal1 >>
rect -481 2819 -435 2831
rect -481 -2757 -475 2819
rect -441 -2757 -435 2819
rect -481 -2769 -435 -2757
rect -23 2819 23 2831
rect -23 -2757 -17 2819
rect 17 -2757 23 2819
rect -23 -2769 23 -2757
rect 435 2819 481 2831
rect 435 -2757 441 2819
rect 475 -2757 481 2819
rect 435 -2769 481 -2757
rect -425 -2807 -33 -2801
rect -425 -2841 -413 -2807
rect -45 -2841 -33 -2807
rect -425 -2847 -33 -2841
rect 33 -2807 425 -2801
rect 33 -2841 45 -2807
rect 413 -2841 425 -2807
rect 33 -2847 425 -2841
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 28.0 l 2.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
