magic
tech sky130A
magscale 1 2
timestamp 1666815934
<< metal3 >>
rect -1150 1072 1149 1100
rect -1150 -1072 1065 1072
rect 1129 -1072 1149 1072
rect -1150 -1100 1149 -1072
<< via3 >>
rect 1065 -1072 1129 1072
<< mimcap >>
rect -1050 960 950 1000
rect -1050 -960 -1010 960
rect 910 -960 950 960
rect -1050 -1000 950 -960
<< mimcapcontact >>
rect -1010 -960 910 960
<< metal4 >>
rect 1049 1072 1145 1088
rect -1011 960 911 961
rect -1011 -960 -1010 960
rect 910 -960 911 960
rect -1011 -961 911 -960
rect 1049 -1072 1065 1072
rect 1129 -1072 1145 1072
rect 1049 -1088 1145 -1072
<< properties >>
string FIXED_BBOX -1150 -1100 1050 1100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 10.0 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
