magic
tech sky130A
magscale 1 2
timestamp 1667951016
<< error_p >>
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect -29 -347 29 -341
<< nmos >>
rect -30 -269 30 331
<< ndiff >>
rect -88 319 -30 331
rect -88 -257 -76 319
rect -42 -257 -30 319
rect -88 -269 -30 -257
rect 30 319 88 331
rect 30 -257 42 319
rect 76 -257 88 319
rect 30 -269 88 -257
<< ndiffc >>
rect -76 -257 -42 319
rect 42 -257 76 319
<< poly >>
rect -30 331 30 357
rect -30 -291 30 -269
rect -33 -307 33 -291
rect -33 -341 -17 -307
rect 17 -341 33 -307
rect -33 -357 33 -341
<< polycont >>
rect -17 -341 17 -307
<< locali >>
rect -76 319 -42 335
rect -76 -273 -42 -257
rect 42 319 76 335
rect 42 -273 76 -257
rect -33 -341 -17 -307
rect 17 -341 33 -307
<< viali >>
rect -76 -257 -42 319
rect 42 -257 76 319
rect -17 -341 17 -307
<< metal1 >>
rect -82 319 -36 331
rect -82 -257 -76 319
rect -42 -257 -36 319
rect -82 -269 -36 -257
rect 36 319 82 331
rect 36 -257 42 319
rect 76 -257 82 319
rect 36 -269 82 -257
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect 17 -341 29 -307
rect -29 -347 29 -341
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
