magic
tech sky130A
magscale 1 2
timestamp 1668017421
<< nmos >>
rect -30 -569 30 631
<< ndiff >>
rect -88 619 -30 631
rect -88 -557 -76 619
rect -42 -557 -30 619
rect -88 -569 -30 -557
rect 30 619 88 631
rect 30 -557 42 619
rect 76 -557 88 619
rect 30 -569 88 -557
<< ndiffc >>
rect -76 -557 -42 619
rect 42 -557 76 619
<< poly >>
rect -30 631 30 657
rect -30 -591 30 -569
rect -33 -607 33 -591
rect -33 -641 -17 -607
rect 17 -641 33 -607
rect -33 -657 33 -641
<< polycont >>
rect -17 -641 17 -607
<< locali >>
rect -76 619 -42 635
rect -76 -573 -42 -557
rect 42 619 76 635
rect 42 -573 76 -557
rect -33 -641 -17 -607
rect 17 -641 33 -607
<< viali >>
rect -76 -557 -42 619
rect 42 -557 76 619
rect -17 -641 17 -607
<< metal1 >>
rect -82 619 -36 631
rect -82 -557 -76 619
rect -42 -557 -36 619
rect -82 -569 -36 -557
rect 36 619 82 631
rect 36 -557 42 619
rect 76 -557 82 619
rect 36 -569 82 -557
rect -29 -607 29 -601
rect -29 -641 -17 -607
rect 17 -641 29 -607
rect -29 -647 29 -641
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
