magic
tech sky130A
magscale 1 2
timestamp 1668223520
<< error_p >>
rect -88 1041 -30 1047
rect 30 1041 88 1047
rect -88 1007 -76 1041
rect 30 1007 42 1041
rect -88 1001 -30 1007
rect 30 1001 88 1007
rect -88 -1007 -30 -1001
rect 30 -1007 88 -1001
rect -88 -1041 -76 -1007
rect 30 -1041 42 -1007
rect -88 -1047 -30 -1041
rect 30 -1047 88 -1041
<< nwell >>
rect -183 -1060 183 1060
<< pmos >>
rect -89 -960 -29 960
rect 29 -960 89 960
<< pdiff >>
rect -147 948 -89 960
rect -147 -948 -135 948
rect -101 -948 -89 948
rect -147 -960 -89 -948
rect -29 948 29 960
rect -29 -948 -17 948
rect 17 -948 29 948
rect -29 -960 29 -948
rect 89 948 147 960
rect 89 -948 101 948
rect 135 -948 147 948
rect 89 -960 147 -948
<< pdiffc >>
rect -135 -948 -101 948
rect -17 -948 17 948
rect 101 -948 135 948
<< poly >>
rect -92 1041 -26 1057
rect -92 1007 -76 1041
rect -42 1007 -26 1041
rect -92 991 -26 1007
rect 26 1041 92 1057
rect 26 1007 42 1041
rect 76 1007 92 1041
rect 26 991 92 1007
rect -89 960 -29 991
rect 29 960 89 991
rect -89 -991 -29 -960
rect 29 -991 89 -960
rect -92 -1007 -26 -991
rect -92 -1041 -76 -1007
rect -42 -1041 -26 -1007
rect -92 -1057 -26 -1041
rect 26 -1007 92 -991
rect 26 -1041 42 -1007
rect 76 -1041 92 -1007
rect 26 -1057 92 -1041
<< polycont >>
rect -76 1007 -42 1041
rect 42 1007 76 1041
rect -76 -1041 -42 -1007
rect 42 -1041 76 -1007
<< locali >>
rect -92 1007 -76 1041
rect -42 1007 -26 1041
rect 26 1007 42 1041
rect 76 1007 92 1041
rect -135 948 -101 964
rect -135 -964 -101 -948
rect -17 948 17 964
rect -17 -964 17 -948
rect 101 948 135 964
rect 101 -964 135 -948
rect -92 -1041 -76 -1007
rect -42 -1041 -26 -1007
rect 26 -1041 42 -1007
rect 76 -1041 92 -1007
<< viali >>
rect -76 1007 -42 1041
rect 42 1007 76 1041
rect -135 -948 -101 948
rect -17 -948 17 948
rect 101 -948 135 948
rect -76 -1041 -42 -1007
rect 42 -1041 76 -1007
<< metal1 >>
rect -88 1041 -30 1047
rect -88 1007 -76 1041
rect -42 1007 -30 1041
rect -88 1001 -30 1007
rect 30 1041 88 1047
rect 30 1007 42 1041
rect 76 1007 88 1041
rect 30 1001 88 1007
rect -141 948 -95 960
rect -141 -948 -135 948
rect -101 -948 -95 948
rect -141 -960 -95 -948
rect -23 948 23 960
rect -23 -948 -17 948
rect 17 -948 23 948
rect -23 -960 23 -948
rect 95 948 141 960
rect 95 -948 101 948
rect 135 -948 141 948
rect 95 -960 141 -948
rect -88 -1007 -30 -1001
rect -88 -1041 -76 -1007
rect -42 -1041 -30 -1007
rect -88 -1047 -30 -1041
rect 30 -1007 88 -1001
rect 30 -1041 42 -1007
rect 76 -1041 88 -1007
rect 30 -1047 88 -1041
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9.6 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
