magic
tech sky130A
magscale 1 2
timestamp 1667322124
<< error_p >>
rect -223 1636 -161 1642
rect -223 1602 -211 1636
rect -223 1596 -161 1602
<< nwell >>
rect -321 -1655 321 1655
<< pmoslvt >>
rect -227 -1555 -157 1555
rect -99 -1555 -29 1555
rect 29 -1555 99 1555
rect 157 -1555 227 1555
<< pdiff >>
rect -285 1543 -227 1555
rect -285 -1543 -273 1543
rect -239 -1543 -227 1543
rect -285 -1555 -227 -1543
rect -157 1543 -99 1555
rect -157 -1543 -145 1543
rect -111 -1543 -99 1543
rect -157 -1555 -99 -1543
rect -29 1543 29 1555
rect -29 -1543 -17 1543
rect 17 -1543 29 1543
rect -29 -1555 29 -1543
rect 99 1543 157 1555
rect 99 -1543 111 1543
rect 145 -1543 157 1543
rect 99 -1555 157 -1543
rect 227 1543 285 1555
rect 227 -1543 239 1543
rect 273 -1543 285 1543
rect 227 -1555 285 -1543
<< pdiffc >>
rect -273 -1543 -239 1543
rect -145 -1543 -111 1543
rect -17 -1543 17 1543
rect 111 -1543 145 1543
rect 239 -1543 273 1543
<< poly >>
rect -227 1636 -157 1652
rect -227 1602 -211 1636
rect -173 1602 -157 1636
rect -227 1555 -157 1602
rect -99 1578 99 1652
rect -99 1555 -29 1578
rect 29 1555 99 1578
rect 157 1555 227 1606
rect -227 -1578 -157 -1555
rect -99 -1578 -29 -1555
rect -227 -1652 -29 -1578
rect 29 -1578 99 -1555
rect 157 -1578 227 -1555
rect 29 -1652 227 -1578
<< polycont >>
rect -211 1602 -173 1636
<< locali >>
rect -227 1602 -211 1636
rect -173 1602 -157 1636
rect -273 1543 -239 1559
rect -273 -1559 -239 -1543
rect -145 1543 -111 1559
rect -145 -1559 -111 -1543
rect -17 1543 17 1559
rect -17 -1559 17 -1543
rect 111 1543 145 1559
rect 111 -1559 145 -1543
rect 239 1543 273 1559
rect 239 -1559 273 -1543
<< viali >>
rect -211 1602 -173 1636
rect -273 -1543 -239 1543
rect -145 -1543 -111 1543
rect -17 -1543 17 1543
rect 111 -1543 145 1543
rect 239 -1543 273 1543
<< metal1 >>
rect -223 1636 -161 1642
rect -223 1602 -211 1636
rect -173 1602 -161 1636
rect -223 1596 -161 1602
rect -279 1543 -233 1555
rect -279 -1543 -273 1543
rect -239 -1543 -233 1543
rect -279 -1555 -233 -1543
rect -151 1543 -105 1555
rect -151 -1543 -145 1543
rect -111 -1543 -105 1543
rect -151 -1555 -105 -1543
rect -23 1543 23 1555
rect -23 -1543 -17 1543
rect 17 -1543 23 1543
rect -23 -1555 23 -1543
rect 105 1543 151 1555
rect 105 -1543 111 1543
rect 145 -1543 151 1543
rect 105 -1555 151 -1543
rect 233 1543 279 1555
rect 233 -1543 239 1543
rect 273 -1543 279 1543
rect 233 -1555 279 -1543
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 15.55 l 0.35 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
