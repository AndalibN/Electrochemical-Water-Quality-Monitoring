magic
tech sky130A
magscale 1 2
timestamp 1666903823
<< nmos >>
rect -1000 -131 1000 69
<< ndiff >>
rect -1058 57 -1000 69
rect -1058 -119 -1046 57
rect -1012 -119 -1000 57
rect -1058 -131 -1000 -119
rect 1000 57 1058 69
rect 1000 -119 1012 57
rect 1046 -119 1058 57
rect 1000 -131 1058 -119
<< ndiffc >>
rect -1046 -119 -1012 57
rect 1012 -119 1046 57
<< poly >>
rect -1000 141 1000 157
rect -1000 107 -984 141
rect 984 107 1000 141
rect -1000 69 1000 107
rect -1000 -157 1000 -131
<< polycont >>
rect -984 107 984 141
<< locali >>
rect -1000 107 -984 141
rect 984 107 1000 141
rect -1046 57 -1012 73
rect -1046 -135 -1012 -119
rect 1012 57 1046 73
rect 1012 -135 1046 -119
<< viali >>
rect -984 107 984 141
rect -1046 -119 -1012 57
rect 1012 -119 1046 57
<< metal1 >>
rect -996 141 996 147
rect -996 107 -984 141
rect 984 107 996 141
rect -996 101 996 107
rect -1052 57 -1006 69
rect -1052 -119 -1046 57
rect -1012 -119 -1006 57
rect -1052 -131 -1006 -119
rect 1006 57 1052 69
rect 1006 -119 1012 57
rect 1046 -119 1052 57
rect 1006 -131 1052 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
