magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -109 -274 109 290
<< pmos >>
rect -15 -156 15 228
<< pdiff >>
rect -73 189 -15 228
rect -73 155 -61 189
rect -27 155 -15 189
rect -73 121 -15 155
rect -73 87 -61 121
rect -27 87 -15 121
rect -73 53 -15 87
rect -73 19 -61 53
rect -27 19 -15 53
rect -73 -15 -15 19
rect -73 -49 -61 -15
rect -27 -49 -15 -15
rect -73 -83 -15 -49
rect -73 -117 -61 -83
rect -27 -117 -15 -83
rect -73 -156 -15 -117
rect 15 189 73 228
rect 15 155 27 189
rect 61 155 73 189
rect 15 121 73 155
rect 15 87 27 121
rect 61 87 73 121
rect 15 53 73 87
rect 15 19 27 53
rect 61 19 73 53
rect 15 -15 73 19
rect 15 -49 27 -15
rect 61 -49 73 -15
rect 15 -83 73 -49
rect 15 -117 27 -83
rect 61 -117 73 -83
rect 15 -156 73 -117
<< pdiffc >>
rect -61 155 -27 189
rect -61 87 -27 121
rect -61 19 -27 53
rect -61 -49 -27 -15
rect -61 -117 -27 -83
rect 27 155 61 189
rect 27 87 61 121
rect 27 19 61 53
rect 27 -49 61 -15
rect 27 -117 61 -83
<< poly >>
rect -15 228 15 254
rect -15 -207 15 -156
rect -33 -223 33 -207
rect -33 -257 -17 -223
rect 17 -257 33 -223
rect -33 -273 33 -257
<< polycont >>
rect -17 -257 17 -223
<< locali >>
rect -61 197 -27 232
rect -61 125 -27 155
rect -61 53 -27 87
rect -61 -15 -27 19
rect -61 -83 -27 -53
rect -61 -160 -27 -125
rect 27 197 61 232
rect 27 125 61 155
rect 27 53 61 87
rect 27 -15 61 19
rect 27 -83 61 -53
rect 27 -160 61 -125
rect -33 -257 -17 -223
rect 17 -257 33 -223
<< viali >>
rect -61 189 -27 197
rect -61 163 -27 189
rect -61 121 -27 125
rect -61 91 -27 121
rect -61 19 -27 53
rect -61 -49 -27 -19
rect -61 -53 -27 -49
rect -61 -117 -27 -91
rect -61 -125 -27 -117
rect 27 189 61 197
rect 27 163 61 189
rect 27 121 61 125
rect 27 91 61 121
rect 27 19 61 53
rect 27 -49 61 -19
rect 27 -53 61 -49
rect 27 -117 61 -91
rect 27 -125 61 -117
rect -17 -257 17 -223
<< metal1 >>
rect -67 197 -21 228
rect -67 163 -61 197
rect -27 163 -21 197
rect -67 125 -21 163
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -156 -21 -125
rect 21 197 67 228
rect 21 163 27 197
rect 61 163 67 197
rect 21 125 67 163
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -156 67 -125
rect -31 -223 31 -213
rect -31 -257 -17 -223
rect 17 -257 31 -223
rect -31 -267 31 -257
<< end >>
