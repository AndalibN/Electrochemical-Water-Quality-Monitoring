magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -134 -1057 134 995
<< nmos >>
rect -50 -1031 50 969
<< ndiff >>
rect -108 938 -50 969
rect -108 904 -96 938
rect -62 904 -50 938
rect -108 870 -50 904
rect -108 836 -96 870
rect -62 836 -50 870
rect -108 802 -50 836
rect -108 768 -96 802
rect -62 768 -50 802
rect -108 734 -50 768
rect -108 700 -96 734
rect -62 700 -50 734
rect -108 666 -50 700
rect -108 632 -96 666
rect -62 632 -50 666
rect -108 598 -50 632
rect -108 564 -96 598
rect -62 564 -50 598
rect -108 530 -50 564
rect -108 496 -96 530
rect -62 496 -50 530
rect -108 462 -50 496
rect -108 428 -96 462
rect -62 428 -50 462
rect -108 394 -50 428
rect -108 360 -96 394
rect -62 360 -50 394
rect -108 326 -50 360
rect -108 292 -96 326
rect -62 292 -50 326
rect -108 258 -50 292
rect -108 224 -96 258
rect -62 224 -50 258
rect -108 190 -50 224
rect -108 156 -96 190
rect -62 156 -50 190
rect -108 122 -50 156
rect -108 88 -96 122
rect -62 88 -50 122
rect -108 54 -50 88
rect -108 20 -96 54
rect -62 20 -50 54
rect -108 -14 -50 20
rect -108 -48 -96 -14
rect -62 -48 -50 -14
rect -108 -82 -50 -48
rect -108 -116 -96 -82
rect -62 -116 -50 -82
rect -108 -150 -50 -116
rect -108 -184 -96 -150
rect -62 -184 -50 -150
rect -108 -218 -50 -184
rect -108 -252 -96 -218
rect -62 -252 -50 -218
rect -108 -286 -50 -252
rect -108 -320 -96 -286
rect -62 -320 -50 -286
rect -108 -354 -50 -320
rect -108 -388 -96 -354
rect -62 -388 -50 -354
rect -108 -422 -50 -388
rect -108 -456 -96 -422
rect -62 -456 -50 -422
rect -108 -490 -50 -456
rect -108 -524 -96 -490
rect -62 -524 -50 -490
rect -108 -558 -50 -524
rect -108 -592 -96 -558
rect -62 -592 -50 -558
rect -108 -626 -50 -592
rect -108 -660 -96 -626
rect -62 -660 -50 -626
rect -108 -694 -50 -660
rect -108 -728 -96 -694
rect -62 -728 -50 -694
rect -108 -762 -50 -728
rect -108 -796 -96 -762
rect -62 -796 -50 -762
rect -108 -830 -50 -796
rect -108 -864 -96 -830
rect -62 -864 -50 -830
rect -108 -898 -50 -864
rect -108 -932 -96 -898
rect -62 -932 -50 -898
rect -108 -966 -50 -932
rect -108 -1000 -96 -966
rect -62 -1000 -50 -966
rect -108 -1031 -50 -1000
rect 50 938 108 969
rect 50 904 62 938
rect 96 904 108 938
rect 50 870 108 904
rect 50 836 62 870
rect 96 836 108 870
rect 50 802 108 836
rect 50 768 62 802
rect 96 768 108 802
rect 50 734 108 768
rect 50 700 62 734
rect 96 700 108 734
rect 50 666 108 700
rect 50 632 62 666
rect 96 632 108 666
rect 50 598 108 632
rect 50 564 62 598
rect 96 564 108 598
rect 50 530 108 564
rect 50 496 62 530
rect 96 496 108 530
rect 50 462 108 496
rect 50 428 62 462
rect 96 428 108 462
rect 50 394 108 428
rect 50 360 62 394
rect 96 360 108 394
rect 50 326 108 360
rect 50 292 62 326
rect 96 292 108 326
rect 50 258 108 292
rect 50 224 62 258
rect 96 224 108 258
rect 50 190 108 224
rect 50 156 62 190
rect 96 156 108 190
rect 50 122 108 156
rect 50 88 62 122
rect 96 88 108 122
rect 50 54 108 88
rect 50 20 62 54
rect 96 20 108 54
rect 50 -14 108 20
rect 50 -48 62 -14
rect 96 -48 108 -14
rect 50 -82 108 -48
rect 50 -116 62 -82
rect 96 -116 108 -82
rect 50 -150 108 -116
rect 50 -184 62 -150
rect 96 -184 108 -150
rect 50 -218 108 -184
rect 50 -252 62 -218
rect 96 -252 108 -218
rect 50 -286 108 -252
rect 50 -320 62 -286
rect 96 -320 108 -286
rect 50 -354 108 -320
rect 50 -388 62 -354
rect 96 -388 108 -354
rect 50 -422 108 -388
rect 50 -456 62 -422
rect 96 -456 108 -422
rect 50 -490 108 -456
rect 50 -524 62 -490
rect 96 -524 108 -490
rect 50 -558 108 -524
rect 50 -592 62 -558
rect 96 -592 108 -558
rect 50 -626 108 -592
rect 50 -660 62 -626
rect 96 -660 108 -626
rect 50 -694 108 -660
rect 50 -728 62 -694
rect 96 -728 108 -694
rect 50 -762 108 -728
rect 50 -796 62 -762
rect 96 -796 108 -762
rect 50 -830 108 -796
rect 50 -864 62 -830
rect 96 -864 108 -830
rect 50 -898 108 -864
rect 50 -932 62 -898
rect 96 -932 108 -898
rect 50 -966 108 -932
rect 50 -1000 62 -966
rect 96 -1000 108 -966
rect 50 -1031 108 -1000
<< ndiffc >>
rect -96 904 -62 938
rect -96 836 -62 870
rect -96 768 -62 802
rect -96 700 -62 734
rect -96 632 -62 666
rect -96 564 -62 598
rect -96 496 -62 530
rect -96 428 -62 462
rect -96 360 -62 394
rect -96 292 -62 326
rect -96 224 -62 258
rect -96 156 -62 190
rect -96 88 -62 122
rect -96 20 -62 54
rect -96 -48 -62 -14
rect -96 -116 -62 -82
rect -96 -184 -62 -150
rect -96 -252 -62 -218
rect -96 -320 -62 -286
rect -96 -388 -62 -354
rect -96 -456 -62 -422
rect -96 -524 -62 -490
rect -96 -592 -62 -558
rect -96 -660 -62 -626
rect -96 -728 -62 -694
rect -96 -796 -62 -762
rect -96 -864 -62 -830
rect -96 -932 -62 -898
rect -96 -1000 -62 -966
rect 62 904 96 938
rect 62 836 96 870
rect 62 768 96 802
rect 62 700 96 734
rect 62 632 96 666
rect 62 564 96 598
rect 62 496 96 530
rect 62 428 96 462
rect 62 360 96 394
rect 62 292 96 326
rect 62 224 96 258
rect 62 156 96 190
rect 62 88 96 122
rect 62 20 96 54
rect 62 -48 96 -14
rect 62 -116 96 -82
rect 62 -184 96 -150
rect 62 -252 96 -218
rect 62 -320 96 -286
rect 62 -388 96 -354
rect 62 -456 96 -422
rect 62 -524 96 -490
rect 62 -592 96 -558
rect 62 -660 96 -626
rect 62 -728 96 -694
rect 62 -796 96 -762
rect 62 -864 96 -830
rect 62 -932 96 -898
rect 62 -1000 96 -966
<< poly >>
rect -50 1041 50 1057
rect -50 1007 -17 1041
rect 17 1007 50 1041
rect -50 969 50 1007
rect -50 -1057 50 -1031
<< polycont >>
rect -17 1007 17 1041
<< locali >>
rect -50 1007 -17 1041
rect 17 1007 50 1041
rect -96 938 -62 973
rect -96 870 -62 888
rect -96 802 -62 816
rect -96 734 -62 744
rect -96 666 -62 672
rect -96 598 -62 600
rect -96 562 -62 564
rect -96 490 -62 496
rect -96 418 -62 428
rect -96 346 -62 360
rect -96 274 -62 292
rect -96 202 -62 224
rect -96 130 -62 156
rect -96 58 -62 88
rect -96 -14 -62 20
rect -96 -82 -62 -48
rect -96 -150 -62 -120
rect -96 -218 -62 -192
rect -96 -286 -62 -264
rect -96 -354 -62 -336
rect -96 -422 -62 -408
rect -96 -490 -62 -480
rect -96 -558 -62 -552
rect -96 -626 -62 -624
rect -96 -662 -62 -660
rect -96 -734 -62 -728
rect -96 -806 -62 -796
rect -96 -878 -62 -864
rect -96 -950 -62 -932
rect -96 -1035 -62 -1000
rect 62 938 96 973
rect 62 870 96 888
rect 62 802 96 816
rect 62 734 96 744
rect 62 666 96 672
rect 62 598 96 600
rect 62 562 96 564
rect 62 490 96 496
rect 62 418 96 428
rect 62 346 96 360
rect 62 274 96 292
rect 62 202 96 224
rect 62 130 96 156
rect 62 58 96 88
rect 62 -14 96 20
rect 62 -82 96 -48
rect 62 -150 96 -120
rect 62 -218 96 -192
rect 62 -286 96 -264
rect 62 -354 96 -336
rect 62 -422 96 -408
rect 62 -490 96 -480
rect 62 -558 96 -552
rect 62 -626 96 -624
rect 62 -662 96 -660
rect 62 -734 96 -728
rect 62 -806 96 -796
rect 62 -878 96 -864
rect 62 -950 96 -932
rect 62 -1035 96 -1000
<< viali >>
rect -17 1007 17 1041
rect -96 904 -62 922
rect -96 888 -62 904
rect -96 836 -62 850
rect -96 816 -62 836
rect -96 768 -62 778
rect -96 744 -62 768
rect -96 700 -62 706
rect -96 672 -62 700
rect -96 632 -62 634
rect -96 600 -62 632
rect -96 530 -62 562
rect -96 528 -62 530
rect -96 462 -62 490
rect -96 456 -62 462
rect -96 394 -62 418
rect -96 384 -62 394
rect -96 326 -62 346
rect -96 312 -62 326
rect -96 258 -62 274
rect -96 240 -62 258
rect -96 190 -62 202
rect -96 168 -62 190
rect -96 122 -62 130
rect -96 96 -62 122
rect -96 54 -62 58
rect -96 24 -62 54
rect -96 -48 -62 -14
rect -96 -116 -62 -86
rect -96 -120 -62 -116
rect -96 -184 -62 -158
rect -96 -192 -62 -184
rect -96 -252 -62 -230
rect -96 -264 -62 -252
rect -96 -320 -62 -302
rect -96 -336 -62 -320
rect -96 -388 -62 -374
rect -96 -408 -62 -388
rect -96 -456 -62 -446
rect -96 -480 -62 -456
rect -96 -524 -62 -518
rect -96 -552 -62 -524
rect -96 -592 -62 -590
rect -96 -624 -62 -592
rect -96 -694 -62 -662
rect -96 -696 -62 -694
rect -96 -762 -62 -734
rect -96 -768 -62 -762
rect -96 -830 -62 -806
rect -96 -840 -62 -830
rect -96 -898 -62 -878
rect -96 -912 -62 -898
rect -96 -966 -62 -950
rect -96 -984 -62 -966
rect 62 904 96 922
rect 62 888 96 904
rect 62 836 96 850
rect 62 816 96 836
rect 62 768 96 778
rect 62 744 96 768
rect 62 700 96 706
rect 62 672 96 700
rect 62 632 96 634
rect 62 600 96 632
rect 62 530 96 562
rect 62 528 96 530
rect 62 462 96 490
rect 62 456 96 462
rect 62 394 96 418
rect 62 384 96 394
rect 62 326 96 346
rect 62 312 96 326
rect 62 258 96 274
rect 62 240 96 258
rect 62 190 96 202
rect 62 168 96 190
rect 62 122 96 130
rect 62 96 96 122
rect 62 54 96 58
rect 62 24 96 54
rect 62 -48 96 -14
rect 62 -116 96 -86
rect 62 -120 96 -116
rect 62 -184 96 -158
rect 62 -192 96 -184
rect 62 -252 96 -230
rect 62 -264 96 -252
rect 62 -320 96 -302
rect 62 -336 96 -320
rect 62 -388 96 -374
rect 62 -408 96 -388
rect 62 -456 96 -446
rect 62 -480 96 -456
rect 62 -524 96 -518
rect 62 -552 96 -524
rect 62 -592 96 -590
rect 62 -624 96 -592
rect 62 -694 96 -662
rect 62 -696 96 -694
rect 62 -762 96 -734
rect 62 -768 96 -762
rect 62 -830 96 -806
rect 62 -840 96 -830
rect 62 -898 96 -878
rect 62 -912 96 -898
rect 62 -966 96 -950
rect 62 -984 96 -966
<< metal1 >>
rect -46 1041 46 1047
rect -46 1007 -17 1041
rect 17 1007 46 1041
rect -46 1001 46 1007
rect -102 922 -56 969
rect -102 888 -96 922
rect -62 888 -56 922
rect -102 850 -56 888
rect -102 816 -96 850
rect -62 816 -56 850
rect -102 778 -56 816
rect -102 744 -96 778
rect -62 744 -56 778
rect -102 706 -56 744
rect -102 672 -96 706
rect -62 672 -56 706
rect -102 634 -56 672
rect -102 600 -96 634
rect -62 600 -56 634
rect -102 562 -56 600
rect -102 528 -96 562
rect -62 528 -56 562
rect -102 490 -56 528
rect -102 456 -96 490
rect -62 456 -56 490
rect -102 418 -56 456
rect -102 384 -96 418
rect -62 384 -56 418
rect -102 346 -56 384
rect -102 312 -96 346
rect -62 312 -56 346
rect -102 274 -56 312
rect -102 240 -96 274
rect -62 240 -56 274
rect -102 202 -56 240
rect -102 168 -96 202
rect -62 168 -56 202
rect -102 130 -56 168
rect -102 96 -96 130
rect -62 96 -56 130
rect -102 58 -56 96
rect -102 24 -96 58
rect -62 24 -56 58
rect -102 -14 -56 24
rect -102 -48 -96 -14
rect -62 -48 -56 -14
rect -102 -86 -56 -48
rect -102 -120 -96 -86
rect -62 -120 -56 -86
rect -102 -158 -56 -120
rect -102 -192 -96 -158
rect -62 -192 -56 -158
rect -102 -230 -56 -192
rect -102 -264 -96 -230
rect -62 -264 -56 -230
rect -102 -302 -56 -264
rect -102 -336 -96 -302
rect -62 -336 -56 -302
rect -102 -374 -56 -336
rect -102 -408 -96 -374
rect -62 -408 -56 -374
rect -102 -446 -56 -408
rect -102 -480 -96 -446
rect -62 -480 -56 -446
rect -102 -518 -56 -480
rect -102 -552 -96 -518
rect -62 -552 -56 -518
rect -102 -590 -56 -552
rect -102 -624 -96 -590
rect -62 -624 -56 -590
rect -102 -662 -56 -624
rect -102 -696 -96 -662
rect -62 -696 -56 -662
rect -102 -734 -56 -696
rect -102 -768 -96 -734
rect -62 -768 -56 -734
rect -102 -806 -56 -768
rect -102 -840 -96 -806
rect -62 -840 -56 -806
rect -102 -878 -56 -840
rect -102 -912 -96 -878
rect -62 -912 -56 -878
rect -102 -950 -56 -912
rect -102 -984 -96 -950
rect -62 -984 -56 -950
rect -102 -1031 -56 -984
rect 56 922 102 969
rect 56 888 62 922
rect 96 888 102 922
rect 56 850 102 888
rect 56 816 62 850
rect 96 816 102 850
rect 56 778 102 816
rect 56 744 62 778
rect 96 744 102 778
rect 56 706 102 744
rect 56 672 62 706
rect 96 672 102 706
rect 56 634 102 672
rect 56 600 62 634
rect 96 600 102 634
rect 56 562 102 600
rect 56 528 62 562
rect 96 528 102 562
rect 56 490 102 528
rect 56 456 62 490
rect 96 456 102 490
rect 56 418 102 456
rect 56 384 62 418
rect 96 384 102 418
rect 56 346 102 384
rect 56 312 62 346
rect 96 312 102 346
rect 56 274 102 312
rect 56 240 62 274
rect 96 240 102 274
rect 56 202 102 240
rect 56 168 62 202
rect 96 168 102 202
rect 56 130 102 168
rect 56 96 62 130
rect 96 96 102 130
rect 56 58 102 96
rect 56 24 62 58
rect 96 24 102 58
rect 56 -14 102 24
rect 56 -48 62 -14
rect 96 -48 102 -14
rect 56 -86 102 -48
rect 56 -120 62 -86
rect 96 -120 102 -86
rect 56 -158 102 -120
rect 56 -192 62 -158
rect 96 -192 102 -158
rect 56 -230 102 -192
rect 56 -264 62 -230
rect 96 -264 102 -230
rect 56 -302 102 -264
rect 56 -336 62 -302
rect 96 -336 102 -302
rect 56 -374 102 -336
rect 56 -408 62 -374
rect 96 -408 102 -374
rect 56 -446 102 -408
rect 56 -480 62 -446
rect 96 -480 102 -446
rect 56 -518 102 -480
rect 56 -552 62 -518
rect 96 -552 102 -518
rect 56 -590 102 -552
rect 56 -624 62 -590
rect 96 -624 102 -590
rect 56 -662 102 -624
rect 56 -696 62 -662
rect 96 -696 102 -662
rect 56 -734 102 -696
rect 56 -768 62 -734
rect 96 -768 102 -734
rect 56 -806 102 -768
rect 56 -840 62 -806
rect 96 -840 102 -806
rect 56 -878 102 -840
rect 56 -912 62 -878
rect 96 -912 102 -878
rect 56 -950 102 -912
rect 56 -984 62 -950
rect 96 -984 102 -950
rect 56 -1031 102 -984
<< end >>
