magic
tech sky130A
magscale 1 2
timestamp 1667325748
<< nwell >>
rect -1099 -741 947 741
<< pmos >>
rect -755 -625 -715 625
rect -657 -625 -617 625
rect -559 -625 -519 625
rect -461 -625 -421 625
rect -363 -625 -323 625
rect -265 -625 -225 625
rect -167 -625 -127 625
rect -69 -625 -29 625
rect 29 -625 69 625
rect 127 -625 167 625
rect 225 -625 265 625
rect 323 -625 363 625
rect 421 -625 461 625
rect 519 -625 559 625
rect 617 -625 657 625
rect 715 -625 755 625
<< pdiff >>
rect -813 613 -755 625
rect -813 -613 -801 613
rect -767 -613 -755 613
rect -813 -625 -755 -613
rect -715 613 -657 625
rect -715 -613 -703 613
rect -669 -613 -657 613
rect -715 -625 -657 -613
rect -617 613 -559 625
rect -617 -613 -605 613
rect -571 -613 -559 613
rect -617 -625 -559 -613
rect -519 613 -461 625
rect -519 -613 -507 613
rect -473 -613 -461 613
rect -519 -625 -461 -613
rect -421 613 -363 625
rect -421 -613 -409 613
rect -375 -613 -363 613
rect -421 -625 -363 -613
rect -323 613 -265 625
rect -323 -613 -311 613
rect -277 -613 -265 613
rect -323 -625 -265 -613
rect -225 613 -167 625
rect -225 -613 -213 613
rect -179 -613 -167 613
rect -225 -625 -167 -613
rect -127 613 -69 625
rect -127 -613 -115 613
rect -81 -613 -69 613
rect -127 -625 -69 -613
rect -29 613 29 625
rect -29 -613 -17 613
rect 17 -613 29 613
rect -29 -625 29 -613
rect 69 613 127 625
rect 69 -613 81 613
rect 115 -613 127 613
rect 69 -625 127 -613
rect 167 613 225 625
rect 167 -613 179 613
rect 213 -613 225 613
rect 167 -625 225 -613
rect 265 613 323 625
rect 265 -613 277 613
rect 311 -613 323 613
rect 265 -625 323 -613
rect 363 613 421 625
rect 363 -613 375 613
rect 409 -613 421 613
rect 363 -625 421 -613
rect 461 613 519 625
rect 461 -613 473 613
rect 507 -613 519 613
rect 461 -625 519 -613
rect 559 613 617 625
rect 559 -613 571 613
rect 605 -613 617 613
rect 559 -625 617 -613
rect 657 613 715 625
rect 657 -613 669 613
rect 703 -613 715 613
rect 657 -625 715 -613
rect 755 613 813 625
rect 755 -613 767 613
rect 801 -613 813 613
rect 755 -625 813 -613
<< pdiffc >>
rect -801 -613 -767 613
rect -703 -613 -669 613
rect -605 -613 -571 613
rect -507 -613 -473 613
rect -409 -613 -375 613
rect -311 -613 -277 613
rect -213 -613 -179 613
rect -115 -613 -81 613
rect -17 -613 17 613
rect 81 -613 115 613
rect 179 -613 213 613
rect 277 -613 311 613
rect 375 -613 409 613
rect 473 -613 507 613
rect 571 -613 605 613
rect 669 -613 703 613
rect 767 -613 801 613
<< poly >>
rect -1089 715 657 731
rect -1089 571 -1071 715
rect -927 693 657 715
rect -927 571 -911 693
rect -1089 555 -911 571
rect -1089 -571 -911 -555
rect -1089 -715 -1071 -571
rect -927 -693 -911 -571
rect -869 -651 -829 651
rect -755 625 -715 651
rect -657 625 -617 693
rect -559 625 -519 693
rect -461 625 -421 651
rect -363 625 -323 651
rect -265 625 -225 693
rect -167 625 -127 693
rect -69 625 -29 651
rect 29 625 69 651
rect 127 625 167 693
rect 225 625 265 693
rect 323 625 363 651
rect 421 625 461 651
rect 519 625 559 693
rect 617 625 657 693
rect 715 625 755 651
rect -755 -693 -715 -625
rect -657 -651 -617 -625
rect -559 -651 -519 -625
rect -461 -693 -421 -625
rect -363 -693 -323 -625
rect -265 -651 -225 -625
rect -167 -651 -127 -625
rect -69 -693 -29 -625
rect 29 -693 69 -625
rect 127 -651 167 -625
rect 225 -651 265 -625
rect 323 -693 363 -625
rect 421 -693 461 -625
rect 519 -651 559 -625
rect 617 -651 657 -625
rect 715 -693 755 -625
rect 829 -651 869 651
rect -927 -715 755 -693
rect -1089 -731 755 -715
<< polycont >>
rect -1071 571 -927 715
rect -1071 -715 -927 -571
<< locali >>
rect -1089 715 -911 731
rect -1089 571 -1071 715
rect -927 571 -911 715
rect -1089 555 -911 571
rect -801 613 -767 629
rect -1089 -571 -911 -555
rect -1089 -715 -1071 -571
rect -927 -715 -911 -571
rect -801 -629 -767 -613
rect -703 613 -669 629
rect -703 -629 -669 -613
rect -605 613 -571 629
rect -605 -629 -571 -613
rect -507 613 -473 629
rect -507 -629 -473 -613
rect -409 613 -375 629
rect -409 -629 -375 -613
rect -311 613 -277 629
rect -311 -629 -277 -613
rect -213 613 -179 629
rect -213 -629 -179 -613
rect -115 613 -81 629
rect -115 -629 -81 -613
rect -17 613 17 629
rect -17 -629 17 -613
rect 81 613 115 629
rect 81 -629 115 -613
rect 179 613 213 629
rect 179 -629 213 -613
rect 277 613 311 629
rect 277 -629 311 -613
rect 375 613 409 629
rect 375 -629 409 -613
rect 473 613 507 629
rect 473 -629 507 -613
rect 571 613 605 629
rect 571 -629 605 -613
rect 669 613 703 629
rect 669 -629 703 -613
rect 767 613 801 629
rect 767 -629 801 -613
rect -1089 -731 -911 -715
<< viali >>
rect -801 -613 -767 613
rect -703 -613 -669 613
rect -605 -613 -571 613
rect -507 -613 -473 613
rect -409 -613 -375 613
rect -311 -613 -277 613
rect -213 -613 -179 613
rect -115 -613 -81 613
rect -17 -613 17 613
rect 81 -613 115 613
rect 179 -613 213 613
rect 277 -613 311 613
rect 375 -613 409 613
rect 473 -613 507 613
rect 571 -613 605 613
rect 669 -613 703 613
rect 767 -613 801 613
<< metal1 >>
rect -1089 555 -911 731
rect -807 613 -761 625
rect -1089 -731 -911 -555
rect -807 -613 -801 613
rect -767 -613 -761 613
rect -807 -625 -761 -613
rect -709 613 -663 625
rect -709 -613 -703 613
rect -669 -613 -663 613
rect -709 -625 -663 -613
rect -611 613 -565 625
rect -611 -613 -605 613
rect -571 -613 -565 613
rect -611 -625 -565 -613
rect -513 613 -467 625
rect -513 -613 -507 613
rect -473 -613 -467 613
rect -513 -625 -467 -613
rect -415 613 -369 625
rect -415 -613 -409 613
rect -375 -613 -369 613
rect -415 -625 -369 -613
rect -317 613 -271 625
rect -317 -613 -311 613
rect -277 -613 -271 613
rect -317 -625 -271 -613
rect -219 613 -173 625
rect -219 -613 -213 613
rect -179 -613 -173 613
rect -219 -625 -173 -613
rect -121 613 -75 625
rect -121 -613 -115 613
rect -81 -613 -75 613
rect -121 -625 -75 -613
rect -23 613 23 625
rect -23 -613 -17 613
rect 17 -613 23 613
rect -23 -625 23 -613
rect 75 613 121 625
rect 75 -613 81 613
rect 115 -613 121 613
rect 75 -625 121 -613
rect 173 613 219 625
rect 173 -613 179 613
rect 213 -613 219 613
rect 173 -625 219 -613
rect 271 613 317 625
rect 271 -613 277 613
rect 311 -613 317 613
rect 271 -625 317 -613
rect 369 613 415 625
rect 369 -613 375 613
rect 409 -613 415 613
rect 369 -625 415 -613
rect 467 613 513 625
rect 467 -613 473 613
rect 507 -613 513 613
rect 467 -625 513 -613
rect 565 613 611 625
rect 565 -613 571 613
rect 605 -613 611 613
rect 565 -625 611 -613
rect 663 613 709 625
rect 663 -613 669 613
rect 703 -613 709 613
rect 663 -625 709 -613
rect 761 613 807 625
rect 761 -613 767 613
rect 801 -613 807 613
rect 761 -625 807 -613
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.25 l 0.2 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
