magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nwell >>
rect -223 -10100 223 10100
<< pmos >>
rect -129 -10000 -29 10000
rect 29 -10000 129 10000
<< pdiff >>
rect -187 9988 -129 10000
rect -187 -9988 -175 9988
rect -141 -9988 -129 9988
rect -187 -10000 -129 -9988
rect -29 9988 29 10000
rect -29 -9988 -17 9988
rect 17 -9988 29 9988
rect -29 -10000 29 -9988
rect 129 9988 187 10000
rect 129 -9988 141 9988
rect 175 -9988 187 9988
rect 129 -10000 187 -9988
<< pdiffc >>
rect -175 -9988 -141 9988
rect -17 -9988 17 9988
rect 141 -9988 175 9988
<< poly >>
rect -129 10081 -29 10097
rect -129 10047 -113 10081
rect -45 10047 -29 10081
rect -129 10000 -29 10047
rect 29 10081 129 10097
rect 29 10047 45 10081
rect 113 10047 129 10081
rect 29 10000 129 10047
rect -129 -10047 -29 -10000
rect -129 -10081 -113 -10047
rect -45 -10081 -29 -10047
rect -129 -10097 -29 -10081
rect 29 -10047 129 -10000
rect 29 -10081 45 -10047
rect 113 -10081 129 -10047
rect 29 -10097 129 -10081
<< polycont >>
rect -113 10047 -45 10081
rect 45 10047 113 10081
rect -113 -10081 -45 -10047
rect 45 -10081 113 -10047
<< locali >>
rect -129 10047 -113 10081
rect -45 10047 -29 10081
rect 29 10047 45 10081
rect 113 10047 129 10081
rect -175 9988 -141 10004
rect -175 -10004 -141 -9988
rect -17 9988 17 10004
rect -17 -10004 17 -9988
rect 141 9988 175 10004
rect 141 -10004 175 -9988
rect -129 -10081 -113 -10047
rect -45 -10081 -29 -10047
rect 29 -10081 45 -10047
rect 113 -10081 129 -10047
<< viali >>
rect -113 10047 -45 10081
rect 45 10047 113 10081
rect -175 -9988 -141 9988
rect -17 -9988 17 9988
rect 141 -9988 175 9988
rect -113 -10081 -45 -10047
rect 45 -10081 113 -10047
<< metal1 >>
rect -125 10081 -33 10087
rect -125 10047 -113 10081
rect -45 10047 -33 10081
rect -125 10041 -33 10047
rect 33 10081 125 10087
rect 33 10047 45 10081
rect 113 10047 125 10081
rect 33 10041 125 10047
rect -181 9988 -135 10000
rect -181 -9988 -175 9988
rect -141 -9988 -135 9988
rect -181 -10000 -135 -9988
rect -23 9988 23 10000
rect -23 -9988 -17 9988
rect 17 -9988 23 9988
rect -23 -10000 23 -9988
rect 135 9988 181 10000
rect 135 -9988 141 9988
rect 175 -9988 181 9988
rect 135 -10000 181 -9988
rect -125 -10047 -33 -10041
rect -125 -10081 -113 -10047
rect -45 -10081 -33 -10047
rect -125 -10087 -33 -10081
rect 33 -10047 125 -10041
rect 33 -10081 45 -10047
rect 113 -10081 125 -10047
rect 33 -10087 125 -10081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 100.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
