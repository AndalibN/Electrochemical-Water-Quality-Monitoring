magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -88 -307 -30 -301
rect 30 -307 88 -301
rect -88 -341 -76 -307
rect 30 -341 42 -307
rect -88 -347 -30 -341
rect 30 -347 88 -341
<< pwell >>
rect -173 -295 173 357
<< nmos >>
rect -89 -269 -29 331
rect 29 -269 89 331
<< ndiff >>
rect -147 286 -89 331
rect -147 252 -135 286
rect -101 252 -89 286
rect -147 218 -89 252
rect -147 184 -135 218
rect -101 184 -89 218
rect -147 150 -89 184
rect -147 116 -135 150
rect -101 116 -89 150
rect -147 82 -89 116
rect -147 48 -135 82
rect -101 48 -89 82
rect -147 14 -89 48
rect -147 -20 -135 14
rect -101 -20 -89 14
rect -147 -54 -89 -20
rect -147 -88 -135 -54
rect -101 -88 -89 -54
rect -147 -122 -89 -88
rect -147 -156 -135 -122
rect -101 -156 -89 -122
rect -147 -190 -89 -156
rect -147 -224 -135 -190
rect -101 -224 -89 -190
rect -147 -269 -89 -224
rect -29 286 29 331
rect -29 252 -17 286
rect 17 252 29 286
rect -29 218 29 252
rect -29 184 -17 218
rect 17 184 29 218
rect -29 150 29 184
rect -29 116 -17 150
rect 17 116 29 150
rect -29 82 29 116
rect -29 48 -17 82
rect 17 48 29 82
rect -29 14 29 48
rect -29 -20 -17 14
rect 17 -20 29 14
rect -29 -54 29 -20
rect -29 -88 -17 -54
rect 17 -88 29 -54
rect -29 -122 29 -88
rect -29 -156 -17 -122
rect 17 -156 29 -122
rect -29 -190 29 -156
rect -29 -224 -17 -190
rect 17 -224 29 -190
rect -29 -269 29 -224
rect 89 286 147 331
rect 89 252 101 286
rect 135 252 147 286
rect 89 218 147 252
rect 89 184 101 218
rect 135 184 147 218
rect 89 150 147 184
rect 89 116 101 150
rect 135 116 147 150
rect 89 82 147 116
rect 89 48 101 82
rect 135 48 147 82
rect 89 14 147 48
rect 89 -20 101 14
rect 135 -20 147 14
rect 89 -54 147 -20
rect 89 -88 101 -54
rect 135 -88 147 -54
rect 89 -122 147 -88
rect 89 -156 101 -122
rect 135 -156 147 -122
rect 89 -190 147 -156
rect 89 -224 101 -190
rect 135 -224 147 -190
rect 89 -269 147 -224
<< ndiffc >>
rect -135 252 -101 286
rect -135 184 -101 218
rect -135 116 -101 150
rect -135 48 -101 82
rect -135 -20 -101 14
rect -135 -88 -101 -54
rect -135 -156 -101 -122
rect -135 -224 -101 -190
rect -17 252 17 286
rect -17 184 17 218
rect -17 116 17 150
rect -17 48 17 82
rect -17 -20 17 14
rect -17 -88 17 -54
rect -17 -156 17 -122
rect -17 -224 17 -190
rect 101 252 135 286
rect 101 184 135 218
rect 101 116 135 150
rect 101 48 135 82
rect 101 -20 135 14
rect 101 -88 135 -54
rect 101 -156 135 -122
rect 101 -224 135 -190
<< poly >>
rect -89 355 89 398
rect -89 331 -29 355
rect 29 331 89 355
rect -89 -291 -29 -269
rect 29 -291 89 -269
rect -92 -307 -26 -291
rect -92 -341 -76 -307
rect -42 -341 -26 -307
rect -92 -357 -26 -341
rect 26 -307 92 -291
rect 26 -341 42 -307
rect 76 -341 92 -307
rect 26 -357 92 -341
<< polycont >>
rect -76 -341 -42 -307
rect 42 -341 76 -307
<< locali >>
rect -135 300 -101 335
rect -135 228 -101 252
rect -135 156 -101 184
rect -135 84 -101 116
rect -135 14 -101 48
rect -135 -54 -101 -22
rect -135 -122 -101 -94
rect -135 -190 -101 -166
rect -135 -273 -101 -238
rect -17 300 17 335
rect -17 228 17 252
rect -17 156 17 184
rect -17 84 17 116
rect -17 14 17 48
rect -17 -54 17 -22
rect -17 -122 17 -94
rect -17 -190 17 -166
rect -17 -273 17 -238
rect 101 300 135 335
rect 101 228 135 252
rect 101 156 135 184
rect 101 84 135 116
rect 101 14 135 48
rect 101 -54 135 -22
rect 101 -122 135 -94
rect 101 -190 135 -166
rect 101 -273 135 -238
rect -92 -341 -76 -307
rect -42 -341 -26 -307
rect 26 -341 42 -307
rect 76 -341 92 -307
<< viali >>
rect -135 286 -101 300
rect -135 266 -101 286
rect -135 218 -101 228
rect -135 194 -101 218
rect -135 150 -101 156
rect -135 122 -101 150
rect -135 82 -101 84
rect -135 50 -101 82
rect -135 -20 -101 12
rect -135 -22 -101 -20
rect -135 -88 -101 -60
rect -135 -94 -101 -88
rect -135 -156 -101 -132
rect -135 -166 -101 -156
rect -135 -224 -101 -204
rect -135 -238 -101 -224
rect -17 286 17 300
rect -17 266 17 286
rect -17 218 17 228
rect -17 194 17 218
rect -17 150 17 156
rect -17 122 17 150
rect -17 82 17 84
rect -17 50 17 82
rect -17 -20 17 12
rect -17 -22 17 -20
rect -17 -88 17 -60
rect -17 -94 17 -88
rect -17 -156 17 -132
rect -17 -166 17 -156
rect -17 -224 17 -204
rect -17 -238 17 -224
rect 101 286 135 300
rect 101 266 135 286
rect 101 218 135 228
rect 101 194 135 218
rect 101 150 135 156
rect 101 122 135 150
rect 101 82 135 84
rect 101 50 135 82
rect 101 -20 135 12
rect 101 -22 135 -20
rect 101 -88 135 -60
rect 101 -94 135 -88
rect 101 -156 135 -132
rect 101 -166 135 -156
rect 101 -224 135 -204
rect 101 -238 135 -224
rect -76 -341 -42 -307
rect 42 -341 76 -307
<< metal1 >>
rect -141 300 -95 331
rect -141 266 -135 300
rect -101 266 -95 300
rect -141 228 -95 266
rect -141 194 -135 228
rect -101 194 -95 228
rect -141 156 -95 194
rect -141 122 -135 156
rect -101 122 -95 156
rect -141 84 -95 122
rect -141 50 -135 84
rect -101 50 -95 84
rect -141 12 -95 50
rect -141 -22 -135 12
rect -101 -22 -95 12
rect -141 -60 -95 -22
rect -141 -94 -135 -60
rect -101 -94 -95 -60
rect -141 -132 -95 -94
rect -141 -166 -135 -132
rect -101 -166 -95 -132
rect -141 -204 -95 -166
rect -141 -238 -135 -204
rect -101 -238 -95 -204
rect -141 -269 -95 -238
rect -23 300 23 331
rect -23 266 -17 300
rect 17 266 23 300
rect -23 228 23 266
rect -23 194 -17 228
rect 17 194 23 228
rect -23 156 23 194
rect -23 122 -17 156
rect 17 122 23 156
rect -23 84 23 122
rect -23 50 -17 84
rect 17 50 23 84
rect -23 12 23 50
rect -23 -22 -17 12
rect 17 -22 23 12
rect -23 -60 23 -22
rect -23 -94 -17 -60
rect 17 -94 23 -60
rect -23 -132 23 -94
rect -23 -166 -17 -132
rect 17 -166 23 -132
rect -23 -204 23 -166
rect -23 -238 -17 -204
rect 17 -238 23 -204
rect -23 -269 23 -238
rect 95 300 141 331
rect 95 266 101 300
rect 135 266 141 300
rect 95 228 141 266
rect 95 194 101 228
rect 135 194 141 228
rect 95 156 141 194
rect 95 122 101 156
rect 135 122 141 156
rect 95 84 141 122
rect 95 50 101 84
rect 135 50 141 84
rect 95 12 141 50
rect 95 -22 101 12
rect 135 -22 141 12
rect 95 -60 141 -22
rect 95 -94 101 -60
rect 135 -94 141 -60
rect 95 -132 141 -94
rect 95 -166 101 -132
rect 135 -166 141 -132
rect 95 -204 141 -166
rect 95 -238 101 -204
rect 135 -238 141 -204
rect 95 -269 141 -238
rect -88 -307 -30 -301
rect -88 -341 -76 -307
rect -42 -341 -30 -307
rect -88 -347 -30 -341
rect 30 -307 88 -301
rect 30 -341 42 -307
rect 76 -341 88 -307
rect 30 -347 88 -341
<< end >>
