magic
tech sky130A
magscale 1 2
timestamp 1667951165
<< metal4 >>
rect -50200 -23712 -33400 -23600
rect -50200 -27088 -50088 -23712
rect -46712 -27088 -36888 -23712
rect -33512 -27088 -33400 -23712
rect -50200 -27200 -33400 -27088
<< via4 >>
rect -50088 -27088 -46712 -23712
rect -36888 -27088 -33512 -23712
<< metal5 >>
tri -37600 1125 -33725 5000 se
rect -33725 1400 -10475 5000
tri -10475 1400 -6875 5000 sw
rect -33725 1125 -32834 1400
tri -38937 -212 -37600 1125 se
rect -37600 800 -32834 1125
tri -32834 800 -32234 1400 nw
tri -11966 800 -11366 1400 ne
rect -11366 800 -6875 1400
rect -37600 -49 -33683 800
tri -33683 -49 -32834 800 nw
tri -32834 -49 -31985 800 se
rect -31985 -49 -12215 800
tri -12215 -49 -11366 800 sw
tri -11366 -49 -10517 800 ne
rect -10517 -49 -6875 800
rect -37600 -212 -33846 -49
tri -33846 -212 -33683 -49 nw
tri -32997 -212 -32834 -49 se
rect -32834 -212 -11366 -49
tri -41800 -3075 -38937 -212 se
rect -38937 -1061 -34695 -212
tri -34695 -1061 -33846 -212 nw
tri -33846 -1061 -32997 -212 se
rect -32997 -898 -11366 -212
tri -11366 -898 -10517 -49 sw
tri -10517 -898 -9668 -49 ne
rect -9668 -898 -6875 -49
rect -32997 -1061 -10517 -898
rect -38937 -1910 -35544 -1061
tri -35544 -1910 -34695 -1061 nw
tri -34695 -1910 -33846 -1061 se
rect -33846 -1102 -10517 -1061
tri -10517 -1102 -10313 -898 sw
tri -9668 -1102 -9464 -898 ne
rect -9464 -1102 -6875 -898
rect -33846 -1910 -10313 -1102
rect -38937 -1951 -35585 -1910
tri -35585 -1951 -35544 -1910 nw
tri -34736 -1951 -34695 -1910 se
rect -34695 -1951 -10313 -1910
tri -10313 -1951 -9464 -1102 sw
tri -9464 -1951 -8615 -1102 ne
rect -8615 -1951 -6875 -1102
rect -38937 -2800 -36434 -1951
tri -36434 -2800 -35585 -1951 nw
tri -35585 -2800 -34736 -1951 se
rect -34736 -2800 -9464 -1951
tri -9464 -2800 -8615 -1951 sw
tri -8615 -2800 -7766 -1951 ne
rect -7766 -2800 -6875 -1951
tri -6875 -2800 -2675 1400 sw
rect -38937 -3075 -37283 -2800
tri -42691 -3966 -41800 -3075 se
rect -41800 -3649 -37283 -3075
tri -37283 -3649 -36434 -2800 nw
tri -36434 -3649 -35585 -2800 se
rect -35585 -3400 -31094 -2800
tri -31094 -3400 -30494 -2800 nw
tri -13706 -3400 -13106 -2800 ne
rect -13106 -3400 -8615 -2800
rect -35585 -3649 -31942 -3400
rect -41800 -3966 -37600 -3649
tri -37600 -3966 -37283 -3649 nw
tri -36751 -3966 -36434 -3649 se
rect -36434 -3966 -31942 -3649
tri -46000 -7275 -42691 -3966 se
rect -42691 -4815 -38449 -3966
tri -38449 -4815 -37600 -3966 nw
tri -37600 -4815 -36751 -3966 se
rect -36751 -4248 -31942 -3966
tri -31942 -4248 -31094 -3400 nw
tri -31094 -4248 -30246 -3400 se
rect -30246 -4248 -13954 -3400
tri -13954 -4248 -13106 -3400 sw
tri -13106 -4248 -12258 -3400 ne
rect -12258 -3649 -8615 -3400
tri -8615 -3649 -7766 -2800 sw
tri -7766 -3649 -6917 -2800 ne
rect -6917 -3649 -2675 -2800
rect -12258 -4248 -7766 -3649
rect -36751 -4815 -32790 -4248
rect -42691 -5664 -39298 -4815
tri -39298 -5664 -38449 -4815 nw
tri -38449 -5664 -37600 -4815 se
rect -37600 -5096 -32790 -4815
tri -32790 -5096 -31942 -4248 nw
tri -31942 -5096 -31094 -4248 se
rect -31094 -5096 -13106 -4248
tri -13106 -5096 -12258 -4248 sw
tri -12258 -5096 -11410 -4248 ne
rect -11410 -4498 -7766 -4248
tri -7766 -4498 -6917 -3649 sw
tri -6917 -4498 -6068 -3649 ne
rect -6068 -4498 -2675 -3649
rect -11410 -5096 -6917 -4498
rect -37600 -5304 -32998 -5096
tri -32998 -5304 -32790 -5096 nw
tri -32150 -5304 -31942 -5096 se
rect -31942 -5304 -12258 -5096
tri -12258 -5304 -12050 -5096 sw
tri -11410 -5304 -11202 -5096 ne
rect -11202 -5302 -6917 -5096
tri -6917 -5302 -6113 -4498 sw
tri -6068 -5302 -5264 -4498 ne
rect -5264 -5302 -2675 -4498
rect -11202 -5304 -6113 -5302
rect -37600 -5664 -33846 -5304
rect -42691 -6152 -39786 -5664
tri -39786 -6152 -39298 -5664 nw
tri -38937 -6152 -38449 -5664 se
rect -38449 -6152 -33846 -5664
tri -33846 -6152 -32998 -5304 nw
tri -32998 -6152 -32150 -5304 se
rect -32150 -6152 -12050 -5304
tri -12050 -6152 -11202 -5304 sw
tri -11202 -6152 -10354 -5304 ne
rect -10354 -6151 -6113 -5304
tri -6113 -6151 -5264 -5302 sw
tri -5264 -6151 -4415 -5302 ne
rect -4415 -6151 -2675 -5302
rect -10354 -6152 -5264 -6151
rect -42691 -7001 -40635 -6152
tri -40635 -7001 -39786 -6152 nw
tri -39786 -7001 -38937 -6152 se
rect -38937 -7000 -34694 -6152
tri -34694 -7000 -33846 -6152 nw
tri -33846 -7000 -32998 -6152 se
rect -32998 -7000 -11202 -6152
tri -11202 -7000 -10354 -6152 sw
tri -10354 -7000 -9506 -6152 ne
rect -9506 -7000 -5264 -6152
tri -5264 -7000 -4415 -6151 sw
tri -4415 -7000 -3566 -6151 ne
rect -3566 -7000 -2675 -6151
tri -2675 -7000 1525 -2800 sw
rect -38937 -7001 -35542 -7000
rect -42691 -7275 -40951 -7001
tri -46891 -8166 -46000 -7275 se
rect -46000 -7317 -40951 -7275
tri -40951 -7317 -40635 -7001 nw
tri -40102 -7317 -39786 -7001 se
rect -39786 -7317 -35542 -7001
rect -46000 -8166 -41800 -7317
tri -41800 -8166 -40951 -7317 nw
tri -40951 -8166 -40102 -7317 se
rect -40102 -7848 -35542 -7317
tri -35542 -7848 -34694 -7000 nw
tri -34694 -7848 -33846 -7000 se
rect -40102 -8166 -36390 -7848
tri -49600 -10875 -46891 -8166 se
rect -46891 -9015 -42649 -8166
tri -42649 -9015 -41800 -8166 nw
tri -41800 -9015 -40951 -8166 se
rect -40951 -8696 -36390 -8166
tri -36390 -8696 -35542 -7848 nw
tri -35542 -8696 -34694 -7848 se
rect -34694 -8696 -33846 -7848
rect -40951 -9015 -36752 -8696
rect -46891 -9864 -43498 -9015
tri -43498 -9864 -42649 -9015 nw
tri -42649 -9864 -41800 -9015 se
rect -41800 -9058 -36752 -9015
tri -36752 -9058 -36390 -8696 nw
tri -35904 -9058 -35542 -8696 se
rect -35542 -9058 -33846 -8696
rect -41800 -9864 -37600 -9058
rect -46891 -9906 -43540 -9864
tri -43540 -9906 -43498 -9864 nw
tri -42691 -9906 -42649 -9864 se
rect -42649 -9906 -37600 -9864
tri -37600 -9906 -36752 -9058 nw
tri -36752 -9906 -35904 -9058 se
rect -35904 -9906 -33846 -9058
rect -46891 -10755 -44389 -9906
tri -44389 -10755 -43540 -9906 nw
tri -43540 -10755 -42691 -9906 se
rect -42691 -10754 -38448 -9906
tri -38448 -10754 -37600 -9906 nw
tri -37600 -10754 -36752 -9906 se
rect -36752 -10754 -33846 -9906
rect -42691 -10755 -39296 -10754
rect -46891 -10875 -44551 -10755
rect -49600 -10917 -44551 -10875
tri -44551 -10917 -44389 -10755 nw
tri -43702 -10917 -43540 -10755 se
rect -43540 -10917 -39296 -10755
rect -49600 -11766 -45400 -10917
tri -45400 -11766 -44551 -10917 nw
tri -44551 -11766 -43702 -10917 se
rect -43702 -11602 -39296 -10917
tri -39296 -11602 -38448 -10754 nw
tri -38448 -11602 -37600 -10754 se
rect -37600 -11602 -33846 -10754
rect -43702 -11766 -39785 -11602
rect -49600 -12800 -46000 -11766
tri -46000 -12366 -45400 -11766 nw
rect -53200 -16400 -46000 -12800
tri -45400 -12615 -44551 -11766 se
rect -44551 -12091 -39785 -11766
tri -39785 -12091 -39296 -11602 nw
tri -38937 -12091 -38448 -11602 se
rect -38448 -12091 -33846 -11602
tri -33846 -12091 -28755 -7000 nw
tri -15445 -12091 -10354 -7000 ne
tri -10354 -7848 -9506 -7000 sw
tri -9506 -7848 -8658 -7000 ne
rect -8658 -7848 -4415 -7000
rect -10354 -8696 -9506 -7848
tri -9506 -8696 -8658 -7848 sw
tri -8658 -8696 -7810 -7848 ne
rect -7810 -7849 -4415 -7848
tri -4415 -7849 -3566 -7000 sw
tri -3566 -7849 -2717 -7000 ne
rect -2717 -7849 1525 -7000
rect -7810 -8696 -3566 -7849
rect -10354 -9058 -8658 -8696
tri -8658 -9058 -8296 -8696 sw
tri -7810 -9058 -7448 -8696 ne
rect -7448 -8698 -3566 -8696
tri -3566 -8698 -2717 -7849 sw
tri -2717 -8698 -1868 -7849 ne
rect -1868 -8698 1525 -7849
rect -7448 -9056 -2717 -8698
tri -2717 -9056 -2359 -8698 sw
tri -1868 -9056 -1510 -8698 ne
rect -1510 -9056 1525 -8698
rect -7448 -9058 -2359 -9056
rect -10354 -9906 -8296 -9058
tri -8296 -9906 -7448 -9058 sw
tri -7448 -9906 -6600 -9058 ne
rect -6600 -9905 -2359 -9058
tri -2359 -9905 -1510 -9056 sw
tri -1510 -9905 -661 -9056 ne
rect -661 -9905 1525 -9056
rect -6600 -9906 -1510 -9905
rect -10354 -10754 -7448 -9906
tri -7448 -10754 -6600 -9906 sw
tri -6600 -10754 -5752 -9906 ne
rect -5752 -10754 -1510 -9906
tri -1510 -10754 -661 -9905 sw
tri -661 -10754 188 -9905 ne
rect 188 -10754 1525 -9905
rect -10354 -11602 -6600 -10754
tri -6600 -11602 -5752 -10754 sw
tri -5752 -11602 -4904 -10754 ne
rect -4904 -11602 -661 -10754
rect -10354 -12091 -5752 -11602
rect -44551 -12615 -40494 -12091
rect -45400 -12800 -40494 -12615
tri -40494 -12800 -39785 -12091 nw
tri -39646 -12800 -38937 -12091 se
rect -38937 -12800 -37600 -12091
rect -45400 -13506 -41200 -12800
tri -41200 -13506 -40494 -12800 nw
tri -40352 -13506 -39646 -12800 se
rect -39646 -13506 -37600 -12800
rect -50200 -23712 -46600 -23600
rect -50200 -27088 -50088 -23712
rect -46712 -27088 -46600 -23712
rect -50200 -27200 -46600 -27088
rect -45400 -29464 -41800 -13506
tri -41800 -14106 -41200 -13506 nw
tri -41200 -14354 -40352 -13506 se
rect -40352 -14354 -37600 -13506
rect -41200 -27724 -37600 -14354
tri -37600 -15845 -33846 -12091 nw
tri -10354 -15845 -6600 -12091 ne
rect -6600 -12450 -5752 -12091
tri -5752 -12450 -4904 -11602 sw
tri -4904 -12450 -4056 -11602 ne
rect -4056 -11603 -661 -11602
tri -661 -11603 188 -10754 sw
tri 188 -11603 1037 -10754 ne
rect 1037 -10875 1525 -10754
tri 1525 -10875 5400 -7000 sw
rect 1037 -11603 5400 -10875
rect -4056 -12366 188 -11603
tri 188 -12366 951 -11603 sw
tri 1037 -12366 1800 -11603 ne
rect -4056 -12450 951 -12366
rect -6600 -12658 -4904 -12450
tri -4904 -12658 -4696 -12450 sw
tri -4056 -12658 -3848 -12450 ne
rect -3848 -12615 951 -12450
tri 951 -12615 1200 -12366 sw
rect -3848 -12658 1200 -12615
rect -6600 -13506 -4696 -12658
tri -4696 -13506 -3848 -12658 sw
tri -3848 -13506 -3000 -12658 ne
rect -3000 -13506 1200 -12658
rect -6600 -14354 -3848 -13506
tri -3848 -14354 -3000 -13506 sw
tri -3000 -14106 -2400 -13506 ne
rect -37000 -23712 -33400 -23600
rect -37000 -27088 -36888 -23712
rect -33512 -27088 -33400 -23712
tri -37600 -27724 -37000 -27124 sw
rect -37000 -27200 -33400 -27088
tri -36676 -27724 -36152 -27200 ne
rect -36152 -27724 -33400 -27200
rect -41200 -28572 -37000 -27724
tri -37000 -28572 -36152 -27724 sw
tri -36152 -28572 -35304 -27724 ne
rect -35304 -28572 -33400 -27724
rect -41200 -28616 -36152 -28572
tri -41800 -29464 -41200 -28864 sw
tri -41200 -29464 -40352 -28616 ne
rect -40352 -28780 -36152 -28616
tri -36152 -28780 -35944 -28572 sw
tri -35304 -28780 -35096 -28572 ne
rect -35096 -28780 -33400 -28572
rect -40352 -29464 -35944 -28780
rect -45400 -29628 -41200 -29464
tri -41200 -29628 -41036 -29464 sw
tri -40352 -29628 -40188 -29464 ne
rect -40188 -29628 -35944 -29464
tri -35944 -29628 -35096 -28780 sw
tri -35096 -29628 -34248 -28780 ne
rect -34248 -29628 -33400 -28780
rect -45400 -30355 -41036 -29628
tri -45400 -33000 -42755 -30355 ne
rect -42755 -30476 -41036 -30355
tri -41036 -30476 -40188 -29628 sw
tri -40188 -30476 -39340 -29628 ne
rect -39340 -30476 -35096 -29628
tri -35096 -30476 -34248 -29628 sw
tri -34248 -30476 -33400 -29628 ne
tri -33400 -30476 -28309 -25385 sw
tri -9124 -27909 -6600 -25385 se
rect -6600 -26876 -3000 -14354
rect -6600 -27724 -3848 -26876
tri -3848 -27724 -3000 -26876 nw
tri -3000 -27724 -2400 -27124 se
rect -2400 -27724 1200 -13506
rect -6600 -27909 -4033 -27724
tri -4033 -27909 -3848 -27724 nw
tri -3185 -27909 -3000 -27724 se
rect -3000 -27909 1200 -27724
tri -11691 -30476 -9124 -27909 se
rect -9124 -28757 -4881 -27909
tri -4881 -28757 -4033 -27909 nw
tri -4033 -28757 -3185 -27909 se
rect -3185 -28616 1200 -27909
rect -3185 -28757 352 -28616
rect -9124 -28780 -4904 -28757
tri -4904 -28780 -4881 -28757 nw
tri -4056 -28780 -4033 -28757 se
rect -4033 -28780 352 -28757
rect -9124 -29628 -5752 -28780
tri -5752 -29628 -4904 -28780 nw
tri -4904 -29628 -4056 -28780 se
rect -4056 -29464 352 -28780
tri 352 -29464 1200 -28616 nw
tri 1200 -29464 1800 -28864 se
rect 1800 -29464 5400 -11603
rect -4056 -29628 -496 -29464
rect -9124 -30476 -6600 -29628
tri -6600 -30476 -5752 -29628 nw
tri -5752 -30476 -4904 -29628 se
rect -4904 -30312 -496 -29628
tri -496 -30312 352 -29464 nw
tri 352 -30312 1200 -29464 se
rect 1200 -30312 5400 -29464
rect -4904 -30476 -660 -30312
tri -660 -30476 -496 -30312 nw
tri 188 -30476 352 -30312 se
rect 352 -30355 5400 -30312
rect 352 -30476 1800 -30355
rect -42755 -31324 -40188 -30476
tri -40188 -31324 -39340 -30476 sw
tri -39340 -31324 -38492 -30476 ne
rect -38492 -31324 -34248 -30476
tri -34248 -31324 -33400 -30476 sw
tri -33400 -31324 -32552 -30476 ne
rect -32552 -31324 -28309 -30476
rect -42755 -32152 -39340 -31324
tri -39340 -32152 -38512 -31324 sw
tri -38492 -32152 -37664 -31324 ne
rect -37664 -32152 -33400 -31324
tri -33400 -32152 -32572 -31324 sw
tri -32552 -32152 -31724 -31324 ne
rect -31724 -32152 -28309 -31324
rect -42755 -33000 -38512 -32152
tri -38512 -33000 -37664 -32152 sw
tri -37664 -33000 -36816 -32152 ne
rect -36816 -33000 -32572 -32152
tri -32572 -33000 -31724 -32152 sw
tri -31724 -33000 -30876 -32152 ne
rect -30876 -33000 -28309 -32152
tri -28309 -33000 -25785 -30476 sw
tri -14215 -33000 -11691 -30476 se
rect -11691 -31324 -7448 -30476
tri -7448 -31324 -6600 -30476 nw
tri -6600 -31324 -5752 -30476 se
rect -5752 -31324 -1508 -30476
tri -1508 -31324 -660 -30476 nw
tri -660 -31324 188 -30476 se
rect 188 -31324 1800 -30476
rect -11691 -32152 -8276 -31324
tri -8276 -32152 -7448 -31324 nw
tri -7428 -32152 -6600 -31324 se
rect -6600 -31368 -1552 -31324
tri -1552 -31368 -1508 -31324 nw
tri -704 -31368 -660 -31324 se
rect -660 -31368 1800 -31324
rect -6600 -32152 -2400 -31368
rect -11691 -33000 -9124 -32152
tri -9124 -33000 -8276 -32152 nw
tri -8276 -33000 -7428 -32152 se
rect -7428 -32216 -2400 -32152
tri -2400 -32216 -1552 -31368 nw
tri -1552 -32216 -704 -31368 se
rect -704 -32216 1800 -31368
rect -7428 -33000 -3248 -32216
tri -42755 -37200 -38555 -33000 ne
rect -38555 -33848 -37664 -33000
tri -37664 -33848 -36816 -33000 sw
tri -36816 -33848 -35968 -33000 ne
rect -35968 -33848 -31724 -33000
tri -31724 -33848 -30876 -33000 sw
tri -30876 -33848 -30028 -33000 ne
rect -30028 -33848 -9972 -33000
tri -9972 -33848 -9124 -33000 nw
tri -9124 -33848 -8276 -33000 se
rect -8276 -33064 -3248 -33000
tri -3248 -33064 -2400 -32216 nw
tri -2400 -33064 -1552 -32216 se
rect -1552 -33064 1800 -32216
rect -8276 -33848 -4032 -33064
tri -4032 -33848 -3248 -33064 nw
tri -3184 -33848 -2400 -33064 se
rect -2400 -33848 1800 -33064
rect -38555 -34696 -36816 -33848
tri -36816 -34696 -35968 -33848 sw
tri -35968 -34696 -35120 -33848 ne
rect -35120 -34696 -30876 -33848
tri -30876 -34696 -30028 -33848 sw
tri -30028 -34696 -29180 -33848 ne
rect -29180 -34696 -10820 -33848
tri -10820 -34696 -9972 -33848 nw
tri -9972 -34696 -9124 -33848 se
rect -9124 -34696 -4880 -33848
tri -4880 -34696 -4032 -33848 nw
tri -4032 -34696 -3184 -33848 se
rect -3184 -33955 1800 -33848
tri 1800 -33955 5400 -30355 nw
rect -3184 -34696 -2400 -33955
rect -38555 -35504 -35968 -34696
tri -35968 -35504 -35160 -34696 sw
tri -35120 -35504 -34312 -34696 ne
rect -34312 -34904 -30028 -34696
tri -30028 -34904 -29820 -34696 sw
tri -29180 -34904 -28972 -34696 ne
rect -28972 -34904 -11028 -34696
tri -11028 -34904 -10820 -34696 nw
tri -10180 -34904 -9972 -34696 se
rect -9972 -34720 -4904 -34696
tri -4904 -34720 -4880 -34696 nw
tri -4056 -34720 -4032 -34696 se
rect -4032 -34720 -2400 -34696
rect -9972 -34904 -5752 -34720
rect -34312 -35504 -29820 -34904
rect -38555 -36352 -35160 -35504
tri -35160 -36352 -34312 -35504 sw
tri -34312 -36352 -33464 -35504 ne
rect -33464 -35752 -29820 -35504
tri -29820 -35752 -28972 -34904 sw
tri -28972 -35752 -28124 -34904 ne
rect -28124 -35752 -11876 -34904
tri -11876 -35752 -11028 -34904 nw
tri -11028 -35752 -10180 -34904 se
rect -10180 -35568 -5752 -34904
tri -5752 -35568 -4904 -34720 nw
tri -4904 -35568 -4056 -34720 se
rect -4056 -35568 -2400 -34720
rect -10180 -35752 -6600 -35568
rect -33464 -36352 -28972 -35752
rect -38555 -37200 -34312 -36352
tri -34312 -37200 -33464 -36352 sw
tri -33464 -37200 -32616 -36352 ne
rect -32616 -36600 -28972 -36352
tri -28972 -36600 -28124 -35752 sw
tri -28124 -36600 -27276 -35752 ne
rect -27276 -36600 -12724 -35752
tri -12724 -36600 -11876 -35752 nw
tri -11876 -36600 -11028 -35752 se
rect -11028 -36416 -6600 -35752
tri -6600 -36416 -5752 -35568 nw
tri -5752 -36416 -4904 -35568 se
rect -4904 -36416 -2400 -35568
rect -11028 -36600 -7448 -36416
rect -32616 -37200 -28124 -36600
tri -28124 -37200 -27524 -36600 sw
tri -12476 -37200 -11876 -36600 se
rect -11876 -37200 -7448 -36600
tri -38555 -41400 -34355 -37200 ne
rect -34355 -38048 -33464 -37200
tri -33464 -38048 -32616 -37200 sw
tri -32616 -38048 -31768 -37200 ne
rect -31768 -37264 -7448 -37200
tri -7448 -37264 -6600 -36416 nw
tri -6600 -37264 -5752 -36416 se
rect -5752 -37264 -2400 -36416
rect -31768 -38048 -8276 -37264
rect -34355 -38896 -32616 -38048
tri -32616 -38896 -31768 -38048 sw
tri -31768 -38896 -30920 -38048 ne
rect -30920 -38092 -8276 -38048
tri -8276 -38092 -7448 -37264 nw
tri -7428 -38092 -6600 -37264 se
rect -6600 -38092 -2400 -37264
rect -30920 -38896 -9124 -38092
rect -34355 -39104 -31768 -38896
tri -31768 -39104 -31560 -38896 sw
tri -30920 -39104 -30712 -38896 ne
rect -30712 -38940 -9124 -38896
tri -9124 -38940 -8276 -38092 nw
tri -8276 -38940 -7428 -38092 se
rect -7428 -38155 -2400 -38092
tri -2400 -38155 1800 -33955 nw
rect -7428 -38940 -6600 -38155
rect -30712 -39104 -9972 -38940
rect -34355 -39952 -31560 -39104
tri -31560 -39952 -30712 -39104 sw
tri -30712 -39952 -29864 -39104 ne
rect -29864 -39788 -9972 -39104
tri -9972 -39788 -9124 -38940 nw
tri -9124 -39788 -8276 -38940 se
rect -8276 -39788 -6600 -38940
rect -29864 -39952 -10136 -39788
tri -10136 -39952 -9972 -39788 nw
tri -9288 -39952 -9124 -39788 se
rect -9124 -39952 -6600 -39788
rect -34355 -40800 -30712 -39952
tri -30712 -40800 -29864 -39952 sw
tri -29864 -40800 -29016 -39952 ne
rect -29016 -40800 -10984 -39952
tri -10984 -40800 -10136 -39952 nw
tri -10136 -40800 -9288 -39952 se
rect -9288 -40800 -6600 -39952
rect -34355 -41400 -29864 -40800
tri -29864 -41400 -29264 -40800 sw
tri -10736 -41400 -10136 -40800 se
rect -10136 -41400 -6600 -40800
tri -34355 -45000 -30755 -41400 ne
rect -30755 -42355 -6600 -41400
tri -6600 -42355 -2400 -38155 nw
rect -30755 -45000 -9245 -42355
tri -9245 -45000 -6600 -42355 nw
<< end >>
