magic
tech sky130A
magscale 1 2
timestamp 1666811438
<< error_p >>
rect -227 3683 -163 3689
rect -97 3683 -33 3689
rect 33 3683 97 3689
rect 163 3683 227 3689
rect -227 3649 -215 3683
rect -97 3649 -85 3683
rect 33 3649 45 3683
rect 163 3649 175 3683
rect -227 3643 -163 3649
rect -97 3643 -33 3649
rect 33 3643 97 3649
rect 163 3643 227 3649
rect -227 -3649 -163 -3643
rect -97 -3649 -33 -3643
rect 33 -3649 97 -3643
rect 163 -3649 227 -3643
rect -227 -3683 -215 -3649
rect -97 -3683 -85 -3649
rect 33 -3683 45 -3649
rect 163 -3683 175 -3649
rect -227 -3689 -163 -3683
rect -97 -3689 -33 -3683
rect 33 -3689 97 -3683
rect 163 -3689 227 -3683
<< nmos >>
rect -231 -3611 -159 3611
rect -101 -3611 -29 3611
rect 29 -3611 101 3611
rect 159 -3611 231 3611
<< ndiff >>
rect -289 3599 -231 3611
rect -289 -3599 -277 3599
rect -243 -3599 -231 3599
rect -289 -3611 -231 -3599
rect -159 3599 -101 3611
rect -159 -3599 -147 3599
rect -113 -3599 -101 3599
rect -159 -3611 -101 -3599
rect -29 3599 29 3611
rect -29 -3599 -17 3599
rect 17 -3599 29 3599
rect -29 -3611 29 -3599
rect 101 3599 159 3611
rect 101 -3599 113 3599
rect 147 -3599 159 3599
rect 101 -3611 159 -3599
rect 231 3599 289 3611
rect 231 -3599 243 3599
rect 277 -3599 289 3599
rect 231 -3611 289 -3599
<< ndiffc >>
rect -277 -3599 -243 3599
rect -147 -3599 -113 3599
rect -17 -3599 17 3599
rect 113 -3599 147 3599
rect 243 -3599 277 3599
<< poly >>
rect -231 3683 -159 3699
rect -231 3649 -215 3683
rect -175 3649 -159 3683
rect -231 3611 -159 3649
rect -101 3683 -29 3699
rect -101 3649 -85 3683
rect -45 3649 -29 3683
rect -101 3611 -29 3649
rect 29 3683 101 3699
rect 29 3649 45 3683
rect 85 3649 101 3683
rect 29 3611 101 3649
rect 159 3683 231 3699
rect 159 3649 175 3683
rect 215 3649 231 3683
rect 159 3611 231 3649
rect -231 -3649 -159 -3611
rect -231 -3683 -215 -3649
rect -175 -3683 -159 -3649
rect -231 -3699 -159 -3683
rect -101 -3649 -29 -3611
rect -101 -3683 -85 -3649
rect -45 -3683 -29 -3649
rect -101 -3699 -29 -3683
rect 29 -3649 101 -3611
rect 29 -3683 45 -3649
rect 85 -3683 101 -3649
rect 29 -3699 101 -3683
rect 159 -3649 231 -3611
rect 159 -3683 175 -3649
rect 215 -3683 231 -3649
rect 159 -3699 231 -3683
<< polycont >>
rect -215 3649 -175 3683
rect -85 3649 -45 3683
rect 45 3649 85 3683
rect 175 3649 215 3683
rect -215 -3683 -175 -3649
rect -85 -3683 -45 -3649
rect 45 -3683 85 -3649
rect 175 -3683 215 -3649
<< locali >>
rect -231 3649 -215 3683
rect -175 3649 -159 3683
rect -101 3649 -85 3683
rect -45 3649 -29 3683
rect 29 3649 45 3683
rect 85 3649 101 3683
rect 159 3649 175 3683
rect 215 3649 231 3683
rect -277 3599 -243 3615
rect -277 -3615 -243 -3599
rect -147 3599 -113 3615
rect -147 -3615 -113 -3599
rect -17 3599 17 3615
rect -17 -3615 17 -3599
rect 113 3599 147 3615
rect 113 -3615 147 -3599
rect 243 3599 277 3615
rect 243 -3615 277 -3599
rect -231 -3683 -215 -3649
rect -175 -3683 -159 -3649
rect -101 -3683 -85 -3649
rect -45 -3683 -29 -3649
rect 29 -3683 45 -3649
rect 85 -3683 101 -3649
rect 159 -3683 175 -3649
rect 215 -3683 231 -3649
<< viali >>
rect -215 3649 -175 3683
rect -85 3649 -45 3683
rect 45 3649 85 3683
rect 175 3649 215 3683
rect -277 -3599 -243 3599
rect -147 -3599 -113 3599
rect -17 -3599 17 3599
rect 113 -3599 147 3599
rect 243 -3599 277 3599
rect -215 -3683 -175 -3649
rect -85 -3683 -45 -3649
rect 45 -3683 85 -3649
rect 175 -3683 215 -3649
<< metal1 >>
rect -227 3683 -163 3689
rect -227 3649 -215 3683
rect -175 3649 -163 3683
rect -227 3643 -163 3649
rect -97 3683 -33 3689
rect -97 3649 -85 3683
rect -45 3649 -33 3683
rect -97 3643 -33 3649
rect 33 3683 97 3689
rect 33 3649 45 3683
rect 85 3649 97 3683
rect 33 3643 97 3649
rect 163 3683 227 3689
rect 163 3649 175 3683
rect 215 3649 227 3683
rect 163 3643 227 3649
rect -283 3599 -237 3611
rect -283 -3599 -277 3599
rect -243 -3599 -237 3599
rect -283 -3611 -237 -3599
rect -153 3599 -107 3611
rect -153 -3599 -147 3599
rect -113 -3599 -107 3599
rect -153 -3611 -107 -3599
rect -23 3599 23 3611
rect -23 -3599 -17 3599
rect 17 -3599 23 3599
rect -23 -3611 23 -3599
rect 107 3599 153 3611
rect 107 -3599 113 3599
rect 147 -3599 153 3599
rect 107 -3611 153 -3599
rect 237 3599 283 3611
rect 237 -3599 243 3599
rect 277 -3599 283 3599
rect 237 -3611 283 -3599
rect -227 -3649 -163 -3643
rect -227 -3683 -215 -3649
rect -175 -3683 -163 -3649
rect -227 -3689 -163 -3683
rect -97 -3649 -33 -3643
rect -97 -3683 -85 -3649
rect -45 -3683 -33 -3649
rect -97 -3689 -33 -3683
rect 33 -3649 97 -3643
rect 33 -3683 45 -3649
rect 85 -3683 97 -3649
rect 33 -3689 97 -3683
rect 163 -3649 227 -3643
rect 163 -3683 175 -3649
rect 215 -3683 227 -3649
rect 163 -3689 227 -3683
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 36.112 l 0.361 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
