magic
tech sky130A
magscale 1 2
timestamp 1666963525
<< nwell >>
rect -396 -1619 396 1619
<< pmos >>
rect -200 -1400 200 1400
<< pdiff >>
rect -258 1388 -200 1400
rect -258 -1388 -246 1388
rect -212 -1388 -200 1388
rect -258 -1400 -200 -1388
rect 200 1388 258 1400
rect 200 -1388 212 1388
rect 246 -1388 258 1388
rect 200 -1400 258 -1388
<< pdiffc >>
rect -246 -1388 -212 1388
rect 212 -1388 246 1388
<< nsubdiff >>
rect -360 1549 -264 1583
rect 264 1549 360 1583
rect -360 1487 -326 1549
rect 326 1487 360 1549
rect -360 -1549 -326 -1487
rect 326 -1549 360 -1487
rect -360 -1583 -264 -1549
rect 264 -1583 360 -1549
<< nsubdiffcont >>
rect -264 1549 264 1583
rect -360 -1487 -326 1487
rect 326 -1487 360 1487
rect -264 -1583 264 -1549
<< poly >>
rect -200 1481 200 1497
rect -200 1447 -184 1481
rect 184 1447 200 1481
rect -200 1400 200 1447
rect -200 -1447 200 -1400
rect -200 -1481 -184 -1447
rect 184 -1481 200 -1447
rect -200 -1497 200 -1481
<< polycont >>
rect -184 1447 184 1481
rect -184 -1481 184 -1447
<< locali >>
rect -360 1549 -264 1583
rect 264 1549 360 1583
rect -360 1487 -326 1549
rect 326 1487 360 1549
rect -200 1447 -184 1481
rect 184 1447 200 1481
rect -246 1388 -212 1404
rect -246 -1404 -212 -1388
rect 212 1388 246 1404
rect 212 -1404 246 -1388
rect -200 -1481 -184 -1447
rect 184 -1481 200 -1447
rect -360 -1549 -326 -1487
rect 326 -1549 360 -1487
rect -360 -1583 -264 -1549
rect 264 -1583 360 -1549
<< viali >>
rect -184 1447 184 1481
rect -246 -1388 -212 1388
rect 212 -1388 246 1388
rect -184 -1481 184 -1447
<< metal1 >>
rect -196 1481 196 1487
rect -196 1447 -184 1481
rect 184 1447 196 1481
rect -196 1441 196 1447
rect -252 1388 -206 1400
rect -252 -1388 -246 1388
rect -212 -1388 -206 1388
rect -252 -1400 -206 -1388
rect 206 1388 252 1400
rect 206 -1388 212 1388
rect 246 -1388 252 1388
rect 206 -1400 252 -1388
rect -196 -1447 196 -1441
rect -196 -1481 -184 -1447
rect 184 -1481 196 -1447
rect -196 -1487 196 -1481
<< properties >>
string FIXED_BBOX -343 -1566 343 1566
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 14.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
