magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 60 35 492
rect -35 -492 35 -60
<< ppolyres >>
rect -35 -60 35 60
<< viali >>
rect -17 438 17 472
rect -17 366 17 400
rect -17 294 17 328
rect -17 222 17 256
rect -17 150 17 184
rect -17 78 17 112
rect -17 -113 17 -79
rect -17 -185 17 -151
rect -17 -257 17 -223
rect -17 -329 17 -295
rect -17 -401 17 -367
rect -17 -473 17 -439
<< metal1 >>
rect -25 472 25 486
rect -25 438 -17 472
rect 17 438 25 472
rect -25 400 25 438
rect -25 366 -17 400
rect 17 366 25 400
rect -25 328 25 366
rect -25 294 -17 328
rect 17 294 25 328
rect -25 256 25 294
rect -25 222 -17 256
rect 17 222 25 256
rect -25 184 25 222
rect -25 150 -17 184
rect 17 150 25 184
rect -25 112 25 150
rect -25 78 -17 112
rect 17 78 25 112
rect -25 65 25 78
rect -25 -79 25 -65
rect -25 -113 -17 -79
rect 17 -113 25 -79
rect -25 -151 25 -113
rect -25 -185 -17 -151
rect 17 -185 25 -151
rect -25 -223 25 -185
rect -25 -257 -17 -223
rect 17 -257 25 -223
rect -25 -295 25 -257
rect -25 -329 -17 -295
rect 17 -329 25 -295
rect -25 -367 25 -329
rect -25 -401 -17 -367
rect 17 -401 25 -367
rect -25 -439 25 -401
rect -25 -473 -17 -439
rect 17 -473 25 -439
rect -25 -486 25 -473
<< end >>
