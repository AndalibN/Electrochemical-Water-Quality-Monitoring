magic
tech sky130A
magscale 1 2
timestamp 1666895121
<< error_p >>
rect -77 512 -31 524
rect 31 512 77 524
rect -77 472 -71 512
rect 31 472 37 512
rect -77 460 -31 472
rect 31 460 77 472
rect -77 108 -31 120
rect 31 108 77 120
rect -77 68 -71 108
rect 31 68 37 108
rect -77 56 -31 68
rect 31 56 77 68
rect -77 -68 -31 -56
rect 31 -68 77 -56
rect -77 -108 -71 -68
rect 31 -108 37 -68
rect -77 -120 -31 -108
rect 31 -120 77 -108
rect -77 -472 -31 -460
rect 31 -472 77 -460
rect -77 -512 -71 -472
rect 31 -512 37 -472
rect -77 -524 -31 -512
rect 31 -524 77 -512
<< pwell >>
rect -253 -694 253 694
<< psubdiff >>
rect -217 624 -121 658
rect 121 624 217 658
rect -217 562 -183 624
rect 183 562 217 624
rect -217 -624 -183 -562
rect 183 -624 217 -562
rect -217 -658 -121 -624
rect 121 -658 217 -624
<< psubdiffcont >>
rect -121 624 121 658
rect -217 -562 -183 562
rect 183 -562 217 562
rect -121 -658 121 -624
<< poly >>
rect -87 512 -21 528
rect -87 478 -71 512
rect -37 478 -21 512
rect -87 455 -21 478
rect -87 102 -21 125
rect -87 68 -71 102
rect -37 68 -21 102
rect -87 52 -21 68
rect 21 512 87 528
rect 21 478 37 512
rect 71 478 87 512
rect 21 455 87 478
rect 21 102 87 125
rect 21 68 37 102
rect 71 68 87 102
rect 21 52 87 68
rect -87 -68 -21 -52
rect -87 -102 -71 -68
rect -37 -102 -21 -68
rect -87 -125 -21 -102
rect -87 -478 -21 -455
rect -87 -512 -71 -478
rect -37 -512 -21 -478
rect -87 -528 -21 -512
rect 21 -68 87 -52
rect 21 -102 37 -68
rect 71 -102 87 -68
rect 21 -125 87 -102
rect 21 -478 87 -455
rect 21 -512 37 -478
rect 71 -512 87 -478
rect 21 -528 87 -512
<< polycont >>
rect -71 478 -37 512
rect -71 68 -37 102
rect 37 478 71 512
rect 37 68 71 102
rect -71 -102 -37 -68
rect -71 -512 -37 -478
rect 37 -102 71 -68
rect 37 -512 71 -478
<< npolyres >>
rect -87 125 -21 455
rect 21 125 87 455
rect -87 -455 -21 -125
rect 21 -455 87 -125
<< locali >>
rect -217 624 -121 658
rect 121 624 217 658
rect -217 562 -183 624
rect 183 562 217 624
rect -87 478 -71 512
rect -37 478 -21 512
rect 21 478 37 512
rect 71 478 87 512
rect -87 68 -71 102
rect -37 68 -21 102
rect 21 68 37 102
rect 71 68 87 102
rect -87 -102 -71 -68
rect -37 -102 -21 -68
rect 21 -102 37 -68
rect 71 -102 87 -68
rect -87 -512 -71 -478
rect -37 -512 -21 -478
rect 21 -512 37 -478
rect 71 -512 87 -478
rect -217 -624 -183 -562
rect 183 -624 217 -562
rect -217 -658 -121 -624
rect 121 -658 217 -624
<< viali >>
rect -71 478 -37 512
rect 37 478 71 512
rect -71 472 -37 478
rect 37 472 71 478
rect -71 102 -37 108
rect 37 102 71 108
rect -71 68 -37 102
rect 37 68 71 102
rect -71 -102 -37 -68
rect 37 -102 71 -68
rect -71 -108 -37 -102
rect 37 -108 71 -102
rect -71 -478 -37 -472
rect 37 -478 71 -472
rect -71 -512 -37 -478
rect 37 -512 71 -478
<< metal1 >>
rect -77 512 -31 524
rect -77 472 -71 512
rect -37 472 -31 512
rect -77 460 -31 472
rect 31 512 77 524
rect 31 472 37 512
rect 71 472 77 512
rect 31 460 77 472
rect -77 108 -31 120
rect -77 68 -71 108
rect -37 68 -31 108
rect -77 56 -31 68
rect 31 108 77 120
rect 31 68 37 108
rect 71 68 77 108
rect 31 56 77 68
rect -77 -68 -31 -56
rect -77 -108 -71 -68
rect -37 -108 -31 -68
rect -77 -120 -31 -108
rect 31 -68 77 -56
rect 31 -108 37 -68
rect 71 -108 77 -68
rect 31 -120 77 -108
rect -77 -472 -31 -460
rect -77 -512 -71 -472
rect -37 -512 -31 -472
rect -77 -524 -31 -512
rect 31 -472 77 -460
rect 31 -512 37 -472
rect 71 -512 77 -472
rect 31 -524 77 -512
<< properties >>
string FIXED_BBOX -200 -641 200 641
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 1.650 m 2 nx 2 wmin 0.330 lmin 1.650 rho 48.2 val 241.0 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
