magic
tech sky130A
magscale 1 2
timestamp 1668702877
<< error_p >>
rect -29 4272 29 4278
rect -29 4238 -17 4272
rect -29 4232 29 4238
rect -29 -4238 29 -4232
rect -29 -4272 -17 -4238
rect -29 -4278 29 -4272
<< pwell >>
rect -226 -4410 226 4410
<< nmos >>
rect -30 -4200 30 4200
<< ndiff >>
rect -88 4188 -30 4200
rect -88 -4188 -76 4188
rect -42 -4188 -30 4188
rect -88 -4200 -30 -4188
rect 30 4188 88 4200
rect 30 -4188 42 4188
rect 76 -4188 88 4188
rect 30 -4200 88 -4188
<< ndiffc >>
rect -76 -4188 -42 4188
rect 42 -4188 76 4188
<< psubdiff >>
rect -190 4340 -94 4374
rect 94 4340 190 4374
rect -190 4278 -156 4340
rect 156 4278 190 4340
rect -190 -4340 -156 -4278
rect 156 -4340 190 -4278
rect -190 -4374 -94 -4340
rect 94 -4374 190 -4340
<< psubdiffcont >>
rect -94 4340 94 4374
rect -190 -4278 -156 4278
rect 156 -4278 190 4278
rect -94 -4374 94 -4340
<< poly >>
rect -33 4272 33 4288
rect -33 4238 -17 4272
rect 17 4238 33 4272
rect -33 4222 33 4238
rect -30 4200 30 4222
rect -30 -4222 30 -4200
rect -33 -4238 33 -4222
rect -33 -4272 -17 -4238
rect 17 -4272 33 -4238
rect -33 -4288 33 -4272
<< polycont >>
rect -17 4238 17 4272
rect -17 -4272 17 -4238
<< locali >>
rect -190 4340 -94 4374
rect 94 4340 190 4374
rect -190 4278 -156 4340
rect 156 4278 190 4340
rect -33 4238 -17 4272
rect 17 4238 33 4272
rect -76 4188 -42 4204
rect -76 -4204 -42 -4188
rect 42 4188 76 4204
rect 42 -4204 76 -4188
rect -33 -4272 -17 -4238
rect 17 -4272 33 -4238
rect -190 -4340 -156 -4278
rect 156 -4340 190 -4278
rect -190 -4374 -94 -4340
rect 94 -4374 190 -4340
<< viali >>
rect -17 4238 17 4272
rect -76 -4188 -42 4188
rect 42 -4188 76 4188
rect -17 -4272 17 -4238
<< metal1 >>
rect -29 4272 29 4278
rect -29 4238 -17 4272
rect 17 4238 29 4272
rect -29 4232 29 4238
rect -82 4188 -36 4200
rect -82 -4188 -76 4188
rect -42 -4188 -36 4188
rect -82 -4200 -36 -4188
rect 36 4188 82 4200
rect 36 -4188 42 4188
rect 76 -4188 82 4188
rect 36 -4200 82 -4188
rect -29 -4238 29 -4232
rect -29 -4272 -17 -4238
rect 17 -4272 29 -4238
rect -29 -4278 29 -4272
<< properties >>
string FIXED_BBOX -173 -4357 173 4357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 42.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
