magic
tech sky130A
magscale 1 2
timestamp 1667977299
<< pwell >>
rect -226 -510 226 510
<< nmos >>
rect -30 -300 30 300
<< ndiff >>
rect -88 288 -30 300
rect -88 -288 -76 288
rect -42 -288 -30 288
rect -88 -300 -30 -288
rect 30 288 88 300
rect 30 -288 42 288
rect 76 -288 88 288
rect 30 -300 88 -288
<< ndiffc >>
rect -76 -288 -42 288
rect 42 -288 76 288
<< psubdiff >>
rect -190 440 -94 474
rect 94 440 190 474
rect -190 378 -156 440
rect 156 378 190 440
rect -190 -440 -156 -378
rect 156 -440 190 -378
rect -190 -474 -94 -440
rect 94 -474 190 -440
<< psubdiffcont >>
rect -94 440 94 474
rect -190 -378 -156 378
rect 156 -378 190 378
rect -94 -474 94 -440
<< poly >>
rect -33 372 33 388
rect -33 338 -17 372
rect 17 338 33 372
rect -33 322 33 338
rect -30 300 30 322
rect -30 -322 30 -300
rect -33 -338 33 -322
rect -33 -372 -17 -338
rect 17 -372 33 -338
rect -33 -388 33 -372
<< polycont >>
rect -17 338 17 372
rect -17 -372 17 -338
<< locali >>
rect -190 440 -94 474
rect 94 440 190 474
rect -190 378 -156 440
rect 156 378 190 440
rect -33 338 -17 372
rect 17 338 33 372
rect -76 288 -42 304
rect -76 -304 -42 -288
rect 42 288 76 304
rect 42 -304 76 -288
rect -33 -372 -17 -338
rect 17 -372 33 -338
rect -190 -440 -156 -378
rect 156 -440 190 -378
rect -190 -474 -94 -440
rect 94 -474 190 -440
<< viali >>
rect -17 338 17 372
rect -76 -288 -42 288
rect 42 -288 76 288
rect -17 -372 17 -338
<< metal1 >>
rect -29 372 29 378
rect -29 338 -17 372
rect 17 338 29 372
rect -29 332 29 338
rect -82 288 -36 300
rect -82 -288 -76 288
rect -42 -288 -36 288
rect -82 -300 -36 -288
rect 36 288 82 300
rect 36 -288 42 288
rect 76 -288 82 288
rect 36 -300 82 -288
rect -29 -338 29 -332
rect -29 -372 -17 -338
rect 17 -372 29 -338
rect -29 -378 29 -372
<< properties >>
string FIXED_BBOX -173 -457 173 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
