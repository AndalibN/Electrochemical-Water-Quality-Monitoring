magic
tech sky130A
magscale 1 2
timestamp 1667937831
<< error_p >>
rect -88 345 -30 351
rect 30 345 88 351
rect -88 311 -76 345
rect 30 311 42 345
rect -88 305 -30 311
rect 30 305 88 311
<< nwell >>
rect -183 -398 183 364
<< pmos >>
rect -89 -336 -29 264
rect 29 -336 89 264
<< pdiff >>
rect -147 252 -89 264
rect -147 -324 -135 252
rect -101 -324 -89 252
rect -147 -336 -89 -324
rect -29 252 29 264
rect -29 -324 -17 252
rect 17 -324 29 252
rect -29 -336 29 -324
rect 89 252 147 264
rect 89 -324 101 252
rect 135 -324 147 252
rect 89 -336 147 -324
<< pdiffc >>
rect -135 -324 -101 252
rect -17 -324 17 252
rect 101 -324 135 252
<< poly >>
rect -92 345 -26 361
rect -92 311 -76 345
rect -42 311 -26 345
rect -92 295 -26 311
rect 26 345 92 361
rect 26 311 42 345
rect 76 311 92 345
rect 26 295 92 311
rect -89 264 -29 295
rect 29 264 89 295
rect -89 -362 -29 -336
rect 29 -362 89 -336
<< polycont >>
rect -76 311 -42 345
rect 42 311 76 345
<< locali >>
rect -92 311 -76 345
rect -42 311 -26 345
rect 26 311 42 345
rect 76 311 92 345
rect -135 252 -101 268
rect -135 -340 -101 -324
rect -17 252 17 268
rect -17 -340 17 -324
rect 101 252 135 268
rect 101 -340 135 -324
<< viali >>
rect -76 311 -42 345
rect 42 311 76 345
rect -135 -324 -101 252
rect -17 -324 17 252
rect 101 -324 135 252
<< metal1 >>
rect -88 345 -30 351
rect -88 311 -76 345
rect -42 311 -30 345
rect -88 305 -30 311
rect 30 345 88 351
rect 30 311 42 345
rect 76 311 88 345
rect 30 305 88 311
rect -141 252 -95 264
rect -141 -324 -135 252
rect -101 -324 -95 252
rect -141 -336 -95 -324
rect -23 252 23 264
rect -23 -324 -17 252
rect 17 -324 23 252
rect -23 -336 23 -324
rect 95 252 141 264
rect 95 -324 101 252
rect 135 -324 141 252
rect 95 -336 141 -324
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3 l 0.30 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
