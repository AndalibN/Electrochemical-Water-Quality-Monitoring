magic
tech sky130A
magscale 1 2
timestamp 1666968066
<< nwell >>
rect -1094 -1064 1094 1098
<< pmos >>
rect -1000 -964 1000 1036
<< pdiff >>
rect -1058 1024 -1000 1036
rect -1058 -952 -1046 1024
rect -1012 -952 -1000 1024
rect -1058 -964 -1000 -952
rect 1000 1024 1058 1036
rect 1000 -952 1012 1024
rect 1046 -952 1058 1024
rect 1000 -964 1058 -952
<< pdiffc >>
rect -1046 -952 -1012 1024
rect 1012 -952 1046 1024
<< poly >>
rect -1000 1036 1000 1062
rect -1000 -1011 1000 -964
rect -1000 -1045 -984 -1011
rect 984 -1045 1000 -1011
rect -1000 -1061 1000 -1045
<< polycont >>
rect -984 -1045 984 -1011
<< locali >>
rect -1046 1024 -1012 1040
rect -1046 -968 -1012 -952
rect 1012 1024 1046 1040
rect 1012 -968 1046 -952
rect -1000 -1045 -984 -1011
rect 984 -1045 1000 -1011
<< viali >>
rect -1046 -952 -1012 1024
rect 1012 -952 1046 1024
rect -984 -1045 984 -1011
<< metal1 >>
rect -1052 1024 -1006 1036
rect -1052 -952 -1046 1024
rect -1012 -952 -1006 1024
rect -1052 -964 -1006 -952
rect 1006 1024 1052 1036
rect 1006 -952 1012 1024
rect 1046 -952 1052 1024
rect 1006 -964 1052 -952
rect -996 -1011 996 -1005
rect -996 -1045 -984 -1011
rect 984 -1045 996 -1011
rect -996 -1051 996 -1045
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
