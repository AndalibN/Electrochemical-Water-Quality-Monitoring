magic
tech sky130A
magscale 1 2
timestamp 1666802529
<< checkpaint >>
rect 96 4395 5491 4927
rect -1260 -660 5491 4395
rect -1260 -2460 1460 -660
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_GDJJ3U  XXM1
timestamp 1666802528
transform 1 0 53 0 1 1800
box -53 -1200 409 1335
use sky130_fd_pr__pfet_01v8_RWVM3U  XXM2
timestamp 1666802528
transform 1 0 515 0 1 1800
box -53 -1200 409 1335
use sky130_fd_pr__nfet_01v8_S4GQ7J  XXM3
timestamp 1666802528
transform 1 0 977 0 1 1800
box -53 -1200 379 1067
use sky130_fd_pr__nfet_01v8_QY8CNP  XXM4
timestamp 1666802528
transform 1 0 1409 0 1 2600
box -53 -2000 758 1067
use sky130_fd_pr__pfet_01v8_79XL75  XXM5
timestamp 1666802529
transform 1 0 2220 0 1 1800
box -53 -1200 409 1335
use sky130_fd_pr__nfet_01v8_Y6ED9L  XXM6
timestamp 1666802529
transform 1 0 2682 0 1 2600
box -53 -2000 758 1067
use sky130_fd_pr__nfet_01v8_75NWZG  XXM7
timestamp 1666802529
transform 1 0 3493 0 1 2600
box -53 -2000 738 1067
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 In
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 GND
port 3 nsew
<< end >>
