magic
tech sky130A
magscale 1 2
timestamp 1667856991
<< error_p >>
rect -2259 2210 -2199 3550
rect -2179 2210 -2119 3550
rect -800 2210 -740 3550
rect -720 2210 -660 3550
rect 659 2210 719 3550
rect 739 2210 799 3550
rect 2118 2210 2178 3550
rect 2198 2210 2258 3550
rect -2259 770 -2199 2110
rect -2179 770 -2119 2110
rect -800 770 -740 2110
rect -720 770 -660 2110
rect 659 770 719 2110
rect 739 770 799 2110
rect 2118 770 2178 2110
rect 2198 770 2258 2110
rect -2259 -670 -2199 670
rect -2179 -670 -2119 670
rect -800 -670 -740 670
rect -720 -670 -660 670
rect 659 -670 719 670
rect 739 -670 799 670
rect 2118 -670 2178 670
rect 2198 -670 2258 670
rect -2259 -2110 -2199 -770
rect -2179 -2110 -2119 -770
rect -800 -2110 -740 -770
rect -720 -2110 -660 -770
rect 659 -2110 719 -770
rect 739 -2110 799 -770
rect 2118 -2110 2178 -770
rect 2198 -2110 2258 -770
rect -2259 -3550 -2199 -2210
rect -2179 -3550 -2119 -2210
rect -800 -3550 -740 -2210
rect -720 -3550 -660 -2210
rect 659 -3550 719 -2210
rect 739 -3550 799 -2210
rect 2118 -3550 2178 -2210
rect 2198 -3550 2258 -2210
<< metal3 >>
rect -3638 3522 -2199 3550
rect -3638 2238 -2283 3522
rect -2219 2238 -2199 3522
rect -3638 2210 -2199 2238
rect -2179 3522 -740 3550
rect -2179 2238 -824 3522
rect -760 2238 -740 3522
rect -2179 2210 -740 2238
rect -720 3522 719 3550
rect -720 2238 635 3522
rect 699 2238 719 3522
rect -720 2210 719 2238
rect 739 3522 2178 3550
rect 739 2238 2094 3522
rect 2158 2238 2178 3522
rect 739 2210 2178 2238
rect 2198 3522 3637 3550
rect 2198 2238 3553 3522
rect 3617 2238 3637 3522
rect 2198 2210 3637 2238
rect -3638 2082 -2199 2110
rect -3638 798 -2283 2082
rect -2219 798 -2199 2082
rect -3638 770 -2199 798
rect -2179 2082 -740 2110
rect -2179 798 -824 2082
rect -760 798 -740 2082
rect -2179 770 -740 798
rect -720 2082 719 2110
rect -720 798 635 2082
rect 699 798 719 2082
rect -720 770 719 798
rect 739 2082 2178 2110
rect 739 798 2094 2082
rect 2158 798 2178 2082
rect 739 770 2178 798
rect 2198 2082 3637 2110
rect 2198 798 3553 2082
rect 3617 798 3637 2082
rect 2198 770 3637 798
rect -3638 642 -2199 670
rect -3638 -642 -2283 642
rect -2219 -642 -2199 642
rect -3638 -670 -2199 -642
rect -2179 642 -740 670
rect -2179 -642 -824 642
rect -760 -642 -740 642
rect -2179 -670 -740 -642
rect -720 642 719 670
rect -720 -642 635 642
rect 699 -642 719 642
rect -720 -670 719 -642
rect 739 642 2178 670
rect 739 -642 2094 642
rect 2158 -642 2178 642
rect 739 -670 2178 -642
rect 2198 642 3637 670
rect 2198 -642 3553 642
rect 3617 -642 3637 642
rect 2198 -670 3637 -642
rect -3638 -798 -2199 -770
rect -3638 -2082 -2283 -798
rect -2219 -2082 -2199 -798
rect -3638 -2110 -2199 -2082
rect -2179 -798 -740 -770
rect -2179 -2082 -824 -798
rect -760 -2082 -740 -798
rect -2179 -2110 -740 -2082
rect -720 -798 719 -770
rect -720 -2082 635 -798
rect 699 -2082 719 -798
rect -720 -2110 719 -2082
rect 739 -798 2178 -770
rect 739 -2082 2094 -798
rect 2158 -2082 2178 -798
rect 739 -2110 2178 -2082
rect 2198 -798 3637 -770
rect 2198 -2082 3553 -798
rect 3617 -2082 3637 -798
rect 2198 -2110 3637 -2082
rect -3638 -2238 -2199 -2210
rect -3638 -3522 -2283 -2238
rect -2219 -3522 -2199 -2238
rect -3638 -3550 -2199 -3522
rect -2179 -2238 -740 -2210
rect -2179 -3522 -824 -2238
rect -760 -3522 -740 -2238
rect -2179 -3550 -740 -3522
rect -720 -2238 719 -2210
rect -720 -3522 635 -2238
rect 699 -3522 719 -2238
rect -720 -3550 719 -3522
rect 739 -2238 2178 -2210
rect 739 -3522 2094 -2238
rect 2158 -3522 2178 -2238
rect 739 -3550 2178 -3522
rect 2198 -2238 3637 -2210
rect 2198 -3522 3553 -2238
rect 3617 -3522 3637 -2238
rect 2198 -3550 3637 -3522
<< via3 >>
rect -2283 2238 -2219 3522
rect -824 2238 -760 3522
rect 635 2238 699 3522
rect 2094 2238 2158 3522
rect 3553 2238 3617 3522
rect -2283 798 -2219 2082
rect -824 798 -760 2082
rect 635 798 699 2082
rect 2094 798 2158 2082
rect 3553 798 3617 2082
rect -2283 -642 -2219 642
rect -824 -642 -760 642
rect 635 -642 699 642
rect 2094 -642 2158 642
rect 3553 -642 3617 642
rect -2283 -2082 -2219 -798
rect -824 -2082 -760 -798
rect 635 -2082 699 -798
rect 2094 -2082 2158 -798
rect 3553 -2082 3617 -798
rect -2283 -3522 -2219 -2238
rect -824 -3522 -760 -2238
rect 635 -3522 699 -2238
rect 2094 -3522 2158 -2238
rect 3553 -3522 3617 -2238
<< mimcap >>
rect -3538 3410 -2398 3450
rect -3538 2350 -3498 3410
rect -2438 2350 -2398 3410
rect -3538 2310 -2398 2350
rect -2079 3410 -939 3450
rect -2079 2350 -2039 3410
rect -979 2350 -939 3410
rect -2079 2310 -939 2350
rect -620 3410 520 3450
rect -620 2350 -580 3410
rect 480 2350 520 3410
rect -620 2310 520 2350
rect 839 3410 1979 3450
rect 839 2350 879 3410
rect 1939 2350 1979 3410
rect 839 2310 1979 2350
rect 2298 3410 3438 3450
rect 2298 2350 2338 3410
rect 3398 2350 3438 3410
rect 2298 2310 3438 2350
rect -3538 1970 -2398 2010
rect -3538 910 -3498 1970
rect -2438 910 -2398 1970
rect -3538 870 -2398 910
rect -2079 1970 -939 2010
rect -2079 910 -2039 1970
rect -979 910 -939 1970
rect -2079 870 -939 910
rect -620 1970 520 2010
rect -620 910 -580 1970
rect 480 910 520 1970
rect -620 870 520 910
rect 839 1970 1979 2010
rect 839 910 879 1970
rect 1939 910 1979 1970
rect 839 870 1979 910
rect 2298 1970 3438 2010
rect 2298 910 2338 1970
rect 3398 910 3438 1970
rect 2298 870 3438 910
rect -3538 530 -2398 570
rect -3538 -530 -3498 530
rect -2438 -530 -2398 530
rect -3538 -570 -2398 -530
rect -2079 530 -939 570
rect -2079 -530 -2039 530
rect -979 -530 -939 530
rect -2079 -570 -939 -530
rect -620 530 520 570
rect -620 -530 -580 530
rect 480 -530 520 530
rect -620 -570 520 -530
rect 839 530 1979 570
rect 839 -530 879 530
rect 1939 -530 1979 530
rect 839 -570 1979 -530
rect 2298 530 3438 570
rect 2298 -530 2338 530
rect 3398 -530 3438 530
rect 2298 -570 3438 -530
rect -3538 -910 -2398 -870
rect -3538 -1970 -3498 -910
rect -2438 -1970 -2398 -910
rect -3538 -2010 -2398 -1970
rect -2079 -910 -939 -870
rect -2079 -1970 -2039 -910
rect -979 -1970 -939 -910
rect -2079 -2010 -939 -1970
rect -620 -910 520 -870
rect -620 -1970 -580 -910
rect 480 -1970 520 -910
rect -620 -2010 520 -1970
rect 839 -910 1979 -870
rect 839 -1970 879 -910
rect 1939 -1970 1979 -910
rect 839 -2010 1979 -1970
rect 2298 -910 3438 -870
rect 2298 -1970 2338 -910
rect 3398 -1970 3438 -910
rect 2298 -2010 3438 -1970
rect -3538 -2350 -2398 -2310
rect -3538 -3410 -3498 -2350
rect -2438 -3410 -2398 -2350
rect -3538 -3450 -2398 -3410
rect -2079 -2350 -939 -2310
rect -2079 -3410 -2039 -2350
rect -979 -3410 -939 -2350
rect -2079 -3450 -939 -3410
rect -620 -2350 520 -2310
rect -620 -3410 -580 -2350
rect 480 -3410 520 -2350
rect -620 -3450 520 -3410
rect 839 -2350 1979 -2310
rect 839 -3410 879 -2350
rect 1939 -3410 1979 -2350
rect 839 -3450 1979 -3410
rect 2298 -2350 3438 -2310
rect 2298 -3410 2338 -2350
rect 3398 -3410 3438 -2350
rect 2298 -3450 3438 -3410
<< mimcapcontact >>
rect -3498 2350 -2438 3410
rect -2039 2350 -979 3410
rect -580 2350 480 3410
rect 879 2350 1939 3410
rect 2338 2350 3398 3410
rect -3498 910 -2438 1970
rect -2039 910 -979 1970
rect -580 910 480 1970
rect 879 910 1939 1970
rect 2338 910 3398 1970
rect -3498 -530 -2438 530
rect -2039 -530 -979 530
rect -580 -530 480 530
rect 879 -530 1939 530
rect 2338 -530 3398 530
rect -3498 -1970 -2438 -910
rect -2039 -1970 -979 -910
rect -580 -1970 480 -910
rect 879 -1970 1939 -910
rect 2338 -1970 3398 -910
rect -3498 -3410 -2438 -2350
rect -2039 -3410 -979 -2350
rect -580 -3410 480 -2350
rect 879 -3410 1939 -2350
rect 2338 -3410 3398 -2350
<< metal4 >>
rect -3020 3411 -2916 3600
rect -2330 3538 -2226 3600
rect -2330 3522 -2203 3538
rect -3499 3410 -2437 3411
rect -3499 2350 -3498 3410
rect -2438 2350 -2437 3410
rect -3499 2349 -2437 2350
rect -3020 1971 -2916 2349
rect -2330 2238 -2283 3522
rect -2219 2238 -2203 3522
rect -1561 3411 -1457 3600
rect -871 3538 -767 3600
rect -871 3522 -744 3538
rect -2040 3410 -978 3411
rect -2040 2350 -2039 3410
rect -979 2350 -978 3410
rect -2040 2349 -978 2350
rect -2330 2222 -2203 2238
rect -2330 2098 -2226 2222
rect -2330 2082 -2203 2098
rect -3499 1970 -2437 1971
rect -3499 910 -3498 1970
rect -2438 910 -2437 1970
rect -3499 909 -2437 910
rect -3020 531 -2916 909
rect -2330 798 -2283 2082
rect -2219 798 -2203 2082
rect -1561 1971 -1457 2349
rect -871 2238 -824 3522
rect -760 2238 -744 3522
rect -102 3411 2 3600
rect 588 3538 692 3600
rect 588 3522 715 3538
rect -581 3410 481 3411
rect -581 2350 -580 3410
rect 480 2350 481 3410
rect -581 2349 481 2350
rect -871 2222 -744 2238
rect -871 2098 -767 2222
rect -871 2082 -744 2098
rect -2040 1970 -978 1971
rect -2040 910 -2039 1970
rect -979 910 -978 1970
rect -2040 909 -978 910
rect -2330 782 -2203 798
rect -2330 658 -2226 782
rect -2330 642 -2203 658
rect -3499 530 -2437 531
rect -3499 -530 -3498 530
rect -2438 -530 -2437 530
rect -3499 -531 -2437 -530
rect -3020 -909 -2916 -531
rect -2330 -642 -2283 642
rect -2219 -642 -2203 642
rect -1561 531 -1457 909
rect -871 798 -824 2082
rect -760 798 -744 2082
rect -102 1971 2 2349
rect 588 2238 635 3522
rect 699 2238 715 3522
rect 1357 3411 1461 3600
rect 2047 3538 2151 3600
rect 2047 3522 2174 3538
rect 878 3410 1940 3411
rect 878 2350 879 3410
rect 1939 2350 1940 3410
rect 878 2349 1940 2350
rect 588 2222 715 2238
rect 588 2098 692 2222
rect 588 2082 715 2098
rect -581 1970 481 1971
rect -581 910 -580 1970
rect 480 910 481 1970
rect -581 909 481 910
rect -871 782 -744 798
rect -871 658 -767 782
rect -871 642 -744 658
rect -2040 530 -978 531
rect -2040 -530 -2039 530
rect -979 -530 -978 530
rect -2040 -531 -978 -530
rect -2330 -658 -2203 -642
rect -2330 -782 -2226 -658
rect -2330 -798 -2203 -782
rect -3499 -910 -2437 -909
rect -3499 -1970 -3498 -910
rect -2438 -1970 -2437 -910
rect -3499 -1971 -2437 -1970
rect -3020 -2349 -2916 -1971
rect -2330 -2082 -2283 -798
rect -2219 -2082 -2203 -798
rect -1561 -909 -1457 -531
rect -871 -642 -824 642
rect -760 -642 -744 642
rect -102 531 2 909
rect 588 798 635 2082
rect 699 798 715 2082
rect 1357 1971 1461 2349
rect 2047 2238 2094 3522
rect 2158 2238 2174 3522
rect 2816 3411 2920 3600
rect 3506 3538 3610 3600
rect 3506 3522 3633 3538
rect 2337 3410 3399 3411
rect 2337 2350 2338 3410
rect 3398 2350 3399 3410
rect 2337 2349 3399 2350
rect 2047 2222 2174 2238
rect 2047 2098 2151 2222
rect 2047 2082 2174 2098
rect 878 1970 1940 1971
rect 878 910 879 1970
rect 1939 910 1940 1970
rect 878 909 1940 910
rect 588 782 715 798
rect 588 658 692 782
rect 588 642 715 658
rect -581 530 481 531
rect -581 -530 -580 530
rect 480 -530 481 530
rect -581 -531 481 -530
rect -871 -658 -744 -642
rect -871 -782 -767 -658
rect -871 -798 -744 -782
rect -2040 -910 -978 -909
rect -2040 -1970 -2039 -910
rect -979 -1970 -978 -910
rect -2040 -1971 -978 -1970
rect -2330 -2098 -2203 -2082
rect -2330 -2222 -2226 -2098
rect -2330 -2238 -2203 -2222
rect -3499 -2350 -2437 -2349
rect -3499 -3410 -3498 -2350
rect -2438 -3410 -2437 -2350
rect -3499 -3411 -2437 -3410
rect -3020 -3600 -2916 -3411
rect -2330 -3522 -2283 -2238
rect -2219 -3522 -2203 -2238
rect -1561 -2349 -1457 -1971
rect -871 -2082 -824 -798
rect -760 -2082 -744 -798
rect -102 -909 2 -531
rect 588 -642 635 642
rect 699 -642 715 642
rect 1357 531 1461 909
rect 2047 798 2094 2082
rect 2158 798 2174 2082
rect 2816 1971 2920 2349
rect 3506 2238 3553 3522
rect 3617 2238 3633 3522
rect 3506 2222 3633 2238
rect 3506 2098 3610 2222
rect 3506 2082 3633 2098
rect 2337 1970 3399 1971
rect 2337 910 2338 1970
rect 3398 910 3399 1970
rect 2337 909 3399 910
rect 2047 782 2174 798
rect 2047 658 2151 782
rect 2047 642 2174 658
rect 878 530 1940 531
rect 878 -530 879 530
rect 1939 -530 1940 530
rect 878 -531 1940 -530
rect 588 -658 715 -642
rect 588 -782 692 -658
rect 588 -798 715 -782
rect -581 -910 481 -909
rect -581 -1970 -580 -910
rect 480 -1970 481 -910
rect -581 -1971 481 -1970
rect -871 -2098 -744 -2082
rect -871 -2222 -767 -2098
rect -871 -2238 -744 -2222
rect -2040 -2350 -978 -2349
rect -2040 -3410 -2039 -2350
rect -979 -3410 -978 -2350
rect -2040 -3411 -978 -3410
rect -2330 -3538 -2203 -3522
rect -2330 -3600 -2226 -3538
rect -1561 -3600 -1457 -3411
rect -871 -3522 -824 -2238
rect -760 -3522 -744 -2238
rect -102 -2349 2 -1971
rect 588 -2082 635 -798
rect 699 -2082 715 -798
rect 1357 -909 1461 -531
rect 2047 -642 2094 642
rect 2158 -642 2174 642
rect 2816 531 2920 909
rect 3506 798 3553 2082
rect 3617 798 3633 2082
rect 3506 782 3633 798
rect 3506 658 3610 782
rect 3506 642 3633 658
rect 2337 530 3399 531
rect 2337 -530 2338 530
rect 3398 -530 3399 530
rect 2337 -531 3399 -530
rect 2047 -658 2174 -642
rect 2047 -782 2151 -658
rect 2047 -798 2174 -782
rect 878 -910 1940 -909
rect 878 -1970 879 -910
rect 1939 -1970 1940 -910
rect 878 -1971 1940 -1970
rect 588 -2098 715 -2082
rect 588 -2222 692 -2098
rect 588 -2238 715 -2222
rect -581 -2350 481 -2349
rect -581 -3410 -580 -2350
rect 480 -3410 481 -2350
rect -581 -3411 481 -3410
rect -871 -3538 -744 -3522
rect -871 -3600 -767 -3538
rect -102 -3600 2 -3411
rect 588 -3522 635 -2238
rect 699 -3522 715 -2238
rect 1357 -2349 1461 -1971
rect 2047 -2082 2094 -798
rect 2158 -2082 2174 -798
rect 2816 -909 2920 -531
rect 3506 -642 3553 642
rect 3617 -642 3633 642
rect 3506 -658 3633 -642
rect 3506 -782 3610 -658
rect 3506 -798 3633 -782
rect 2337 -910 3399 -909
rect 2337 -1970 2338 -910
rect 3398 -1970 3399 -910
rect 2337 -1971 3399 -1970
rect 2047 -2098 2174 -2082
rect 2047 -2222 2151 -2098
rect 2047 -2238 2174 -2222
rect 878 -2350 1940 -2349
rect 878 -3410 879 -2350
rect 1939 -3410 1940 -2350
rect 878 -3411 1940 -3410
rect 588 -3538 715 -3522
rect 588 -3600 692 -3538
rect 1357 -3600 1461 -3411
rect 2047 -3522 2094 -2238
rect 2158 -3522 2174 -2238
rect 2816 -2349 2920 -1971
rect 3506 -2082 3553 -798
rect 3617 -2082 3633 -798
rect 3506 -2098 3633 -2082
rect 3506 -2222 3610 -2098
rect 3506 -2238 3633 -2222
rect 2337 -2350 3399 -2349
rect 2337 -3410 2338 -2350
rect 3398 -3410 3399 -2350
rect 2337 -3411 3399 -3410
rect 2047 -3538 2174 -3522
rect 2047 -3600 2151 -3538
rect 2816 -3600 2920 -3411
rect 3506 -3522 3553 -2238
rect 3617 -3522 3633 -2238
rect 3506 -3538 3633 -3522
rect 3506 -3600 3610 -3538
<< properties >>
string FIXED_BBOX 2198 2210 3538 3550
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5.7 l 5.7 val 69.312 carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
