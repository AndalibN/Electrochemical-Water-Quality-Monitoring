magic
tech sky130A
magscale 1 2
timestamp 1669223049
<< error_s >>
rect 5536 2572 41834 2606
rect 5440 520 5474 2510
rect 5536 424 41834 458
<< nwell >>
rect 15505 14880 20461 15135
rect 15504 14810 20461 14880
rect 15504 12624 20455 14810
rect 5395 10446 10351 10701
rect 10738 10558 10843 10560
rect 11140 10558 11310 10597
rect 10724 10468 10725 10558
rect 10736 10470 11310 10558
rect 10736 10468 10843 10470
rect 5395 10376 10352 10446
rect 5401 8190 10352 10376
rect 10724 8625 10843 10468
rect 11140 10443 11310 10470
rect 11151 10437 11261 10443
rect 11151 8625 11260 10437
rect 16402 8710 17024 9416
rect 10724 8547 11261 8625
rect 10739 8544 11261 8547
rect 10703 6261 11317 7604
rect 16396 7314 17018 8020
rect 17368 7809 18302 9465
rect 19869 8705 20491 9411
rect 19865 7374 20487 8080
rect 10764 5647 11317 6261
rect 19883 6132 20505 6838
rect 10703 5507 11317 5647
rect 12956 5388 15053 6002
rect 15026 2643 16162 2647
rect 15024 2642 16162 2643
<< psubdiff >>
rect 11788 14794 14530 15044
rect 11788 14792 12164 14794
rect 11788 12961 12152 14792
rect 11788 12375 12151 12961
rect 11788 12374 12164 12375
rect 14218 12374 14530 14794
rect 11788 12046 14530 12374
rect 15681 11953 20257 11990
rect 10751 11159 11240 11180
rect 10751 10687 10776 11159
rect 10836 11092 11155 11110
rect 10836 10756 10860 11092
rect 11131 10756 11155 11092
rect 10836 10736 11155 10756
rect 11215 10687 11240 11159
rect 15681 10808 15716 11953
rect 15828 11804 20114 11840
rect 15828 10967 15855 11804
rect 20090 10967 20114 11804
rect 15828 10934 20114 10967
rect 20230 10808 20257 11953
rect 15681 10781 20257 10808
rect 10751 10668 11240 10687
rect 16348 9878 16980 9908
rect 16348 9843 16381 9878
rect 16348 9464 16382 9843
rect 16443 9821 16882 9843
rect 16443 9524 16480 9821
rect 16848 9524 16882 9821
rect 16443 9505 16882 9524
rect 16943 9464 16980 9878
rect 16348 9442 16980 9464
rect 19815 9874 20447 9904
rect 19815 9839 19848 9874
rect 19815 9460 19849 9839
rect 19910 9817 20349 9839
rect 19910 9520 19947 9817
rect 20315 9520 20349 9817
rect 19910 9501 20349 9520
rect 20410 9460 20447 9874
rect 19815 9438 20447 9460
rect 16344 8483 16976 8513
rect 16344 8448 16377 8483
rect 10753 8162 11242 8183
rect 10753 7690 10778 8162
rect 10838 8095 11157 8113
rect 10838 7759 10862 8095
rect 11133 7759 11157 8095
rect 10838 7739 11157 7759
rect 11217 7690 11242 8162
rect 16344 8069 16378 8448
rect 16439 8426 16878 8448
rect 16439 8129 16476 8426
rect 16844 8129 16878 8426
rect 16439 8110 16878 8129
rect 16939 8069 16976 8483
rect 16344 8047 16976 8069
rect 10753 7671 11242 7690
rect 5602 7519 10178 7556
rect 5602 6374 5629 7519
rect 5745 7370 10031 7406
rect 5745 6533 5769 7370
rect 10004 6533 10031 7370
rect 5745 6500 10031 6533
rect 10143 6374 10178 7519
rect 5602 6347 10178 6374
rect 18529 9408 19439 9428
rect 18529 7956 18553 9408
rect 18589 9407 19379 9408
rect 18528 7872 18553 7956
rect 18589 9323 19379 9343
rect 18589 7956 18614 9323
rect 19354 7956 19379 9323
rect 18589 7937 19379 7956
rect 19415 7872 19439 9408
rect 19812 8543 20444 8573
rect 19812 8508 19845 8543
rect 19812 8129 19846 8508
rect 19907 8486 20346 8508
rect 19907 8189 19944 8486
rect 20312 8189 20346 8486
rect 19907 8170 20346 8189
rect 20407 8129 20444 8543
rect 19812 8107 20444 8129
rect 18528 7851 19439 7872
rect 18529 7850 18614 7851
rect 19354 7850 19439 7851
rect 19826 7301 20458 7331
rect 19826 7266 19859 7301
rect 19826 6887 19860 7266
rect 19921 7244 20360 7266
rect 19921 6947 19958 7244
rect 20326 6947 20360 7244
rect 19921 6928 20360 6947
rect 20421 6887 20458 7301
rect 19826 6865 20458 6887
rect 12377 5920 12889 5945
rect 12377 5481 12398 5920
rect 12447 5836 12821 5860
rect 12447 5565 12465 5836
rect 12801 5565 12821 5836
rect 12447 5541 12821 5565
rect 12870 5481 12889 5920
rect 12377 5456 12889 5481
<< nsubdiff >>
rect 15679 15056 20254 15086
rect 15679 12841 15716 15056
rect 15821 14954 20120 14973
rect 20218 14962 20254 15056
rect 15821 14397 15855 14954
rect 15820 14394 15855 14397
rect 17454 14619 17629 14661
rect 15820 12990 15854 14394
rect 17454 14272 17492 14619
rect 17453 13154 17492 14272
rect 17593 14226 17629 14619
rect 17592 13154 17629 14226
rect 17453 13126 17629 13154
rect 19230 14604 19407 14657
rect 19230 13161 19273 14604
rect 19369 14209 19407 14604
rect 19369 13161 19405 14209
rect 19230 13128 19405 13161
rect 20078 12990 20120 14954
rect 20219 14402 20254 14962
rect 15820 12954 20120 12990
rect 20218 12841 20254 14402
rect 15679 12805 20254 12841
rect 5602 10622 10177 10652
rect 5602 10528 5638 10622
rect 5602 9968 5637 10528
rect 5736 10520 10035 10539
rect 5602 8407 5638 9968
rect 5736 8556 5778 10520
rect 6449 10170 6626 10223
rect 6449 9775 6487 10170
rect 6451 8727 6487 9775
rect 6583 8727 6626 10170
rect 6451 8694 6626 8727
rect 8227 10185 8402 10227
rect 8227 9792 8263 10185
rect 8364 9838 8402 10185
rect 10001 9963 10035 10520
rect 10001 9960 10036 9963
rect 8227 8720 8264 9792
rect 8364 8720 8403 9838
rect 8227 8692 8403 8720
rect 10002 8556 10036 9960
rect 5736 8520 10036 8556
rect 10140 8407 10177 10622
rect 10738 10558 10843 10560
rect 10736 10543 11261 10558
rect 10736 10542 10764 10543
rect 10823 10542 11261 10543
rect 10736 10490 10760 10542
rect 10736 10470 10764 10490
rect 10738 8570 10764 10470
rect 10823 10470 11174 10490
rect 10823 8625 10843 10470
rect 11151 8625 11174 10470
rect 10823 8604 11174 8625
rect 11234 10437 11261 10542
rect 11234 8625 11260 10437
rect 17411 9407 18264 9426
rect 16441 9359 16977 9380
rect 16441 8770 16468 9359
rect 16546 9303 16868 9322
rect 16546 8825 16574 9303
rect 16839 8825 16868 9303
rect 16546 8807 16868 8825
rect 16946 8770 16977 9359
rect 16441 8747 16977 8770
rect 17411 9373 17438 9407
rect 11234 8604 11261 8625
rect 11235 8570 11261 8604
rect 10738 8549 11261 8570
rect 10739 8544 11261 8549
rect 5602 8371 10177 8407
rect 16435 7963 16971 7984
rect 10745 7565 10850 7567
rect 10743 7550 11268 7565
rect 10743 7549 10771 7550
rect 10830 7549 11268 7550
rect 10743 7497 10767 7549
rect 10743 7477 10771 7497
rect 10745 5577 10771 7477
rect 10830 7477 11181 7497
rect 10830 5632 10850 7477
rect 11158 5632 11181 7477
rect 10830 5611 11181 5632
rect 11241 7444 11268 7549
rect 11241 5632 11267 7444
rect 16435 7374 16462 7963
rect 16540 7907 16862 7926
rect 16540 7429 16568 7907
rect 16833 7429 16862 7907
rect 16540 7411 16862 7429
rect 16940 7374 16971 7963
rect 17411 7879 17439 9373
rect 17481 9359 18203 9373
rect 17481 7955 17509 9359
rect 17566 8939 18083 8959
rect 17566 8904 17591 8939
rect 18055 8904 18083 8939
rect 17566 8883 18083 8904
rect 18179 7955 18203 9359
rect 17481 7926 18203 7955
rect 18238 7879 18264 9407
rect 17411 7850 18264 7879
rect 19908 9354 20444 9375
rect 19908 8765 19935 9354
rect 20013 9298 20335 9317
rect 20013 8820 20041 9298
rect 20306 8820 20335 9298
rect 20013 8802 20335 8820
rect 20413 8765 20444 9354
rect 19908 8742 20444 8765
rect 19904 8023 20440 8044
rect 19904 7434 19931 8023
rect 20009 7967 20331 7986
rect 20009 7489 20037 7967
rect 20302 7489 20331 7967
rect 20009 7471 20331 7489
rect 20409 7434 20440 8023
rect 19904 7411 20440 7434
rect 16435 7351 16971 7374
rect 19922 6781 20458 6802
rect 19922 6192 19949 6781
rect 20027 6725 20349 6744
rect 20027 6247 20055 6725
rect 20320 6247 20349 6725
rect 20027 6229 20349 6247
rect 20427 6192 20458 6781
rect 19922 6169 20458 6192
rect 12995 5952 13116 5953
rect 14928 5952 15009 5953
rect 11241 5611 11268 5632
rect 11242 5577 11268 5611
rect 10745 5556 11268 5577
rect 10746 5551 11268 5556
rect 12995 5927 15009 5952
rect 12995 5926 14949 5927
rect 12995 5535 13011 5926
rect 12993 5515 13011 5535
rect 13063 5843 14949 5866
rect 13063 5535 13083 5843
rect 14928 5535 14949 5843
rect 13063 5515 14949 5535
rect 12993 5456 13010 5515
rect 14983 5456 15009 5927
rect 12993 5452 13011 5456
rect 13063 5452 15009 5456
rect 12993 5431 15009 5452
rect 12993 5430 15004 5431
rect 12995 5428 13083 5430
rect 5440 2572 5536 2606
rect 41834 2572 41896 2606
rect 5440 2510 5474 2572
rect 5440 458 5474 520
rect 5440 424 5536 458
rect 41834 424 41896 458
<< psubdiffcont >>
rect 12164 14792 14218 14794
rect 12152 12961 14218 14792
rect 12151 12375 14218 12961
rect 12164 12374 14218 12375
rect 10776 11110 11215 11159
rect 10776 10736 10836 11110
rect 11155 10736 11215 11110
rect 10776 10687 11215 10736
rect 15716 11840 20230 11953
rect 15716 10934 15828 11840
rect 20114 10934 20230 11840
rect 15716 10808 20230 10934
rect 16381 9843 16943 9878
rect 16382 9505 16443 9843
rect 16882 9505 16943 9843
rect 16382 9464 16943 9505
rect 19848 9839 20410 9874
rect 19849 9501 19910 9839
rect 20349 9501 20410 9839
rect 19849 9460 20410 9501
rect 16377 8448 16939 8483
rect 10778 8113 11217 8162
rect 10778 7739 10838 8113
rect 11157 7739 11217 8113
rect 10778 7690 11217 7739
rect 16378 8110 16439 8448
rect 16878 8110 16939 8448
rect 16378 8069 16939 8110
rect 5629 7406 10143 7519
rect 5629 6500 5745 7406
rect 10031 6500 10143 7406
rect 5629 6374 10143 6500
rect 18553 9407 18589 9408
rect 19379 9407 19415 9408
rect 18553 9343 19415 9407
rect 18553 7937 18589 9343
rect 19379 7937 19415 9343
rect 18553 7872 19415 7937
rect 19845 8508 20407 8543
rect 19846 8170 19907 8508
rect 20346 8170 20407 8508
rect 19846 8129 20407 8170
rect 19859 7266 20421 7301
rect 19860 6928 19921 7266
rect 20360 6928 20421 7266
rect 19860 6887 20421 6928
rect 12398 5860 12870 5920
rect 12398 5541 12447 5860
rect 12821 5541 12870 5860
rect 12398 5481 12870 5541
<< nsubdiffcont >>
rect 15716 14973 20218 15056
rect 15716 14397 15821 14973
rect 20120 14962 20218 14973
rect 15716 12954 15820 14397
rect 17492 14226 17593 14619
rect 17492 13154 17592 14226
rect 19273 13161 19369 14604
rect 20120 14402 20219 14962
rect 20120 12954 20218 14402
rect 15716 12841 20218 12954
rect 5638 10539 10140 10622
rect 5638 10528 5736 10539
rect 5637 9968 5736 10528
rect 5638 8520 5736 9968
rect 6487 8727 6583 10170
rect 8263 9792 8364 10185
rect 10035 9963 10140 10539
rect 8264 8720 8364 9792
rect 10036 8520 10140 9963
rect 5638 8407 10140 8520
rect 10764 10542 10823 10543
rect 10760 10490 11234 10542
rect 10764 8604 10823 10490
rect 11174 8604 11234 10490
rect 16468 9322 16946 9359
rect 16468 8807 16546 9322
rect 16868 8807 16946 9322
rect 16468 8770 16946 8807
rect 17438 9373 18238 9407
rect 10764 8570 11235 8604
rect 10771 7549 10830 7550
rect 10767 7497 11241 7549
rect 10771 5611 10830 7497
rect 11181 5611 11241 7497
rect 16462 7926 16940 7963
rect 16462 7411 16540 7926
rect 16862 7411 16940 7926
rect 16462 7374 16940 7411
rect 17439 7926 17481 9373
rect 17591 8904 18055 8939
rect 18203 7926 18238 9373
rect 17439 7879 18238 7926
rect 19935 9317 20413 9354
rect 19935 8802 20013 9317
rect 20335 8802 20413 9317
rect 19935 8765 20413 8802
rect 19931 7986 20409 8023
rect 19931 7471 20009 7986
rect 20331 7471 20409 7986
rect 19931 7434 20409 7471
rect 19949 6744 20427 6781
rect 19949 6229 20027 6744
rect 20349 6229 20427 6744
rect 19949 6192 20427 6229
rect 10771 5577 11242 5611
rect 14949 5926 14983 5927
rect 13011 5866 14983 5926
rect 13011 5515 13063 5866
rect 14949 5515 14983 5866
rect 13010 5456 14983 5515
rect 13011 5452 13063 5456
rect 5536 2572 41834 2606
rect 5440 520 5474 2510
rect 5536 424 41834 458
<< locali >>
rect 15694 15056 20241 15073
rect 11930 14794 14414 14936
rect 11930 14792 12164 14794
rect 11930 12961 12152 14792
rect 11930 12375 12151 12961
rect 11930 12374 12164 12375
rect 14218 12374 14414 14794
rect 15694 12841 15716 15056
rect 15821 14964 20120 14973
rect 15821 14397 15841 14964
rect 15820 12973 15841 14397
rect 17468 14619 17615 14641
rect 17468 13154 17492 14619
rect 17593 14226 17615 14619
rect 17592 13154 17615 14226
rect 17468 13136 17615 13154
rect 19247 14604 19391 14635
rect 19247 13161 19273 14604
rect 19369 13161 19391 14604
rect 19247 13139 19391 13161
rect 20095 12973 20120 14964
rect 20218 14962 20241 15056
rect 20219 14959 20241 14962
rect 20219 14402 20242 14959
rect 15820 12954 20120 12973
rect 20218 12841 20241 14402
rect 15694 12840 15850 12841
rect 15972 12840 20241 12841
rect 15694 12821 20241 12840
rect 11930 12218 14414 12374
rect 15700 11953 20246 11971
rect 10755 11159 11235 11172
rect 10755 10687 10776 11159
rect 10836 11096 11155 11110
rect 10836 10750 10856 11096
rect 11134 10750 11155 11096
rect 10836 10736 11155 10750
rect 11215 10954 11235 11159
rect 11215 10874 11236 10954
rect 11215 10687 11235 10874
rect 15700 10808 15716 11953
rect 15828 11822 20114 11840
rect 15828 10950 15838 11822
rect 20106 10950 20114 11822
rect 15828 10934 20114 10950
rect 20230 10808 20246 11953
rect 15700 10791 20246 10808
rect 10755 10671 11235 10687
rect 5615 10622 10162 10639
rect 5615 10528 5638 10622
rect 5736 10530 10035 10539
rect 5615 10525 5637 10528
rect 5614 9968 5637 10525
rect 5615 8407 5638 9968
rect 5736 8539 5761 10530
rect 6465 10170 6609 10201
rect 6465 8727 6487 10170
rect 6583 8727 6609 10170
rect 6465 8705 6609 8727
rect 8241 10185 8388 10207
rect 8241 9792 8263 10185
rect 8241 8720 8264 9792
rect 8364 8720 8388 10185
rect 8241 8702 8388 8720
rect 10015 9963 10035 10530
rect 10015 8539 10036 9963
rect 5736 8520 10036 8539
rect 10140 8407 10162 10622
rect 10741 10543 11253 10553
rect 10741 10542 10764 10543
rect 10823 10542 11253 10543
rect 10741 10490 10760 10542
rect 10741 10476 10764 10490
rect 10747 8570 10764 10476
rect 10823 10476 11174 10490
rect 10823 8616 10833 10476
rect 11158 8616 11174 10476
rect 10823 8604 11174 8616
rect 11234 8604 11253 10542
rect 16361 9878 16965 9896
rect 16361 9843 16381 9878
rect 16361 9464 16382 9843
rect 16443 9830 16882 9843
rect 16443 9516 16465 9830
rect 16859 9516 16882 9830
rect 16443 9505 16882 9516
rect 16943 9464 16965 9878
rect 16361 9449 16965 9464
rect 19828 9874 20432 9892
rect 19828 9839 19848 9874
rect 19828 9460 19849 9839
rect 19910 9826 20349 9839
rect 19910 9512 19932 9826
rect 20326 9512 20349 9826
rect 19910 9501 20349 9512
rect 20410 9460 20432 9874
rect 19828 9445 20432 9460
rect 17420 9407 18253 9423
rect 17420 9373 17438 9407
rect 16452 9359 16966 9371
rect 16452 8770 16468 9359
rect 16546 9312 16868 9322
rect 16546 8818 16563 9312
rect 16846 8818 16868 9312
rect 16546 8807 16868 8818
rect 16946 8770 16966 9359
rect 16452 8755 16966 8770
rect 11235 8570 11253 8604
rect 10747 8553 11253 8570
rect 5615 8387 10162 8407
rect 16357 8484 16961 8501
rect 16357 8483 16886 8484
rect 16926 8483 16961 8484
rect 16357 8448 16377 8483
rect 10757 8162 11237 8175
rect 10757 7690 10778 8162
rect 10838 8099 11157 8113
rect 10838 7753 10858 8099
rect 11136 7753 11157 8099
rect 10838 7739 11157 7753
rect 11217 7957 11237 8162
rect 16357 8069 16378 8448
rect 16439 8435 16878 8448
rect 16439 8121 16461 8435
rect 16855 8121 16878 8435
rect 16439 8110 16878 8121
rect 16939 8069 16961 8483
rect 16357 8054 16961 8069
rect 16446 7963 16960 7975
rect 11217 7877 11238 7957
rect 11217 7690 11237 7877
rect 10757 7674 11237 7690
rect 10748 7550 11260 7560
rect 10748 7549 10771 7550
rect 10830 7549 11260 7550
rect 5613 7519 10159 7537
rect 5613 6374 5629 7519
rect 5745 7388 10031 7406
rect 5745 6516 5753 7388
rect 10021 6516 10031 7388
rect 5745 6500 10031 6516
rect 10143 6374 10159 7519
rect 10748 7497 10767 7549
rect 10748 7483 10771 7497
rect 5613 6357 10159 6374
rect 10754 5577 10771 7483
rect 10830 7483 11181 7497
rect 10830 5623 10840 7483
rect 11165 5623 11181 7483
rect 10830 5611 11181 5623
rect 11241 5611 11260 7549
rect 16446 7374 16462 7963
rect 16540 7916 16862 7926
rect 16540 7422 16557 7916
rect 16840 7422 16862 7916
rect 16540 7411 16862 7422
rect 16940 7374 16960 7963
rect 17420 7879 17439 9373
rect 17481 9366 18203 9373
rect 17481 7944 17498 9366
rect 17570 8939 18075 8954
rect 17570 8904 17591 8939
rect 18055 8904 18075 8939
rect 17570 8888 18075 8904
rect 18189 7944 18203 9366
rect 17481 7926 18203 7944
rect 18238 7879 18253 9407
rect 18539 9408 19429 9424
rect 18539 7951 18553 9408
rect 18589 9407 19379 9408
rect 17420 7858 18253 7879
rect 18537 7872 18553 7951
rect 18589 9330 19379 9343
rect 18589 7951 18603 9330
rect 19365 7951 19379 9330
rect 18589 7937 19379 7951
rect 19415 7950 19429 9408
rect 19919 9354 20433 9366
rect 19919 8765 19935 9354
rect 20013 9307 20335 9317
rect 20013 9050 20030 9307
rect 20014 8948 20030 9050
rect 20013 8813 20030 8948
rect 20313 8813 20335 9307
rect 20013 8802 20335 8813
rect 20413 8765 20433 9354
rect 19919 8750 20433 8765
rect 19825 8543 20429 8561
rect 19825 8508 19845 8543
rect 19825 8129 19846 8508
rect 19907 8495 20346 8508
rect 19907 8181 19929 8495
rect 20323 8181 20346 8495
rect 19907 8170 20346 8181
rect 20407 8129 20429 8543
rect 19825 8114 20429 8129
rect 19915 8023 20429 8035
rect 19415 7872 19435 7950
rect 18537 7858 19435 7872
rect 18537 7857 19429 7858
rect 19915 7434 19931 8023
rect 20009 7976 20331 7986
rect 20009 7482 20026 7976
rect 20309 7482 20331 7976
rect 20009 7471 20331 7482
rect 20409 7434 20429 8023
rect 19915 7419 20429 7434
rect 16446 7359 16960 7374
rect 19839 7301 20443 7319
rect 19839 7266 19859 7301
rect 19839 6887 19860 7266
rect 19921 7253 20360 7266
rect 19921 6939 19943 7253
rect 20337 6939 20360 7253
rect 19921 6928 20360 6939
rect 20421 6887 20443 7301
rect 19839 6872 20443 6887
rect 19933 6781 20447 6793
rect 19933 6288 19949 6781
rect 20027 6734 20349 6744
rect 19933 6194 19948 6288
rect 20027 6240 20044 6734
rect 20327 6240 20349 6734
rect 20027 6229 20349 6240
rect 19933 6192 19949 6194
rect 20427 6192 20447 6781
rect 19933 6177 20447 6192
rect 12603 5940 12683 5941
rect 11242 5577 11260 5611
rect 10754 5560 11260 5577
rect 12385 5920 12886 5940
rect 12385 5481 12398 5920
rect 12447 5839 12821 5860
rect 12447 5561 12461 5839
rect 12807 5561 12821 5839
rect 12447 5541 12821 5561
rect 12870 5481 12886 5920
rect 12385 5460 12886 5481
rect 13000 5927 15000 5945
rect 13000 5926 14949 5927
rect 13000 5548 13011 5926
rect 13063 5850 14949 5866
rect 13000 5460 13008 5548
rect 13063 5525 13077 5850
rect 14937 5525 14949 5850
rect 13063 5515 14949 5525
rect 13000 5456 13010 5460
rect 14983 5456 15000 5927
rect 13000 5452 13011 5456
rect 13063 5452 15000 5456
rect 13000 5439 15000 5452
rect 13000 5433 13077 5439
rect 5440 2572 5536 2606
rect 41834 2572 41896 2606
rect 5440 2510 5474 2572
rect 5440 458 5474 520
rect 5440 424 5536 458
rect 41834 424 41896 458
<< viali >>
rect 12376 12482 14054 12774
rect 15850 12841 15972 12928
rect 15850 12840 15972 12841
rect 10786 10752 10826 11094
rect 15740 10830 16170 10916
rect 5644 8422 5718 8556
rect 11176 8604 11228 8692
rect 16892 9602 16932 9712
rect 20362 9600 20406 9670
rect 16480 9238 16532 9344
rect 16886 8483 16926 8484
rect 10782 7846 10832 7974
rect 16886 8358 16926 8483
rect 9712 6398 10120 6482
rect 11188 5604 11240 5692
rect 16470 7822 16522 7928
rect 17442 7884 17768 7920
rect 19272 9362 19402 9396
rect 19938 8948 20013 9050
rect 20013 8948 20014 9050
rect 20358 8248 20402 8318
rect 19932 7876 20008 7978
rect 20364 7022 20416 7114
rect 19948 6194 19949 6288
rect 19949 6194 20004 6288
rect 12426 5490 12650 5532
rect 13008 5515 13011 5548
rect 13011 5515 13060 5548
rect 13008 5460 13010 5515
rect 13010 5460 13060 5515
rect 11401 458 12487 463
rect 15028 458 16114 461
rect 18681 458 19767 460
rect 22324 458 23410 470
rect 25949 458 27035 465
rect 29580 458 30666 460
rect 33227 458 34313 465
rect 36856 458 37942 467
rect 40551 458 41637 461
rect 7750 424 8836 458
rect 11401 424 12487 458
rect 15028 424 16114 458
rect 18681 424 19767 458
rect 22324 427 23410 458
rect 25949 424 27035 458
rect 29580 424 30666 458
rect 33227 424 34313 458
rect 36856 424 37942 458
rect 40551 424 41637 458
rect 7750 415 8836 424
rect 11401 420 12487 424
rect 15028 418 16114 424
rect 18681 417 19767 424
rect 25949 422 27035 424
rect 29580 417 30666 424
rect 33227 422 34313 424
rect 40551 418 41637 424
<< metal1 >>
rect 15842 12950 15994 12960
rect 10425 12902 12152 12906
rect 10425 12774 14210 12902
rect 15842 12840 15850 12950
rect 15982 12840 15994 12950
rect 15842 12826 15994 12840
rect 10425 12482 12376 12774
rect 14054 12482 14210 12774
rect 10425 12380 14210 12482
rect 10425 11478 10595 12380
rect 12156 12370 14210 12380
rect 19709 12278 19810 12363
rect 15398 11478 15573 11482
rect 10425 11255 15576 11478
rect 10425 10964 10595 11255
rect 10774 11094 10838 11110
rect 10774 10964 10786 11094
rect 10425 10810 10786 10964
rect 4417 8586 5486 8587
rect 4417 8556 5746 8586
rect 4417 8422 5644 8556
rect 5718 8422 5746 8556
rect 4417 8398 5746 8422
rect 4417 5140 5153 8398
rect 10425 7987 10595 10810
rect 10774 10752 10786 10810
rect 10826 10752 10838 11094
rect 10983 11024 11086 11034
rect 10983 10972 10994 11024
rect 11076 10972 11086 11024
rect 10983 10967 11086 10972
rect 15398 10937 15573 11255
rect 15398 10916 16519 10937
rect 15398 10830 15740 10916
rect 16170 10830 16519 10916
rect 15398 10817 16519 10830
rect 15398 10815 15573 10817
rect 10774 10736 10838 10752
rect 16333 10111 16519 10817
rect 16333 10109 17650 10111
rect 16333 10107 18381 10109
rect 16333 10103 19462 10107
rect 16333 9985 20702 10103
rect 16339 9983 20702 9985
rect 17070 9981 20702 9983
rect 16671 9803 16761 9813
rect 16671 9739 16680 9803
rect 16750 9739 16761 9803
rect 16671 9732 16761 9739
rect 16882 9712 16944 9724
rect 16882 9647 16892 9712
rect 16880 9602 16892 9647
rect 16932 9647 16944 9712
rect 17078 9647 17179 9981
rect 18151 9979 20702 9981
rect 19255 9976 20702 9979
rect 16932 9602 17179 9647
rect 16880 9591 17179 9602
rect 17078 9572 17179 9591
rect 16442 9348 16554 9360
rect 16442 9226 16466 9348
rect 16546 9226 16554 9348
rect 16442 9216 16554 9226
rect 16648 8905 16758 8914
rect 16648 8852 16665 8905
rect 16740 8852 16758 8905
rect 16648 8842 16758 8852
rect 10966 8752 11073 8760
rect 10966 8695 10971 8752
rect 11047 8695 11073 8752
rect 10966 8688 11073 8695
rect 11160 8692 11634 8710
rect 11160 8604 11176 8692
rect 11228 8604 11634 8692
rect 11160 8584 11634 8604
rect 10967 8026 11073 8033
rect 10425 7974 10842 7987
rect 6050 7863 6163 7937
rect 10425 7846 10782 7974
rect 10832 7846 10842 7974
rect 10967 7972 10973 8026
rect 11065 7972 11073 8026
rect 10967 7967 11073 7972
rect 10425 7833 10842 7846
rect 10425 6861 10595 7833
rect 10425 6860 10592 6861
rect 10422 6678 10592 6860
rect 10422 6677 10587 6678
rect 10420 6503 10587 6677
rect 9679 6482 10587 6503
rect 9679 6398 9712 6482
rect 10120 6398 10587 6482
rect 9679 6374 10587 6398
rect 10420 5346 10587 6374
rect 10943 5759 11058 5768
rect 10943 5706 10959 5759
rect 11043 5706 11058 5759
rect 11508 5717 11634 8584
rect 17081 8491 17177 9572
rect 19256 9410 19387 9976
rect 20589 9974 20702 9976
rect 20589 9904 20703 9974
rect 20139 9805 20221 9813
rect 20139 9740 20150 9805
rect 20210 9740 20221 9805
rect 20139 9732 20221 9740
rect 20589 9683 20704 9904
rect 20343 9670 20704 9683
rect 20343 9600 20362 9670
rect 20406 9600 20704 9670
rect 20343 9587 20704 9600
rect 17438 9372 18239 9408
rect 17438 9130 17482 9372
rect 17595 9304 17731 9313
rect 17595 9240 17605 9304
rect 17720 9240 17731 9304
rect 17595 9232 17731 9240
rect 17759 9299 17837 9301
rect 17759 9246 17766 9299
rect 17829 9246 17837 9299
rect 17759 9240 17837 9246
rect 17759 9212 17821 9240
rect 17759 9068 17820 9212
rect 18202 8948 18239 9372
rect 19256 9396 19414 9410
rect 19256 9362 19272 9396
rect 19402 9362 19414 9396
rect 19256 9345 19414 9362
rect 18942 9296 19099 9312
rect 18942 9224 18954 9296
rect 19082 9224 19099 9296
rect 18942 9212 19099 9224
rect 17591 8905 18239 8948
rect 19377 8943 19414 9345
rect 19590 9050 20033 9064
rect 19590 8948 19938 9050
rect 20014 8948 20033 9050
rect 17591 8904 18061 8905
rect 16874 8484 17177 8491
rect 16641 8417 16737 8425
rect 16641 8348 16651 8417
rect 16729 8348 16737 8417
rect 16641 8340 16737 8348
rect 16874 8358 16886 8484
rect 16926 8428 17177 8484
rect 16926 8358 16940 8428
rect 17081 8427 17177 8428
rect 17538 8718 17686 8720
rect 17538 8702 17689 8718
rect 17538 8384 17560 8702
rect 17673 8384 17689 8702
rect 17538 8365 17689 8384
rect 17538 8359 17686 8365
rect 16874 8344 16940 8358
rect 16446 7954 16548 7964
rect 16446 7810 16460 7954
rect 16534 7810 16548 7954
rect 16446 7798 16548 7810
rect 17399 7929 17623 7942
rect 18202 7929 18238 8905
rect 18995 8903 19416 8943
rect 19590 8921 20033 8948
rect 19590 8847 19782 8921
rect 20133 8907 20217 8914
rect 19591 8001 19781 8847
rect 20133 8846 20146 8907
rect 20209 8846 20217 8907
rect 20133 8839 20217 8846
rect 20137 8456 20214 8466
rect 20137 8400 20143 8456
rect 20207 8400 20214 8456
rect 20137 8395 20214 8400
rect 20589 8334 20704 9587
rect 20339 8318 20704 8334
rect 20339 8248 20358 8318
rect 20402 8248 20704 8318
rect 20339 8238 20704 8248
rect 19591 7978 20033 8001
rect 17399 7920 18241 7929
rect 17399 7884 17442 7920
rect 17768 7884 18241 7920
rect 17399 7879 18241 7884
rect 17399 7870 18240 7879
rect 19591 7876 19932 7978
rect 20008 7876 20033 7978
rect 16636 7510 16766 7520
rect 16636 7443 16645 7510
rect 16753 7443 16766 7510
rect 16636 7435 16766 7443
rect 12514 5769 12591 5770
rect 12507 5762 12591 5769
rect 10943 5697 11058 5706
rect 11174 5692 11636 5717
rect 12507 5703 12528 5762
rect 12582 5703 12591 5762
rect 12507 5697 12591 5703
rect 14797 5722 14882 5738
rect 11174 5604 11188 5692
rect 11240 5604 11636 5692
rect 14797 5670 14803 5722
rect 14856 5670 14882 5722
rect 14797 5656 14882 5670
rect 11174 5591 11636 5604
rect 10420 5262 10450 5346
rect 10559 5262 10587 5346
rect 10420 5246 10587 5262
rect 11508 5140 11634 5591
rect 12985 5548 13088 5566
rect 12416 5544 12512 5546
rect 12414 5534 12666 5544
rect 12414 5480 12426 5534
rect 12499 5532 12666 5534
rect 12650 5490 12666 5532
rect 12416 5479 12426 5480
rect 12499 5480 12666 5490
rect 12499 5479 12512 5480
rect 12985 5460 13008 5548
rect 13060 5460 13088 5548
rect 4412 5138 11676 5140
rect 12985 5139 13088 5460
rect 17399 5163 17623 7870
rect 19591 7858 20033 7876
rect 19591 6304 19781 7858
rect 20132 7569 20222 7577
rect 20132 7497 20140 7569
rect 20212 7497 20222 7569
rect 20132 7487 20222 7497
rect 20152 7216 20231 7223
rect 20152 7159 20159 7216
rect 20223 7159 20231 7216
rect 20152 7152 20231 7159
rect 20354 7120 20426 7122
rect 20589 7120 20704 8238
rect 20351 7114 20704 7120
rect 20351 7041 20364 7114
rect 20354 7022 20364 7041
rect 20416 7042 20704 7114
rect 20416 7041 20692 7042
rect 20416 7022 20426 7041
rect 20354 7010 20426 7022
rect 20146 6323 20231 6331
rect 19591 6288 20025 6304
rect 19591 6194 19948 6288
rect 20004 6194 20025 6288
rect 20146 6256 20155 6323
rect 20224 6256 20231 6323
rect 20146 6248 20231 6256
rect 19591 6161 20025 6194
rect 19591 5163 19781 6161
rect 27240 5395 27403 5404
rect 22419 5337 22547 5350
rect 22419 5246 22433 5337
rect 22531 5246 22547 5337
rect 23408 5328 23517 5337
rect 22846 5266 23087 5311
rect 22419 5233 22547 5246
rect 23408 5246 23417 5328
rect 23510 5246 23517 5328
rect 23408 5235 23517 5246
rect 27240 5241 27251 5395
rect 27390 5241 27403 5395
rect 15841 5142 15999 5147
rect 17399 5142 19781 5163
rect 15841 5140 19781 5142
rect 14520 5139 19781 5140
rect 12985 5138 19781 5139
rect 4412 5130 19781 5138
rect 4412 5018 15860 5130
rect 15980 5018 19781 5130
rect 27240 5093 27403 5241
rect 4412 5013 19781 5018
rect 4412 5008 19743 5013
rect 4417 -474 5153 5008
rect 11508 5006 19743 5008
rect 11508 5004 17457 5006
rect 11508 5002 15999 5004
rect 11508 5001 14552 5002
rect 11594 5000 13088 5001
rect 15841 4998 15999 5002
rect 27239 569 27403 5093
rect 4417 -528 5171 -474
rect 4417 -1121 4485 -528
rect 5107 -1121 5171 -528
rect 4417 -1169 5171 -1121
<< via1 >>
rect 15850 12928 15982 12950
rect 15850 12840 15972 12928
rect 15972 12840 15982 12928
rect 10994 10972 11076 11024
rect 16680 9739 16750 9803
rect 16466 9344 16546 9348
rect 16466 9238 16480 9344
rect 16480 9238 16532 9344
rect 16532 9238 16546 9344
rect 16466 9226 16546 9238
rect 16665 8852 16740 8905
rect 10971 8695 11047 8752
rect 10973 7972 11065 8026
rect 10959 5706 11043 5759
rect 20150 9740 20210 9805
rect 17605 9240 17720 9304
rect 17766 9246 17829 9299
rect 18954 9224 19082 9296
rect 16651 8348 16729 8417
rect 17560 8384 17673 8702
rect 16460 7928 16534 7954
rect 16460 7822 16470 7928
rect 16470 7822 16522 7928
rect 16522 7822 16534 7928
rect 16460 7810 16534 7822
rect 20146 8846 20209 8907
rect 20143 8400 20207 8456
rect 16645 7443 16753 7510
rect 12528 5703 12582 5762
rect 14803 5670 14856 5722
rect 10450 5262 10559 5346
rect 12426 5532 12499 5534
rect 12426 5490 12499 5532
rect 12426 5479 12499 5490
rect 20140 7497 20212 7569
rect 20159 7159 20223 7216
rect 20155 6256 20224 6323
rect 22433 5246 22531 5337
rect 23417 5246 23510 5328
rect 27251 5241 27390 5395
rect 15860 5018 15980 5130
rect 4485 -1121 5107 -528
<< metal2 >>
rect 15842 12950 15994 12960
rect 15842 12840 15850 12950
rect 15982 12840 15994 12950
rect 10983 11028 11086 11034
rect 10983 10972 10994 11028
rect 11076 10972 11086 11028
rect 10983 10967 11086 10972
rect 11033 10380 11114 10400
rect 10918 9168 10966 9228
rect 11092 8842 11114 10380
rect 15842 9360 15994 12840
rect 16192 11625 16327 11643
rect 16192 11546 16207 11625
rect 16309 11546 16327 11625
rect 16192 11531 16327 11546
rect 16801 11625 16904 11637
rect 16801 11502 16814 11625
rect 16894 11502 16904 11625
rect 16801 11487 16904 11502
rect 18943 10574 19099 10591
rect 18943 10476 18958 10574
rect 19081 10476 19099 10574
rect 16671 9803 16761 9813
rect 16671 9739 16680 9803
rect 16750 9739 16761 9803
rect 16671 9732 16761 9739
rect 17759 9804 17837 9813
rect 17759 9739 17767 9804
rect 17828 9739 17837 9804
rect 15842 9348 16554 9360
rect 15842 9226 16466 9348
rect 16546 9226 16554 9348
rect 17595 9304 17731 9313
rect 17595 9241 17604 9304
rect 17721 9241 17731 9304
rect 17595 9240 17605 9241
rect 17720 9240 17731 9241
rect 17759 9299 17837 9739
rect 18943 9313 19099 10476
rect 20139 9805 20221 9813
rect 20139 9740 20150 9805
rect 20210 9740 20221 9805
rect 20139 9732 20221 9740
rect 19626 9314 19703 9315
rect 19543 9313 19704 9314
rect 17759 9246 17766 9299
rect 17829 9246 17837 9299
rect 17759 9240 17837 9246
rect 18941 9296 19704 9313
rect 17595 9232 17731 9240
rect 15842 9216 16554 9226
rect 18941 9224 18954 9296
rect 19082 9224 19704 9296
rect 11076 8799 11114 8842
rect 10966 8752 11073 8760
rect 10966 8695 10971 8752
rect 11047 8750 11073 8752
rect 10966 8688 10974 8695
rect 11063 8688 11073 8750
rect 10966 8679 11073 8688
rect 10967 8041 11073 8051
rect 15844 8047 16002 9216
rect 18941 9214 19704 9224
rect 18941 9213 19548 9214
rect 18943 9212 19099 9213
rect 16609 9137 16692 9147
rect 16609 8954 16626 9137
rect 16682 8954 16692 9137
rect 16609 8946 16692 8954
rect 16726 9141 16826 9149
rect 16726 8953 16759 9141
rect 16815 8953 16826 9141
rect 16726 8946 16826 8953
rect 19626 8914 19703 9214
rect 20196 9147 20326 9162
rect 20076 9131 20095 9140
rect 20076 9006 20088 9131
rect 20076 8997 20095 9006
rect 20196 8974 20234 9147
rect 20313 8974 20326 9147
rect 20196 8962 20326 8974
rect 16648 8905 16758 8914
rect 16648 8852 16665 8905
rect 16740 8852 16758 8905
rect 19626 8907 20217 8914
rect 16648 8820 16758 8852
rect 16648 8754 16664 8820
rect 16739 8754 16758 8820
rect 17974 8863 18099 8876
rect 17974 8775 17988 8863
rect 18080 8775 18099 8863
rect 17974 8763 18099 8775
rect 18770 8849 18887 8864
rect 18770 8770 18782 8849
rect 18870 8770 18887 8849
rect 19626 8846 20146 8907
rect 20209 8846 20217 8907
rect 18770 8758 18887 8770
rect 19136 8834 19244 8846
rect 19136 8764 19148 8834
rect 19228 8764 19244 8834
rect 16648 8734 16758 8754
rect 19136 8753 19244 8764
rect 19626 8839 20217 8846
rect 17538 8718 17686 8720
rect 17538 8702 17689 8718
rect 16641 8417 16737 8425
rect 16641 8348 16651 8417
rect 16729 8348 16737 8417
rect 17538 8384 17560 8702
rect 17673 8384 17689 8702
rect 18354 8553 18395 8597
rect 17538 8365 17689 8384
rect 17538 8359 17686 8365
rect 16641 8340 16737 8348
rect 10967 7972 10973 8041
rect 11066 7977 11073 8041
rect 11065 7972 11073 7977
rect 10967 7967 11073 7972
rect 15843 7964 16002 8047
rect 15843 7954 16548 7964
rect 15843 7810 16460 7954
rect 16534 7810 16548 7954
rect 15843 7798 16548 7810
rect 10909 7386 10986 7396
rect 10909 5838 10919 7386
rect 10976 5838 10986 7386
rect 10909 5829 10986 5838
rect 11049 6472 11140 6491
rect 11049 5851 11064 6472
rect 11122 5851 11140 6472
rect 11049 5837 11140 5851
rect 10943 5762 11058 5768
rect 10943 5702 10953 5762
rect 11048 5702 11058 5762
rect 10943 5697 11058 5702
rect 12507 5762 12591 5770
rect 12507 5705 12516 5762
rect 12507 5703 12528 5705
rect 12582 5703 12591 5762
rect 14797 5722 14882 5738
rect 12507 5697 12591 5703
rect 14797 5670 14803 5722
rect 14856 5721 14882 5722
rect 14797 5663 14806 5670
rect 14864 5663 14882 5721
rect 14797 5656 14882 5663
rect 13159 5556 14759 5618
rect 12415 5534 12512 5545
rect 12415 5479 12426 5534
rect 12499 5479 12512 5534
rect 12415 5366 12512 5479
rect 13159 5485 13181 5556
rect 14738 5485 14759 5556
rect 13159 5467 14759 5485
rect 10428 5346 12512 5366
rect 10428 5262 10450 5346
rect 10559 5262 12512 5346
rect 10428 5246 12512 5262
rect 15843 5147 16000 7798
rect 16612 7743 16686 7752
rect 16612 7560 16622 7743
rect 16678 7560 16686 7743
rect 16612 7550 16686 7560
rect 16722 7746 16825 7754
rect 16722 7558 16757 7746
rect 16813 7558 16825 7746
rect 16722 7551 16825 7558
rect 19626 7577 19702 8839
rect 20137 8458 20214 8466
rect 20137 8456 20146 8458
rect 20204 8456 20214 8458
rect 20137 8400 20143 8456
rect 20207 8400 20214 8456
rect 20137 8395 20214 8400
rect 20028 7792 20146 7800
rect 20028 7615 20037 7792
rect 20139 7615 20146 7792
rect 20196 7668 20228 7698
rect 20028 7606 20146 7615
rect 19626 7569 20222 7577
rect 16636 7510 16766 7520
rect 16636 7443 16645 7510
rect 16753 7443 16766 7510
rect 16636 7427 16766 7443
rect 16636 7353 16645 7427
rect 16755 7353 16766 7427
rect 16636 7343 16766 7353
rect 19626 7497 20140 7569
rect 20212 7497 20222 7569
rect 19626 7467 20222 7497
rect 19626 6331 19702 7467
rect 20152 7220 20231 7231
rect 20152 7159 20159 7220
rect 20223 7159 20231 7220
rect 20152 7154 20231 7159
rect 20056 6560 20162 6566
rect 20056 6375 20065 6560
rect 20155 6375 20162 6560
rect 20218 6472 20234 6490
rect 20056 6369 20162 6375
rect 19626 6323 20231 6331
rect 19626 6256 20155 6323
rect 20224 6256 20231 6323
rect 19626 6244 20231 6256
rect 27240 5395 27403 5405
rect 22419 5337 22547 5350
rect 22419 5246 22433 5337
rect 22531 5246 22547 5337
rect 22419 5233 22547 5246
rect 23408 5328 23517 5337
rect 23408 5246 23417 5328
rect 23510 5246 23517 5328
rect 23408 5235 23517 5246
rect 27240 5241 27251 5395
rect 27390 5241 27403 5395
rect 27240 5229 27403 5241
rect 15841 5130 16000 5147
rect 15841 5018 15860 5130
rect 15980 5023 16000 5130
rect 15980 5018 15999 5023
rect 15841 4998 15999 5018
rect 4417 -528 5171 -474
rect 4417 -1121 4485 -528
rect 5107 -1121 5171 -528
rect 4417 -1169 5171 -1121
<< via2 >>
rect 10994 11024 11076 11028
rect 10994 10972 11076 11024
rect 11033 8842 11092 10380
rect 16207 11546 16309 11625
rect 16814 11502 16894 11625
rect 18958 10476 19081 10574
rect 16680 9739 16750 9803
rect 17767 9739 17828 9804
rect 17604 9241 17605 9304
rect 17605 9241 17720 9304
rect 17720 9241 17721 9304
rect 20150 9740 20210 9805
rect 10974 8695 11047 8750
rect 11047 8695 11063 8750
rect 10974 8688 11063 8695
rect 16626 8954 16682 9137
rect 16759 8953 16815 9141
rect 17631 8956 17713 9033
rect 20088 9006 20150 9131
rect 20234 8974 20313 9147
rect 16664 8754 16739 8820
rect 17988 8775 18080 8863
rect 18782 8770 18870 8849
rect 19148 8764 19228 8834
rect 16651 8348 16726 8416
rect 17560 8384 17673 8702
rect 10973 8026 11066 8041
rect 10973 7977 11065 8026
rect 11065 7977 11066 8026
rect 8973 7124 9030 7202
rect 9555 7121 9633 7191
rect 10919 5838 10976 7386
rect 11064 5851 11122 6472
rect 10953 5759 11048 5762
rect 10953 5706 10959 5759
rect 10959 5706 11043 5759
rect 11043 5706 11048 5759
rect 10953 5702 11048 5706
rect 12516 5705 12528 5762
rect 12528 5705 12580 5762
rect 13169 5719 14726 5775
rect 14806 5670 14856 5721
rect 14856 5670 14864 5721
rect 14806 5663 14864 5670
rect 13181 5485 14738 5556
rect 16622 7560 16678 7743
rect 16757 7558 16813 7746
rect 20146 8456 20204 8458
rect 20146 8402 20204 8456
rect 20037 7615 20139 7792
rect 16645 7353 16755 7427
rect 20159 7216 20223 7220
rect 20159 7163 20223 7216
rect 20065 6375 20155 6560
rect 22433 5246 22531 5337
rect 23417 5246 23510 5328
rect 27251 5241 27390 5395
rect 4485 -1121 5107 -528
<< metal3 >>
rect 16192 11625 16327 11643
rect 16192 11546 16207 11625
rect 16309 11546 16327 11625
rect 10738 11028 11086 11034
rect 10738 10972 10994 11028
rect 11076 10972 11086 11028
rect 10738 10957 11086 10972
rect 10738 10862 10843 10957
rect 8944 7209 9069 7215
rect 8944 7124 8973 7209
rect 9044 7124 9069 7209
rect 10737 7208 10843 10862
rect 16192 10662 16327 11546
rect 16801 11625 16904 11637
rect 16801 11502 16814 11625
rect 16894 11502 16904 11625
rect 16801 11487 16904 11502
rect 16191 10553 16327 10662
rect 18943 10574 19098 10594
rect 11028 10380 11099 10388
rect 11028 8841 11033 10380
rect 11092 10379 11099 10380
rect 11098 8841 11099 10379
rect 16191 10345 16326 10553
rect 18943 10476 18958 10574
rect 19081 10476 19098 10574
rect 18943 10460 19098 10476
rect 16190 10145 16326 10345
rect 16190 9813 16325 10145
rect 16190 9805 20529 9813
rect 16190 9804 20150 9805
rect 16190 9803 17767 9804
rect 16190 9739 16680 9803
rect 16750 9739 17767 9803
rect 17828 9740 20150 9804
rect 20210 9740 20529 9805
rect 17828 9739 20529 9740
rect 16190 9732 20529 9739
rect 16190 9051 16325 9732
rect 17594 9410 20326 9498
rect 17594 9304 17731 9410
rect 17594 9241 17604 9304
rect 17721 9241 17731 9304
rect 17594 9232 17731 9241
rect 11028 8835 11099 8841
rect 10967 8750 11073 8769
rect 10967 8688 10974 8750
rect 11063 8688 11073 8750
rect 10967 8387 11073 8688
rect 16189 8579 16325 9051
rect 16609 9138 16692 9147
rect 16609 8957 16616 9138
rect 16685 8957 16692 9138
rect 16609 8954 16626 8957
rect 16682 8954 16692 8957
rect 16609 8946 16692 8954
rect 16752 9141 16850 9150
rect 16752 8953 16759 9141
rect 16815 9048 16850 9141
rect 20224 9149 20326 9410
rect 18596 9131 20158 9140
rect 16815 9033 17725 9048
rect 16815 8956 17631 9033
rect 17713 8956 17725 9033
rect 16815 8953 17725 8956
rect 16752 8946 17725 8953
rect 18596 9006 20088 9131
rect 20150 9006 20158 9131
rect 20224 9027 20233 9149
rect 18596 8997 20158 9006
rect 17974 8863 18099 8876
rect 16648 8820 16758 8842
rect 16648 8754 16664 8820
rect 16739 8754 16758 8820
rect 17974 8775 17988 8863
rect 18080 8775 18099 8863
rect 17974 8763 18099 8775
rect 16648 8734 16758 8754
rect 17538 8718 17686 8720
rect 17538 8702 17689 8718
rect 18596 8714 18703 8997
rect 20225 8972 20233 9027
rect 20314 8972 20326 9149
rect 20225 8962 20326 8972
rect 18770 8849 18887 8864
rect 18770 8770 18782 8849
rect 18870 8770 18887 8849
rect 18770 8758 18887 8770
rect 19136 8834 19277 8846
rect 19136 8764 19148 8834
rect 19228 8764 19277 8834
rect 19136 8753 19277 8764
rect 16189 8425 16324 8579
rect 16189 8416 16737 8425
rect 10967 8377 11349 8387
rect 10967 8268 10972 8377
rect 11065 8268 11349 8377
rect 16189 8348 16651 8416
rect 16726 8348 16737 8416
rect 17538 8384 17560 8702
rect 17673 8384 17689 8702
rect 18594 8397 18703 8714
rect 17538 8365 17689 8384
rect 17538 8359 17686 8365
rect 16189 8339 16737 8348
rect 10967 8261 11349 8268
rect 10967 8041 11073 8261
rect 10967 7977 10973 8041
rect 11066 7977 11073 8041
rect 10967 7957 11073 7977
rect 10909 7389 10986 7396
rect 8944 7114 9069 7124
rect 9547 7191 10842 7208
rect 9547 7121 9555 7191
rect 9633 7121 10842 7191
rect 9547 7108 10842 7121
rect 10736 5769 10842 7108
rect 10909 5835 10914 7389
rect 10981 5835 10986 7389
rect 11049 6473 11140 6491
rect 11049 5851 11064 6473
rect 11128 5851 11140 6473
rect 11248 5980 11349 8261
rect 19165 7757 19277 8753
rect 20137 8462 20214 8466
rect 20460 8462 20529 9732
rect 20137 8458 20529 8462
rect 20137 8402 20146 8458
rect 20204 8402 20529 8458
rect 20137 8392 20529 8402
rect 20460 8168 20529 8392
rect 20459 7930 20529 8168
rect 18528 7756 19277 7757
rect 17963 7755 19277 7756
rect 17401 7754 19277 7755
rect 16599 7743 16686 7753
rect 16599 7741 16622 7743
rect 16678 7741 16686 7743
rect 16599 7560 16610 7741
rect 16679 7560 16686 7741
rect 16599 7550 16686 7560
rect 16748 7746 19277 7754
rect 16748 7558 16757 7746
rect 16813 7558 19277 7746
rect 20028 7792 20146 7800
rect 20028 7615 20037 7792
rect 20139 7615 20146 7792
rect 20028 7606 20146 7615
rect 16748 7554 19277 7558
rect 16748 7553 18556 7554
rect 19081 7553 19244 7554
rect 16748 7552 17994 7553
rect 16748 7551 17417 7552
rect 16636 7427 16766 7435
rect 16636 7353 16645 7427
rect 16755 7353 16766 7427
rect 16636 7343 16766 7353
rect 20459 7227 20528 7930
rect 20152 7220 20528 7227
rect 20152 7163 20159 7220
rect 20223 7163 20528 7220
rect 20152 7152 20528 7163
rect 20056 6560 20162 6566
rect 20056 6375 20065 6560
rect 20155 6375 20162 6560
rect 20056 6369 20162 6375
rect 11248 5867 14882 5980
rect 11049 5837 11140 5851
rect 10909 5829 10986 5835
rect 13158 5789 14735 5799
rect 10736 5762 12599 5769
rect 10736 5702 10953 5762
rect 11048 5705 12516 5762
rect 12580 5705 12599 5762
rect 13158 5719 13169 5789
rect 14727 5776 14735 5789
rect 14727 5719 14736 5776
rect 13158 5710 14736 5719
rect 14797 5721 14882 5867
rect 13158 5709 14735 5710
rect 11048 5702 12599 5705
rect 10736 5697 12599 5702
rect 14797 5663 14806 5721
rect 14864 5663 14882 5721
rect 14797 5656 14882 5663
rect 13159 5556 14759 5578
rect 13159 5485 13181 5556
rect 14738 5485 14759 5556
rect 13159 5467 14759 5485
rect 27240 5395 27403 5405
rect 22419 5337 22547 5350
rect 22419 5246 22433 5337
rect 22531 5246 22547 5337
rect 22419 5233 22547 5246
rect 23402 5335 23525 5343
rect 23402 5237 23412 5335
rect 23515 5237 23525 5335
rect 23402 5230 23525 5237
rect 27240 5241 27251 5395
rect 27390 5241 27403 5395
rect 27240 5229 27403 5241
rect 4417 -476 5171 -474
rect 4417 -528 6104 -476
rect 4417 -1121 4485 -528
rect 5107 -1121 6104 -528
rect 4417 -1169 6104 -1121
rect 5136 -1170 6104 -1169
<< via3 >>
rect 8973 7202 9044 7209
rect 8973 7124 9030 7202
rect 9030 7124 9044 7202
rect 16814 11502 16894 11625
rect 11033 8842 11092 10379
rect 11092 8842 11098 10379
rect 11033 8841 11098 8842
rect 18958 10476 19081 10574
rect 16616 9137 16685 9138
rect 16616 8957 16626 9137
rect 16626 8957 16682 9137
rect 16682 8957 16685 9137
rect 20233 9147 20314 9149
rect 16664 8754 16739 8820
rect 17988 8775 18080 8863
rect 20233 8974 20234 9147
rect 20234 8974 20313 9147
rect 20313 8974 20314 9147
rect 20233 8972 20314 8974
rect 18782 8770 18870 8849
rect 10972 8268 11065 8377
rect 17560 8384 17673 8702
rect 10914 7386 10981 7389
rect 10914 5838 10919 7386
rect 10919 5838 10976 7386
rect 10976 5838 10981 7386
rect 10914 5835 10981 5838
rect 11064 6472 11128 6473
rect 11064 5851 11122 6472
rect 11122 5851 11128 6472
rect 16610 7560 16622 7741
rect 16622 7560 16678 7741
rect 16678 7560 16679 7741
rect 20037 7615 20139 7792
rect 16645 7353 16755 7427
rect 20065 6375 20155 6560
rect 13169 5775 14727 5789
rect 13169 5719 14726 5775
rect 14726 5719 14727 5775
rect 13181 5485 14738 5556
rect 22433 5246 22531 5337
rect 23412 5328 23515 5335
rect 23412 5246 23417 5328
rect 23417 5246 23510 5328
rect 23510 5246 23515 5328
rect 23412 5237 23515 5246
rect 27251 5241 27390 5395
<< metal4 >>
rect 16801 11625 16904 11637
rect 16801 11502 16814 11625
rect 16894 11502 16904 11625
rect 16801 11487 16904 11502
rect 16802 10592 16881 11487
rect 17581 10592 19099 10593
rect 16802 10574 19099 10592
rect 16802 10476 18958 10574
rect 19081 10476 19099 10574
rect 16802 10460 19099 10476
rect 16802 10459 17623 10460
rect 11028 10379 12098 10388
rect 11028 8841 11033 10379
rect 11098 8841 12098 10379
rect 16211 9138 16692 9147
rect 16211 8957 16616 9138
rect 16685 8957 16692 9138
rect 16211 8947 16692 8957
rect 11028 8811 12098 8841
rect 10534 8377 11098 8386
rect 10534 8268 10972 8377
rect 11065 8268 11098 8377
rect 10534 8262 11098 8268
rect 10534 7342 10653 8262
rect 16212 7753 16329 8947
rect 16803 8842 16882 10459
rect 20225 9149 21793 9170
rect 20225 8972 20233 9149
rect 20314 8972 21793 9149
rect 20225 8962 21793 8972
rect 16648 8820 16882 8842
rect 16648 8754 16664 8820
rect 16739 8754 16882 8820
rect 16648 8734 16882 8754
rect 16212 7741 16687 7753
rect 16212 7560 16610 7741
rect 16679 7560 16687 7741
rect 16212 7550 16687 7560
rect 8959 7253 10653 7342
rect 10909 7390 10986 7396
rect 10909 7389 12051 7390
rect 8959 7209 9049 7253
rect 8959 7124 8973 7209
rect 9044 7124 9049 7209
rect 8959 7114 9049 7124
rect 10909 5835 10914 7389
rect 10981 6572 12051 7389
rect 10981 5835 10986 6572
rect 10909 5829 10986 5835
rect 11049 6473 11140 6491
rect 11049 5851 11064 6473
rect 11128 5851 11140 6473
rect 16212 6423 16329 7550
rect 16803 7435 16882 8734
rect 17969 8863 18102 8880
rect 18881 8864 18979 8865
rect 17969 8775 17988 8863
rect 18080 8775 18102 8863
rect 16636 7427 16882 7435
rect 16636 7353 16645 7427
rect 16755 7353 16882 7427
rect 16636 7343 16882 7353
rect 17538 8718 17686 8720
rect 17538 8702 17689 8718
rect 17538 8384 17560 8702
rect 17673 8384 17689 8702
rect 11049 5752 11140 5851
rect 11048 5349 11140 5752
rect 13158 5789 14757 6418
rect 15785 6327 16329 6423
rect 15785 6326 16323 6327
rect 13158 5719 13169 5789
rect 14727 5719 14757 5789
rect 13158 5710 14757 5719
rect 17538 5579 17689 8384
rect 17969 8185 18102 8775
rect 18770 8849 18979 8864
rect 18770 8770 18782 8849
rect 18870 8770 18979 8849
rect 18770 8758 18979 8770
rect 18881 8600 18979 8758
rect 17968 7170 18102 8185
rect 18880 7909 18979 8600
rect 18880 7800 18978 7909
rect 18880 7792 20147 7800
rect 18880 7615 20037 7792
rect 20139 7615 20147 7792
rect 18880 7596 20147 7615
rect 17968 6566 18101 7170
rect 17968 6560 20162 6566
rect 17968 6375 20065 6560
rect 20155 6375 20162 6560
rect 17968 6369 20162 6375
rect 26109 6157 27403 6368
rect 13159 5556 17689 5579
rect 13159 5485 13181 5556
rect 14738 5485 17689 5556
rect 13159 5467 17689 5485
rect 11048 5337 22547 5349
rect 11048 5246 22433 5337
rect 22531 5246 22547 5337
rect 11048 5234 22547 5246
rect 11048 5233 13123 5234
rect 13309 5233 22547 5234
rect 23402 5335 23527 5718
rect 23402 5237 23412 5335
rect 23515 5237 23527 5335
rect 19120 4266 20674 5233
rect 23402 5230 23527 5237
rect 27240 5395 27403 6157
rect 27240 5241 27251 5395
rect 27390 5241 27403 5395
rect 27240 5229 27403 5241
use pseudolayout  CLKgenerator /research/mlab/chipathon/Final_layout
timestamp 1669223049
transform 1 0 5266 0 1 6298
box 356 74 4887 4325
use pseudolayout  ENgenerator
timestamp 1669223049
transform -1 0 20592 0 1 10732
box 356 74 4887 4325
use Liza_Tgate  amplify /research/mlab/chipathon/Final_layout
timestamp 1669223049
transform 0 -1 15126 1 0 5215
box 173 68 787 2594
use Liza_Tgate  autozero
timestamp 1669223049
transform 1 0 10524 0 1 5429
box 173 68 787 2594
use Liza_enable  bottomleft_enable /research/mlab/chipathon/Final_layout
timestamp 1669223049
transform 1 0 16070 0 1 7094
box 434 356 744 1300
use Liza_enable  n_enable
timestamp 1669223049
transform 1 0 19540 0 1 7153
box 434 356 744 1300
use Liza_enable  p_enable
timestamp 1669223049
transform 1 0 19556 0 1 5912
box 434 356 744 1300
use sky130_fd_pr__pfet_01v8_J2H2S6  pass
timestamp 1669223049
transform 0 1 23685 1 0 1515
box -3371 -18281 3401 18341
use rldo  rldo_0
timestamp 1669223049
transform 1 0 12335 0 1 4667
box 5103 3281 6955 4741
use Liza_Tgate  sample
timestamp 1669223049
transform 1 0 10523 0 1 8432
box 173 68 787 2594
use sky130_fd_pr__cap_mim_m3_1_3RKQ3N  sky130_fd_pr__cap_mim_m3_1_3RKQ3N_0
timestamp 1669223049
transform 0 1 23906 -1 0 7783
box -2150 -2600 2149 2600
use sky130_fd_pr__cap_mim_m3_1_BSSJ5K  sky130_fd_pr__cap_mim_m3_1_BSSJ5K_0
timestamp 1669223049
transform 0 1 13844 -1 0 8471
box -2150 -2100 2149 2100
use sky130_fd_pr__res_generic_po_B4RDC6  sky130_fd_pr__res_generic_po_B4RDC6_0
timestamp 1669223049
transform 0 -1 22968 1 0 5288
box -33 -528 33 528
use Liza_enable  topleft_enable
timestamp 1669223049
transform 1 0 16074 0 1 8490
box 434 356 744 1300
use Liza_enable  topright_enable
timestamp 1669223049
transform 1 0 19544 0 1 8486
box 434 356 744 1300
<< labels >>
rlabel metal3 9688 7158 9688 7158 7 CLK
rlabel metal4 9688 7306 9690 7306 7 CLKinverted
rlabel metal3 16261 10599 16262 10600 7 EN
rlabel metal4 16826 11045 16826 11045 7 ENinverted
rlabel metal4 22086 5298 22086 5298 7 Vout
port 5 w
rlabel metal2 10940 9192 10940 9192 7 Vref
port 2 w
rlabel metal2 20212 7682 20212 7682 7 NMOS_DZ
port 6 w
rlabel metal2 20224 6482 20224 6482 7 PMOS_DZ
port 7 w
rlabel metal4 11552 9160 11552 9174 7 net5
rlabel metal4 16168 6370 16168 6370 7 net6
rlabel metal3 17190 8974 17190 8974 7 net7
rlabel metal3 17238 7620 17238 7620 7 net8
rlabel metal4 15660 5518 15660 5518 7 net1
rlabel metal3 18662 8786 18662 8786 7 net2
rlabel metal4 20644 9030 20644 9030 7 net4
rlabel metal2 18373 8572 18373 8572 7 net3
rlabel metal1 4811 0 4811 0 7 Vin
port 1 w
rlabel nsubdiffcont 11204 7519 11204 7519 7 Vin
rlabel nsubdiffcont 13041 5889 13041 5889 5 Vin
rlabel nsubdiffcont 11197 10512 11197 10512 7 Vin
rlabel nsubdiffcont 16887 9284 16921 9357 7 Vin
rlabel metal1 6105 7900 6105 7900 7 CLKin
port 3 w
rlabel metal1 19753 12322 19753 12322 7 ENPin
port 4 w
rlabel metal1 10510 11916 10510 11916 7 GND
<< end >>
