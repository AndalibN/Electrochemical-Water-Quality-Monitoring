magic
tech sky130A
timestamp 1667977299
<< pwell >>
rect -128 -255 128 255
<< nmos >>
rect -30 -150 30 150
<< ndiff >>
rect -59 144 -30 150
rect -59 -144 -53 144
rect -36 -144 -30 144
rect -59 -150 -30 -144
rect 30 144 59 150
rect 30 -144 36 144
rect 53 -144 59 144
rect 30 -150 59 -144
<< ndiffc >>
rect -53 -144 -36 144
rect 36 -144 53 144
<< psubdiff >>
rect -110 220 -62 237
rect 62 220 110 237
rect -110 189 -93 220
rect 93 189 110 220
rect -110 -220 -93 -189
rect 93 -220 110 -189
rect -110 -237 -62 -220
rect 62 -237 110 -220
<< psubdiffcont >>
rect -62 220 62 237
rect -110 -189 -93 189
rect 93 -189 110 189
rect -62 -237 62 -220
<< poly >>
rect -30 186 30 194
rect -30 169 -22 186
rect 22 169 30 186
rect -30 150 30 169
rect -30 -169 30 -150
rect -30 -186 -22 -169
rect 22 -186 30 -169
rect -30 -194 30 -186
<< polycont >>
rect -22 169 22 186
rect -22 -186 22 -169
<< locali >>
rect -110 220 -62 237
rect 62 220 110 237
rect -110 189 -93 220
rect 93 189 110 220
rect -30 169 -22 186
rect 22 169 30 186
rect -53 144 -36 152
rect -53 -152 -36 -144
rect 36 144 53 152
rect 36 -152 53 -144
rect -30 -186 -22 -169
rect 22 -186 30 -169
rect -110 -220 -93 -189
rect 93 -220 110 -189
rect -110 -237 -62 -220
rect 62 -237 110 -220
<< viali >>
rect -22 169 22 186
rect -53 -144 -36 144
rect 36 -144 53 144
rect -22 -186 22 -169
<< metal1 >>
rect -28 186 28 189
rect -28 169 -22 186
rect 22 169 28 186
rect -28 166 28 169
rect -56 144 -33 150
rect -56 -144 -53 144
rect -36 -144 -33 144
rect -56 -150 -33 -144
rect 33 144 56 150
rect 33 -144 36 144
rect 53 -144 56 144
rect 33 -150 56 -144
rect -28 -169 28 -166
rect -28 -186 -22 -169
rect 22 -186 28 -169
rect -28 -189 28 -186
<< properties >>
string FIXED_BBOX -101 -228 101 228
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
