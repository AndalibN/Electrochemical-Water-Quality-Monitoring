magic
tech sky130A
magscale 1 2
timestamp 1665001199
<< nmos >>
rect -229 -1400 -29 1400
rect 29 -1400 229 1400
<< ndiff >>
rect -287 1388 -229 1400
rect -287 -1388 -275 1388
rect -241 -1388 -229 1388
rect -287 -1400 -229 -1388
rect -29 1388 29 1400
rect -29 -1388 -17 1388
rect 17 -1388 29 1388
rect -29 -1400 29 -1388
rect 229 1388 287 1400
rect 229 -1388 241 1388
rect 275 -1388 287 1388
rect 229 -1400 287 -1388
<< ndiffc >>
rect -275 -1388 -241 1388
rect -17 -1388 17 1388
rect 241 -1388 275 1388
<< poly >>
rect -229 1472 -29 1488
rect -229 1438 -213 1472
rect -45 1438 -29 1472
rect -229 1400 -29 1438
rect 29 1472 229 1488
rect 29 1438 45 1472
rect 213 1438 229 1472
rect 29 1400 229 1438
rect -229 -1438 -29 -1400
rect -229 -1472 -213 -1438
rect -45 -1472 -29 -1438
rect -229 -1488 -29 -1472
rect 29 -1438 229 -1400
rect 29 -1472 45 -1438
rect 213 -1472 229 -1438
rect 29 -1488 229 -1472
<< polycont >>
rect -213 1438 -45 1472
rect 45 1438 213 1472
rect -213 -1472 -45 -1438
rect 45 -1472 213 -1438
<< locali >>
rect -229 1438 -213 1472
rect -45 1438 -29 1472
rect 29 1438 45 1472
rect 213 1438 229 1472
rect -275 1388 -241 1404
rect -275 -1404 -241 -1388
rect -17 1388 17 1404
rect -17 -1404 17 -1388
rect 241 1388 275 1404
rect 241 -1404 275 -1388
rect -229 -1472 -213 -1438
rect -45 -1472 -29 -1438
rect 29 -1472 45 -1438
rect 213 -1472 229 -1438
<< viali >>
rect -213 1438 -45 1472
rect 45 1438 213 1472
rect -275 -1388 -241 1388
rect -17 -1388 17 1388
rect 241 -1388 275 1388
rect -213 -1472 -45 -1438
rect 45 -1472 213 -1438
<< metal1 >>
rect -225 1472 -33 1478
rect -225 1438 -213 1472
rect -45 1438 -33 1472
rect -225 1432 -33 1438
rect 33 1472 225 1478
rect 33 1438 45 1472
rect 213 1438 225 1472
rect 33 1432 225 1438
rect -281 1388 -235 1400
rect -281 -1388 -275 1388
rect -241 -1388 -235 1388
rect -281 -1400 -235 -1388
rect -23 1388 23 1400
rect -23 -1388 -17 1388
rect 17 -1388 23 1388
rect -23 -1400 23 -1388
rect 235 1388 281 1400
rect 235 -1388 241 1388
rect 275 -1388 281 1388
rect 235 -1400 281 -1388
rect -225 -1438 -33 -1432
rect -225 -1472 -213 -1438
rect -45 -1472 -33 -1438
rect -225 -1478 -33 -1472
rect 33 -1438 225 -1432
rect 33 -1472 45 -1438
rect 213 -1472 225 -1438
rect 33 -1478 225 -1472
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 14 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
