magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect 15505 14880 20461 15135
rect 15504 14810 20461 14880
rect 15504 12624 20455 14810
rect 5395 10446 10351 10701
rect 10738 10558 10843 10560
rect 11140 10558 11310 10597
rect 10724 10468 10725 10558
rect 10736 10470 11310 10558
rect 10736 10468 10843 10470
rect 5395 10376 10352 10446
rect 5401 8190 10352 10376
rect 10724 8625 10843 10468
rect 11140 10443 11310 10470
rect 11151 10437 11261 10443
rect 11151 8625 11260 10437
rect 16402 8710 17024 9416
rect 10724 8547 11261 8625
rect 10739 8544 11261 8547
rect 10703 6261 11317 7604
rect 16396 7314 17018 8020
rect 17368 7809 18302 9465
rect 19869 8705 20491 9411
rect 19865 7374 20487 8080
rect 10764 5647 11317 6261
rect 19883 6132 20505 6838
rect 10703 5507 11317 5647
rect 12956 5388 15053 6002
rect 15026 2643 16162 2647
rect 15024 2642 16162 2643
<< pwell >>
rect 11762 12020 14556 15070
rect 15655 11778 20283 12016
rect 10725 11066 11266 11206
rect 10725 10782 10886 11066
rect 11105 10782 11266 11066
rect 10725 10642 11266 10782
rect 15655 10993 15881 11778
rect 20064 10993 20283 11778
rect 15655 10755 20283 10993
rect 16322 9795 17006 9934
rect 16322 9550 16506 9795
rect 16822 9550 17006 9795
rect 16322 9416 17006 9550
rect 19789 9791 20473 9930
rect 19789 9546 19973 9791
rect 20289 9546 20473 9791
rect 16318 8400 17002 8539
rect 10727 8069 11268 8209
rect 10727 7785 10888 8069
rect 11107 7785 11268 8069
rect 16318 8155 16502 8400
rect 16818 8155 17002 8400
rect 16318 8021 17002 8155
rect 10727 7645 11268 7785
rect 5576 7344 10204 7582
rect 5576 6559 5795 7344
rect 9978 6559 10204 7344
rect 5576 6321 10204 6559
rect 18503 9297 19465 9454
rect 19789 9412 20473 9546
rect 18503 7982 18640 9297
rect 19328 7982 19465 9297
rect 19786 8460 20470 8599
rect 19786 8215 19970 8460
rect 20286 8215 20470 8460
rect 19786 8081 20470 8215
rect 18502 7825 19465 7982
rect 18503 7824 18640 7825
rect 19328 7824 19465 7825
rect 19800 7218 20484 7357
rect 19800 6973 19984 7218
rect 20300 6973 20484 7218
rect 19800 6839 20484 6973
rect 12351 5810 12915 5971
rect 12351 5591 12491 5810
rect 12775 5591 12915 5810
rect 12351 5430 12915 5591
<< psubdiff >>
rect 11788 14791 14530 15044
rect 11788 12377 12181 14791
rect 14187 12377 14530 14791
rect 11788 12046 14530 12377
rect 15681 11941 20257 11990
rect 15681 11907 15746 11941
rect 15780 11907 15814 11941
rect 15848 11907 15882 11941
rect 15916 11907 15950 11941
rect 15984 11907 16018 11941
rect 16052 11907 16086 11941
rect 16120 11907 16154 11941
rect 16188 11907 16222 11941
rect 16256 11907 16290 11941
rect 16324 11907 16358 11941
rect 16392 11907 16426 11941
rect 16460 11907 16494 11941
rect 16528 11907 16562 11941
rect 16596 11907 16630 11941
rect 16664 11907 16698 11941
rect 16732 11907 16766 11941
rect 16800 11907 16834 11941
rect 16868 11907 16902 11941
rect 16936 11907 16970 11941
rect 17004 11907 17038 11941
rect 17072 11907 17106 11941
rect 17140 11907 17174 11941
rect 17208 11907 17242 11941
rect 17276 11907 17310 11941
rect 17344 11907 17378 11941
rect 17412 11907 17446 11941
rect 17480 11907 17514 11941
rect 17548 11907 17582 11941
rect 17616 11907 17650 11941
rect 17684 11907 17718 11941
rect 17752 11907 17786 11941
rect 17820 11907 17854 11941
rect 17888 11907 17922 11941
rect 17956 11907 17990 11941
rect 18024 11907 18058 11941
rect 18092 11907 18126 11941
rect 18160 11907 18194 11941
rect 18228 11907 18262 11941
rect 18296 11907 18330 11941
rect 18364 11907 18398 11941
rect 18432 11907 18466 11941
rect 18500 11907 18534 11941
rect 18568 11907 18602 11941
rect 18636 11907 18670 11941
rect 18704 11907 18738 11941
rect 18772 11907 18806 11941
rect 18840 11907 18874 11941
rect 18908 11907 18942 11941
rect 18976 11907 19010 11941
rect 19044 11907 19078 11941
rect 19112 11907 19146 11941
rect 19180 11907 19214 11941
rect 19248 11907 19282 11941
rect 19316 11907 19350 11941
rect 19384 11907 19418 11941
rect 19452 11907 19486 11941
rect 19520 11907 19554 11941
rect 19588 11907 19622 11941
rect 19656 11907 19690 11941
rect 19724 11907 19758 11941
rect 19792 11907 19826 11941
rect 19860 11907 19894 11941
rect 19928 11907 19962 11941
rect 19996 11907 20030 11941
rect 20064 11907 20098 11941
rect 20132 11907 20166 11941
rect 20200 11907 20257 11941
rect 15681 11873 20257 11907
rect 15681 11839 15746 11873
rect 15780 11839 20166 11873
rect 20200 11839 20257 11873
rect 15681 11805 20257 11839
rect 15681 11771 15746 11805
rect 15780 11804 20166 11805
rect 15780 11771 15855 11804
rect 15681 11737 15855 11771
rect 15681 11703 15746 11737
rect 15780 11703 15855 11737
rect 15681 11669 15855 11703
rect 15681 11635 15746 11669
rect 15780 11635 15855 11669
rect 15681 11601 15855 11635
rect 15681 11567 15746 11601
rect 15780 11567 15855 11601
rect 15681 11533 15855 11567
rect 15681 11499 15746 11533
rect 15780 11499 15855 11533
rect 15681 11465 15855 11499
rect 15681 11431 15746 11465
rect 15780 11431 15855 11465
rect 15681 11397 15855 11431
rect 15681 11363 15746 11397
rect 15780 11363 15855 11397
rect 15681 11329 15855 11363
rect 15681 11295 15746 11329
rect 15780 11295 15855 11329
rect 15681 11261 15855 11295
rect 15681 11227 15746 11261
rect 15780 11227 15855 11261
rect 15681 11193 15855 11227
rect 10751 11151 11240 11180
rect 10751 11117 10789 11151
rect 10823 11117 10876 11151
rect 10910 11117 10944 11151
rect 10978 11117 11012 11151
rect 11046 11117 11080 11151
rect 11114 11117 11168 11151
rect 11202 11117 11240 11151
rect 10751 11092 11240 11117
rect 10751 11076 10860 11092
rect 10751 11042 10789 11076
rect 10823 11042 10860 11076
rect 10751 11008 10860 11042
rect 10751 10974 10789 11008
rect 10823 10974 10860 11008
rect 10751 10940 10860 10974
rect 10751 10906 10789 10940
rect 10823 10906 10860 10940
rect 10751 10872 10860 10906
rect 10751 10838 10789 10872
rect 10823 10838 10860 10872
rect 10751 10804 10860 10838
rect 10751 10770 10789 10804
rect 10823 10770 10860 10804
rect 10751 10756 10860 10770
rect 11131 11076 11240 11092
rect 11131 11042 11168 11076
rect 11202 11042 11240 11076
rect 11131 11008 11240 11042
rect 11131 10974 11168 11008
rect 11202 10974 11240 11008
rect 11131 10940 11240 10974
rect 11131 10906 11168 10940
rect 11202 10906 11240 10940
rect 11131 10872 11240 10906
rect 11131 10838 11168 10872
rect 11202 10838 11240 10872
rect 11131 10804 11240 10838
rect 11131 10770 11168 10804
rect 11202 10770 11240 10804
rect 15681 11159 15746 11193
rect 15780 11159 15855 11193
rect 15681 11125 15855 11159
rect 15681 11091 15746 11125
rect 15780 11091 15855 11125
rect 15681 11057 15855 11091
rect 15681 11023 15746 11057
rect 15780 11023 15855 11057
rect 15681 10989 15855 11023
rect 15681 10955 15746 10989
rect 15780 10967 15855 10989
rect 20090 11771 20166 11804
rect 20200 11771 20257 11805
rect 20090 11737 20257 11771
rect 20090 11703 20166 11737
rect 20200 11703 20257 11737
rect 20090 11669 20257 11703
rect 20090 11635 20166 11669
rect 20200 11635 20257 11669
rect 20090 11601 20257 11635
rect 20090 11567 20166 11601
rect 20200 11567 20257 11601
rect 20090 11533 20257 11567
rect 20090 11499 20166 11533
rect 20200 11499 20257 11533
rect 20090 11465 20257 11499
rect 20090 11431 20166 11465
rect 20200 11431 20257 11465
rect 20090 11397 20257 11431
rect 20090 11363 20166 11397
rect 20200 11363 20257 11397
rect 20090 11329 20257 11363
rect 20090 11295 20166 11329
rect 20200 11295 20257 11329
rect 20090 11261 20257 11295
rect 20090 11227 20166 11261
rect 20200 11227 20257 11261
rect 20090 11193 20257 11227
rect 20090 11159 20166 11193
rect 20200 11159 20257 11193
rect 20090 11125 20257 11159
rect 20090 11091 20166 11125
rect 20200 11091 20257 11125
rect 20090 11057 20257 11091
rect 20090 11023 20166 11057
rect 20200 11023 20257 11057
rect 20090 10989 20257 11023
rect 20090 10967 20166 10989
rect 15780 10955 20166 10967
rect 20200 10955 20257 10989
rect 15681 10921 20257 10955
rect 15681 10819 15746 10921
rect 20200 10819 20257 10921
rect 15681 10781 20257 10819
rect 11131 10756 11240 10770
rect 10751 10728 11240 10756
rect 10751 10694 10789 10728
rect 10823 10694 10876 10728
rect 10910 10694 10944 10728
rect 10978 10694 11012 10728
rect 11046 10694 11080 10728
rect 11114 10694 11168 10728
rect 11202 10694 11240 10728
rect 10751 10668 11240 10694
rect 16348 9877 16980 9908
rect 16348 9843 16395 9877
rect 16429 9843 16509 9877
rect 16543 9843 16577 9877
rect 16611 9843 16645 9877
rect 16679 9843 16713 9877
rect 16747 9843 16781 9877
rect 16815 9843 16895 9877
rect 16929 9843 16980 9877
rect 16348 9821 16980 9843
rect 16348 9793 16480 9821
rect 16348 9759 16395 9793
rect 16429 9759 16480 9793
rect 16348 9725 16480 9759
rect 16348 9691 16395 9725
rect 16429 9691 16480 9725
rect 16348 9657 16480 9691
rect 16348 9623 16395 9657
rect 16429 9623 16480 9657
rect 16348 9589 16480 9623
rect 16348 9555 16395 9589
rect 16429 9555 16480 9589
rect 16348 9524 16480 9555
rect 16848 9793 16980 9821
rect 16848 9759 16895 9793
rect 16929 9759 16980 9793
rect 16848 9725 16980 9759
rect 16848 9691 16895 9725
rect 16929 9691 16980 9725
rect 16848 9657 16980 9691
rect 16848 9623 16895 9657
rect 16929 9623 16980 9657
rect 16848 9589 16980 9623
rect 16848 9555 16895 9589
rect 16929 9555 16980 9589
rect 16848 9524 16980 9555
rect 16348 9501 16980 9524
rect 16348 9467 16395 9501
rect 16429 9467 16509 9501
rect 16543 9467 16577 9501
rect 16611 9467 16645 9501
rect 16679 9467 16713 9501
rect 16747 9467 16781 9501
rect 16815 9467 16895 9501
rect 16929 9467 16980 9501
rect 16348 9442 16980 9467
rect 19815 9873 20447 9904
rect 19815 9839 19862 9873
rect 19896 9839 19976 9873
rect 20010 9839 20044 9873
rect 20078 9839 20112 9873
rect 20146 9839 20180 9873
rect 20214 9839 20248 9873
rect 20282 9839 20362 9873
rect 20396 9839 20447 9873
rect 19815 9817 20447 9839
rect 19815 9789 19947 9817
rect 19815 9755 19862 9789
rect 19896 9755 19947 9789
rect 19815 9721 19947 9755
rect 19815 9687 19862 9721
rect 19896 9687 19947 9721
rect 19815 9653 19947 9687
rect 19815 9619 19862 9653
rect 19896 9619 19947 9653
rect 19815 9585 19947 9619
rect 19815 9551 19862 9585
rect 19896 9551 19947 9585
rect 19815 9520 19947 9551
rect 20315 9789 20447 9817
rect 20315 9755 20362 9789
rect 20396 9755 20447 9789
rect 20315 9721 20447 9755
rect 20315 9687 20362 9721
rect 20396 9687 20447 9721
rect 20315 9653 20447 9687
rect 20315 9619 20362 9653
rect 20396 9619 20447 9653
rect 20315 9585 20447 9619
rect 20315 9551 20362 9585
rect 20396 9551 20447 9585
rect 20315 9520 20447 9551
rect 19815 9497 20447 9520
rect 19815 9463 19862 9497
rect 19896 9463 19976 9497
rect 20010 9463 20044 9497
rect 20078 9463 20112 9497
rect 20146 9463 20180 9497
rect 20214 9463 20248 9497
rect 20282 9463 20362 9497
rect 20396 9463 20447 9497
rect 19815 9438 20447 9463
rect 16344 8482 16976 8513
rect 16344 8448 16391 8482
rect 16425 8448 16505 8482
rect 16539 8448 16573 8482
rect 16607 8448 16641 8482
rect 16675 8448 16709 8482
rect 16743 8448 16777 8482
rect 16811 8448 16891 8482
rect 16925 8448 16976 8482
rect 16344 8426 16976 8448
rect 16344 8398 16476 8426
rect 16344 8364 16391 8398
rect 16425 8364 16476 8398
rect 16344 8330 16476 8364
rect 16344 8296 16391 8330
rect 16425 8296 16476 8330
rect 16344 8262 16476 8296
rect 16344 8228 16391 8262
rect 16425 8228 16476 8262
rect 16344 8194 16476 8228
rect 10753 8154 11242 8183
rect 10753 8120 10791 8154
rect 10825 8120 10878 8154
rect 10912 8120 10946 8154
rect 10980 8120 11014 8154
rect 11048 8120 11082 8154
rect 11116 8120 11170 8154
rect 11204 8120 11242 8154
rect 10753 8095 11242 8120
rect 10753 8079 10862 8095
rect 10753 8045 10791 8079
rect 10825 8045 10862 8079
rect 10753 8011 10862 8045
rect 10753 7977 10791 8011
rect 10825 7977 10862 8011
rect 10753 7943 10862 7977
rect 10753 7909 10791 7943
rect 10825 7909 10862 7943
rect 10753 7875 10862 7909
rect 10753 7841 10791 7875
rect 10825 7841 10862 7875
rect 10753 7807 10862 7841
rect 10753 7773 10791 7807
rect 10825 7773 10862 7807
rect 10753 7759 10862 7773
rect 11133 8079 11242 8095
rect 11133 8045 11170 8079
rect 11204 8045 11242 8079
rect 16344 8160 16391 8194
rect 16425 8160 16476 8194
rect 16344 8129 16476 8160
rect 16844 8398 16976 8426
rect 16844 8364 16891 8398
rect 16925 8364 16976 8398
rect 16844 8330 16976 8364
rect 16844 8296 16891 8330
rect 16925 8296 16976 8330
rect 16844 8262 16976 8296
rect 16844 8228 16891 8262
rect 16925 8228 16976 8262
rect 16844 8194 16976 8228
rect 16844 8160 16891 8194
rect 16925 8160 16976 8194
rect 16844 8129 16976 8160
rect 16344 8106 16976 8129
rect 16344 8072 16391 8106
rect 16425 8072 16505 8106
rect 16539 8072 16573 8106
rect 16607 8072 16641 8106
rect 16675 8072 16709 8106
rect 16743 8072 16777 8106
rect 16811 8072 16891 8106
rect 16925 8072 16976 8106
rect 16344 8047 16976 8072
rect 11133 8011 11242 8045
rect 11133 7977 11170 8011
rect 11204 7977 11242 8011
rect 11133 7943 11242 7977
rect 11133 7909 11170 7943
rect 11204 7909 11242 7943
rect 11133 7875 11242 7909
rect 11133 7841 11170 7875
rect 11204 7841 11242 7875
rect 11133 7807 11242 7841
rect 11133 7773 11170 7807
rect 11204 7773 11242 7807
rect 11133 7759 11242 7773
rect 10753 7731 11242 7759
rect 10753 7697 10791 7731
rect 10825 7697 10878 7731
rect 10912 7697 10946 7731
rect 10980 7697 11014 7731
rect 11048 7697 11082 7731
rect 11116 7697 11170 7731
rect 11204 7697 11242 7731
rect 10753 7671 11242 7697
rect 5602 7507 10178 7556
rect 5602 7473 5659 7507
rect 5693 7473 5727 7507
rect 5761 7473 5795 7507
rect 5829 7473 5863 7507
rect 5897 7473 5931 7507
rect 5965 7473 5999 7507
rect 6033 7473 6067 7507
rect 6101 7473 6135 7507
rect 6169 7473 6203 7507
rect 6237 7473 6271 7507
rect 6305 7473 6339 7507
rect 6373 7473 6407 7507
rect 6441 7473 6475 7507
rect 6509 7473 6543 7507
rect 6577 7473 6611 7507
rect 6645 7473 6679 7507
rect 6713 7473 6747 7507
rect 6781 7473 6815 7507
rect 6849 7473 6883 7507
rect 6917 7473 6951 7507
rect 6985 7473 7019 7507
rect 7053 7473 7087 7507
rect 7121 7473 7155 7507
rect 7189 7473 7223 7507
rect 7257 7473 7291 7507
rect 7325 7473 7359 7507
rect 7393 7473 7427 7507
rect 7461 7473 7495 7507
rect 7529 7473 7563 7507
rect 7597 7473 7631 7507
rect 7665 7473 7699 7507
rect 7733 7473 7767 7507
rect 7801 7473 7835 7507
rect 7869 7473 7903 7507
rect 7937 7473 7971 7507
rect 8005 7473 8039 7507
rect 8073 7473 8107 7507
rect 8141 7473 8175 7507
rect 8209 7473 8243 7507
rect 8277 7473 8311 7507
rect 8345 7473 8379 7507
rect 8413 7473 8447 7507
rect 8481 7473 8515 7507
rect 8549 7473 8583 7507
rect 8617 7473 8651 7507
rect 8685 7473 8719 7507
rect 8753 7473 8787 7507
rect 8821 7473 8855 7507
rect 8889 7473 8923 7507
rect 8957 7473 8991 7507
rect 9025 7473 9059 7507
rect 9093 7473 9127 7507
rect 9161 7473 9195 7507
rect 9229 7473 9263 7507
rect 9297 7473 9331 7507
rect 9365 7473 9399 7507
rect 9433 7473 9467 7507
rect 9501 7473 9535 7507
rect 9569 7473 9603 7507
rect 9637 7473 9671 7507
rect 9705 7473 9739 7507
rect 9773 7473 9807 7507
rect 9841 7473 9875 7507
rect 9909 7473 9943 7507
rect 9977 7473 10011 7507
rect 10045 7473 10079 7507
rect 10113 7473 10178 7507
rect 5602 7439 10178 7473
rect 5602 7405 5659 7439
rect 5693 7405 10079 7439
rect 10113 7405 10178 7439
rect 5602 7371 10178 7405
rect 5602 7337 5659 7371
rect 5693 7370 10079 7371
rect 5693 7337 5769 7370
rect 5602 7303 5769 7337
rect 5602 7269 5659 7303
rect 5693 7269 5769 7303
rect 5602 7235 5769 7269
rect 5602 7201 5659 7235
rect 5693 7201 5769 7235
rect 5602 7167 5769 7201
rect 5602 7133 5659 7167
rect 5693 7133 5769 7167
rect 5602 7099 5769 7133
rect 5602 7065 5659 7099
rect 5693 7065 5769 7099
rect 5602 7031 5769 7065
rect 5602 6997 5659 7031
rect 5693 6997 5769 7031
rect 5602 6963 5769 6997
rect 5602 6929 5659 6963
rect 5693 6929 5769 6963
rect 5602 6895 5769 6929
rect 5602 6861 5659 6895
rect 5693 6861 5769 6895
rect 5602 6827 5769 6861
rect 5602 6793 5659 6827
rect 5693 6793 5769 6827
rect 5602 6759 5769 6793
rect 5602 6725 5659 6759
rect 5693 6725 5769 6759
rect 5602 6691 5769 6725
rect 5602 6657 5659 6691
rect 5693 6657 5769 6691
rect 5602 6623 5769 6657
rect 5602 6589 5659 6623
rect 5693 6589 5769 6623
rect 5602 6555 5769 6589
rect 5602 6521 5659 6555
rect 5693 6533 5769 6555
rect 10004 7337 10079 7370
rect 10113 7337 10178 7371
rect 10004 7303 10178 7337
rect 10004 7269 10079 7303
rect 10113 7269 10178 7303
rect 10004 7235 10178 7269
rect 10004 7201 10079 7235
rect 10113 7201 10178 7235
rect 10004 7167 10178 7201
rect 10004 7133 10079 7167
rect 10113 7133 10178 7167
rect 10004 7099 10178 7133
rect 10004 7065 10079 7099
rect 10113 7065 10178 7099
rect 10004 7031 10178 7065
rect 10004 6997 10079 7031
rect 10113 6997 10178 7031
rect 10004 6963 10178 6997
rect 10004 6929 10079 6963
rect 10113 6929 10178 6963
rect 10004 6895 10178 6929
rect 10004 6861 10079 6895
rect 10113 6861 10178 6895
rect 10004 6827 10178 6861
rect 10004 6793 10079 6827
rect 10113 6793 10178 6827
rect 10004 6759 10178 6793
rect 10004 6725 10079 6759
rect 10113 6725 10178 6759
rect 10004 6691 10178 6725
rect 10004 6657 10079 6691
rect 10113 6657 10178 6691
rect 10004 6623 10178 6657
rect 10004 6589 10079 6623
rect 10113 6589 10178 6623
rect 10004 6555 10178 6589
rect 10004 6533 10079 6555
rect 5693 6521 10079 6533
rect 10113 6521 10178 6555
rect 5602 6487 10178 6521
rect 5602 6385 5659 6487
rect 10113 6385 10178 6487
rect 5602 6347 10178 6385
rect 18529 9392 19439 9428
rect 18529 9358 18554 9392
rect 18588 9358 18627 9392
rect 18661 9358 18695 9392
rect 18729 9358 18763 9392
rect 18797 9358 18831 9392
rect 18865 9358 18899 9392
rect 18933 9358 18967 9392
rect 19001 9358 19035 9392
rect 19069 9358 19103 9392
rect 19137 9358 19171 9392
rect 19205 9358 19239 9392
rect 19273 9358 19307 9392
rect 19341 9358 19380 9392
rect 19414 9358 19439 9392
rect 18529 9323 19439 9358
rect 18529 9303 18614 9323
rect 18529 9269 18554 9303
rect 18588 9269 18614 9303
rect 18529 9235 18614 9269
rect 18529 9201 18554 9235
rect 18588 9201 18614 9235
rect 18529 9167 18614 9201
rect 18529 9133 18554 9167
rect 18588 9133 18614 9167
rect 18529 9099 18614 9133
rect 18529 9065 18554 9099
rect 18588 9065 18614 9099
rect 18529 9031 18614 9065
rect 18529 8997 18554 9031
rect 18588 8997 18614 9031
rect 18529 8963 18614 8997
rect 18529 8929 18554 8963
rect 18588 8929 18614 8963
rect 18529 8895 18614 8929
rect 18529 8861 18554 8895
rect 18588 8861 18614 8895
rect 18529 8827 18614 8861
rect 18529 8793 18554 8827
rect 18588 8793 18614 8827
rect 18529 8759 18614 8793
rect 18529 8725 18554 8759
rect 18588 8725 18614 8759
rect 18529 8691 18614 8725
rect 18529 8657 18554 8691
rect 18588 8657 18614 8691
rect 18529 8623 18614 8657
rect 18529 8589 18554 8623
rect 18588 8589 18614 8623
rect 18529 8555 18614 8589
rect 18529 8521 18554 8555
rect 18588 8521 18614 8555
rect 18529 8487 18614 8521
rect 18529 8453 18554 8487
rect 18588 8453 18614 8487
rect 18529 8419 18614 8453
rect 18529 8385 18554 8419
rect 18588 8385 18614 8419
rect 18529 8351 18614 8385
rect 18529 8317 18554 8351
rect 18588 8317 18614 8351
rect 18529 8283 18614 8317
rect 18529 8249 18554 8283
rect 18588 8249 18614 8283
rect 18529 8215 18614 8249
rect 18529 8181 18554 8215
rect 18588 8181 18614 8215
rect 18529 8147 18614 8181
rect 18529 8113 18554 8147
rect 18588 8113 18614 8147
rect 18529 8079 18614 8113
rect 18529 8045 18554 8079
rect 18588 8045 18614 8079
rect 18529 8011 18614 8045
rect 18529 7977 18554 8011
rect 18588 7977 18614 8011
rect 18529 7956 18614 7977
rect 19354 9303 19439 9323
rect 19354 9269 19380 9303
rect 19414 9269 19439 9303
rect 19354 9235 19439 9269
rect 19354 9201 19380 9235
rect 19414 9201 19439 9235
rect 19354 9167 19439 9201
rect 19354 9133 19380 9167
rect 19414 9133 19439 9167
rect 19354 9099 19439 9133
rect 19354 9065 19380 9099
rect 19414 9065 19439 9099
rect 19354 9031 19439 9065
rect 19354 8997 19380 9031
rect 19414 8997 19439 9031
rect 19354 8963 19439 8997
rect 19354 8929 19380 8963
rect 19414 8929 19439 8963
rect 19354 8895 19439 8929
rect 19354 8861 19380 8895
rect 19414 8861 19439 8895
rect 19354 8827 19439 8861
rect 19354 8793 19380 8827
rect 19414 8793 19439 8827
rect 19354 8759 19439 8793
rect 19354 8725 19380 8759
rect 19414 8725 19439 8759
rect 19354 8691 19439 8725
rect 19354 8657 19380 8691
rect 19414 8657 19439 8691
rect 19354 8623 19439 8657
rect 19354 8589 19380 8623
rect 19414 8589 19439 8623
rect 19354 8555 19439 8589
rect 19354 8521 19380 8555
rect 19414 8521 19439 8555
rect 19354 8487 19439 8521
rect 19354 8453 19380 8487
rect 19414 8453 19439 8487
rect 19354 8419 19439 8453
rect 19354 8385 19380 8419
rect 19414 8385 19439 8419
rect 19354 8351 19439 8385
rect 19354 8317 19380 8351
rect 19414 8317 19439 8351
rect 19354 8283 19439 8317
rect 19354 8249 19380 8283
rect 19414 8249 19439 8283
rect 19354 8215 19439 8249
rect 19354 8181 19380 8215
rect 19414 8181 19439 8215
rect 19354 8147 19439 8181
rect 19354 8113 19380 8147
rect 19414 8113 19439 8147
rect 19354 8079 19439 8113
rect 19812 8542 20444 8573
rect 19812 8508 19859 8542
rect 19893 8508 19973 8542
rect 20007 8508 20041 8542
rect 20075 8508 20109 8542
rect 20143 8508 20177 8542
rect 20211 8508 20245 8542
rect 20279 8508 20359 8542
rect 20393 8508 20444 8542
rect 19812 8486 20444 8508
rect 19812 8458 19944 8486
rect 19812 8424 19859 8458
rect 19893 8424 19944 8458
rect 19812 8390 19944 8424
rect 19812 8356 19859 8390
rect 19893 8356 19944 8390
rect 19812 8322 19944 8356
rect 19812 8288 19859 8322
rect 19893 8288 19944 8322
rect 19812 8254 19944 8288
rect 19812 8220 19859 8254
rect 19893 8220 19944 8254
rect 19812 8189 19944 8220
rect 20312 8458 20444 8486
rect 20312 8424 20359 8458
rect 20393 8424 20444 8458
rect 20312 8390 20444 8424
rect 20312 8356 20359 8390
rect 20393 8356 20444 8390
rect 20312 8322 20444 8356
rect 20312 8288 20359 8322
rect 20393 8288 20444 8322
rect 20312 8254 20444 8288
rect 20312 8220 20359 8254
rect 20393 8220 20444 8254
rect 20312 8189 20444 8220
rect 19812 8166 20444 8189
rect 19812 8132 19859 8166
rect 19893 8132 19973 8166
rect 20007 8132 20041 8166
rect 20075 8132 20109 8166
rect 20143 8132 20177 8166
rect 20211 8132 20245 8166
rect 20279 8132 20359 8166
rect 20393 8132 20444 8166
rect 19812 8107 20444 8132
rect 19354 8045 19380 8079
rect 19414 8045 19439 8079
rect 19354 8011 19439 8045
rect 19354 7977 19380 8011
rect 19414 7977 19439 8011
rect 19354 7956 19439 7977
rect 18528 7921 19439 7956
rect 18528 7887 18554 7921
rect 18588 7887 18627 7921
rect 18661 7887 18695 7921
rect 18729 7887 18763 7921
rect 18797 7887 18831 7921
rect 18865 7887 18899 7921
rect 18933 7887 18967 7921
rect 19001 7887 19035 7921
rect 19069 7887 19103 7921
rect 19137 7887 19171 7921
rect 19205 7887 19239 7921
rect 19273 7887 19307 7921
rect 19341 7887 19380 7921
rect 19414 7887 19439 7921
rect 18528 7851 19439 7887
rect 18529 7850 18614 7851
rect 19354 7850 19439 7851
rect 19826 7300 20458 7331
rect 19826 7266 19873 7300
rect 19907 7266 19987 7300
rect 20021 7266 20055 7300
rect 20089 7266 20123 7300
rect 20157 7266 20191 7300
rect 20225 7266 20259 7300
rect 20293 7266 20373 7300
rect 20407 7266 20458 7300
rect 19826 7244 20458 7266
rect 19826 7216 19958 7244
rect 19826 7182 19873 7216
rect 19907 7182 19958 7216
rect 19826 7148 19958 7182
rect 19826 7114 19873 7148
rect 19907 7114 19958 7148
rect 19826 7080 19958 7114
rect 19826 7046 19873 7080
rect 19907 7046 19958 7080
rect 19826 7012 19958 7046
rect 19826 6978 19873 7012
rect 19907 6978 19958 7012
rect 19826 6947 19958 6978
rect 20326 7216 20458 7244
rect 20326 7182 20373 7216
rect 20407 7182 20458 7216
rect 20326 7148 20458 7182
rect 20326 7114 20373 7148
rect 20407 7114 20458 7148
rect 20326 7080 20458 7114
rect 20326 7046 20373 7080
rect 20407 7046 20458 7080
rect 20326 7012 20458 7046
rect 20326 6978 20373 7012
rect 20407 6978 20458 7012
rect 20326 6947 20458 6978
rect 19826 6924 20458 6947
rect 19826 6890 19873 6924
rect 19907 6890 19987 6924
rect 20021 6890 20055 6924
rect 20089 6890 20123 6924
rect 20157 6890 20191 6924
rect 20225 6890 20259 6924
rect 20293 6890 20373 6924
rect 20407 6890 20458 6924
rect 19826 6865 20458 6890
rect 12377 5907 12889 5945
rect 12377 5873 12405 5907
rect 12439 5873 12481 5907
rect 12515 5873 12549 5907
rect 12583 5873 12617 5907
rect 12651 5873 12685 5907
rect 12719 5873 12753 5907
rect 12787 5873 12828 5907
rect 12862 5873 12889 5907
rect 12377 5836 12889 5873
rect 12377 5819 12465 5836
rect 12377 5785 12405 5819
rect 12439 5785 12465 5819
rect 12377 5751 12465 5785
rect 12377 5717 12405 5751
rect 12439 5717 12465 5751
rect 12377 5683 12465 5717
rect 12377 5649 12405 5683
rect 12439 5649 12465 5683
rect 12377 5615 12465 5649
rect 12377 5581 12405 5615
rect 12439 5581 12465 5615
rect 12377 5565 12465 5581
rect 12801 5819 12889 5836
rect 12801 5785 12828 5819
rect 12862 5785 12889 5819
rect 12801 5751 12889 5785
rect 12801 5717 12828 5751
rect 12862 5717 12889 5751
rect 12801 5683 12889 5717
rect 12801 5649 12828 5683
rect 12862 5649 12889 5683
rect 12801 5615 12889 5649
rect 12801 5581 12828 5615
rect 12862 5581 12889 5615
rect 12801 5565 12889 5581
rect 12377 5528 12889 5565
rect 12377 5494 12405 5528
rect 12439 5494 12481 5528
rect 12515 5494 12549 5528
rect 12583 5494 12617 5528
rect 12651 5494 12685 5528
rect 12719 5494 12753 5528
rect 12787 5494 12828 5528
rect 12862 5494 12889 5528
rect 12377 5456 12889 5494
<< nsubdiff >>
rect 15679 15053 20254 15086
rect 15679 15019 15740 15053
rect 15774 15031 20254 15053
rect 15774 15019 15879 15031
rect 15679 14997 15879 15019
rect 15913 14997 15947 15031
rect 15981 14997 16015 15031
rect 16049 14997 16083 15031
rect 16117 14997 16151 15031
rect 16185 14997 16219 15031
rect 16253 14997 16287 15031
rect 16321 14997 16355 15031
rect 16389 14997 16423 15031
rect 16457 14997 16491 15031
rect 16525 14997 16559 15031
rect 16593 14997 16627 15031
rect 16661 14997 16695 15031
rect 16729 14997 16763 15031
rect 16797 14997 16831 15031
rect 16865 14997 16899 15031
rect 16933 14997 16967 15031
rect 17001 14997 17035 15031
rect 17069 14997 17103 15031
rect 17137 14997 17171 15031
rect 17205 14997 17239 15031
rect 17273 14997 17307 15031
rect 17341 14997 17375 15031
rect 17409 14997 17443 15031
rect 17477 14997 17511 15031
rect 17545 14997 17579 15031
rect 17613 14997 17647 15031
rect 17681 14997 17715 15031
rect 17749 14997 17783 15031
rect 17817 14997 17851 15031
rect 17885 14997 17919 15031
rect 17953 14997 17987 15031
rect 18021 14997 18055 15031
rect 18089 14997 18123 15031
rect 18157 14997 18191 15031
rect 18225 14997 18259 15031
rect 18293 14997 18327 15031
rect 18361 14997 18395 15031
rect 18429 14997 18463 15031
rect 18497 14997 18531 15031
rect 18565 14997 18599 15031
rect 18633 14997 18667 15031
rect 18701 14997 18735 15031
rect 18769 14997 18803 15031
rect 18837 14997 18871 15031
rect 18905 14997 18939 15031
rect 18973 14997 19007 15031
rect 19041 14997 19075 15031
rect 19109 14997 19143 15031
rect 19177 14997 19211 15031
rect 19245 14997 19279 15031
rect 19313 14997 19347 15031
rect 19381 14997 19415 15031
rect 19449 14997 19483 15031
rect 19517 14997 19551 15031
rect 19585 14997 19619 15031
rect 19653 14997 19687 15031
rect 19721 14997 19755 15031
rect 19789 14997 19823 15031
rect 19857 14997 19891 15031
rect 19925 14997 19959 15031
rect 19993 14997 20027 15031
rect 20061 15026 20254 15031
rect 20061 14997 20152 15026
rect 15679 14992 20152 14997
rect 20186 14992 20254 15026
rect 15679 14985 20254 14992
rect 15679 14951 15740 14985
rect 15774 14954 20254 14985
rect 15774 14951 15855 14954
rect 15679 14917 15855 14951
rect 15679 14883 15740 14917
rect 15774 14883 15855 14917
rect 15679 14849 15855 14883
rect 15679 14815 15740 14849
rect 15774 14815 15855 14849
rect 15679 14781 15855 14815
rect 15679 14747 15740 14781
rect 15774 14747 15855 14781
rect 15679 14713 15855 14747
rect 15679 14679 15740 14713
rect 15774 14679 15855 14713
rect 15679 14645 15855 14679
rect 20078 14920 20152 14954
rect 20186 14920 20254 14954
rect 20078 14886 20254 14920
rect 20078 14852 20152 14886
rect 20186 14852 20254 14886
rect 20078 14818 20254 14852
rect 20078 14784 20152 14818
rect 20186 14784 20254 14818
rect 20078 14750 20254 14784
rect 20078 14716 20152 14750
rect 20186 14716 20254 14750
rect 20078 14682 20254 14716
rect 15679 14611 15740 14645
rect 15774 14611 15855 14645
rect 15679 14577 15855 14611
rect 15679 14543 15740 14577
rect 15774 14543 15855 14577
rect 15679 14509 15855 14543
rect 15679 14475 15740 14509
rect 15774 14475 15855 14509
rect 15679 14441 15855 14475
rect 15679 14407 15740 14441
rect 15774 14407 15855 14441
rect 15679 14394 15855 14407
rect 17454 14592 17629 14661
rect 17454 14558 17525 14592
rect 17559 14558 17629 14592
rect 17454 14524 17629 14558
rect 17454 14490 17525 14524
rect 17559 14490 17629 14524
rect 17454 14456 17629 14490
rect 17454 14422 17525 14456
rect 17559 14422 17629 14456
rect 15679 14373 15854 14394
rect 15679 14339 15740 14373
rect 15774 14339 15854 14373
rect 15679 14305 15854 14339
rect 15679 14271 15740 14305
rect 15774 14271 15854 14305
rect 17454 14388 17629 14422
rect 17454 14354 17525 14388
rect 17559 14354 17629 14388
rect 17454 14320 17629 14354
rect 17454 14286 17525 14320
rect 17559 14286 17629 14320
rect 17454 14272 17629 14286
rect 15679 14237 15854 14271
rect 15679 14203 15740 14237
rect 15774 14203 15854 14237
rect 15679 14169 15854 14203
rect 15679 14135 15740 14169
rect 15774 14135 15854 14169
rect 15679 14101 15854 14135
rect 15679 14067 15740 14101
rect 15774 14067 15854 14101
rect 15679 14033 15854 14067
rect 15679 13999 15740 14033
rect 15774 13999 15854 14033
rect 15679 13965 15854 13999
rect 15679 13931 15740 13965
rect 15774 13931 15854 13965
rect 15679 13897 15854 13931
rect 15679 13863 15740 13897
rect 15774 13863 15854 13897
rect 15679 13829 15854 13863
rect 15679 13795 15740 13829
rect 15774 13795 15854 13829
rect 15679 13761 15854 13795
rect 15679 13727 15740 13761
rect 15774 13727 15854 13761
rect 15679 13693 15854 13727
rect 15679 13659 15740 13693
rect 15774 13659 15854 13693
rect 15679 13625 15854 13659
rect 15679 13591 15740 13625
rect 15774 13591 15854 13625
rect 15679 13557 15854 13591
rect 15679 13523 15740 13557
rect 15774 13523 15854 13557
rect 15679 13489 15854 13523
rect 15679 13455 15740 13489
rect 15774 13455 15854 13489
rect 15679 13421 15854 13455
rect 15679 13387 15740 13421
rect 15774 13387 15854 13421
rect 15679 13353 15854 13387
rect 15679 13319 15740 13353
rect 15774 13319 15854 13353
rect 15679 13285 15854 13319
rect 15679 13251 15740 13285
rect 15774 13251 15854 13285
rect 15679 13217 15854 13251
rect 15679 13183 15740 13217
rect 15774 13183 15854 13217
rect 15679 13149 15854 13183
rect 15679 13115 15740 13149
rect 15774 13115 15854 13149
rect 17453 14166 17629 14272
rect 17453 14132 17525 14166
rect 17559 14132 17629 14166
rect 17453 14098 17629 14132
rect 17453 14064 17525 14098
rect 17559 14064 17629 14098
rect 17453 14030 17629 14064
rect 17453 13996 17525 14030
rect 17559 13996 17629 14030
rect 17453 13962 17629 13996
rect 17453 13928 17525 13962
rect 17559 13928 17629 13962
rect 17453 13894 17629 13928
rect 17453 13860 17525 13894
rect 17559 13860 17629 13894
rect 17453 13826 17629 13860
rect 17453 13792 17525 13826
rect 17559 13792 17629 13826
rect 17453 13758 17629 13792
rect 17453 13724 17525 13758
rect 17559 13724 17629 13758
rect 17453 13690 17629 13724
rect 17453 13656 17525 13690
rect 17559 13656 17629 13690
rect 17453 13622 17629 13656
rect 17453 13588 17525 13622
rect 17559 13588 17629 13622
rect 17453 13554 17629 13588
rect 17453 13520 17525 13554
rect 17559 13520 17629 13554
rect 17453 13486 17629 13520
rect 17453 13452 17525 13486
rect 17559 13452 17629 13486
rect 17453 13418 17629 13452
rect 17453 13384 17525 13418
rect 17559 13384 17629 13418
rect 17453 13350 17629 13384
rect 17453 13316 17525 13350
rect 17559 13316 17629 13350
rect 17453 13282 17629 13316
rect 17453 13248 17525 13282
rect 17559 13248 17629 13282
rect 17453 13214 17629 13248
rect 17453 13180 17525 13214
rect 17559 13180 17629 13214
rect 17453 13126 17629 13180
rect 19230 14579 19407 14657
rect 19230 14545 19304 14579
rect 19338 14545 19407 14579
rect 19230 14511 19407 14545
rect 19230 14477 19304 14511
rect 19338 14477 19407 14511
rect 19230 14443 19407 14477
rect 19230 14409 19304 14443
rect 19338 14409 19407 14443
rect 19230 14375 19407 14409
rect 19230 14341 19304 14375
rect 19338 14341 19407 14375
rect 19230 14307 19407 14341
rect 19230 14273 19304 14307
rect 19338 14273 19407 14307
rect 19230 14239 19407 14273
rect 19230 14205 19304 14239
rect 19338 14209 19407 14239
rect 20078 14648 20152 14682
rect 20186 14648 20254 14682
rect 20078 14614 20254 14648
rect 20078 14580 20152 14614
rect 20186 14580 20254 14614
rect 20078 14546 20254 14580
rect 20078 14512 20152 14546
rect 20186 14512 20254 14546
rect 20078 14478 20254 14512
rect 20078 14444 20152 14478
rect 20186 14444 20254 14478
rect 20078 14341 20254 14444
rect 20078 14307 20152 14341
rect 20186 14307 20254 14341
rect 20078 14273 20254 14307
rect 20078 14239 20152 14273
rect 20186 14239 20254 14273
rect 19338 14205 19405 14209
rect 19230 14171 19405 14205
rect 19230 14137 19304 14171
rect 19338 14137 19405 14171
rect 19230 14103 19405 14137
rect 19230 14069 19304 14103
rect 19338 14069 19405 14103
rect 19230 14035 19405 14069
rect 19230 14001 19304 14035
rect 19338 14001 19405 14035
rect 19230 13967 19405 14001
rect 19230 13933 19304 13967
rect 19338 13933 19405 13967
rect 19230 13899 19405 13933
rect 19230 13865 19304 13899
rect 19338 13865 19405 13899
rect 19230 13831 19405 13865
rect 19230 13797 19304 13831
rect 19338 13797 19405 13831
rect 19230 13763 19405 13797
rect 19230 13729 19304 13763
rect 19338 13729 19405 13763
rect 19230 13695 19405 13729
rect 19230 13661 19304 13695
rect 19338 13661 19405 13695
rect 19230 13627 19405 13661
rect 19230 13593 19304 13627
rect 19338 13593 19405 13627
rect 19230 13559 19405 13593
rect 19230 13525 19304 13559
rect 19338 13525 19405 13559
rect 19230 13491 19405 13525
rect 19230 13457 19304 13491
rect 19338 13457 19405 13491
rect 19230 13423 19405 13457
rect 19230 13389 19304 13423
rect 19338 13389 19405 13423
rect 19230 13355 19405 13389
rect 19230 13321 19304 13355
rect 19338 13321 19405 13355
rect 19230 13287 19405 13321
rect 19230 13253 19304 13287
rect 19338 13253 19405 13287
rect 19230 13219 19405 13253
rect 19230 13185 19304 13219
rect 19338 13185 19405 13219
rect 19230 13128 19405 13185
rect 20078 14205 20254 14239
rect 20078 14171 20152 14205
rect 20186 14171 20254 14205
rect 20078 14137 20254 14171
rect 20078 14103 20152 14137
rect 20186 14103 20254 14137
rect 20078 14069 20254 14103
rect 20078 14035 20152 14069
rect 20186 14035 20254 14069
rect 20078 14001 20254 14035
rect 20078 13967 20152 14001
rect 20186 13967 20254 14001
rect 20078 13933 20254 13967
rect 20078 13899 20152 13933
rect 20186 13899 20254 13933
rect 20078 13865 20254 13899
rect 20078 13831 20152 13865
rect 20186 13831 20254 13865
rect 20078 13797 20254 13831
rect 20078 13763 20152 13797
rect 20186 13763 20254 13797
rect 20078 13729 20254 13763
rect 20078 13695 20152 13729
rect 20186 13695 20254 13729
rect 20078 13661 20254 13695
rect 20078 13627 20152 13661
rect 20186 13627 20254 13661
rect 20078 13593 20254 13627
rect 20078 13559 20152 13593
rect 20186 13559 20254 13593
rect 20078 13525 20254 13559
rect 20078 13491 20152 13525
rect 20186 13491 20254 13525
rect 20078 13457 20254 13491
rect 20078 13423 20152 13457
rect 20186 13423 20254 13457
rect 20078 13389 20254 13423
rect 20078 13355 20152 13389
rect 20186 13355 20254 13389
rect 20078 13321 20254 13355
rect 20078 13287 20152 13321
rect 20186 13287 20254 13321
rect 20078 13253 20254 13287
rect 20078 13219 20152 13253
rect 20186 13219 20254 13253
rect 20078 13185 20254 13219
rect 20078 13151 20152 13185
rect 20186 13151 20254 13185
rect 15679 13081 15854 13115
rect 15679 13047 15740 13081
rect 15774 13047 15854 13081
rect 15679 13013 15854 13047
rect 15679 12979 15740 13013
rect 15774 12990 15854 13013
rect 20078 13117 20254 13151
rect 20078 13083 20152 13117
rect 20186 13083 20254 13117
rect 20078 13049 20254 13083
rect 20078 13015 20152 13049
rect 20186 13015 20254 13049
rect 20078 12990 20254 13015
rect 15774 12979 20254 12990
rect 15679 12945 20254 12979
rect 15679 12843 15740 12945
rect 20194 12843 20254 12945
rect 15679 12805 20254 12843
rect 5602 10619 10177 10652
rect 5602 10597 10082 10619
rect 5602 10592 5794 10597
rect 5602 10558 5670 10592
rect 5704 10563 5794 10592
rect 5828 10563 5862 10597
rect 5896 10563 5930 10597
rect 5964 10563 5998 10597
rect 6032 10563 6066 10597
rect 6100 10563 6134 10597
rect 6168 10563 6202 10597
rect 6236 10563 6270 10597
rect 6304 10563 6338 10597
rect 6372 10563 6406 10597
rect 6440 10563 6474 10597
rect 6508 10563 6542 10597
rect 6576 10563 6610 10597
rect 6644 10563 6678 10597
rect 6712 10563 6746 10597
rect 6780 10563 6814 10597
rect 6848 10563 6882 10597
rect 6916 10563 6950 10597
rect 6984 10563 7018 10597
rect 7052 10563 7086 10597
rect 7120 10563 7154 10597
rect 7188 10563 7222 10597
rect 7256 10563 7290 10597
rect 7324 10563 7358 10597
rect 7392 10563 7426 10597
rect 7460 10563 7494 10597
rect 7528 10563 7562 10597
rect 7596 10563 7630 10597
rect 7664 10563 7698 10597
rect 7732 10563 7766 10597
rect 7800 10563 7834 10597
rect 7868 10563 7902 10597
rect 7936 10563 7970 10597
rect 8004 10563 8038 10597
rect 8072 10563 8106 10597
rect 8140 10563 8174 10597
rect 8208 10563 8242 10597
rect 8276 10563 8310 10597
rect 8344 10563 8378 10597
rect 8412 10563 8446 10597
rect 8480 10563 8514 10597
rect 8548 10563 8582 10597
rect 8616 10563 8650 10597
rect 8684 10563 8718 10597
rect 8752 10563 8786 10597
rect 8820 10563 8854 10597
rect 8888 10563 8922 10597
rect 8956 10563 8990 10597
rect 9024 10563 9058 10597
rect 9092 10563 9126 10597
rect 9160 10563 9194 10597
rect 9228 10563 9262 10597
rect 9296 10563 9330 10597
rect 9364 10563 9398 10597
rect 9432 10563 9466 10597
rect 9500 10563 9534 10597
rect 9568 10563 9602 10597
rect 9636 10563 9670 10597
rect 9704 10563 9738 10597
rect 9772 10563 9806 10597
rect 9840 10563 9874 10597
rect 9908 10563 9942 10597
rect 9976 10585 10082 10597
rect 10116 10585 10177 10619
rect 9976 10563 10177 10585
rect 5704 10558 10177 10563
rect 10738 10558 10843 10560
rect 5602 10551 10177 10558
rect 5602 10520 10082 10551
rect 5602 10486 5778 10520
rect 5602 10452 5669 10486
rect 5703 10452 5778 10486
rect 5602 10418 5778 10452
rect 5602 10384 5669 10418
rect 5703 10384 5778 10418
rect 5602 10350 5778 10384
rect 5602 10316 5669 10350
rect 5703 10316 5778 10350
rect 5602 10282 5778 10316
rect 5602 10248 5669 10282
rect 5703 10248 5778 10282
rect 5602 10214 5778 10248
rect 10001 10517 10082 10520
rect 10116 10517 10177 10551
rect 10001 10483 10177 10517
rect 10001 10449 10082 10483
rect 10116 10449 10177 10483
rect 10736 10533 11261 10558
rect 10736 10499 10776 10533
rect 10810 10499 10879 10533
rect 10913 10499 10947 10533
rect 10981 10499 11015 10533
rect 11049 10499 11083 10533
rect 11117 10499 11187 10533
rect 11221 10499 11261 10533
rect 10736 10470 11261 10499
rect 10001 10415 10177 10449
rect 10001 10381 10082 10415
rect 10116 10381 10177 10415
rect 10001 10347 10177 10381
rect 10001 10313 10082 10347
rect 10116 10313 10177 10347
rect 10001 10279 10177 10313
rect 10001 10245 10082 10279
rect 10116 10245 10177 10279
rect 5602 10180 5669 10214
rect 5703 10180 5778 10214
rect 5602 10146 5778 10180
rect 5602 10112 5669 10146
rect 5703 10112 5778 10146
rect 5602 10078 5778 10112
rect 5602 10044 5669 10078
rect 5703 10044 5778 10078
rect 5602 10010 5778 10044
rect 5602 9976 5669 10010
rect 5703 9976 5778 10010
rect 5602 9907 5778 9976
rect 5602 9873 5670 9907
rect 5704 9873 5778 9907
rect 5602 9839 5778 9873
rect 5602 9805 5670 9839
rect 5704 9805 5778 9839
rect 5602 9771 5778 9805
rect 6449 10145 6626 10223
rect 6449 10111 6518 10145
rect 6552 10111 6626 10145
rect 6449 10077 6626 10111
rect 6449 10043 6518 10077
rect 6552 10043 6626 10077
rect 6449 10009 6626 10043
rect 6449 9975 6518 10009
rect 6552 9975 6626 10009
rect 6449 9941 6626 9975
rect 6449 9907 6518 9941
rect 6552 9907 6626 9941
rect 6449 9873 6626 9907
rect 6449 9839 6518 9873
rect 6552 9839 6626 9873
rect 6449 9805 6626 9839
rect 6449 9775 6518 9805
rect 5602 9737 5670 9771
rect 5704 9737 5778 9771
rect 5602 9703 5778 9737
rect 5602 9669 5670 9703
rect 5704 9669 5778 9703
rect 5602 9635 5778 9669
rect 5602 9601 5670 9635
rect 5704 9601 5778 9635
rect 5602 9567 5778 9601
rect 5602 9533 5670 9567
rect 5704 9533 5778 9567
rect 5602 9499 5778 9533
rect 5602 9465 5670 9499
rect 5704 9465 5778 9499
rect 5602 9431 5778 9465
rect 5602 9397 5670 9431
rect 5704 9397 5778 9431
rect 5602 9363 5778 9397
rect 5602 9329 5670 9363
rect 5704 9329 5778 9363
rect 5602 9295 5778 9329
rect 5602 9261 5670 9295
rect 5704 9261 5778 9295
rect 5602 9227 5778 9261
rect 5602 9193 5670 9227
rect 5704 9193 5778 9227
rect 5602 9159 5778 9193
rect 5602 9125 5670 9159
rect 5704 9125 5778 9159
rect 5602 9091 5778 9125
rect 5602 9057 5670 9091
rect 5704 9057 5778 9091
rect 5602 9023 5778 9057
rect 5602 8989 5670 9023
rect 5704 8989 5778 9023
rect 5602 8955 5778 8989
rect 5602 8921 5670 8955
rect 5704 8921 5778 8955
rect 5602 8887 5778 8921
rect 5602 8853 5670 8887
rect 5704 8853 5778 8887
rect 5602 8819 5778 8853
rect 5602 8785 5670 8819
rect 5704 8785 5778 8819
rect 5602 8751 5778 8785
rect 5602 8717 5670 8751
rect 5704 8717 5778 8751
rect 5602 8683 5778 8717
rect 6451 9771 6518 9775
rect 6552 9771 6626 9805
rect 6451 9737 6626 9771
rect 6451 9703 6518 9737
rect 6552 9703 6626 9737
rect 6451 9669 6626 9703
rect 6451 9635 6518 9669
rect 6552 9635 6626 9669
rect 6451 9601 6626 9635
rect 6451 9567 6518 9601
rect 6552 9567 6626 9601
rect 6451 9533 6626 9567
rect 6451 9499 6518 9533
rect 6552 9499 6626 9533
rect 6451 9465 6626 9499
rect 6451 9431 6518 9465
rect 6552 9431 6626 9465
rect 6451 9397 6626 9431
rect 6451 9363 6518 9397
rect 6552 9363 6626 9397
rect 6451 9329 6626 9363
rect 6451 9295 6518 9329
rect 6552 9295 6626 9329
rect 6451 9261 6626 9295
rect 6451 9227 6518 9261
rect 6552 9227 6626 9261
rect 6451 9193 6626 9227
rect 6451 9159 6518 9193
rect 6552 9159 6626 9193
rect 6451 9125 6626 9159
rect 6451 9091 6518 9125
rect 6552 9091 6626 9125
rect 6451 9057 6626 9091
rect 6451 9023 6518 9057
rect 6552 9023 6626 9057
rect 6451 8989 6626 9023
rect 6451 8955 6518 8989
rect 6552 8955 6626 8989
rect 6451 8921 6626 8955
rect 6451 8887 6518 8921
rect 6552 8887 6626 8921
rect 6451 8853 6626 8887
rect 6451 8819 6518 8853
rect 6552 8819 6626 8853
rect 6451 8785 6626 8819
rect 6451 8751 6518 8785
rect 6552 8751 6626 8785
rect 6451 8694 6626 8751
rect 8227 10175 8402 10227
rect 8227 10141 8296 10175
rect 8330 10141 8402 10175
rect 8227 10107 8402 10141
rect 8227 10073 8296 10107
rect 8330 10073 8402 10107
rect 8227 10039 8402 10073
rect 8227 10005 8296 10039
rect 8330 10005 8402 10039
rect 8227 9971 8402 10005
rect 8227 9937 8296 9971
rect 8330 9937 8402 9971
rect 10001 10211 10177 10245
rect 10001 10177 10082 10211
rect 10116 10177 10177 10211
rect 10001 10143 10177 10177
rect 10001 10109 10082 10143
rect 10116 10109 10177 10143
rect 10001 10075 10177 10109
rect 10001 10041 10082 10075
rect 10116 10041 10177 10075
rect 10001 10007 10177 10041
rect 10001 9973 10082 10007
rect 10116 9973 10177 10007
rect 10001 9960 10177 9973
rect 8227 9903 8402 9937
rect 8227 9869 8296 9903
rect 8330 9869 8402 9903
rect 8227 9838 8402 9869
rect 10002 9939 10177 9960
rect 10002 9905 10082 9939
rect 10116 9905 10177 9939
rect 10002 9871 10177 9905
rect 8227 9835 8403 9838
rect 8227 9801 8296 9835
rect 8330 9801 8403 9835
rect 8227 9732 8403 9801
rect 8227 9698 8297 9732
rect 8331 9698 8403 9732
rect 8227 9664 8403 9698
rect 8227 9630 8297 9664
rect 8331 9630 8403 9664
rect 8227 9596 8403 9630
rect 8227 9562 8297 9596
rect 8331 9562 8403 9596
rect 8227 9528 8403 9562
rect 8227 9494 8297 9528
rect 8331 9494 8403 9528
rect 8227 9460 8403 9494
rect 8227 9426 8297 9460
rect 8331 9426 8403 9460
rect 8227 9392 8403 9426
rect 8227 9358 8297 9392
rect 8331 9358 8403 9392
rect 8227 9324 8403 9358
rect 8227 9290 8297 9324
rect 8331 9290 8403 9324
rect 8227 9256 8403 9290
rect 8227 9222 8297 9256
rect 8331 9222 8403 9256
rect 8227 9188 8403 9222
rect 8227 9154 8297 9188
rect 8331 9154 8403 9188
rect 8227 9120 8403 9154
rect 8227 9086 8297 9120
rect 8331 9086 8403 9120
rect 8227 9052 8403 9086
rect 8227 9018 8297 9052
rect 8331 9018 8403 9052
rect 8227 8984 8403 9018
rect 8227 8950 8297 8984
rect 8331 8950 8403 8984
rect 8227 8916 8403 8950
rect 8227 8882 8297 8916
rect 8331 8882 8403 8916
rect 8227 8848 8403 8882
rect 8227 8814 8297 8848
rect 8331 8814 8403 8848
rect 8227 8780 8403 8814
rect 8227 8746 8297 8780
rect 8331 8746 8403 8780
rect 8227 8692 8403 8746
rect 10002 9837 10082 9871
rect 10116 9837 10177 9871
rect 10002 9803 10177 9837
rect 10002 9769 10082 9803
rect 10116 9769 10177 9803
rect 10002 9735 10177 9769
rect 10002 9701 10082 9735
rect 10116 9701 10177 9735
rect 10002 9667 10177 9701
rect 10002 9633 10082 9667
rect 10116 9633 10177 9667
rect 10002 9599 10177 9633
rect 10002 9565 10082 9599
rect 10116 9565 10177 9599
rect 10002 9531 10177 9565
rect 10002 9497 10082 9531
rect 10116 9497 10177 9531
rect 10002 9463 10177 9497
rect 10002 9429 10082 9463
rect 10116 9429 10177 9463
rect 10002 9395 10177 9429
rect 10002 9361 10082 9395
rect 10116 9361 10177 9395
rect 10002 9327 10177 9361
rect 10002 9293 10082 9327
rect 10116 9293 10177 9327
rect 10002 9259 10177 9293
rect 10002 9225 10082 9259
rect 10116 9225 10177 9259
rect 10002 9191 10177 9225
rect 10002 9157 10082 9191
rect 10116 9157 10177 9191
rect 10002 9123 10177 9157
rect 10002 9089 10082 9123
rect 10116 9089 10177 9123
rect 10002 9055 10177 9089
rect 10002 9021 10082 9055
rect 10116 9021 10177 9055
rect 10002 8987 10177 9021
rect 10002 8953 10082 8987
rect 10116 8953 10177 8987
rect 10002 8919 10177 8953
rect 10002 8885 10082 8919
rect 10116 8885 10177 8919
rect 10002 8851 10177 8885
rect 10002 8817 10082 8851
rect 10116 8817 10177 8851
rect 10002 8783 10177 8817
rect 10002 8749 10082 8783
rect 10116 8749 10177 8783
rect 10002 8715 10177 8749
rect 5602 8649 5670 8683
rect 5704 8649 5778 8683
rect 5602 8615 5778 8649
rect 5602 8581 5670 8615
rect 5704 8581 5778 8615
rect 5602 8556 5778 8581
rect 10002 8681 10082 8715
rect 10116 8681 10177 8715
rect 10002 8647 10177 8681
rect 10002 8613 10082 8647
rect 10116 8613 10177 8647
rect 10002 8579 10177 8613
rect 10002 8556 10082 8579
rect 5602 8545 10082 8556
rect 10116 8545 10177 8579
rect 10738 10448 10843 10470
rect 10738 10414 10776 10448
rect 10810 10414 10843 10448
rect 10738 10380 10843 10414
rect 10738 10346 10776 10380
rect 10810 10346 10843 10380
rect 10738 10312 10843 10346
rect 10738 10278 10776 10312
rect 10810 10278 10843 10312
rect 10738 10244 10843 10278
rect 10738 10210 10776 10244
rect 10810 10210 10843 10244
rect 10738 10176 10843 10210
rect 10738 10142 10776 10176
rect 10810 10142 10843 10176
rect 10738 10108 10843 10142
rect 10738 10074 10776 10108
rect 10810 10074 10843 10108
rect 10738 10040 10843 10074
rect 10738 10006 10776 10040
rect 10810 10006 10843 10040
rect 10738 9972 10843 10006
rect 10738 9938 10776 9972
rect 10810 9938 10843 9972
rect 10738 9904 10843 9938
rect 10738 9870 10776 9904
rect 10810 9870 10843 9904
rect 10738 9836 10843 9870
rect 10738 9802 10776 9836
rect 10810 9802 10843 9836
rect 10738 9768 10843 9802
rect 10738 9734 10776 9768
rect 10810 9734 10843 9768
rect 10738 9700 10843 9734
rect 10738 9666 10776 9700
rect 10810 9666 10843 9700
rect 10738 9632 10843 9666
rect 10738 9598 10776 9632
rect 10810 9598 10843 9632
rect 10738 9564 10843 9598
rect 10738 9530 10776 9564
rect 10810 9530 10843 9564
rect 10738 9496 10843 9530
rect 10738 9462 10776 9496
rect 10810 9462 10843 9496
rect 10738 9428 10843 9462
rect 10738 9394 10776 9428
rect 10810 9394 10843 9428
rect 10738 9360 10843 9394
rect 10738 9326 10776 9360
rect 10810 9326 10843 9360
rect 10738 9292 10843 9326
rect 10738 9258 10776 9292
rect 10810 9258 10843 9292
rect 10738 9224 10843 9258
rect 10738 9190 10776 9224
rect 10810 9190 10843 9224
rect 10738 9156 10843 9190
rect 10738 9122 10776 9156
rect 10810 9122 10843 9156
rect 10738 9088 10843 9122
rect 10738 9054 10776 9088
rect 10810 9054 10843 9088
rect 10738 9020 10843 9054
rect 10738 8986 10776 9020
rect 10810 8986 10843 9020
rect 10738 8952 10843 8986
rect 10738 8918 10776 8952
rect 10810 8918 10843 8952
rect 10738 8884 10843 8918
rect 10738 8850 10776 8884
rect 10810 8850 10843 8884
rect 10738 8816 10843 8850
rect 10738 8782 10776 8816
rect 10810 8782 10843 8816
rect 10738 8748 10843 8782
rect 10738 8714 10776 8748
rect 10810 8714 10843 8748
rect 10738 8680 10843 8714
rect 10738 8646 10776 8680
rect 10810 8646 10843 8680
rect 10738 8625 10843 8646
rect 11151 10448 11261 10470
rect 11151 10414 11187 10448
rect 11221 10437 11261 10448
rect 11221 10414 11260 10437
rect 11151 10380 11260 10414
rect 11151 10346 11187 10380
rect 11221 10346 11260 10380
rect 11151 10312 11260 10346
rect 11151 10278 11187 10312
rect 11221 10278 11260 10312
rect 11151 10244 11260 10278
rect 11151 10210 11187 10244
rect 11221 10210 11260 10244
rect 11151 10176 11260 10210
rect 11151 10142 11187 10176
rect 11221 10142 11260 10176
rect 11151 10108 11260 10142
rect 11151 10074 11187 10108
rect 11221 10074 11260 10108
rect 11151 10040 11260 10074
rect 11151 10006 11187 10040
rect 11221 10006 11260 10040
rect 11151 9972 11260 10006
rect 11151 9938 11187 9972
rect 11221 9938 11260 9972
rect 11151 9904 11260 9938
rect 11151 9870 11187 9904
rect 11221 9870 11260 9904
rect 11151 9836 11260 9870
rect 11151 9802 11187 9836
rect 11221 9802 11260 9836
rect 11151 9768 11260 9802
rect 11151 9734 11187 9768
rect 11221 9734 11260 9768
rect 11151 9700 11260 9734
rect 11151 9666 11187 9700
rect 11221 9666 11260 9700
rect 11151 9632 11260 9666
rect 11151 9598 11187 9632
rect 11221 9598 11260 9632
rect 11151 9564 11260 9598
rect 11151 9530 11187 9564
rect 11221 9530 11260 9564
rect 11151 9496 11260 9530
rect 11151 9462 11187 9496
rect 11221 9462 11260 9496
rect 11151 9428 11260 9462
rect 11151 9394 11187 9428
rect 11221 9394 11260 9428
rect 11151 9360 11260 9394
rect 17411 9407 18264 9426
rect 11151 9326 11187 9360
rect 11221 9326 11260 9360
rect 11151 9292 11260 9326
rect 11151 9258 11187 9292
rect 11221 9258 11260 9292
rect 11151 9224 11260 9258
rect 11151 9190 11187 9224
rect 11221 9190 11260 9224
rect 11151 9156 11260 9190
rect 11151 9122 11187 9156
rect 11221 9122 11260 9156
rect 11151 9088 11260 9122
rect 11151 9054 11187 9088
rect 11221 9054 11260 9088
rect 11151 9020 11260 9054
rect 11151 8986 11187 9020
rect 11221 8986 11260 9020
rect 11151 8952 11260 8986
rect 11151 8918 11187 8952
rect 11221 8918 11260 8952
rect 11151 8884 11260 8918
rect 11151 8850 11187 8884
rect 11221 8850 11260 8884
rect 11151 8816 11260 8850
rect 11151 8782 11187 8816
rect 11221 8782 11260 8816
rect 11151 8748 11260 8782
rect 11151 8714 11187 8748
rect 11221 8714 11260 8748
rect 16441 9357 16977 9380
rect 16441 9323 16490 9357
rect 16524 9323 16588 9357
rect 16622 9323 16656 9357
rect 16690 9323 16724 9357
rect 16758 9323 16792 9357
rect 16826 9323 16890 9357
rect 16924 9323 16977 9357
rect 16441 9303 16977 9323
rect 16441 9285 16574 9303
rect 16441 9251 16490 9285
rect 16524 9251 16574 9285
rect 16441 9217 16574 9251
rect 16441 9183 16490 9217
rect 16524 9183 16574 9217
rect 16441 9149 16574 9183
rect 16441 9115 16490 9149
rect 16524 9115 16574 9149
rect 16441 9081 16574 9115
rect 16441 9047 16490 9081
rect 16524 9047 16574 9081
rect 16441 9013 16574 9047
rect 16441 8979 16490 9013
rect 16524 8979 16574 9013
rect 16441 8945 16574 8979
rect 16441 8911 16490 8945
rect 16524 8911 16574 8945
rect 16441 8877 16574 8911
rect 16441 8843 16490 8877
rect 16524 8843 16574 8877
rect 16441 8825 16574 8843
rect 16839 9285 16977 9303
rect 16839 9251 16890 9285
rect 16924 9251 16977 9285
rect 16839 9217 16977 9251
rect 16839 9183 16890 9217
rect 16924 9183 16977 9217
rect 16839 9149 16977 9183
rect 16839 9115 16890 9149
rect 16924 9115 16977 9149
rect 16839 9081 16977 9115
rect 16839 9047 16890 9081
rect 16924 9047 16977 9081
rect 16839 9013 16977 9047
rect 16839 8979 16890 9013
rect 16924 8979 16977 9013
rect 16839 8945 16977 8979
rect 16839 8911 16890 8945
rect 16924 8911 16977 8945
rect 16839 8877 16977 8911
rect 16839 8843 16890 8877
rect 16924 8843 16977 8877
rect 16839 8825 16977 8843
rect 16441 8805 16977 8825
rect 16441 8771 16490 8805
rect 16524 8771 16588 8805
rect 16622 8771 16656 8805
rect 16690 8771 16724 8805
rect 16758 8771 16792 8805
rect 16826 8771 16890 8805
rect 16924 8771 16977 8805
rect 16441 8747 16977 8771
rect 17411 9373 17443 9407
rect 17477 9373 17519 9407
rect 17553 9373 17587 9407
rect 17621 9373 17655 9407
rect 17689 9373 17723 9407
rect 17757 9373 17791 9407
rect 17825 9373 17859 9407
rect 17893 9373 17927 9407
rect 17961 9373 17995 9407
rect 18029 9373 18063 9407
rect 18097 9373 18131 9407
rect 18165 9373 18203 9407
rect 18237 9373 18264 9407
rect 17411 9359 18264 9373
rect 17411 9312 17509 9359
rect 17411 9278 17443 9312
rect 17477 9278 17509 9312
rect 17411 9244 17509 9278
rect 17411 9210 17443 9244
rect 17477 9210 17509 9244
rect 17411 9176 17509 9210
rect 17411 9142 17443 9176
rect 17477 9142 17509 9176
rect 17411 9108 17509 9142
rect 17411 9074 17443 9108
rect 17477 9074 17509 9108
rect 17411 9040 17509 9074
rect 17411 9006 17443 9040
rect 17477 9006 17509 9040
rect 17411 8972 17509 9006
rect 17411 8938 17443 8972
rect 17477 8938 17509 8972
rect 18179 9312 18264 9359
rect 18179 9278 18203 9312
rect 18237 9278 18264 9312
rect 18179 9244 18264 9278
rect 18179 9210 18203 9244
rect 18237 9210 18264 9244
rect 18179 9176 18264 9210
rect 18179 9142 18203 9176
rect 18237 9142 18264 9176
rect 18179 9108 18264 9142
rect 18179 9074 18203 9108
rect 18237 9074 18264 9108
rect 18179 9040 18264 9074
rect 18179 9006 18203 9040
rect 18237 9006 18264 9040
rect 18179 8972 18264 9006
rect 17411 8904 17509 8938
rect 17411 8870 17443 8904
rect 17477 8870 17509 8904
rect 17566 8938 18083 8959
rect 17566 8904 17602 8938
rect 17636 8904 17670 8938
rect 17704 8904 17738 8938
rect 17772 8904 17806 8938
rect 17840 8904 17874 8938
rect 17908 8904 17942 8938
rect 17976 8904 18010 8938
rect 18044 8904 18083 8938
rect 17566 8883 18083 8904
rect 18179 8938 18203 8972
rect 18237 8938 18264 8972
rect 18179 8904 18264 8938
rect 17411 8836 17509 8870
rect 17411 8802 17443 8836
rect 17477 8802 17509 8836
rect 17411 8768 17509 8802
rect 11151 8680 11260 8714
rect 11151 8646 11187 8680
rect 11221 8646 11260 8680
rect 11151 8625 11260 8646
rect 17411 8734 17443 8768
rect 17477 8734 17509 8768
rect 17411 8700 17509 8734
rect 17411 8666 17443 8700
rect 17477 8666 17509 8700
rect 17411 8632 17509 8666
rect 10738 8604 11261 8625
rect 10738 8570 10776 8604
rect 10810 8570 10879 8604
rect 10913 8570 10947 8604
rect 10981 8570 11015 8604
rect 11049 8570 11083 8604
rect 11117 8570 11187 8604
rect 11221 8570 11261 8604
rect 10738 8549 11261 8570
rect 5602 8511 10177 8545
rect 10739 8544 11261 8549
rect 17411 8598 17443 8632
rect 17477 8598 17509 8632
rect 17411 8564 17509 8598
rect 17411 8530 17443 8564
rect 17477 8530 17509 8564
rect 5602 8409 5662 8511
rect 10116 8409 10177 8511
rect 5602 8371 10177 8409
rect 17411 8496 17509 8530
rect 17411 8462 17443 8496
rect 17477 8462 17509 8496
rect 17411 8428 17509 8462
rect 17411 8394 17443 8428
rect 17477 8394 17509 8428
rect 17411 8360 17509 8394
rect 17411 8326 17443 8360
rect 17477 8326 17509 8360
rect 17411 8292 17509 8326
rect 17411 8258 17443 8292
rect 17477 8258 17509 8292
rect 17411 8224 17509 8258
rect 17411 8190 17443 8224
rect 17477 8190 17509 8224
rect 17411 8156 17509 8190
rect 17411 8122 17443 8156
rect 17477 8122 17509 8156
rect 17411 8088 17509 8122
rect 17411 8054 17443 8088
rect 17477 8054 17509 8088
rect 17411 8020 17509 8054
rect 17411 7986 17443 8020
rect 17477 7986 17509 8020
rect 16435 7961 16971 7984
rect 16435 7927 16484 7961
rect 16518 7927 16582 7961
rect 16616 7927 16650 7961
rect 16684 7927 16718 7961
rect 16752 7927 16786 7961
rect 16820 7927 16884 7961
rect 16918 7927 16971 7961
rect 16435 7907 16971 7927
rect 16435 7889 16568 7907
rect 16435 7855 16484 7889
rect 16518 7855 16568 7889
rect 16435 7821 16568 7855
rect 16435 7787 16484 7821
rect 16518 7787 16568 7821
rect 16435 7753 16568 7787
rect 16435 7719 16484 7753
rect 16518 7719 16568 7753
rect 16435 7685 16568 7719
rect 16435 7651 16484 7685
rect 16518 7651 16568 7685
rect 16435 7617 16568 7651
rect 16435 7583 16484 7617
rect 16518 7583 16568 7617
rect 10745 7565 10850 7567
rect 10743 7540 11268 7565
rect 10743 7506 10783 7540
rect 10817 7506 10886 7540
rect 10920 7506 10954 7540
rect 10988 7506 11022 7540
rect 11056 7506 11090 7540
rect 11124 7506 11194 7540
rect 11228 7506 11268 7540
rect 10743 7477 11268 7506
rect 10745 7455 10850 7477
rect 10745 7421 10783 7455
rect 10817 7421 10850 7455
rect 10745 7387 10850 7421
rect 10745 7353 10783 7387
rect 10817 7353 10850 7387
rect 10745 7319 10850 7353
rect 10745 7285 10783 7319
rect 10817 7285 10850 7319
rect 10745 7251 10850 7285
rect 10745 7217 10783 7251
rect 10817 7217 10850 7251
rect 10745 7183 10850 7217
rect 10745 7149 10783 7183
rect 10817 7149 10850 7183
rect 10745 7115 10850 7149
rect 10745 7081 10783 7115
rect 10817 7081 10850 7115
rect 10745 7047 10850 7081
rect 10745 7013 10783 7047
rect 10817 7013 10850 7047
rect 10745 6979 10850 7013
rect 10745 6945 10783 6979
rect 10817 6945 10850 6979
rect 10745 6911 10850 6945
rect 10745 6877 10783 6911
rect 10817 6877 10850 6911
rect 10745 6843 10850 6877
rect 10745 6809 10783 6843
rect 10817 6809 10850 6843
rect 10745 6775 10850 6809
rect 10745 6741 10783 6775
rect 10817 6741 10850 6775
rect 10745 6707 10850 6741
rect 10745 6673 10783 6707
rect 10817 6673 10850 6707
rect 10745 6639 10850 6673
rect 10745 6605 10783 6639
rect 10817 6605 10850 6639
rect 10745 6571 10850 6605
rect 10745 6537 10783 6571
rect 10817 6537 10850 6571
rect 10745 6503 10850 6537
rect 10745 6469 10783 6503
rect 10817 6469 10850 6503
rect 10745 6435 10850 6469
rect 10745 6401 10783 6435
rect 10817 6401 10850 6435
rect 10745 6367 10850 6401
rect 10745 6333 10783 6367
rect 10817 6333 10850 6367
rect 10745 6299 10850 6333
rect 10745 6265 10783 6299
rect 10817 6265 10850 6299
rect 10745 6231 10850 6265
rect 10745 6197 10783 6231
rect 10817 6197 10850 6231
rect 10745 6163 10850 6197
rect 10745 6129 10783 6163
rect 10817 6129 10850 6163
rect 10745 6095 10850 6129
rect 10745 6061 10783 6095
rect 10817 6061 10850 6095
rect 10745 6027 10850 6061
rect 10745 5993 10783 6027
rect 10817 5993 10850 6027
rect 10745 5959 10850 5993
rect 10745 5925 10783 5959
rect 10817 5925 10850 5959
rect 10745 5891 10850 5925
rect 10745 5857 10783 5891
rect 10817 5857 10850 5891
rect 10745 5823 10850 5857
rect 10745 5789 10783 5823
rect 10817 5789 10850 5823
rect 10745 5755 10850 5789
rect 10745 5721 10783 5755
rect 10817 5721 10850 5755
rect 10745 5687 10850 5721
rect 10745 5653 10783 5687
rect 10817 5653 10850 5687
rect 10745 5632 10850 5653
rect 11158 7455 11268 7477
rect 11158 7421 11194 7455
rect 11228 7444 11268 7455
rect 16435 7549 16568 7583
rect 16435 7515 16484 7549
rect 16518 7515 16568 7549
rect 16435 7481 16568 7515
rect 16435 7447 16484 7481
rect 16518 7447 16568 7481
rect 11228 7421 11267 7444
rect 11158 7387 11267 7421
rect 11158 7353 11194 7387
rect 11228 7353 11267 7387
rect 11158 7319 11267 7353
rect 16435 7429 16568 7447
rect 16833 7889 16971 7907
rect 16833 7855 16884 7889
rect 16918 7855 16971 7889
rect 16833 7821 16971 7855
rect 17411 7955 17509 7986
rect 18179 8870 18203 8904
rect 18237 8870 18264 8904
rect 18179 8836 18264 8870
rect 18179 8802 18203 8836
rect 18237 8802 18264 8836
rect 18179 8768 18264 8802
rect 18179 8734 18203 8768
rect 18237 8734 18264 8768
rect 18179 8700 18264 8734
rect 18179 8666 18203 8700
rect 18237 8666 18264 8700
rect 18179 8632 18264 8666
rect 18179 8598 18203 8632
rect 18237 8598 18264 8632
rect 18179 8564 18264 8598
rect 18179 8530 18203 8564
rect 18237 8530 18264 8564
rect 18179 8496 18264 8530
rect 18179 8462 18203 8496
rect 18237 8462 18264 8496
rect 18179 8428 18264 8462
rect 18179 8394 18203 8428
rect 18237 8394 18264 8428
rect 18179 8360 18264 8394
rect 18179 8326 18203 8360
rect 18237 8326 18264 8360
rect 18179 8292 18264 8326
rect 18179 8258 18203 8292
rect 18237 8258 18264 8292
rect 18179 8224 18264 8258
rect 18179 8190 18203 8224
rect 18237 8190 18264 8224
rect 18179 8156 18264 8190
rect 18179 8122 18203 8156
rect 18237 8122 18264 8156
rect 18179 8088 18264 8122
rect 18179 8054 18203 8088
rect 18237 8054 18264 8088
rect 18179 8020 18264 8054
rect 18179 7986 18203 8020
rect 18237 7986 18264 8020
rect 18179 7955 18264 7986
rect 19908 9352 20444 9375
rect 19908 9318 19957 9352
rect 19991 9318 20055 9352
rect 20089 9318 20123 9352
rect 20157 9318 20191 9352
rect 20225 9318 20259 9352
rect 20293 9318 20357 9352
rect 20391 9318 20444 9352
rect 19908 9298 20444 9318
rect 19908 9280 20041 9298
rect 19908 9246 19957 9280
rect 19991 9246 20041 9280
rect 19908 9212 20041 9246
rect 19908 9178 19957 9212
rect 19991 9178 20041 9212
rect 19908 9144 20041 9178
rect 19908 9110 19957 9144
rect 19991 9110 20041 9144
rect 19908 9076 20041 9110
rect 19908 9042 19957 9076
rect 19991 9042 20041 9076
rect 19908 9008 20041 9042
rect 19908 8974 19957 9008
rect 19991 8974 20041 9008
rect 19908 8940 20041 8974
rect 19908 8906 19957 8940
rect 19991 8906 20041 8940
rect 19908 8872 20041 8906
rect 19908 8838 19957 8872
rect 19991 8838 20041 8872
rect 19908 8820 20041 8838
rect 20306 9280 20444 9298
rect 20306 9246 20357 9280
rect 20391 9246 20444 9280
rect 20306 9212 20444 9246
rect 20306 9178 20357 9212
rect 20391 9178 20444 9212
rect 20306 9144 20444 9178
rect 20306 9110 20357 9144
rect 20391 9110 20444 9144
rect 20306 9076 20444 9110
rect 20306 9042 20357 9076
rect 20391 9042 20444 9076
rect 20306 9008 20444 9042
rect 20306 8974 20357 9008
rect 20391 8974 20444 9008
rect 20306 8940 20444 8974
rect 20306 8906 20357 8940
rect 20391 8906 20444 8940
rect 20306 8872 20444 8906
rect 20306 8838 20357 8872
rect 20391 8838 20444 8872
rect 20306 8820 20444 8838
rect 19908 8800 20444 8820
rect 19908 8766 19957 8800
rect 19991 8766 20055 8800
rect 20089 8766 20123 8800
rect 20157 8766 20191 8800
rect 20225 8766 20259 8800
rect 20293 8766 20357 8800
rect 20391 8766 20444 8800
rect 19908 8742 20444 8766
rect 17411 7919 18264 7955
rect 17411 7885 17443 7919
rect 17477 7885 17519 7919
rect 17553 7885 17587 7919
rect 17621 7885 17655 7919
rect 17689 7885 17723 7919
rect 17757 7885 17791 7919
rect 17825 7885 17859 7919
rect 17893 7885 17927 7919
rect 17961 7885 17995 7919
rect 18029 7885 18063 7919
rect 18097 7885 18131 7919
rect 18165 7885 18203 7919
rect 18237 7885 18264 7919
rect 17411 7850 18264 7885
rect 19904 8021 20440 8044
rect 19904 7987 19953 8021
rect 19987 7987 20051 8021
rect 20085 7987 20119 8021
rect 20153 7987 20187 8021
rect 20221 7987 20255 8021
rect 20289 7987 20353 8021
rect 20387 7987 20440 8021
rect 19904 7967 20440 7987
rect 19904 7949 20037 7967
rect 19904 7915 19953 7949
rect 19987 7915 20037 7949
rect 19904 7881 20037 7915
rect 16833 7787 16884 7821
rect 16918 7787 16971 7821
rect 16833 7753 16971 7787
rect 16833 7719 16884 7753
rect 16918 7719 16971 7753
rect 16833 7685 16971 7719
rect 16833 7651 16884 7685
rect 16918 7651 16971 7685
rect 16833 7617 16971 7651
rect 16833 7583 16884 7617
rect 16918 7583 16971 7617
rect 16833 7549 16971 7583
rect 16833 7515 16884 7549
rect 16918 7515 16971 7549
rect 16833 7481 16971 7515
rect 16833 7447 16884 7481
rect 16918 7447 16971 7481
rect 16833 7429 16971 7447
rect 16435 7409 16971 7429
rect 19904 7847 19953 7881
rect 19987 7847 20037 7881
rect 19904 7813 20037 7847
rect 19904 7779 19953 7813
rect 19987 7779 20037 7813
rect 19904 7745 20037 7779
rect 19904 7711 19953 7745
rect 19987 7711 20037 7745
rect 19904 7677 20037 7711
rect 19904 7643 19953 7677
rect 19987 7643 20037 7677
rect 19904 7609 20037 7643
rect 19904 7575 19953 7609
rect 19987 7575 20037 7609
rect 19904 7541 20037 7575
rect 19904 7507 19953 7541
rect 19987 7507 20037 7541
rect 19904 7489 20037 7507
rect 20302 7949 20440 7967
rect 20302 7915 20353 7949
rect 20387 7915 20440 7949
rect 20302 7881 20440 7915
rect 20302 7847 20353 7881
rect 20387 7847 20440 7881
rect 20302 7813 20440 7847
rect 20302 7779 20353 7813
rect 20387 7779 20440 7813
rect 20302 7745 20440 7779
rect 20302 7711 20353 7745
rect 20387 7711 20440 7745
rect 20302 7677 20440 7711
rect 20302 7643 20353 7677
rect 20387 7643 20440 7677
rect 20302 7609 20440 7643
rect 20302 7575 20353 7609
rect 20387 7575 20440 7609
rect 20302 7541 20440 7575
rect 20302 7507 20353 7541
rect 20387 7507 20440 7541
rect 20302 7489 20440 7507
rect 19904 7469 20440 7489
rect 19904 7435 19953 7469
rect 19987 7435 20051 7469
rect 20085 7435 20119 7469
rect 20153 7435 20187 7469
rect 20221 7435 20255 7469
rect 20289 7435 20353 7469
rect 20387 7435 20440 7469
rect 19904 7411 20440 7435
rect 16435 7375 16484 7409
rect 16518 7375 16582 7409
rect 16616 7375 16650 7409
rect 16684 7375 16718 7409
rect 16752 7375 16786 7409
rect 16820 7375 16884 7409
rect 16918 7375 16971 7409
rect 16435 7351 16971 7375
rect 11158 7285 11194 7319
rect 11228 7285 11267 7319
rect 11158 7251 11267 7285
rect 11158 7217 11194 7251
rect 11228 7217 11267 7251
rect 11158 7183 11267 7217
rect 11158 7149 11194 7183
rect 11228 7149 11267 7183
rect 11158 7115 11267 7149
rect 11158 7081 11194 7115
rect 11228 7081 11267 7115
rect 11158 7047 11267 7081
rect 11158 7013 11194 7047
rect 11228 7013 11267 7047
rect 11158 6979 11267 7013
rect 11158 6945 11194 6979
rect 11228 6945 11267 6979
rect 11158 6911 11267 6945
rect 11158 6877 11194 6911
rect 11228 6877 11267 6911
rect 11158 6843 11267 6877
rect 11158 6809 11194 6843
rect 11228 6809 11267 6843
rect 11158 6775 11267 6809
rect 11158 6741 11194 6775
rect 11228 6741 11267 6775
rect 11158 6707 11267 6741
rect 11158 6673 11194 6707
rect 11228 6673 11267 6707
rect 11158 6639 11267 6673
rect 11158 6605 11194 6639
rect 11228 6605 11267 6639
rect 11158 6571 11267 6605
rect 11158 6537 11194 6571
rect 11228 6537 11267 6571
rect 11158 6503 11267 6537
rect 11158 6469 11194 6503
rect 11228 6469 11267 6503
rect 11158 6435 11267 6469
rect 11158 6401 11194 6435
rect 11228 6401 11267 6435
rect 11158 6367 11267 6401
rect 11158 6333 11194 6367
rect 11228 6333 11267 6367
rect 11158 6299 11267 6333
rect 11158 6265 11194 6299
rect 11228 6265 11267 6299
rect 11158 6231 11267 6265
rect 11158 6197 11194 6231
rect 11228 6197 11267 6231
rect 11158 6163 11267 6197
rect 19922 6779 20458 6802
rect 19922 6745 19971 6779
rect 20005 6745 20069 6779
rect 20103 6745 20137 6779
rect 20171 6745 20205 6779
rect 20239 6745 20273 6779
rect 20307 6745 20371 6779
rect 20405 6745 20458 6779
rect 19922 6725 20458 6745
rect 19922 6707 20055 6725
rect 19922 6673 19971 6707
rect 20005 6673 20055 6707
rect 19922 6639 20055 6673
rect 19922 6605 19971 6639
rect 20005 6605 20055 6639
rect 19922 6571 20055 6605
rect 19922 6537 19971 6571
rect 20005 6537 20055 6571
rect 19922 6503 20055 6537
rect 19922 6469 19971 6503
rect 20005 6469 20055 6503
rect 19922 6435 20055 6469
rect 19922 6401 19971 6435
rect 20005 6401 20055 6435
rect 19922 6367 20055 6401
rect 19922 6333 19971 6367
rect 20005 6333 20055 6367
rect 19922 6299 20055 6333
rect 19922 6265 19971 6299
rect 20005 6265 20055 6299
rect 19922 6247 20055 6265
rect 20320 6707 20458 6725
rect 20320 6673 20371 6707
rect 20405 6673 20458 6707
rect 20320 6639 20458 6673
rect 20320 6605 20371 6639
rect 20405 6605 20458 6639
rect 20320 6571 20458 6605
rect 20320 6537 20371 6571
rect 20405 6537 20458 6571
rect 20320 6503 20458 6537
rect 20320 6469 20371 6503
rect 20405 6469 20458 6503
rect 20320 6435 20458 6469
rect 20320 6401 20371 6435
rect 20405 6401 20458 6435
rect 20320 6367 20458 6401
rect 20320 6333 20371 6367
rect 20405 6333 20458 6367
rect 20320 6299 20458 6333
rect 20320 6265 20371 6299
rect 20405 6265 20458 6299
rect 20320 6247 20458 6265
rect 19922 6227 20458 6247
rect 19922 6193 19971 6227
rect 20005 6193 20069 6227
rect 20103 6193 20137 6227
rect 20171 6193 20205 6227
rect 20239 6193 20273 6227
rect 20307 6193 20371 6227
rect 20405 6193 20458 6227
rect 19922 6169 20458 6193
rect 11158 6129 11194 6163
rect 11228 6129 11267 6163
rect 11158 6095 11267 6129
rect 11158 6061 11194 6095
rect 11228 6061 11267 6095
rect 11158 6027 11267 6061
rect 11158 5993 11194 6027
rect 11228 5993 11267 6027
rect 11158 5959 11267 5993
rect 11158 5925 11194 5959
rect 11228 5925 11267 5959
rect 12995 5952 13116 5953
rect 14928 5952 15009 5953
rect 11158 5891 11267 5925
rect 11158 5857 11194 5891
rect 11228 5857 11267 5891
rect 11158 5823 11267 5857
rect 11158 5789 11194 5823
rect 11228 5789 11267 5823
rect 11158 5755 11267 5789
rect 11158 5721 11194 5755
rect 11228 5721 11267 5755
rect 11158 5687 11267 5721
rect 11158 5653 11194 5687
rect 11228 5653 11267 5687
rect 11158 5632 11267 5653
rect 10745 5611 11268 5632
rect 10745 5577 10783 5611
rect 10817 5577 10886 5611
rect 10920 5577 10954 5611
rect 10988 5577 11022 5611
rect 11056 5577 11090 5611
rect 11124 5577 11194 5611
rect 11228 5577 11268 5611
rect 10745 5556 11268 5577
rect 10746 5551 11268 5556
rect 12995 5913 15009 5952
rect 12995 5879 13020 5913
rect 13054 5879 13105 5913
rect 13139 5879 13173 5913
rect 13207 5879 13241 5913
rect 13275 5879 13309 5913
rect 13343 5879 13377 5913
rect 13411 5879 13445 5913
rect 13479 5879 13513 5913
rect 13547 5879 13581 5913
rect 13615 5879 13649 5913
rect 13683 5879 13717 5913
rect 13751 5879 13785 5913
rect 13819 5879 13853 5913
rect 13887 5879 13921 5913
rect 13955 5879 13989 5913
rect 14023 5879 14057 5913
rect 14091 5879 14125 5913
rect 14159 5879 14193 5913
rect 14227 5879 14261 5913
rect 14295 5879 14329 5913
rect 14363 5879 14397 5913
rect 14431 5879 14465 5913
rect 14499 5879 14533 5913
rect 14567 5879 14601 5913
rect 14635 5879 14669 5913
rect 14703 5879 14737 5913
rect 14771 5879 14805 5913
rect 14839 5879 14873 5913
rect 14907 5879 14949 5913
rect 14983 5879 15009 5913
rect 12995 5843 15009 5879
rect 12995 5809 13083 5843
rect 12995 5775 13020 5809
rect 13054 5775 13083 5809
rect 12995 5741 13083 5775
rect 12995 5707 13020 5741
rect 13054 5707 13083 5741
rect 12995 5673 13083 5707
rect 12995 5639 13020 5673
rect 13054 5639 13083 5673
rect 12995 5605 13083 5639
rect 12995 5571 13020 5605
rect 13054 5571 13083 5605
rect 12995 5535 13083 5571
rect 14928 5809 15009 5843
rect 14928 5775 14949 5809
rect 14983 5775 15009 5809
rect 14928 5741 15009 5775
rect 14928 5707 14949 5741
rect 14983 5707 15009 5741
rect 14928 5673 15009 5707
rect 14928 5639 14949 5673
rect 14983 5639 15009 5673
rect 14928 5605 15009 5639
rect 14928 5571 14949 5605
rect 14983 5571 15009 5605
rect 14928 5535 15009 5571
rect 12993 5502 15009 5535
rect 12993 5500 13105 5502
rect 12993 5466 13020 5500
rect 13054 5468 13105 5500
rect 13139 5468 13173 5502
rect 13207 5468 13241 5502
rect 13275 5468 13309 5502
rect 13343 5468 13377 5502
rect 13411 5468 13445 5502
rect 13479 5468 13513 5502
rect 13547 5468 13581 5502
rect 13615 5468 13649 5502
rect 13683 5468 13717 5502
rect 13751 5468 13785 5502
rect 13819 5468 13853 5502
rect 13887 5468 13921 5502
rect 13955 5468 13989 5502
rect 14023 5468 14057 5502
rect 14091 5468 14125 5502
rect 14159 5468 14193 5502
rect 14227 5468 14261 5502
rect 14295 5468 14329 5502
rect 14363 5468 14397 5502
rect 14431 5468 14465 5502
rect 14499 5468 14533 5502
rect 14567 5468 14601 5502
rect 14635 5468 14669 5502
rect 14703 5468 14737 5502
rect 14771 5468 14805 5502
rect 14839 5468 14873 5502
rect 14907 5468 14949 5502
rect 14983 5468 15009 5502
rect 13054 5466 15009 5468
rect 12993 5431 15009 5466
rect 12993 5430 15004 5431
rect 12995 5428 13083 5430
rect 5440 2572 5546 2606
rect 5580 2572 5614 2606
rect 5648 2572 5682 2606
rect 5716 2572 5750 2606
rect 5784 2572 5818 2606
rect 5852 2572 5886 2606
rect 5920 2572 5954 2606
rect 5988 2572 6022 2606
rect 6056 2572 6090 2606
rect 6124 2572 6158 2606
rect 6192 2572 6226 2606
rect 6260 2572 6294 2606
rect 6328 2572 6362 2606
rect 6396 2572 6430 2606
rect 6464 2572 6498 2606
rect 6532 2572 6566 2606
rect 6600 2572 6634 2606
rect 6668 2572 6702 2606
rect 6736 2572 6770 2606
rect 6804 2572 6838 2606
rect 6872 2572 6906 2606
rect 6940 2572 6974 2606
rect 7008 2572 7042 2606
rect 7076 2572 7110 2606
rect 7144 2572 7178 2606
rect 7212 2572 7246 2606
rect 7280 2572 7314 2606
rect 7348 2572 7382 2606
rect 7416 2572 7450 2606
rect 7484 2572 7518 2606
rect 7552 2572 7586 2606
rect 7620 2572 7654 2606
rect 7688 2572 7722 2606
rect 7756 2572 7790 2606
rect 7824 2572 7858 2606
rect 7892 2572 7926 2606
rect 7960 2572 7994 2606
rect 8028 2572 8062 2606
rect 8096 2572 8130 2606
rect 8164 2572 8198 2606
rect 8232 2572 8266 2606
rect 8300 2572 8334 2606
rect 8368 2572 8402 2606
rect 8436 2572 8470 2606
rect 8504 2572 8538 2606
rect 8572 2572 8606 2606
rect 8640 2572 8674 2606
rect 8708 2572 8742 2606
rect 8776 2572 8810 2606
rect 8844 2572 8878 2606
rect 8912 2572 8946 2606
rect 8980 2572 9014 2606
rect 9048 2572 9082 2606
rect 9116 2572 9150 2606
rect 9184 2572 9218 2606
rect 9252 2572 9286 2606
rect 9320 2572 9354 2606
rect 9388 2572 9422 2606
rect 9456 2572 9490 2606
rect 9524 2572 9558 2606
rect 9592 2572 9626 2606
rect 9660 2572 9694 2606
rect 9728 2572 9762 2606
rect 9796 2572 9830 2606
rect 9864 2572 9898 2606
rect 9932 2572 9966 2606
rect 10000 2572 10034 2606
rect 10068 2572 10102 2606
rect 10136 2572 10170 2606
rect 10204 2572 10238 2606
rect 10272 2572 10306 2606
rect 10340 2572 10374 2606
rect 10408 2572 10442 2606
rect 10476 2572 10510 2606
rect 10544 2572 10578 2606
rect 10612 2572 10646 2606
rect 10680 2572 10714 2606
rect 10748 2572 10782 2606
rect 10816 2572 10850 2606
rect 10884 2572 10918 2606
rect 10952 2572 10986 2606
rect 11020 2572 11054 2606
rect 11088 2572 11122 2606
rect 11156 2572 11190 2606
rect 11224 2572 11258 2606
rect 11292 2572 11326 2606
rect 11360 2572 11394 2606
rect 11428 2572 11462 2606
rect 11496 2572 11530 2606
rect 11564 2572 11598 2606
rect 11632 2572 11666 2606
rect 11700 2572 11734 2606
rect 11768 2572 11802 2606
rect 11836 2572 11870 2606
rect 11904 2572 11938 2606
rect 11972 2572 12006 2606
rect 12040 2572 12074 2606
rect 12108 2572 12142 2606
rect 12176 2572 12210 2606
rect 12244 2572 12278 2606
rect 12312 2572 12346 2606
rect 12380 2572 12414 2606
rect 12448 2572 12482 2606
rect 12516 2572 12550 2606
rect 12584 2572 12618 2606
rect 12652 2572 12686 2606
rect 12720 2572 12754 2606
rect 12788 2572 12822 2606
rect 12856 2572 12890 2606
rect 12924 2572 12958 2606
rect 12992 2572 13026 2606
rect 13060 2572 13094 2606
rect 13128 2572 13162 2606
rect 13196 2572 13230 2606
rect 13264 2572 13298 2606
rect 13332 2572 13366 2606
rect 13400 2572 13434 2606
rect 13468 2572 13502 2606
rect 13536 2572 13570 2606
rect 13604 2572 13638 2606
rect 13672 2572 13706 2606
rect 13740 2572 13774 2606
rect 13808 2572 13842 2606
rect 13876 2572 13910 2606
rect 13944 2572 13978 2606
rect 14012 2572 14046 2606
rect 14080 2572 14114 2606
rect 14148 2572 14182 2606
rect 14216 2572 14250 2606
rect 14284 2572 14318 2606
rect 14352 2572 14386 2606
rect 14420 2572 14454 2606
rect 14488 2572 14522 2606
rect 14556 2572 14590 2606
rect 14624 2572 14658 2606
rect 14692 2572 14726 2606
rect 14760 2572 14794 2606
rect 14828 2572 14862 2606
rect 14896 2572 14930 2606
rect 14964 2572 14998 2606
rect 15032 2572 15066 2606
rect 15100 2572 15134 2606
rect 15168 2572 15202 2606
rect 15236 2572 15270 2606
rect 15304 2572 15338 2606
rect 15372 2572 15406 2606
rect 15440 2572 15474 2606
rect 15508 2572 15542 2606
rect 15576 2572 15610 2606
rect 15644 2572 15678 2606
rect 15712 2572 15746 2606
rect 15780 2572 15814 2606
rect 15848 2572 15882 2606
rect 15916 2572 15950 2606
rect 15984 2572 16018 2606
rect 16052 2572 16086 2606
rect 16120 2572 16154 2606
rect 16188 2572 16222 2606
rect 16256 2572 16290 2606
rect 16324 2572 16358 2606
rect 16392 2572 16426 2606
rect 16460 2572 16494 2606
rect 16528 2572 16562 2606
rect 16596 2572 16630 2606
rect 16664 2572 16698 2606
rect 16732 2572 16766 2606
rect 16800 2572 16834 2606
rect 16868 2572 16902 2606
rect 16936 2572 16970 2606
rect 17004 2572 17038 2606
rect 17072 2572 17106 2606
rect 17140 2572 17174 2606
rect 17208 2572 17242 2606
rect 17276 2572 17310 2606
rect 17344 2572 17378 2606
rect 17412 2572 17446 2606
rect 17480 2572 17514 2606
rect 17548 2572 17582 2606
rect 17616 2572 17650 2606
rect 17684 2572 17718 2606
rect 17752 2572 17786 2606
rect 17820 2572 17854 2606
rect 17888 2572 17922 2606
rect 17956 2572 17990 2606
rect 18024 2572 18058 2606
rect 18092 2572 18126 2606
rect 18160 2572 18194 2606
rect 18228 2572 18262 2606
rect 18296 2572 18330 2606
rect 18364 2572 18398 2606
rect 18432 2572 18466 2606
rect 18500 2572 18534 2606
rect 18568 2572 18602 2606
rect 18636 2572 18670 2606
rect 18704 2572 18738 2606
rect 18772 2572 18806 2606
rect 18840 2572 18874 2606
rect 18908 2572 18942 2606
rect 18976 2572 19010 2606
rect 19044 2572 19078 2606
rect 19112 2572 19146 2606
rect 19180 2572 19214 2606
rect 19248 2572 19282 2606
rect 19316 2572 19350 2606
rect 19384 2572 19418 2606
rect 19452 2572 19486 2606
rect 19520 2572 19554 2606
rect 19588 2572 19622 2606
rect 19656 2572 19690 2606
rect 19724 2572 19758 2606
rect 19792 2572 19826 2606
rect 19860 2572 19894 2606
rect 19928 2572 19962 2606
rect 19996 2572 20030 2606
rect 20064 2572 20098 2606
rect 20132 2572 20166 2606
rect 20200 2572 20234 2606
rect 20268 2572 20302 2606
rect 20336 2572 20370 2606
rect 20404 2572 20438 2606
rect 20472 2572 20506 2606
rect 20540 2572 20574 2606
rect 20608 2572 20642 2606
rect 20676 2572 20710 2606
rect 20744 2572 20778 2606
rect 20812 2572 20846 2606
rect 20880 2572 20914 2606
rect 20948 2572 20982 2606
rect 21016 2572 21050 2606
rect 21084 2572 21118 2606
rect 21152 2572 21186 2606
rect 21220 2572 21254 2606
rect 21288 2572 21322 2606
rect 21356 2572 21390 2606
rect 21424 2572 21458 2606
rect 21492 2572 21526 2606
rect 21560 2572 21594 2606
rect 21628 2572 21662 2606
rect 21696 2572 21730 2606
rect 21764 2572 21798 2606
rect 21832 2572 21866 2606
rect 21900 2572 21934 2606
rect 21968 2572 22002 2606
rect 22036 2572 22070 2606
rect 22104 2572 22138 2606
rect 22172 2572 22206 2606
rect 22240 2572 22274 2606
rect 22308 2572 22342 2606
rect 22376 2572 22410 2606
rect 22444 2572 22478 2606
rect 22512 2572 22546 2606
rect 22580 2572 22614 2606
rect 22648 2572 22682 2606
rect 22716 2572 22750 2606
rect 22784 2572 22818 2606
rect 22852 2572 22886 2606
rect 22920 2572 22954 2606
rect 22988 2572 23022 2606
rect 23056 2572 23090 2606
rect 23124 2572 23158 2606
rect 23192 2572 23226 2606
rect 23260 2572 23294 2606
rect 23328 2572 23362 2606
rect 23396 2572 23430 2606
rect 23464 2572 23498 2606
rect 23532 2572 23566 2606
rect 23600 2572 23634 2606
rect 23668 2572 23702 2606
rect 23736 2572 23770 2606
rect 23804 2572 23838 2606
rect 23872 2572 23906 2606
rect 23940 2572 23974 2606
rect 24008 2572 24042 2606
rect 24076 2572 24110 2606
rect 24144 2572 24178 2606
rect 24212 2572 24246 2606
rect 24280 2572 24314 2606
rect 24348 2572 24382 2606
rect 24416 2572 24450 2606
rect 24484 2572 24518 2606
rect 24552 2572 24586 2606
rect 24620 2572 24654 2606
rect 24688 2572 24722 2606
rect 24756 2572 24790 2606
rect 24824 2572 24858 2606
rect 24892 2572 24926 2606
rect 24960 2572 24994 2606
rect 25028 2572 25062 2606
rect 25096 2572 25130 2606
rect 25164 2572 25198 2606
rect 25232 2572 25266 2606
rect 25300 2572 25334 2606
rect 25368 2572 25402 2606
rect 25436 2572 25470 2606
rect 25504 2572 25538 2606
rect 25572 2572 25606 2606
rect 25640 2572 25674 2606
rect 25708 2572 25742 2606
rect 25776 2572 25810 2606
rect 25844 2572 25878 2606
rect 25912 2572 25946 2606
rect 25980 2572 26014 2606
rect 26048 2572 26082 2606
rect 26116 2572 26150 2606
rect 26184 2572 26218 2606
rect 26252 2572 26286 2606
rect 26320 2572 26354 2606
rect 26388 2572 26422 2606
rect 26456 2572 26490 2606
rect 26524 2572 26558 2606
rect 26592 2572 26626 2606
rect 26660 2572 26694 2606
rect 26728 2572 26762 2606
rect 26796 2572 26830 2606
rect 26864 2572 26898 2606
rect 26932 2572 26966 2606
rect 27000 2572 27034 2606
rect 27068 2572 27102 2606
rect 27136 2572 27170 2606
rect 27204 2572 27238 2606
rect 27272 2572 27306 2606
rect 27340 2572 27374 2606
rect 27408 2572 27442 2606
rect 27476 2572 27510 2606
rect 27544 2572 27578 2606
rect 27612 2572 27646 2606
rect 27680 2572 27714 2606
rect 27748 2572 27782 2606
rect 27816 2572 27850 2606
rect 27884 2572 27918 2606
rect 27952 2572 27986 2606
rect 28020 2572 28054 2606
rect 28088 2572 28122 2606
rect 28156 2572 28190 2606
rect 28224 2572 28258 2606
rect 28292 2572 28326 2606
rect 28360 2572 28394 2606
rect 28428 2572 28462 2606
rect 28496 2572 28530 2606
rect 28564 2572 28598 2606
rect 28632 2572 28666 2606
rect 28700 2572 28734 2606
rect 28768 2572 28802 2606
rect 28836 2572 28870 2606
rect 28904 2572 28938 2606
rect 28972 2572 29006 2606
rect 29040 2572 29074 2606
rect 29108 2572 29142 2606
rect 29176 2572 29210 2606
rect 29244 2572 29278 2606
rect 29312 2572 29346 2606
rect 29380 2572 29414 2606
rect 29448 2572 29482 2606
rect 29516 2572 29550 2606
rect 29584 2572 29618 2606
rect 29652 2572 29686 2606
rect 29720 2572 29754 2606
rect 29788 2572 29822 2606
rect 29856 2572 29890 2606
rect 29924 2572 29958 2606
rect 29992 2572 30026 2606
rect 30060 2572 30094 2606
rect 30128 2572 30162 2606
rect 30196 2572 30230 2606
rect 30264 2572 30298 2606
rect 30332 2572 30366 2606
rect 30400 2572 30434 2606
rect 30468 2572 30502 2606
rect 30536 2572 30570 2606
rect 30604 2572 30638 2606
rect 30672 2572 30706 2606
rect 30740 2572 30774 2606
rect 30808 2572 30842 2606
rect 30876 2572 30910 2606
rect 30944 2572 30978 2606
rect 31012 2572 31046 2606
rect 31080 2572 31114 2606
rect 31148 2572 31182 2606
rect 31216 2572 31250 2606
rect 31284 2572 31318 2606
rect 31352 2572 31386 2606
rect 31420 2572 31454 2606
rect 31488 2572 31522 2606
rect 31556 2572 31590 2606
rect 31624 2572 31658 2606
rect 31692 2572 31726 2606
rect 31760 2572 31794 2606
rect 31828 2572 31862 2606
rect 31896 2572 31930 2606
rect 31964 2572 31998 2606
rect 32032 2572 32066 2606
rect 32100 2572 32134 2606
rect 32168 2572 32202 2606
rect 32236 2572 32270 2606
rect 32304 2572 32338 2606
rect 32372 2572 32406 2606
rect 32440 2572 32474 2606
rect 32508 2572 32542 2606
rect 32576 2572 32610 2606
rect 32644 2572 32678 2606
rect 32712 2572 32746 2606
rect 32780 2572 32814 2606
rect 32848 2572 32882 2606
rect 32916 2572 32950 2606
rect 32984 2572 33018 2606
rect 33052 2572 33086 2606
rect 33120 2572 33154 2606
rect 33188 2572 33222 2606
rect 33256 2572 33290 2606
rect 33324 2572 33358 2606
rect 33392 2572 33426 2606
rect 33460 2572 33494 2606
rect 33528 2572 33562 2606
rect 33596 2572 33630 2606
rect 33664 2572 33698 2606
rect 33732 2572 33766 2606
rect 33800 2572 33834 2606
rect 33868 2572 33902 2606
rect 33936 2572 33970 2606
rect 34004 2572 34038 2606
rect 34072 2572 34106 2606
rect 34140 2572 34174 2606
rect 34208 2572 34242 2606
rect 34276 2572 34310 2606
rect 34344 2572 34378 2606
rect 34412 2572 34446 2606
rect 34480 2572 34514 2606
rect 34548 2572 34582 2606
rect 34616 2572 34650 2606
rect 34684 2572 34718 2606
rect 34752 2572 34786 2606
rect 34820 2572 34854 2606
rect 34888 2572 34922 2606
rect 34956 2572 34990 2606
rect 35024 2572 35058 2606
rect 35092 2572 35126 2606
rect 35160 2572 35194 2606
rect 35228 2572 35262 2606
rect 35296 2572 35330 2606
rect 35364 2572 35398 2606
rect 35432 2572 35466 2606
rect 35500 2572 35534 2606
rect 35568 2572 35602 2606
rect 35636 2572 35670 2606
rect 35704 2572 35738 2606
rect 35772 2572 35806 2606
rect 35840 2572 35874 2606
rect 35908 2572 35942 2606
rect 35976 2572 36010 2606
rect 36044 2572 36078 2606
rect 36112 2572 36146 2606
rect 36180 2572 36214 2606
rect 36248 2572 36282 2606
rect 36316 2572 36350 2606
rect 36384 2572 36418 2606
rect 36452 2572 36486 2606
rect 36520 2572 36554 2606
rect 36588 2572 36622 2606
rect 36656 2572 36690 2606
rect 36724 2572 36758 2606
rect 36792 2572 36826 2606
rect 36860 2572 36894 2606
rect 36928 2572 36962 2606
rect 36996 2572 37030 2606
rect 37064 2572 37098 2606
rect 37132 2572 37166 2606
rect 37200 2572 37234 2606
rect 37268 2572 37302 2606
rect 37336 2572 37370 2606
rect 37404 2572 37438 2606
rect 37472 2572 37506 2606
rect 37540 2572 37574 2606
rect 37608 2572 37642 2606
rect 37676 2572 37710 2606
rect 37744 2572 37778 2606
rect 37812 2572 37846 2606
rect 37880 2572 37914 2606
rect 37948 2572 37982 2606
rect 38016 2572 38050 2606
rect 38084 2572 38118 2606
rect 38152 2572 38186 2606
rect 38220 2572 38254 2606
rect 38288 2572 38322 2606
rect 38356 2572 38390 2606
rect 38424 2572 38458 2606
rect 38492 2572 38526 2606
rect 38560 2572 38594 2606
rect 38628 2572 38662 2606
rect 38696 2572 38730 2606
rect 38764 2572 38798 2606
rect 38832 2572 38866 2606
rect 38900 2572 38934 2606
rect 38968 2572 39002 2606
rect 39036 2572 39070 2606
rect 39104 2572 39138 2606
rect 39172 2572 39206 2606
rect 39240 2572 39274 2606
rect 39308 2572 39342 2606
rect 39376 2572 39410 2606
rect 39444 2572 39478 2606
rect 39512 2572 39546 2606
rect 39580 2572 39614 2606
rect 39648 2572 39682 2606
rect 39716 2572 39750 2606
rect 39784 2572 39818 2606
rect 39852 2572 39886 2606
rect 39920 2572 39954 2606
rect 39988 2572 40022 2606
rect 40056 2572 40090 2606
rect 40124 2572 40158 2606
rect 40192 2572 40226 2606
rect 40260 2572 40294 2606
rect 40328 2572 40362 2606
rect 40396 2572 40430 2606
rect 40464 2572 40498 2606
rect 40532 2572 40566 2606
rect 40600 2572 40634 2606
rect 40668 2572 40702 2606
rect 40736 2572 40770 2606
rect 40804 2572 40838 2606
rect 40872 2572 40906 2606
rect 40940 2572 40974 2606
rect 41008 2572 41042 2606
rect 41076 2572 41110 2606
rect 41144 2572 41178 2606
rect 41212 2572 41246 2606
rect 41280 2572 41314 2606
rect 41348 2572 41382 2606
rect 41416 2572 41450 2606
rect 41484 2572 41518 2606
rect 41552 2572 41586 2606
rect 41620 2572 41654 2606
rect 41688 2572 41722 2606
rect 41756 2572 41790 2606
rect 41824 2572 41896 2606
rect 5440 2484 5474 2572
rect 5440 2416 5474 2450
rect 5440 2348 5474 2382
rect 5440 2280 5474 2314
rect 5440 2212 5474 2246
rect 5440 2144 5474 2178
rect 5440 2076 5474 2110
rect 5440 2008 5474 2042
rect 5440 1940 5474 1974
rect 5440 1872 5474 1906
rect 5440 1804 5474 1838
rect 5440 1736 5474 1770
rect 5440 1668 5474 1702
rect 5440 1600 5474 1634
rect 5440 1532 5474 1566
rect 5440 1464 5474 1498
rect 5440 1396 5474 1430
rect 5440 1328 5474 1362
rect 5440 1260 5474 1294
rect 5440 1192 5474 1226
rect 5440 1124 5474 1158
rect 5440 1056 5474 1090
rect 5440 988 5474 1022
rect 5440 920 5474 954
rect 5440 852 5474 886
rect 5440 784 5474 818
rect 5440 716 5474 750
rect 5440 648 5474 682
rect 5440 580 5474 614
rect 5440 458 5474 546
rect 5440 424 5546 458
rect 5580 424 5614 458
rect 5648 424 5682 458
rect 5716 424 5750 458
rect 5784 424 5818 458
rect 5852 424 5886 458
rect 5920 424 5954 458
rect 5988 424 6022 458
rect 6056 424 6090 458
rect 6124 424 6158 458
rect 6192 424 6226 458
rect 6260 424 6294 458
rect 6328 424 6362 458
rect 6396 424 6430 458
rect 6464 424 6498 458
rect 6532 424 6566 458
rect 6600 424 6634 458
rect 6668 424 6702 458
rect 6736 424 6770 458
rect 6804 424 6838 458
rect 6872 424 6906 458
rect 6940 424 6974 458
rect 7008 424 7042 458
rect 7076 424 7110 458
rect 7144 424 7178 458
rect 7212 424 7246 458
rect 7280 424 7314 458
rect 7348 424 7382 458
rect 7416 424 7450 458
rect 7484 424 7518 458
rect 7552 424 7586 458
rect 7620 424 7654 458
rect 7688 424 7722 458
rect 7756 424 7790 458
rect 7824 424 7858 458
rect 7892 424 7926 458
rect 7960 424 7994 458
rect 8028 424 8062 458
rect 8096 424 8130 458
rect 8164 424 8198 458
rect 8232 424 8266 458
rect 8300 424 8334 458
rect 8368 424 8402 458
rect 8436 424 8470 458
rect 8504 424 8538 458
rect 8572 424 8606 458
rect 8640 424 8674 458
rect 8708 424 8742 458
rect 8776 424 8810 458
rect 8844 424 8878 458
rect 8912 424 8946 458
rect 8980 424 9014 458
rect 9048 424 9082 458
rect 9116 424 9150 458
rect 9184 424 9218 458
rect 9252 424 9286 458
rect 9320 424 9354 458
rect 9388 424 9422 458
rect 9456 424 9490 458
rect 9524 424 9558 458
rect 9592 424 9626 458
rect 9660 424 9694 458
rect 9728 424 9762 458
rect 9796 424 9830 458
rect 9864 424 9898 458
rect 9932 424 9966 458
rect 10000 424 10034 458
rect 10068 424 10102 458
rect 10136 424 10170 458
rect 10204 424 10238 458
rect 10272 424 10306 458
rect 10340 424 10374 458
rect 10408 424 10442 458
rect 10476 424 10510 458
rect 10544 424 10578 458
rect 10612 424 10646 458
rect 10680 424 10714 458
rect 10748 424 10782 458
rect 10816 424 10850 458
rect 10884 424 10918 458
rect 10952 424 10986 458
rect 11020 424 11054 458
rect 11088 424 11122 458
rect 11156 424 11190 458
rect 11224 424 11258 458
rect 11292 424 11326 458
rect 11360 424 11394 458
rect 11428 424 11462 458
rect 11496 424 11530 458
rect 11564 424 11598 458
rect 11632 424 11666 458
rect 11700 424 11734 458
rect 11768 424 11802 458
rect 11836 424 11870 458
rect 11904 424 11938 458
rect 11972 424 12006 458
rect 12040 424 12074 458
rect 12108 424 12142 458
rect 12176 424 12210 458
rect 12244 424 12278 458
rect 12312 424 12346 458
rect 12380 424 12414 458
rect 12448 424 12482 458
rect 12516 424 12550 458
rect 12584 424 12618 458
rect 12652 424 12686 458
rect 12720 424 12754 458
rect 12788 424 12822 458
rect 12856 424 12890 458
rect 12924 424 12958 458
rect 12992 424 13026 458
rect 13060 424 13094 458
rect 13128 424 13162 458
rect 13196 424 13230 458
rect 13264 424 13298 458
rect 13332 424 13366 458
rect 13400 424 13434 458
rect 13468 424 13502 458
rect 13536 424 13570 458
rect 13604 424 13638 458
rect 13672 424 13706 458
rect 13740 424 13774 458
rect 13808 424 13842 458
rect 13876 424 13910 458
rect 13944 424 13978 458
rect 14012 424 14046 458
rect 14080 424 14114 458
rect 14148 424 14182 458
rect 14216 424 14250 458
rect 14284 424 14318 458
rect 14352 424 14386 458
rect 14420 424 14454 458
rect 14488 424 14522 458
rect 14556 424 14590 458
rect 14624 424 14658 458
rect 14692 424 14726 458
rect 14760 424 14794 458
rect 14828 424 14862 458
rect 14896 424 14930 458
rect 14964 424 14998 458
rect 15032 424 15066 458
rect 15100 424 15134 458
rect 15168 424 15202 458
rect 15236 424 15270 458
rect 15304 424 15338 458
rect 15372 424 15406 458
rect 15440 424 15474 458
rect 15508 424 15542 458
rect 15576 424 15610 458
rect 15644 424 15678 458
rect 15712 424 15746 458
rect 15780 424 15814 458
rect 15848 424 15882 458
rect 15916 424 15950 458
rect 15984 424 16018 458
rect 16052 424 16086 458
rect 16120 424 16154 458
rect 16188 424 16222 458
rect 16256 424 16290 458
rect 16324 424 16358 458
rect 16392 424 16426 458
rect 16460 424 16494 458
rect 16528 424 16562 458
rect 16596 424 16630 458
rect 16664 424 16698 458
rect 16732 424 16766 458
rect 16800 424 16834 458
rect 16868 424 16902 458
rect 16936 424 16970 458
rect 17004 424 17038 458
rect 17072 424 17106 458
rect 17140 424 17174 458
rect 17208 424 17242 458
rect 17276 424 17310 458
rect 17344 424 17378 458
rect 17412 424 17446 458
rect 17480 424 17514 458
rect 17548 424 17582 458
rect 17616 424 17650 458
rect 17684 424 17718 458
rect 17752 424 17786 458
rect 17820 424 17854 458
rect 17888 424 17922 458
rect 17956 424 17990 458
rect 18024 424 18058 458
rect 18092 424 18126 458
rect 18160 424 18194 458
rect 18228 424 18262 458
rect 18296 424 18330 458
rect 18364 424 18398 458
rect 18432 424 18466 458
rect 18500 424 18534 458
rect 18568 424 18602 458
rect 18636 424 18670 458
rect 18704 424 18738 458
rect 18772 424 18806 458
rect 18840 424 18874 458
rect 18908 424 18942 458
rect 18976 424 19010 458
rect 19044 424 19078 458
rect 19112 424 19146 458
rect 19180 424 19214 458
rect 19248 424 19282 458
rect 19316 424 19350 458
rect 19384 424 19418 458
rect 19452 424 19486 458
rect 19520 424 19554 458
rect 19588 424 19622 458
rect 19656 424 19690 458
rect 19724 424 19758 458
rect 19792 424 19826 458
rect 19860 424 19894 458
rect 19928 424 19962 458
rect 19996 424 20030 458
rect 20064 424 20098 458
rect 20132 424 20166 458
rect 20200 424 20234 458
rect 20268 424 20302 458
rect 20336 424 20370 458
rect 20404 424 20438 458
rect 20472 424 20506 458
rect 20540 424 20574 458
rect 20608 424 20642 458
rect 20676 424 20710 458
rect 20744 424 20778 458
rect 20812 424 20846 458
rect 20880 424 20914 458
rect 20948 424 20982 458
rect 21016 424 21050 458
rect 21084 424 21118 458
rect 21152 424 21186 458
rect 21220 424 21254 458
rect 21288 424 21322 458
rect 21356 424 21390 458
rect 21424 424 21458 458
rect 21492 424 21526 458
rect 21560 424 21594 458
rect 21628 424 21662 458
rect 21696 424 21730 458
rect 21764 424 21798 458
rect 21832 424 21866 458
rect 21900 424 21934 458
rect 21968 424 22002 458
rect 22036 424 22070 458
rect 22104 424 22138 458
rect 22172 424 22206 458
rect 22240 424 22274 458
rect 22308 424 22342 458
rect 22376 424 22410 458
rect 22444 424 22478 458
rect 22512 424 22546 458
rect 22580 424 22614 458
rect 22648 424 22682 458
rect 22716 424 22750 458
rect 22784 424 22818 458
rect 22852 424 22886 458
rect 22920 424 22954 458
rect 22988 424 23022 458
rect 23056 424 23090 458
rect 23124 424 23158 458
rect 23192 424 23226 458
rect 23260 424 23294 458
rect 23328 424 23362 458
rect 23396 424 23430 458
rect 23464 424 23498 458
rect 23532 424 23566 458
rect 23600 424 23634 458
rect 23668 424 23702 458
rect 23736 424 23770 458
rect 23804 424 23838 458
rect 23872 424 23906 458
rect 23940 424 23974 458
rect 24008 424 24042 458
rect 24076 424 24110 458
rect 24144 424 24178 458
rect 24212 424 24246 458
rect 24280 424 24314 458
rect 24348 424 24382 458
rect 24416 424 24450 458
rect 24484 424 24518 458
rect 24552 424 24586 458
rect 24620 424 24654 458
rect 24688 424 24722 458
rect 24756 424 24790 458
rect 24824 424 24858 458
rect 24892 424 24926 458
rect 24960 424 24994 458
rect 25028 424 25062 458
rect 25096 424 25130 458
rect 25164 424 25198 458
rect 25232 424 25266 458
rect 25300 424 25334 458
rect 25368 424 25402 458
rect 25436 424 25470 458
rect 25504 424 25538 458
rect 25572 424 25606 458
rect 25640 424 25674 458
rect 25708 424 25742 458
rect 25776 424 25810 458
rect 25844 424 25878 458
rect 25912 424 25946 458
rect 25980 424 26014 458
rect 26048 424 26082 458
rect 26116 424 26150 458
rect 26184 424 26218 458
rect 26252 424 26286 458
rect 26320 424 26354 458
rect 26388 424 26422 458
rect 26456 424 26490 458
rect 26524 424 26558 458
rect 26592 424 26626 458
rect 26660 424 26694 458
rect 26728 424 26762 458
rect 26796 424 26830 458
rect 26864 424 26898 458
rect 26932 424 26966 458
rect 27000 424 27034 458
rect 27068 424 27102 458
rect 27136 424 27170 458
rect 27204 424 27238 458
rect 27272 424 27306 458
rect 27340 424 27374 458
rect 27408 424 27442 458
rect 27476 424 27510 458
rect 27544 424 27578 458
rect 27612 424 27646 458
rect 27680 424 27714 458
rect 27748 424 27782 458
rect 27816 424 27850 458
rect 27884 424 27918 458
rect 27952 424 27986 458
rect 28020 424 28054 458
rect 28088 424 28122 458
rect 28156 424 28190 458
rect 28224 424 28258 458
rect 28292 424 28326 458
rect 28360 424 28394 458
rect 28428 424 28462 458
rect 28496 424 28530 458
rect 28564 424 28598 458
rect 28632 424 28666 458
rect 28700 424 28734 458
rect 28768 424 28802 458
rect 28836 424 28870 458
rect 28904 424 28938 458
rect 28972 424 29006 458
rect 29040 424 29074 458
rect 29108 424 29142 458
rect 29176 424 29210 458
rect 29244 424 29278 458
rect 29312 424 29346 458
rect 29380 424 29414 458
rect 29448 424 29482 458
rect 29516 424 29550 458
rect 29584 424 29618 458
rect 29652 424 29686 458
rect 29720 424 29754 458
rect 29788 424 29822 458
rect 29856 424 29890 458
rect 29924 424 29958 458
rect 29992 424 30026 458
rect 30060 424 30094 458
rect 30128 424 30162 458
rect 30196 424 30230 458
rect 30264 424 30298 458
rect 30332 424 30366 458
rect 30400 424 30434 458
rect 30468 424 30502 458
rect 30536 424 30570 458
rect 30604 424 30638 458
rect 30672 424 30706 458
rect 30740 424 30774 458
rect 30808 424 30842 458
rect 30876 424 30910 458
rect 30944 424 30978 458
rect 31012 424 31046 458
rect 31080 424 31114 458
rect 31148 424 31182 458
rect 31216 424 31250 458
rect 31284 424 31318 458
rect 31352 424 31386 458
rect 31420 424 31454 458
rect 31488 424 31522 458
rect 31556 424 31590 458
rect 31624 424 31658 458
rect 31692 424 31726 458
rect 31760 424 31794 458
rect 31828 424 31862 458
rect 31896 424 31930 458
rect 31964 424 31998 458
rect 32032 424 32066 458
rect 32100 424 32134 458
rect 32168 424 32202 458
rect 32236 424 32270 458
rect 32304 424 32338 458
rect 32372 424 32406 458
rect 32440 424 32474 458
rect 32508 424 32542 458
rect 32576 424 32610 458
rect 32644 424 32678 458
rect 32712 424 32746 458
rect 32780 424 32814 458
rect 32848 424 32882 458
rect 32916 424 32950 458
rect 32984 424 33018 458
rect 33052 424 33086 458
rect 33120 424 33154 458
rect 33188 424 33222 458
rect 33256 424 33290 458
rect 33324 424 33358 458
rect 33392 424 33426 458
rect 33460 424 33494 458
rect 33528 424 33562 458
rect 33596 424 33630 458
rect 33664 424 33698 458
rect 33732 424 33766 458
rect 33800 424 33834 458
rect 33868 424 33902 458
rect 33936 424 33970 458
rect 34004 424 34038 458
rect 34072 424 34106 458
rect 34140 424 34174 458
rect 34208 424 34242 458
rect 34276 424 34310 458
rect 34344 424 34378 458
rect 34412 424 34446 458
rect 34480 424 34514 458
rect 34548 424 34582 458
rect 34616 424 34650 458
rect 34684 424 34718 458
rect 34752 424 34786 458
rect 34820 424 34854 458
rect 34888 424 34922 458
rect 34956 424 34990 458
rect 35024 424 35058 458
rect 35092 424 35126 458
rect 35160 424 35194 458
rect 35228 424 35262 458
rect 35296 424 35330 458
rect 35364 424 35398 458
rect 35432 424 35466 458
rect 35500 424 35534 458
rect 35568 424 35602 458
rect 35636 424 35670 458
rect 35704 424 35738 458
rect 35772 424 35806 458
rect 35840 424 35874 458
rect 35908 424 35942 458
rect 35976 424 36010 458
rect 36044 424 36078 458
rect 36112 424 36146 458
rect 36180 424 36214 458
rect 36248 424 36282 458
rect 36316 424 36350 458
rect 36384 424 36418 458
rect 36452 424 36486 458
rect 36520 424 36554 458
rect 36588 424 36622 458
rect 36656 424 36690 458
rect 36724 424 36758 458
rect 36792 424 36826 458
rect 36860 424 36894 458
rect 36928 424 36962 458
rect 36996 424 37030 458
rect 37064 424 37098 458
rect 37132 424 37166 458
rect 37200 424 37234 458
rect 37268 424 37302 458
rect 37336 424 37370 458
rect 37404 424 37438 458
rect 37472 424 37506 458
rect 37540 424 37574 458
rect 37608 424 37642 458
rect 37676 424 37710 458
rect 37744 424 37778 458
rect 37812 424 37846 458
rect 37880 424 37914 458
rect 37948 424 37982 458
rect 38016 424 38050 458
rect 38084 424 38118 458
rect 38152 424 38186 458
rect 38220 424 38254 458
rect 38288 424 38322 458
rect 38356 424 38390 458
rect 38424 424 38458 458
rect 38492 424 38526 458
rect 38560 424 38594 458
rect 38628 424 38662 458
rect 38696 424 38730 458
rect 38764 424 38798 458
rect 38832 424 38866 458
rect 38900 424 38934 458
rect 38968 424 39002 458
rect 39036 424 39070 458
rect 39104 424 39138 458
rect 39172 424 39206 458
rect 39240 424 39274 458
rect 39308 424 39342 458
rect 39376 424 39410 458
rect 39444 424 39478 458
rect 39512 424 39546 458
rect 39580 424 39614 458
rect 39648 424 39682 458
rect 39716 424 39750 458
rect 39784 424 39818 458
rect 39852 424 39886 458
rect 39920 424 39954 458
rect 39988 424 40022 458
rect 40056 424 40090 458
rect 40124 424 40158 458
rect 40192 424 40226 458
rect 40260 424 40294 458
rect 40328 424 40362 458
rect 40396 424 40430 458
rect 40464 424 40498 458
rect 40532 424 40566 458
rect 40600 424 40634 458
rect 40668 424 40702 458
rect 40736 424 40770 458
rect 40804 424 40838 458
rect 40872 424 40906 458
rect 40940 424 40974 458
rect 41008 424 41042 458
rect 41076 424 41110 458
rect 41144 424 41178 458
rect 41212 424 41246 458
rect 41280 424 41314 458
rect 41348 424 41382 458
rect 41416 424 41450 458
rect 41484 424 41518 458
rect 41552 424 41586 458
rect 41620 424 41654 458
rect 41688 424 41722 458
rect 41756 424 41790 458
rect 41824 424 41896 458
<< psubdiffcont >>
rect 12181 12377 14187 14791
rect 15746 11907 15780 11941
rect 15814 11907 15848 11941
rect 15882 11907 15916 11941
rect 15950 11907 15984 11941
rect 16018 11907 16052 11941
rect 16086 11907 16120 11941
rect 16154 11907 16188 11941
rect 16222 11907 16256 11941
rect 16290 11907 16324 11941
rect 16358 11907 16392 11941
rect 16426 11907 16460 11941
rect 16494 11907 16528 11941
rect 16562 11907 16596 11941
rect 16630 11907 16664 11941
rect 16698 11907 16732 11941
rect 16766 11907 16800 11941
rect 16834 11907 16868 11941
rect 16902 11907 16936 11941
rect 16970 11907 17004 11941
rect 17038 11907 17072 11941
rect 17106 11907 17140 11941
rect 17174 11907 17208 11941
rect 17242 11907 17276 11941
rect 17310 11907 17344 11941
rect 17378 11907 17412 11941
rect 17446 11907 17480 11941
rect 17514 11907 17548 11941
rect 17582 11907 17616 11941
rect 17650 11907 17684 11941
rect 17718 11907 17752 11941
rect 17786 11907 17820 11941
rect 17854 11907 17888 11941
rect 17922 11907 17956 11941
rect 17990 11907 18024 11941
rect 18058 11907 18092 11941
rect 18126 11907 18160 11941
rect 18194 11907 18228 11941
rect 18262 11907 18296 11941
rect 18330 11907 18364 11941
rect 18398 11907 18432 11941
rect 18466 11907 18500 11941
rect 18534 11907 18568 11941
rect 18602 11907 18636 11941
rect 18670 11907 18704 11941
rect 18738 11907 18772 11941
rect 18806 11907 18840 11941
rect 18874 11907 18908 11941
rect 18942 11907 18976 11941
rect 19010 11907 19044 11941
rect 19078 11907 19112 11941
rect 19146 11907 19180 11941
rect 19214 11907 19248 11941
rect 19282 11907 19316 11941
rect 19350 11907 19384 11941
rect 19418 11907 19452 11941
rect 19486 11907 19520 11941
rect 19554 11907 19588 11941
rect 19622 11907 19656 11941
rect 19690 11907 19724 11941
rect 19758 11907 19792 11941
rect 19826 11907 19860 11941
rect 19894 11907 19928 11941
rect 19962 11907 19996 11941
rect 20030 11907 20064 11941
rect 20098 11907 20132 11941
rect 20166 11907 20200 11941
rect 15746 11839 15780 11873
rect 20166 11839 20200 11873
rect 15746 11771 15780 11805
rect 15746 11703 15780 11737
rect 15746 11635 15780 11669
rect 15746 11567 15780 11601
rect 15746 11499 15780 11533
rect 15746 11431 15780 11465
rect 15746 11363 15780 11397
rect 15746 11295 15780 11329
rect 15746 11227 15780 11261
rect 10789 11117 10823 11151
rect 10876 11117 10910 11151
rect 10944 11117 10978 11151
rect 11012 11117 11046 11151
rect 11080 11117 11114 11151
rect 11168 11117 11202 11151
rect 10789 11042 10823 11076
rect 10789 10974 10823 11008
rect 10789 10906 10823 10940
rect 10789 10838 10823 10872
rect 10789 10770 10823 10804
rect 11168 11042 11202 11076
rect 11168 10974 11202 11008
rect 11168 10906 11202 10940
rect 11168 10838 11202 10872
rect 11168 10770 11202 10804
rect 15746 11159 15780 11193
rect 15746 11091 15780 11125
rect 15746 11023 15780 11057
rect 15746 10955 15780 10989
rect 20166 11771 20200 11805
rect 20166 11703 20200 11737
rect 20166 11635 20200 11669
rect 20166 11567 20200 11601
rect 20166 11499 20200 11533
rect 20166 11431 20200 11465
rect 20166 11363 20200 11397
rect 20166 11295 20200 11329
rect 20166 11227 20200 11261
rect 20166 11159 20200 11193
rect 20166 11091 20200 11125
rect 20166 11023 20200 11057
rect 20166 10955 20200 10989
rect 15746 10819 20200 10921
rect 10789 10694 10823 10728
rect 10876 10694 10910 10728
rect 10944 10694 10978 10728
rect 11012 10694 11046 10728
rect 11080 10694 11114 10728
rect 11168 10694 11202 10728
rect 16395 9843 16429 9877
rect 16509 9843 16543 9877
rect 16577 9843 16611 9877
rect 16645 9843 16679 9877
rect 16713 9843 16747 9877
rect 16781 9843 16815 9877
rect 16895 9843 16929 9877
rect 16395 9759 16429 9793
rect 16395 9691 16429 9725
rect 16395 9623 16429 9657
rect 16395 9555 16429 9589
rect 16895 9759 16929 9793
rect 16895 9691 16929 9725
rect 16895 9623 16929 9657
rect 16895 9555 16929 9589
rect 16395 9467 16429 9501
rect 16509 9467 16543 9501
rect 16577 9467 16611 9501
rect 16645 9467 16679 9501
rect 16713 9467 16747 9501
rect 16781 9467 16815 9501
rect 16895 9467 16929 9501
rect 19862 9839 19896 9873
rect 19976 9839 20010 9873
rect 20044 9839 20078 9873
rect 20112 9839 20146 9873
rect 20180 9839 20214 9873
rect 20248 9839 20282 9873
rect 20362 9839 20396 9873
rect 19862 9755 19896 9789
rect 19862 9687 19896 9721
rect 19862 9619 19896 9653
rect 19862 9551 19896 9585
rect 20362 9755 20396 9789
rect 20362 9687 20396 9721
rect 20362 9619 20396 9653
rect 20362 9551 20396 9585
rect 19862 9463 19896 9497
rect 19976 9463 20010 9497
rect 20044 9463 20078 9497
rect 20112 9463 20146 9497
rect 20180 9463 20214 9497
rect 20248 9463 20282 9497
rect 20362 9463 20396 9497
rect 16391 8448 16425 8482
rect 16505 8448 16539 8482
rect 16573 8448 16607 8482
rect 16641 8448 16675 8482
rect 16709 8448 16743 8482
rect 16777 8448 16811 8482
rect 16891 8448 16925 8482
rect 16391 8364 16425 8398
rect 16391 8296 16425 8330
rect 16391 8228 16425 8262
rect 10791 8120 10825 8154
rect 10878 8120 10912 8154
rect 10946 8120 10980 8154
rect 11014 8120 11048 8154
rect 11082 8120 11116 8154
rect 11170 8120 11204 8154
rect 10791 8045 10825 8079
rect 10791 7977 10825 8011
rect 10791 7909 10825 7943
rect 10791 7841 10825 7875
rect 10791 7773 10825 7807
rect 11170 8045 11204 8079
rect 16391 8160 16425 8194
rect 16891 8364 16925 8398
rect 16891 8296 16925 8330
rect 16891 8228 16925 8262
rect 16891 8160 16925 8194
rect 16391 8072 16425 8106
rect 16505 8072 16539 8106
rect 16573 8072 16607 8106
rect 16641 8072 16675 8106
rect 16709 8072 16743 8106
rect 16777 8072 16811 8106
rect 16891 8072 16925 8106
rect 11170 7977 11204 8011
rect 11170 7909 11204 7943
rect 11170 7841 11204 7875
rect 11170 7773 11204 7807
rect 10791 7697 10825 7731
rect 10878 7697 10912 7731
rect 10946 7697 10980 7731
rect 11014 7697 11048 7731
rect 11082 7697 11116 7731
rect 11170 7697 11204 7731
rect 5659 7473 5693 7507
rect 5727 7473 5761 7507
rect 5795 7473 5829 7507
rect 5863 7473 5897 7507
rect 5931 7473 5965 7507
rect 5999 7473 6033 7507
rect 6067 7473 6101 7507
rect 6135 7473 6169 7507
rect 6203 7473 6237 7507
rect 6271 7473 6305 7507
rect 6339 7473 6373 7507
rect 6407 7473 6441 7507
rect 6475 7473 6509 7507
rect 6543 7473 6577 7507
rect 6611 7473 6645 7507
rect 6679 7473 6713 7507
rect 6747 7473 6781 7507
rect 6815 7473 6849 7507
rect 6883 7473 6917 7507
rect 6951 7473 6985 7507
rect 7019 7473 7053 7507
rect 7087 7473 7121 7507
rect 7155 7473 7189 7507
rect 7223 7473 7257 7507
rect 7291 7473 7325 7507
rect 7359 7473 7393 7507
rect 7427 7473 7461 7507
rect 7495 7473 7529 7507
rect 7563 7473 7597 7507
rect 7631 7473 7665 7507
rect 7699 7473 7733 7507
rect 7767 7473 7801 7507
rect 7835 7473 7869 7507
rect 7903 7473 7937 7507
rect 7971 7473 8005 7507
rect 8039 7473 8073 7507
rect 8107 7473 8141 7507
rect 8175 7473 8209 7507
rect 8243 7473 8277 7507
rect 8311 7473 8345 7507
rect 8379 7473 8413 7507
rect 8447 7473 8481 7507
rect 8515 7473 8549 7507
rect 8583 7473 8617 7507
rect 8651 7473 8685 7507
rect 8719 7473 8753 7507
rect 8787 7473 8821 7507
rect 8855 7473 8889 7507
rect 8923 7473 8957 7507
rect 8991 7473 9025 7507
rect 9059 7473 9093 7507
rect 9127 7473 9161 7507
rect 9195 7473 9229 7507
rect 9263 7473 9297 7507
rect 9331 7473 9365 7507
rect 9399 7473 9433 7507
rect 9467 7473 9501 7507
rect 9535 7473 9569 7507
rect 9603 7473 9637 7507
rect 9671 7473 9705 7507
rect 9739 7473 9773 7507
rect 9807 7473 9841 7507
rect 9875 7473 9909 7507
rect 9943 7473 9977 7507
rect 10011 7473 10045 7507
rect 10079 7473 10113 7507
rect 5659 7405 5693 7439
rect 10079 7405 10113 7439
rect 5659 7337 5693 7371
rect 5659 7269 5693 7303
rect 5659 7201 5693 7235
rect 5659 7133 5693 7167
rect 5659 7065 5693 7099
rect 5659 6997 5693 7031
rect 5659 6929 5693 6963
rect 5659 6861 5693 6895
rect 5659 6793 5693 6827
rect 5659 6725 5693 6759
rect 5659 6657 5693 6691
rect 5659 6589 5693 6623
rect 5659 6521 5693 6555
rect 10079 7337 10113 7371
rect 10079 7269 10113 7303
rect 10079 7201 10113 7235
rect 10079 7133 10113 7167
rect 10079 7065 10113 7099
rect 10079 6997 10113 7031
rect 10079 6929 10113 6963
rect 10079 6861 10113 6895
rect 10079 6793 10113 6827
rect 10079 6725 10113 6759
rect 10079 6657 10113 6691
rect 10079 6589 10113 6623
rect 10079 6521 10113 6555
rect 5659 6385 10113 6487
rect 18554 9358 18588 9392
rect 18627 9358 18661 9392
rect 18695 9358 18729 9392
rect 18763 9358 18797 9392
rect 18831 9358 18865 9392
rect 18899 9358 18933 9392
rect 18967 9358 19001 9392
rect 19035 9358 19069 9392
rect 19103 9358 19137 9392
rect 19171 9358 19205 9392
rect 19239 9358 19273 9392
rect 19307 9358 19341 9392
rect 19380 9358 19414 9392
rect 18554 9269 18588 9303
rect 18554 9201 18588 9235
rect 18554 9133 18588 9167
rect 18554 9065 18588 9099
rect 18554 8997 18588 9031
rect 18554 8929 18588 8963
rect 18554 8861 18588 8895
rect 18554 8793 18588 8827
rect 18554 8725 18588 8759
rect 18554 8657 18588 8691
rect 18554 8589 18588 8623
rect 18554 8521 18588 8555
rect 18554 8453 18588 8487
rect 18554 8385 18588 8419
rect 18554 8317 18588 8351
rect 18554 8249 18588 8283
rect 18554 8181 18588 8215
rect 18554 8113 18588 8147
rect 18554 8045 18588 8079
rect 18554 7977 18588 8011
rect 19380 9269 19414 9303
rect 19380 9201 19414 9235
rect 19380 9133 19414 9167
rect 19380 9065 19414 9099
rect 19380 8997 19414 9031
rect 19380 8929 19414 8963
rect 19380 8861 19414 8895
rect 19380 8793 19414 8827
rect 19380 8725 19414 8759
rect 19380 8657 19414 8691
rect 19380 8589 19414 8623
rect 19380 8521 19414 8555
rect 19380 8453 19414 8487
rect 19380 8385 19414 8419
rect 19380 8317 19414 8351
rect 19380 8249 19414 8283
rect 19380 8181 19414 8215
rect 19380 8113 19414 8147
rect 19859 8508 19893 8542
rect 19973 8508 20007 8542
rect 20041 8508 20075 8542
rect 20109 8508 20143 8542
rect 20177 8508 20211 8542
rect 20245 8508 20279 8542
rect 20359 8508 20393 8542
rect 19859 8424 19893 8458
rect 19859 8356 19893 8390
rect 19859 8288 19893 8322
rect 19859 8220 19893 8254
rect 20359 8424 20393 8458
rect 20359 8356 20393 8390
rect 20359 8288 20393 8322
rect 20359 8220 20393 8254
rect 19859 8132 19893 8166
rect 19973 8132 20007 8166
rect 20041 8132 20075 8166
rect 20109 8132 20143 8166
rect 20177 8132 20211 8166
rect 20245 8132 20279 8166
rect 20359 8132 20393 8166
rect 19380 8045 19414 8079
rect 19380 7977 19414 8011
rect 18554 7887 18588 7921
rect 18627 7887 18661 7921
rect 18695 7887 18729 7921
rect 18763 7887 18797 7921
rect 18831 7887 18865 7921
rect 18899 7887 18933 7921
rect 18967 7887 19001 7921
rect 19035 7887 19069 7921
rect 19103 7887 19137 7921
rect 19171 7887 19205 7921
rect 19239 7887 19273 7921
rect 19307 7887 19341 7921
rect 19380 7887 19414 7921
rect 19873 7266 19907 7300
rect 19987 7266 20021 7300
rect 20055 7266 20089 7300
rect 20123 7266 20157 7300
rect 20191 7266 20225 7300
rect 20259 7266 20293 7300
rect 20373 7266 20407 7300
rect 19873 7182 19907 7216
rect 19873 7114 19907 7148
rect 19873 7046 19907 7080
rect 19873 6978 19907 7012
rect 20373 7182 20407 7216
rect 20373 7114 20407 7148
rect 20373 7046 20407 7080
rect 20373 6978 20407 7012
rect 19873 6890 19907 6924
rect 19987 6890 20021 6924
rect 20055 6890 20089 6924
rect 20123 6890 20157 6924
rect 20191 6890 20225 6924
rect 20259 6890 20293 6924
rect 20373 6890 20407 6924
rect 12405 5873 12439 5907
rect 12481 5873 12515 5907
rect 12549 5873 12583 5907
rect 12617 5873 12651 5907
rect 12685 5873 12719 5907
rect 12753 5873 12787 5907
rect 12828 5873 12862 5907
rect 12405 5785 12439 5819
rect 12405 5717 12439 5751
rect 12405 5649 12439 5683
rect 12405 5581 12439 5615
rect 12828 5785 12862 5819
rect 12828 5717 12862 5751
rect 12828 5649 12862 5683
rect 12828 5581 12862 5615
rect 12405 5494 12439 5528
rect 12481 5494 12515 5528
rect 12549 5494 12583 5528
rect 12617 5494 12651 5528
rect 12685 5494 12719 5528
rect 12753 5494 12787 5528
rect 12828 5494 12862 5528
<< nsubdiffcont >>
rect 15740 15019 15774 15053
rect 15879 14997 15913 15031
rect 15947 14997 15981 15031
rect 16015 14997 16049 15031
rect 16083 14997 16117 15031
rect 16151 14997 16185 15031
rect 16219 14997 16253 15031
rect 16287 14997 16321 15031
rect 16355 14997 16389 15031
rect 16423 14997 16457 15031
rect 16491 14997 16525 15031
rect 16559 14997 16593 15031
rect 16627 14997 16661 15031
rect 16695 14997 16729 15031
rect 16763 14997 16797 15031
rect 16831 14997 16865 15031
rect 16899 14997 16933 15031
rect 16967 14997 17001 15031
rect 17035 14997 17069 15031
rect 17103 14997 17137 15031
rect 17171 14997 17205 15031
rect 17239 14997 17273 15031
rect 17307 14997 17341 15031
rect 17375 14997 17409 15031
rect 17443 14997 17477 15031
rect 17511 14997 17545 15031
rect 17579 14997 17613 15031
rect 17647 14997 17681 15031
rect 17715 14997 17749 15031
rect 17783 14997 17817 15031
rect 17851 14997 17885 15031
rect 17919 14997 17953 15031
rect 17987 14997 18021 15031
rect 18055 14997 18089 15031
rect 18123 14997 18157 15031
rect 18191 14997 18225 15031
rect 18259 14997 18293 15031
rect 18327 14997 18361 15031
rect 18395 14997 18429 15031
rect 18463 14997 18497 15031
rect 18531 14997 18565 15031
rect 18599 14997 18633 15031
rect 18667 14997 18701 15031
rect 18735 14997 18769 15031
rect 18803 14997 18837 15031
rect 18871 14997 18905 15031
rect 18939 14997 18973 15031
rect 19007 14997 19041 15031
rect 19075 14997 19109 15031
rect 19143 14997 19177 15031
rect 19211 14997 19245 15031
rect 19279 14997 19313 15031
rect 19347 14997 19381 15031
rect 19415 14997 19449 15031
rect 19483 14997 19517 15031
rect 19551 14997 19585 15031
rect 19619 14997 19653 15031
rect 19687 14997 19721 15031
rect 19755 14997 19789 15031
rect 19823 14997 19857 15031
rect 19891 14997 19925 15031
rect 19959 14997 19993 15031
rect 20027 14997 20061 15031
rect 20152 14992 20186 15026
rect 15740 14951 15774 14985
rect 15740 14883 15774 14917
rect 15740 14815 15774 14849
rect 15740 14747 15774 14781
rect 15740 14679 15774 14713
rect 20152 14920 20186 14954
rect 20152 14852 20186 14886
rect 20152 14784 20186 14818
rect 20152 14716 20186 14750
rect 15740 14611 15774 14645
rect 15740 14543 15774 14577
rect 15740 14475 15774 14509
rect 15740 14407 15774 14441
rect 17525 14558 17559 14592
rect 17525 14490 17559 14524
rect 17525 14422 17559 14456
rect 15740 14339 15774 14373
rect 15740 14271 15774 14305
rect 17525 14354 17559 14388
rect 17525 14286 17559 14320
rect 15740 14203 15774 14237
rect 15740 14135 15774 14169
rect 15740 14067 15774 14101
rect 15740 13999 15774 14033
rect 15740 13931 15774 13965
rect 15740 13863 15774 13897
rect 15740 13795 15774 13829
rect 15740 13727 15774 13761
rect 15740 13659 15774 13693
rect 15740 13591 15774 13625
rect 15740 13523 15774 13557
rect 15740 13455 15774 13489
rect 15740 13387 15774 13421
rect 15740 13319 15774 13353
rect 15740 13251 15774 13285
rect 15740 13183 15774 13217
rect 15740 13115 15774 13149
rect 17525 14132 17559 14166
rect 17525 14064 17559 14098
rect 17525 13996 17559 14030
rect 17525 13928 17559 13962
rect 17525 13860 17559 13894
rect 17525 13792 17559 13826
rect 17525 13724 17559 13758
rect 17525 13656 17559 13690
rect 17525 13588 17559 13622
rect 17525 13520 17559 13554
rect 17525 13452 17559 13486
rect 17525 13384 17559 13418
rect 17525 13316 17559 13350
rect 17525 13248 17559 13282
rect 17525 13180 17559 13214
rect 19304 14545 19338 14579
rect 19304 14477 19338 14511
rect 19304 14409 19338 14443
rect 19304 14341 19338 14375
rect 19304 14273 19338 14307
rect 19304 14205 19338 14239
rect 20152 14648 20186 14682
rect 20152 14580 20186 14614
rect 20152 14512 20186 14546
rect 20152 14444 20186 14478
rect 20152 14307 20186 14341
rect 20152 14239 20186 14273
rect 19304 14137 19338 14171
rect 19304 14069 19338 14103
rect 19304 14001 19338 14035
rect 19304 13933 19338 13967
rect 19304 13865 19338 13899
rect 19304 13797 19338 13831
rect 19304 13729 19338 13763
rect 19304 13661 19338 13695
rect 19304 13593 19338 13627
rect 19304 13525 19338 13559
rect 19304 13457 19338 13491
rect 19304 13389 19338 13423
rect 19304 13321 19338 13355
rect 19304 13253 19338 13287
rect 19304 13185 19338 13219
rect 20152 14171 20186 14205
rect 20152 14103 20186 14137
rect 20152 14035 20186 14069
rect 20152 13967 20186 14001
rect 20152 13899 20186 13933
rect 20152 13831 20186 13865
rect 20152 13763 20186 13797
rect 20152 13695 20186 13729
rect 20152 13627 20186 13661
rect 20152 13559 20186 13593
rect 20152 13491 20186 13525
rect 20152 13423 20186 13457
rect 20152 13355 20186 13389
rect 20152 13287 20186 13321
rect 20152 13219 20186 13253
rect 20152 13151 20186 13185
rect 15740 13047 15774 13081
rect 15740 12979 15774 13013
rect 20152 13083 20186 13117
rect 20152 13015 20186 13049
rect 15740 12843 20194 12945
rect 5670 10558 5704 10592
rect 5794 10563 5828 10597
rect 5862 10563 5896 10597
rect 5930 10563 5964 10597
rect 5998 10563 6032 10597
rect 6066 10563 6100 10597
rect 6134 10563 6168 10597
rect 6202 10563 6236 10597
rect 6270 10563 6304 10597
rect 6338 10563 6372 10597
rect 6406 10563 6440 10597
rect 6474 10563 6508 10597
rect 6542 10563 6576 10597
rect 6610 10563 6644 10597
rect 6678 10563 6712 10597
rect 6746 10563 6780 10597
rect 6814 10563 6848 10597
rect 6882 10563 6916 10597
rect 6950 10563 6984 10597
rect 7018 10563 7052 10597
rect 7086 10563 7120 10597
rect 7154 10563 7188 10597
rect 7222 10563 7256 10597
rect 7290 10563 7324 10597
rect 7358 10563 7392 10597
rect 7426 10563 7460 10597
rect 7494 10563 7528 10597
rect 7562 10563 7596 10597
rect 7630 10563 7664 10597
rect 7698 10563 7732 10597
rect 7766 10563 7800 10597
rect 7834 10563 7868 10597
rect 7902 10563 7936 10597
rect 7970 10563 8004 10597
rect 8038 10563 8072 10597
rect 8106 10563 8140 10597
rect 8174 10563 8208 10597
rect 8242 10563 8276 10597
rect 8310 10563 8344 10597
rect 8378 10563 8412 10597
rect 8446 10563 8480 10597
rect 8514 10563 8548 10597
rect 8582 10563 8616 10597
rect 8650 10563 8684 10597
rect 8718 10563 8752 10597
rect 8786 10563 8820 10597
rect 8854 10563 8888 10597
rect 8922 10563 8956 10597
rect 8990 10563 9024 10597
rect 9058 10563 9092 10597
rect 9126 10563 9160 10597
rect 9194 10563 9228 10597
rect 9262 10563 9296 10597
rect 9330 10563 9364 10597
rect 9398 10563 9432 10597
rect 9466 10563 9500 10597
rect 9534 10563 9568 10597
rect 9602 10563 9636 10597
rect 9670 10563 9704 10597
rect 9738 10563 9772 10597
rect 9806 10563 9840 10597
rect 9874 10563 9908 10597
rect 9942 10563 9976 10597
rect 10082 10585 10116 10619
rect 5669 10452 5703 10486
rect 5669 10384 5703 10418
rect 5669 10316 5703 10350
rect 5669 10248 5703 10282
rect 10082 10517 10116 10551
rect 10082 10449 10116 10483
rect 10776 10499 10810 10533
rect 10879 10499 10913 10533
rect 10947 10499 10981 10533
rect 11015 10499 11049 10533
rect 11083 10499 11117 10533
rect 11187 10499 11221 10533
rect 10082 10381 10116 10415
rect 10082 10313 10116 10347
rect 10082 10245 10116 10279
rect 5669 10180 5703 10214
rect 5669 10112 5703 10146
rect 5669 10044 5703 10078
rect 5669 9976 5703 10010
rect 5670 9873 5704 9907
rect 5670 9805 5704 9839
rect 6518 10111 6552 10145
rect 6518 10043 6552 10077
rect 6518 9975 6552 10009
rect 6518 9907 6552 9941
rect 6518 9839 6552 9873
rect 5670 9737 5704 9771
rect 5670 9669 5704 9703
rect 5670 9601 5704 9635
rect 5670 9533 5704 9567
rect 5670 9465 5704 9499
rect 5670 9397 5704 9431
rect 5670 9329 5704 9363
rect 5670 9261 5704 9295
rect 5670 9193 5704 9227
rect 5670 9125 5704 9159
rect 5670 9057 5704 9091
rect 5670 8989 5704 9023
rect 5670 8921 5704 8955
rect 5670 8853 5704 8887
rect 5670 8785 5704 8819
rect 5670 8717 5704 8751
rect 6518 9771 6552 9805
rect 6518 9703 6552 9737
rect 6518 9635 6552 9669
rect 6518 9567 6552 9601
rect 6518 9499 6552 9533
rect 6518 9431 6552 9465
rect 6518 9363 6552 9397
rect 6518 9295 6552 9329
rect 6518 9227 6552 9261
rect 6518 9159 6552 9193
rect 6518 9091 6552 9125
rect 6518 9023 6552 9057
rect 6518 8955 6552 8989
rect 6518 8887 6552 8921
rect 6518 8819 6552 8853
rect 6518 8751 6552 8785
rect 8296 10141 8330 10175
rect 8296 10073 8330 10107
rect 8296 10005 8330 10039
rect 8296 9937 8330 9971
rect 10082 10177 10116 10211
rect 10082 10109 10116 10143
rect 10082 10041 10116 10075
rect 10082 9973 10116 10007
rect 8296 9869 8330 9903
rect 10082 9905 10116 9939
rect 8296 9801 8330 9835
rect 8297 9698 8331 9732
rect 8297 9630 8331 9664
rect 8297 9562 8331 9596
rect 8297 9494 8331 9528
rect 8297 9426 8331 9460
rect 8297 9358 8331 9392
rect 8297 9290 8331 9324
rect 8297 9222 8331 9256
rect 8297 9154 8331 9188
rect 8297 9086 8331 9120
rect 8297 9018 8331 9052
rect 8297 8950 8331 8984
rect 8297 8882 8331 8916
rect 8297 8814 8331 8848
rect 8297 8746 8331 8780
rect 10082 9837 10116 9871
rect 10082 9769 10116 9803
rect 10082 9701 10116 9735
rect 10082 9633 10116 9667
rect 10082 9565 10116 9599
rect 10082 9497 10116 9531
rect 10082 9429 10116 9463
rect 10082 9361 10116 9395
rect 10082 9293 10116 9327
rect 10082 9225 10116 9259
rect 10082 9157 10116 9191
rect 10082 9089 10116 9123
rect 10082 9021 10116 9055
rect 10082 8953 10116 8987
rect 10082 8885 10116 8919
rect 10082 8817 10116 8851
rect 10082 8749 10116 8783
rect 5670 8649 5704 8683
rect 5670 8581 5704 8615
rect 10082 8681 10116 8715
rect 10082 8613 10116 8647
rect 10082 8545 10116 8579
rect 10776 10414 10810 10448
rect 10776 10346 10810 10380
rect 10776 10278 10810 10312
rect 10776 10210 10810 10244
rect 10776 10142 10810 10176
rect 10776 10074 10810 10108
rect 10776 10006 10810 10040
rect 10776 9938 10810 9972
rect 10776 9870 10810 9904
rect 10776 9802 10810 9836
rect 10776 9734 10810 9768
rect 10776 9666 10810 9700
rect 10776 9598 10810 9632
rect 10776 9530 10810 9564
rect 10776 9462 10810 9496
rect 10776 9394 10810 9428
rect 10776 9326 10810 9360
rect 10776 9258 10810 9292
rect 10776 9190 10810 9224
rect 10776 9122 10810 9156
rect 10776 9054 10810 9088
rect 10776 8986 10810 9020
rect 10776 8918 10810 8952
rect 10776 8850 10810 8884
rect 10776 8782 10810 8816
rect 10776 8714 10810 8748
rect 10776 8646 10810 8680
rect 11187 10414 11221 10448
rect 11187 10346 11221 10380
rect 11187 10278 11221 10312
rect 11187 10210 11221 10244
rect 11187 10142 11221 10176
rect 11187 10074 11221 10108
rect 11187 10006 11221 10040
rect 11187 9938 11221 9972
rect 11187 9870 11221 9904
rect 11187 9802 11221 9836
rect 11187 9734 11221 9768
rect 11187 9666 11221 9700
rect 11187 9598 11221 9632
rect 11187 9530 11221 9564
rect 11187 9462 11221 9496
rect 11187 9394 11221 9428
rect 11187 9326 11221 9360
rect 11187 9258 11221 9292
rect 11187 9190 11221 9224
rect 11187 9122 11221 9156
rect 11187 9054 11221 9088
rect 11187 8986 11221 9020
rect 11187 8918 11221 8952
rect 11187 8850 11221 8884
rect 11187 8782 11221 8816
rect 11187 8714 11221 8748
rect 16490 9323 16524 9357
rect 16588 9323 16622 9357
rect 16656 9323 16690 9357
rect 16724 9323 16758 9357
rect 16792 9323 16826 9357
rect 16890 9323 16924 9357
rect 16490 9251 16524 9285
rect 16490 9183 16524 9217
rect 16490 9115 16524 9149
rect 16490 9047 16524 9081
rect 16490 8979 16524 9013
rect 16490 8911 16524 8945
rect 16490 8843 16524 8877
rect 16890 9251 16924 9285
rect 16890 9183 16924 9217
rect 16890 9115 16924 9149
rect 16890 9047 16924 9081
rect 16890 8979 16924 9013
rect 16890 8911 16924 8945
rect 16890 8843 16924 8877
rect 16490 8771 16524 8805
rect 16588 8771 16622 8805
rect 16656 8771 16690 8805
rect 16724 8771 16758 8805
rect 16792 8771 16826 8805
rect 16890 8771 16924 8805
rect 17443 9373 17477 9407
rect 17519 9373 17553 9407
rect 17587 9373 17621 9407
rect 17655 9373 17689 9407
rect 17723 9373 17757 9407
rect 17791 9373 17825 9407
rect 17859 9373 17893 9407
rect 17927 9373 17961 9407
rect 17995 9373 18029 9407
rect 18063 9373 18097 9407
rect 18131 9373 18165 9407
rect 18203 9373 18237 9407
rect 17443 9278 17477 9312
rect 17443 9210 17477 9244
rect 17443 9142 17477 9176
rect 17443 9074 17477 9108
rect 17443 9006 17477 9040
rect 17443 8938 17477 8972
rect 18203 9278 18237 9312
rect 18203 9210 18237 9244
rect 18203 9142 18237 9176
rect 18203 9074 18237 9108
rect 18203 9006 18237 9040
rect 17443 8870 17477 8904
rect 17602 8904 17636 8938
rect 17670 8904 17704 8938
rect 17738 8904 17772 8938
rect 17806 8904 17840 8938
rect 17874 8904 17908 8938
rect 17942 8904 17976 8938
rect 18010 8904 18044 8938
rect 18203 8938 18237 8972
rect 17443 8802 17477 8836
rect 11187 8646 11221 8680
rect 17443 8734 17477 8768
rect 17443 8666 17477 8700
rect 10776 8570 10810 8604
rect 10879 8570 10913 8604
rect 10947 8570 10981 8604
rect 11015 8570 11049 8604
rect 11083 8570 11117 8604
rect 11187 8570 11221 8604
rect 17443 8598 17477 8632
rect 17443 8530 17477 8564
rect 5662 8409 10116 8511
rect 17443 8462 17477 8496
rect 17443 8394 17477 8428
rect 17443 8326 17477 8360
rect 17443 8258 17477 8292
rect 17443 8190 17477 8224
rect 17443 8122 17477 8156
rect 17443 8054 17477 8088
rect 17443 7986 17477 8020
rect 16484 7927 16518 7961
rect 16582 7927 16616 7961
rect 16650 7927 16684 7961
rect 16718 7927 16752 7961
rect 16786 7927 16820 7961
rect 16884 7927 16918 7961
rect 16484 7855 16518 7889
rect 16484 7787 16518 7821
rect 16484 7719 16518 7753
rect 16484 7651 16518 7685
rect 16484 7583 16518 7617
rect 10783 7506 10817 7540
rect 10886 7506 10920 7540
rect 10954 7506 10988 7540
rect 11022 7506 11056 7540
rect 11090 7506 11124 7540
rect 11194 7506 11228 7540
rect 10783 7421 10817 7455
rect 10783 7353 10817 7387
rect 10783 7285 10817 7319
rect 10783 7217 10817 7251
rect 10783 7149 10817 7183
rect 10783 7081 10817 7115
rect 10783 7013 10817 7047
rect 10783 6945 10817 6979
rect 10783 6877 10817 6911
rect 10783 6809 10817 6843
rect 10783 6741 10817 6775
rect 10783 6673 10817 6707
rect 10783 6605 10817 6639
rect 10783 6537 10817 6571
rect 10783 6469 10817 6503
rect 10783 6401 10817 6435
rect 10783 6333 10817 6367
rect 10783 6265 10817 6299
rect 10783 6197 10817 6231
rect 10783 6129 10817 6163
rect 10783 6061 10817 6095
rect 10783 5993 10817 6027
rect 10783 5925 10817 5959
rect 10783 5857 10817 5891
rect 10783 5789 10817 5823
rect 10783 5721 10817 5755
rect 10783 5653 10817 5687
rect 11194 7421 11228 7455
rect 16484 7515 16518 7549
rect 16484 7447 16518 7481
rect 11194 7353 11228 7387
rect 16884 7855 16918 7889
rect 18203 8870 18237 8904
rect 18203 8802 18237 8836
rect 18203 8734 18237 8768
rect 18203 8666 18237 8700
rect 18203 8598 18237 8632
rect 18203 8530 18237 8564
rect 18203 8462 18237 8496
rect 18203 8394 18237 8428
rect 18203 8326 18237 8360
rect 18203 8258 18237 8292
rect 18203 8190 18237 8224
rect 18203 8122 18237 8156
rect 18203 8054 18237 8088
rect 18203 7986 18237 8020
rect 19957 9318 19991 9352
rect 20055 9318 20089 9352
rect 20123 9318 20157 9352
rect 20191 9318 20225 9352
rect 20259 9318 20293 9352
rect 20357 9318 20391 9352
rect 19957 9246 19991 9280
rect 19957 9178 19991 9212
rect 19957 9110 19991 9144
rect 19957 9042 19991 9076
rect 19957 8974 19991 9008
rect 19957 8906 19991 8940
rect 19957 8838 19991 8872
rect 20357 9246 20391 9280
rect 20357 9178 20391 9212
rect 20357 9110 20391 9144
rect 20357 9042 20391 9076
rect 20357 8974 20391 9008
rect 20357 8906 20391 8940
rect 20357 8838 20391 8872
rect 19957 8766 19991 8800
rect 20055 8766 20089 8800
rect 20123 8766 20157 8800
rect 20191 8766 20225 8800
rect 20259 8766 20293 8800
rect 20357 8766 20391 8800
rect 17443 7885 17477 7919
rect 17519 7885 17553 7919
rect 17587 7885 17621 7919
rect 17655 7885 17689 7919
rect 17723 7885 17757 7919
rect 17791 7885 17825 7919
rect 17859 7885 17893 7919
rect 17927 7885 17961 7919
rect 17995 7885 18029 7919
rect 18063 7885 18097 7919
rect 18131 7885 18165 7919
rect 18203 7885 18237 7919
rect 19953 7987 19987 8021
rect 20051 7987 20085 8021
rect 20119 7987 20153 8021
rect 20187 7987 20221 8021
rect 20255 7987 20289 8021
rect 20353 7987 20387 8021
rect 19953 7915 19987 7949
rect 16884 7787 16918 7821
rect 16884 7719 16918 7753
rect 16884 7651 16918 7685
rect 16884 7583 16918 7617
rect 16884 7515 16918 7549
rect 16884 7447 16918 7481
rect 19953 7847 19987 7881
rect 19953 7779 19987 7813
rect 19953 7711 19987 7745
rect 19953 7643 19987 7677
rect 19953 7575 19987 7609
rect 19953 7507 19987 7541
rect 20353 7915 20387 7949
rect 20353 7847 20387 7881
rect 20353 7779 20387 7813
rect 20353 7711 20387 7745
rect 20353 7643 20387 7677
rect 20353 7575 20387 7609
rect 20353 7507 20387 7541
rect 19953 7435 19987 7469
rect 20051 7435 20085 7469
rect 20119 7435 20153 7469
rect 20187 7435 20221 7469
rect 20255 7435 20289 7469
rect 20353 7435 20387 7469
rect 16484 7375 16518 7409
rect 16582 7375 16616 7409
rect 16650 7375 16684 7409
rect 16718 7375 16752 7409
rect 16786 7375 16820 7409
rect 16884 7375 16918 7409
rect 11194 7285 11228 7319
rect 11194 7217 11228 7251
rect 11194 7149 11228 7183
rect 11194 7081 11228 7115
rect 11194 7013 11228 7047
rect 11194 6945 11228 6979
rect 11194 6877 11228 6911
rect 11194 6809 11228 6843
rect 11194 6741 11228 6775
rect 11194 6673 11228 6707
rect 11194 6605 11228 6639
rect 11194 6537 11228 6571
rect 11194 6469 11228 6503
rect 11194 6401 11228 6435
rect 11194 6333 11228 6367
rect 11194 6265 11228 6299
rect 11194 6197 11228 6231
rect 19971 6745 20005 6779
rect 20069 6745 20103 6779
rect 20137 6745 20171 6779
rect 20205 6745 20239 6779
rect 20273 6745 20307 6779
rect 20371 6745 20405 6779
rect 19971 6673 20005 6707
rect 19971 6605 20005 6639
rect 19971 6537 20005 6571
rect 19971 6469 20005 6503
rect 19971 6401 20005 6435
rect 19971 6333 20005 6367
rect 19971 6265 20005 6299
rect 20371 6673 20405 6707
rect 20371 6605 20405 6639
rect 20371 6537 20405 6571
rect 20371 6469 20405 6503
rect 20371 6401 20405 6435
rect 20371 6333 20405 6367
rect 20371 6265 20405 6299
rect 19971 6193 20005 6227
rect 20069 6193 20103 6227
rect 20137 6193 20171 6227
rect 20205 6193 20239 6227
rect 20273 6193 20307 6227
rect 20371 6193 20405 6227
rect 11194 6129 11228 6163
rect 11194 6061 11228 6095
rect 11194 5993 11228 6027
rect 11194 5925 11228 5959
rect 11194 5857 11228 5891
rect 11194 5789 11228 5823
rect 11194 5721 11228 5755
rect 11194 5653 11228 5687
rect 10783 5577 10817 5611
rect 10886 5577 10920 5611
rect 10954 5577 10988 5611
rect 11022 5577 11056 5611
rect 11090 5577 11124 5611
rect 11194 5577 11228 5611
rect 13020 5879 13054 5913
rect 13105 5879 13139 5913
rect 13173 5879 13207 5913
rect 13241 5879 13275 5913
rect 13309 5879 13343 5913
rect 13377 5879 13411 5913
rect 13445 5879 13479 5913
rect 13513 5879 13547 5913
rect 13581 5879 13615 5913
rect 13649 5879 13683 5913
rect 13717 5879 13751 5913
rect 13785 5879 13819 5913
rect 13853 5879 13887 5913
rect 13921 5879 13955 5913
rect 13989 5879 14023 5913
rect 14057 5879 14091 5913
rect 14125 5879 14159 5913
rect 14193 5879 14227 5913
rect 14261 5879 14295 5913
rect 14329 5879 14363 5913
rect 14397 5879 14431 5913
rect 14465 5879 14499 5913
rect 14533 5879 14567 5913
rect 14601 5879 14635 5913
rect 14669 5879 14703 5913
rect 14737 5879 14771 5913
rect 14805 5879 14839 5913
rect 14873 5879 14907 5913
rect 14949 5879 14983 5913
rect 13020 5775 13054 5809
rect 13020 5707 13054 5741
rect 13020 5639 13054 5673
rect 13020 5571 13054 5605
rect 14949 5775 14983 5809
rect 14949 5707 14983 5741
rect 14949 5639 14983 5673
rect 14949 5571 14983 5605
rect 13020 5466 13054 5500
rect 13105 5468 13139 5502
rect 13173 5468 13207 5502
rect 13241 5468 13275 5502
rect 13309 5468 13343 5502
rect 13377 5468 13411 5502
rect 13445 5468 13479 5502
rect 13513 5468 13547 5502
rect 13581 5468 13615 5502
rect 13649 5468 13683 5502
rect 13717 5468 13751 5502
rect 13785 5468 13819 5502
rect 13853 5468 13887 5502
rect 13921 5468 13955 5502
rect 13989 5468 14023 5502
rect 14057 5468 14091 5502
rect 14125 5468 14159 5502
rect 14193 5468 14227 5502
rect 14261 5468 14295 5502
rect 14329 5468 14363 5502
rect 14397 5468 14431 5502
rect 14465 5468 14499 5502
rect 14533 5468 14567 5502
rect 14601 5468 14635 5502
rect 14669 5468 14703 5502
rect 14737 5468 14771 5502
rect 14805 5468 14839 5502
rect 14873 5468 14907 5502
rect 14949 5468 14983 5502
rect 5546 2572 5580 2606
rect 5614 2572 5648 2606
rect 5682 2572 5716 2606
rect 5750 2572 5784 2606
rect 5818 2572 5852 2606
rect 5886 2572 5920 2606
rect 5954 2572 5988 2606
rect 6022 2572 6056 2606
rect 6090 2572 6124 2606
rect 6158 2572 6192 2606
rect 6226 2572 6260 2606
rect 6294 2572 6328 2606
rect 6362 2572 6396 2606
rect 6430 2572 6464 2606
rect 6498 2572 6532 2606
rect 6566 2572 6600 2606
rect 6634 2572 6668 2606
rect 6702 2572 6736 2606
rect 6770 2572 6804 2606
rect 6838 2572 6872 2606
rect 6906 2572 6940 2606
rect 6974 2572 7008 2606
rect 7042 2572 7076 2606
rect 7110 2572 7144 2606
rect 7178 2572 7212 2606
rect 7246 2572 7280 2606
rect 7314 2572 7348 2606
rect 7382 2572 7416 2606
rect 7450 2572 7484 2606
rect 7518 2572 7552 2606
rect 7586 2572 7620 2606
rect 7654 2572 7688 2606
rect 7722 2572 7756 2606
rect 7790 2572 7824 2606
rect 7858 2572 7892 2606
rect 7926 2572 7960 2606
rect 7994 2572 8028 2606
rect 8062 2572 8096 2606
rect 8130 2572 8164 2606
rect 8198 2572 8232 2606
rect 8266 2572 8300 2606
rect 8334 2572 8368 2606
rect 8402 2572 8436 2606
rect 8470 2572 8504 2606
rect 8538 2572 8572 2606
rect 8606 2572 8640 2606
rect 8674 2572 8708 2606
rect 8742 2572 8776 2606
rect 8810 2572 8844 2606
rect 8878 2572 8912 2606
rect 8946 2572 8980 2606
rect 9014 2572 9048 2606
rect 9082 2572 9116 2606
rect 9150 2572 9184 2606
rect 9218 2572 9252 2606
rect 9286 2572 9320 2606
rect 9354 2572 9388 2606
rect 9422 2572 9456 2606
rect 9490 2572 9524 2606
rect 9558 2572 9592 2606
rect 9626 2572 9660 2606
rect 9694 2572 9728 2606
rect 9762 2572 9796 2606
rect 9830 2572 9864 2606
rect 9898 2572 9932 2606
rect 9966 2572 10000 2606
rect 10034 2572 10068 2606
rect 10102 2572 10136 2606
rect 10170 2572 10204 2606
rect 10238 2572 10272 2606
rect 10306 2572 10340 2606
rect 10374 2572 10408 2606
rect 10442 2572 10476 2606
rect 10510 2572 10544 2606
rect 10578 2572 10612 2606
rect 10646 2572 10680 2606
rect 10714 2572 10748 2606
rect 10782 2572 10816 2606
rect 10850 2572 10884 2606
rect 10918 2572 10952 2606
rect 10986 2572 11020 2606
rect 11054 2572 11088 2606
rect 11122 2572 11156 2606
rect 11190 2572 11224 2606
rect 11258 2572 11292 2606
rect 11326 2572 11360 2606
rect 11394 2572 11428 2606
rect 11462 2572 11496 2606
rect 11530 2572 11564 2606
rect 11598 2572 11632 2606
rect 11666 2572 11700 2606
rect 11734 2572 11768 2606
rect 11802 2572 11836 2606
rect 11870 2572 11904 2606
rect 11938 2572 11972 2606
rect 12006 2572 12040 2606
rect 12074 2572 12108 2606
rect 12142 2572 12176 2606
rect 12210 2572 12244 2606
rect 12278 2572 12312 2606
rect 12346 2572 12380 2606
rect 12414 2572 12448 2606
rect 12482 2572 12516 2606
rect 12550 2572 12584 2606
rect 12618 2572 12652 2606
rect 12686 2572 12720 2606
rect 12754 2572 12788 2606
rect 12822 2572 12856 2606
rect 12890 2572 12924 2606
rect 12958 2572 12992 2606
rect 13026 2572 13060 2606
rect 13094 2572 13128 2606
rect 13162 2572 13196 2606
rect 13230 2572 13264 2606
rect 13298 2572 13332 2606
rect 13366 2572 13400 2606
rect 13434 2572 13468 2606
rect 13502 2572 13536 2606
rect 13570 2572 13604 2606
rect 13638 2572 13672 2606
rect 13706 2572 13740 2606
rect 13774 2572 13808 2606
rect 13842 2572 13876 2606
rect 13910 2572 13944 2606
rect 13978 2572 14012 2606
rect 14046 2572 14080 2606
rect 14114 2572 14148 2606
rect 14182 2572 14216 2606
rect 14250 2572 14284 2606
rect 14318 2572 14352 2606
rect 14386 2572 14420 2606
rect 14454 2572 14488 2606
rect 14522 2572 14556 2606
rect 14590 2572 14624 2606
rect 14658 2572 14692 2606
rect 14726 2572 14760 2606
rect 14794 2572 14828 2606
rect 14862 2572 14896 2606
rect 14930 2572 14964 2606
rect 14998 2572 15032 2606
rect 15066 2572 15100 2606
rect 15134 2572 15168 2606
rect 15202 2572 15236 2606
rect 15270 2572 15304 2606
rect 15338 2572 15372 2606
rect 15406 2572 15440 2606
rect 15474 2572 15508 2606
rect 15542 2572 15576 2606
rect 15610 2572 15644 2606
rect 15678 2572 15712 2606
rect 15746 2572 15780 2606
rect 15814 2572 15848 2606
rect 15882 2572 15916 2606
rect 15950 2572 15984 2606
rect 16018 2572 16052 2606
rect 16086 2572 16120 2606
rect 16154 2572 16188 2606
rect 16222 2572 16256 2606
rect 16290 2572 16324 2606
rect 16358 2572 16392 2606
rect 16426 2572 16460 2606
rect 16494 2572 16528 2606
rect 16562 2572 16596 2606
rect 16630 2572 16664 2606
rect 16698 2572 16732 2606
rect 16766 2572 16800 2606
rect 16834 2572 16868 2606
rect 16902 2572 16936 2606
rect 16970 2572 17004 2606
rect 17038 2572 17072 2606
rect 17106 2572 17140 2606
rect 17174 2572 17208 2606
rect 17242 2572 17276 2606
rect 17310 2572 17344 2606
rect 17378 2572 17412 2606
rect 17446 2572 17480 2606
rect 17514 2572 17548 2606
rect 17582 2572 17616 2606
rect 17650 2572 17684 2606
rect 17718 2572 17752 2606
rect 17786 2572 17820 2606
rect 17854 2572 17888 2606
rect 17922 2572 17956 2606
rect 17990 2572 18024 2606
rect 18058 2572 18092 2606
rect 18126 2572 18160 2606
rect 18194 2572 18228 2606
rect 18262 2572 18296 2606
rect 18330 2572 18364 2606
rect 18398 2572 18432 2606
rect 18466 2572 18500 2606
rect 18534 2572 18568 2606
rect 18602 2572 18636 2606
rect 18670 2572 18704 2606
rect 18738 2572 18772 2606
rect 18806 2572 18840 2606
rect 18874 2572 18908 2606
rect 18942 2572 18976 2606
rect 19010 2572 19044 2606
rect 19078 2572 19112 2606
rect 19146 2572 19180 2606
rect 19214 2572 19248 2606
rect 19282 2572 19316 2606
rect 19350 2572 19384 2606
rect 19418 2572 19452 2606
rect 19486 2572 19520 2606
rect 19554 2572 19588 2606
rect 19622 2572 19656 2606
rect 19690 2572 19724 2606
rect 19758 2572 19792 2606
rect 19826 2572 19860 2606
rect 19894 2572 19928 2606
rect 19962 2572 19996 2606
rect 20030 2572 20064 2606
rect 20098 2572 20132 2606
rect 20166 2572 20200 2606
rect 20234 2572 20268 2606
rect 20302 2572 20336 2606
rect 20370 2572 20404 2606
rect 20438 2572 20472 2606
rect 20506 2572 20540 2606
rect 20574 2572 20608 2606
rect 20642 2572 20676 2606
rect 20710 2572 20744 2606
rect 20778 2572 20812 2606
rect 20846 2572 20880 2606
rect 20914 2572 20948 2606
rect 20982 2572 21016 2606
rect 21050 2572 21084 2606
rect 21118 2572 21152 2606
rect 21186 2572 21220 2606
rect 21254 2572 21288 2606
rect 21322 2572 21356 2606
rect 21390 2572 21424 2606
rect 21458 2572 21492 2606
rect 21526 2572 21560 2606
rect 21594 2572 21628 2606
rect 21662 2572 21696 2606
rect 21730 2572 21764 2606
rect 21798 2572 21832 2606
rect 21866 2572 21900 2606
rect 21934 2572 21968 2606
rect 22002 2572 22036 2606
rect 22070 2572 22104 2606
rect 22138 2572 22172 2606
rect 22206 2572 22240 2606
rect 22274 2572 22308 2606
rect 22342 2572 22376 2606
rect 22410 2572 22444 2606
rect 22478 2572 22512 2606
rect 22546 2572 22580 2606
rect 22614 2572 22648 2606
rect 22682 2572 22716 2606
rect 22750 2572 22784 2606
rect 22818 2572 22852 2606
rect 22886 2572 22920 2606
rect 22954 2572 22988 2606
rect 23022 2572 23056 2606
rect 23090 2572 23124 2606
rect 23158 2572 23192 2606
rect 23226 2572 23260 2606
rect 23294 2572 23328 2606
rect 23362 2572 23396 2606
rect 23430 2572 23464 2606
rect 23498 2572 23532 2606
rect 23566 2572 23600 2606
rect 23634 2572 23668 2606
rect 23702 2572 23736 2606
rect 23770 2572 23804 2606
rect 23838 2572 23872 2606
rect 23906 2572 23940 2606
rect 23974 2572 24008 2606
rect 24042 2572 24076 2606
rect 24110 2572 24144 2606
rect 24178 2572 24212 2606
rect 24246 2572 24280 2606
rect 24314 2572 24348 2606
rect 24382 2572 24416 2606
rect 24450 2572 24484 2606
rect 24518 2572 24552 2606
rect 24586 2572 24620 2606
rect 24654 2572 24688 2606
rect 24722 2572 24756 2606
rect 24790 2572 24824 2606
rect 24858 2572 24892 2606
rect 24926 2572 24960 2606
rect 24994 2572 25028 2606
rect 25062 2572 25096 2606
rect 25130 2572 25164 2606
rect 25198 2572 25232 2606
rect 25266 2572 25300 2606
rect 25334 2572 25368 2606
rect 25402 2572 25436 2606
rect 25470 2572 25504 2606
rect 25538 2572 25572 2606
rect 25606 2572 25640 2606
rect 25674 2572 25708 2606
rect 25742 2572 25776 2606
rect 25810 2572 25844 2606
rect 25878 2572 25912 2606
rect 25946 2572 25980 2606
rect 26014 2572 26048 2606
rect 26082 2572 26116 2606
rect 26150 2572 26184 2606
rect 26218 2572 26252 2606
rect 26286 2572 26320 2606
rect 26354 2572 26388 2606
rect 26422 2572 26456 2606
rect 26490 2572 26524 2606
rect 26558 2572 26592 2606
rect 26626 2572 26660 2606
rect 26694 2572 26728 2606
rect 26762 2572 26796 2606
rect 26830 2572 26864 2606
rect 26898 2572 26932 2606
rect 26966 2572 27000 2606
rect 27034 2572 27068 2606
rect 27102 2572 27136 2606
rect 27170 2572 27204 2606
rect 27238 2572 27272 2606
rect 27306 2572 27340 2606
rect 27374 2572 27408 2606
rect 27442 2572 27476 2606
rect 27510 2572 27544 2606
rect 27578 2572 27612 2606
rect 27646 2572 27680 2606
rect 27714 2572 27748 2606
rect 27782 2572 27816 2606
rect 27850 2572 27884 2606
rect 27918 2572 27952 2606
rect 27986 2572 28020 2606
rect 28054 2572 28088 2606
rect 28122 2572 28156 2606
rect 28190 2572 28224 2606
rect 28258 2572 28292 2606
rect 28326 2572 28360 2606
rect 28394 2572 28428 2606
rect 28462 2572 28496 2606
rect 28530 2572 28564 2606
rect 28598 2572 28632 2606
rect 28666 2572 28700 2606
rect 28734 2572 28768 2606
rect 28802 2572 28836 2606
rect 28870 2572 28904 2606
rect 28938 2572 28972 2606
rect 29006 2572 29040 2606
rect 29074 2572 29108 2606
rect 29142 2572 29176 2606
rect 29210 2572 29244 2606
rect 29278 2572 29312 2606
rect 29346 2572 29380 2606
rect 29414 2572 29448 2606
rect 29482 2572 29516 2606
rect 29550 2572 29584 2606
rect 29618 2572 29652 2606
rect 29686 2572 29720 2606
rect 29754 2572 29788 2606
rect 29822 2572 29856 2606
rect 29890 2572 29924 2606
rect 29958 2572 29992 2606
rect 30026 2572 30060 2606
rect 30094 2572 30128 2606
rect 30162 2572 30196 2606
rect 30230 2572 30264 2606
rect 30298 2572 30332 2606
rect 30366 2572 30400 2606
rect 30434 2572 30468 2606
rect 30502 2572 30536 2606
rect 30570 2572 30604 2606
rect 30638 2572 30672 2606
rect 30706 2572 30740 2606
rect 30774 2572 30808 2606
rect 30842 2572 30876 2606
rect 30910 2572 30944 2606
rect 30978 2572 31012 2606
rect 31046 2572 31080 2606
rect 31114 2572 31148 2606
rect 31182 2572 31216 2606
rect 31250 2572 31284 2606
rect 31318 2572 31352 2606
rect 31386 2572 31420 2606
rect 31454 2572 31488 2606
rect 31522 2572 31556 2606
rect 31590 2572 31624 2606
rect 31658 2572 31692 2606
rect 31726 2572 31760 2606
rect 31794 2572 31828 2606
rect 31862 2572 31896 2606
rect 31930 2572 31964 2606
rect 31998 2572 32032 2606
rect 32066 2572 32100 2606
rect 32134 2572 32168 2606
rect 32202 2572 32236 2606
rect 32270 2572 32304 2606
rect 32338 2572 32372 2606
rect 32406 2572 32440 2606
rect 32474 2572 32508 2606
rect 32542 2572 32576 2606
rect 32610 2572 32644 2606
rect 32678 2572 32712 2606
rect 32746 2572 32780 2606
rect 32814 2572 32848 2606
rect 32882 2572 32916 2606
rect 32950 2572 32984 2606
rect 33018 2572 33052 2606
rect 33086 2572 33120 2606
rect 33154 2572 33188 2606
rect 33222 2572 33256 2606
rect 33290 2572 33324 2606
rect 33358 2572 33392 2606
rect 33426 2572 33460 2606
rect 33494 2572 33528 2606
rect 33562 2572 33596 2606
rect 33630 2572 33664 2606
rect 33698 2572 33732 2606
rect 33766 2572 33800 2606
rect 33834 2572 33868 2606
rect 33902 2572 33936 2606
rect 33970 2572 34004 2606
rect 34038 2572 34072 2606
rect 34106 2572 34140 2606
rect 34174 2572 34208 2606
rect 34242 2572 34276 2606
rect 34310 2572 34344 2606
rect 34378 2572 34412 2606
rect 34446 2572 34480 2606
rect 34514 2572 34548 2606
rect 34582 2572 34616 2606
rect 34650 2572 34684 2606
rect 34718 2572 34752 2606
rect 34786 2572 34820 2606
rect 34854 2572 34888 2606
rect 34922 2572 34956 2606
rect 34990 2572 35024 2606
rect 35058 2572 35092 2606
rect 35126 2572 35160 2606
rect 35194 2572 35228 2606
rect 35262 2572 35296 2606
rect 35330 2572 35364 2606
rect 35398 2572 35432 2606
rect 35466 2572 35500 2606
rect 35534 2572 35568 2606
rect 35602 2572 35636 2606
rect 35670 2572 35704 2606
rect 35738 2572 35772 2606
rect 35806 2572 35840 2606
rect 35874 2572 35908 2606
rect 35942 2572 35976 2606
rect 36010 2572 36044 2606
rect 36078 2572 36112 2606
rect 36146 2572 36180 2606
rect 36214 2572 36248 2606
rect 36282 2572 36316 2606
rect 36350 2572 36384 2606
rect 36418 2572 36452 2606
rect 36486 2572 36520 2606
rect 36554 2572 36588 2606
rect 36622 2572 36656 2606
rect 36690 2572 36724 2606
rect 36758 2572 36792 2606
rect 36826 2572 36860 2606
rect 36894 2572 36928 2606
rect 36962 2572 36996 2606
rect 37030 2572 37064 2606
rect 37098 2572 37132 2606
rect 37166 2572 37200 2606
rect 37234 2572 37268 2606
rect 37302 2572 37336 2606
rect 37370 2572 37404 2606
rect 37438 2572 37472 2606
rect 37506 2572 37540 2606
rect 37574 2572 37608 2606
rect 37642 2572 37676 2606
rect 37710 2572 37744 2606
rect 37778 2572 37812 2606
rect 37846 2572 37880 2606
rect 37914 2572 37948 2606
rect 37982 2572 38016 2606
rect 38050 2572 38084 2606
rect 38118 2572 38152 2606
rect 38186 2572 38220 2606
rect 38254 2572 38288 2606
rect 38322 2572 38356 2606
rect 38390 2572 38424 2606
rect 38458 2572 38492 2606
rect 38526 2572 38560 2606
rect 38594 2572 38628 2606
rect 38662 2572 38696 2606
rect 38730 2572 38764 2606
rect 38798 2572 38832 2606
rect 38866 2572 38900 2606
rect 38934 2572 38968 2606
rect 39002 2572 39036 2606
rect 39070 2572 39104 2606
rect 39138 2572 39172 2606
rect 39206 2572 39240 2606
rect 39274 2572 39308 2606
rect 39342 2572 39376 2606
rect 39410 2572 39444 2606
rect 39478 2572 39512 2606
rect 39546 2572 39580 2606
rect 39614 2572 39648 2606
rect 39682 2572 39716 2606
rect 39750 2572 39784 2606
rect 39818 2572 39852 2606
rect 39886 2572 39920 2606
rect 39954 2572 39988 2606
rect 40022 2572 40056 2606
rect 40090 2572 40124 2606
rect 40158 2572 40192 2606
rect 40226 2572 40260 2606
rect 40294 2572 40328 2606
rect 40362 2572 40396 2606
rect 40430 2572 40464 2606
rect 40498 2572 40532 2606
rect 40566 2572 40600 2606
rect 40634 2572 40668 2606
rect 40702 2572 40736 2606
rect 40770 2572 40804 2606
rect 40838 2572 40872 2606
rect 40906 2572 40940 2606
rect 40974 2572 41008 2606
rect 41042 2572 41076 2606
rect 41110 2572 41144 2606
rect 41178 2572 41212 2606
rect 41246 2572 41280 2606
rect 41314 2572 41348 2606
rect 41382 2572 41416 2606
rect 41450 2572 41484 2606
rect 41518 2572 41552 2606
rect 41586 2572 41620 2606
rect 41654 2572 41688 2606
rect 41722 2572 41756 2606
rect 41790 2572 41824 2606
rect 5440 2450 5474 2484
rect 5440 2382 5474 2416
rect 5440 2314 5474 2348
rect 5440 2246 5474 2280
rect 5440 2178 5474 2212
rect 5440 2110 5474 2144
rect 5440 2042 5474 2076
rect 5440 1974 5474 2008
rect 5440 1906 5474 1940
rect 5440 1838 5474 1872
rect 5440 1770 5474 1804
rect 5440 1702 5474 1736
rect 5440 1634 5474 1668
rect 5440 1566 5474 1600
rect 5440 1498 5474 1532
rect 5440 1430 5474 1464
rect 5440 1362 5474 1396
rect 5440 1294 5474 1328
rect 5440 1226 5474 1260
rect 5440 1158 5474 1192
rect 5440 1090 5474 1124
rect 5440 1022 5474 1056
rect 5440 954 5474 988
rect 5440 886 5474 920
rect 5440 818 5474 852
rect 5440 750 5474 784
rect 5440 682 5474 716
rect 5440 614 5474 648
rect 5440 546 5474 580
rect 5546 424 5580 458
rect 5614 424 5648 458
rect 5682 424 5716 458
rect 5750 424 5784 458
rect 5818 424 5852 458
rect 5886 424 5920 458
rect 5954 424 5988 458
rect 6022 424 6056 458
rect 6090 424 6124 458
rect 6158 424 6192 458
rect 6226 424 6260 458
rect 6294 424 6328 458
rect 6362 424 6396 458
rect 6430 424 6464 458
rect 6498 424 6532 458
rect 6566 424 6600 458
rect 6634 424 6668 458
rect 6702 424 6736 458
rect 6770 424 6804 458
rect 6838 424 6872 458
rect 6906 424 6940 458
rect 6974 424 7008 458
rect 7042 424 7076 458
rect 7110 424 7144 458
rect 7178 424 7212 458
rect 7246 424 7280 458
rect 7314 424 7348 458
rect 7382 424 7416 458
rect 7450 424 7484 458
rect 7518 424 7552 458
rect 7586 424 7620 458
rect 7654 424 7688 458
rect 7722 424 7756 458
rect 7790 424 7824 458
rect 7858 424 7892 458
rect 7926 424 7960 458
rect 7994 424 8028 458
rect 8062 424 8096 458
rect 8130 424 8164 458
rect 8198 424 8232 458
rect 8266 424 8300 458
rect 8334 424 8368 458
rect 8402 424 8436 458
rect 8470 424 8504 458
rect 8538 424 8572 458
rect 8606 424 8640 458
rect 8674 424 8708 458
rect 8742 424 8776 458
rect 8810 424 8844 458
rect 8878 424 8912 458
rect 8946 424 8980 458
rect 9014 424 9048 458
rect 9082 424 9116 458
rect 9150 424 9184 458
rect 9218 424 9252 458
rect 9286 424 9320 458
rect 9354 424 9388 458
rect 9422 424 9456 458
rect 9490 424 9524 458
rect 9558 424 9592 458
rect 9626 424 9660 458
rect 9694 424 9728 458
rect 9762 424 9796 458
rect 9830 424 9864 458
rect 9898 424 9932 458
rect 9966 424 10000 458
rect 10034 424 10068 458
rect 10102 424 10136 458
rect 10170 424 10204 458
rect 10238 424 10272 458
rect 10306 424 10340 458
rect 10374 424 10408 458
rect 10442 424 10476 458
rect 10510 424 10544 458
rect 10578 424 10612 458
rect 10646 424 10680 458
rect 10714 424 10748 458
rect 10782 424 10816 458
rect 10850 424 10884 458
rect 10918 424 10952 458
rect 10986 424 11020 458
rect 11054 424 11088 458
rect 11122 424 11156 458
rect 11190 424 11224 458
rect 11258 424 11292 458
rect 11326 424 11360 458
rect 11394 424 11428 458
rect 11462 424 11496 458
rect 11530 424 11564 458
rect 11598 424 11632 458
rect 11666 424 11700 458
rect 11734 424 11768 458
rect 11802 424 11836 458
rect 11870 424 11904 458
rect 11938 424 11972 458
rect 12006 424 12040 458
rect 12074 424 12108 458
rect 12142 424 12176 458
rect 12210 424 12244 458
rect 12278 424 12312 458
rect 12346 424 12380 458
rect 12414 424 12448 458
rect 12482 424 12516 458
rect 12550 424 12584 458
rect 12618 424 12652 458
rect 12686 424 12720 458
rect 12754 424 12788 458
rect 12822 424 12856 458
rect 12890 424 12924 458
rect 12958 424 12992 458
rect 13026 424 13060 458
rect 13094 424 13128 458
rect 13162 424 13196 458
rect 13230 424 13264 458
rect 13298 424 13332 458
rect 13366 424 13400 458
rect 13434 424 13468 458
rect 13502 424 13536 458
rect 13570 424 13604 458
rect 13638 424 13672 458
rect 13706 424 13740 458
rect 13774 424 13808 458
rect 13842 424 13876 458
rect 13910 424 13944 458
rect 13978 424 14012 458
rect 14046 424 14080 458
rect 14114 424 14148 458
rect 14182 424 14216 458
rect 14250 424 14284 458
rect 14318 424 14352 458
rect 14386 424 14420 458
rect 14454 424 14488 458
rect 14522 424 14556 458
rect 14590 424 14624 458
rect 14658 424 14692 458
rect 14726 424 14760 458
rect 14794 424 14828 458
rect 14862 424 14896 458
rect 14930 424 14964 458
rect 14998 424 15032 458
rect 15066 424 15100 458
rect 15134 424 15168 458
rect 15202 424 15236 458
rect 15270 424 15304 458
rect 15338 424 15372 458
rect 15406 424 15440 458
rect 15474 424 15508 458
rect 15542 424 15576 458
rect 15610 424 15644 458
rect 15678 424 15712 458
rect 15746 424 15780 458
rect 15814 424 15848 458
rect 15882 424 15916 458
rect 15950 424 15984 458
rect 16018 424 16052 458
rect 16086 424 16120 458
rect 16154 424 16188 458
rect 16222 424 16256 458
rect 16290 424 16324 458
rect 16358 424 16392 458
rect 16426 424 16460 458
rect 16494 424 16528 458
rect 16562 424 16596 458
rect 16630 424 16664 458
rect 16698 424 16732 458
rect 16766 424 16800 458
rect 16834 424 16868 458
rect 16902 424 16936 458
rect 16970 424 17004 458
rect 17038 424 17072 458
rect 17106 424 17140 458
rect 17174 424 17208 458
rect 17242 424 17276 458
rect 17310 424 17344 458
rect 17378 424 17412 458
rect 17446 424 17480 458
rect 17514 424 17548 458
rect 17582 424 17616 458
rect 17650 424 17684 458
rect 17718 424 17752 458
rect 17786 424 17820 458
rect 17854 424 17888 458
rect 17922 424 17956 458
rect 17990 424 18024 458
rect 18058 424 18092 458
rect 18126 424 18160 458
rect 18194 424 18228 458
rect 18262 424 18296 458
rect 18330 424 18364 458
rect 18398 424 18432 458
rect 18466 424 18500 458
rect 18534 424 18568 458
rect 18602 424 18636 458
rect 18670 424 18704 458
rect 18738 424 18772 458
rect 18806 424 18840 458
rect 18874 424 18908 458
rect 18942 424 18976 458
rect 19010 424 19044 458
rect 19078 424 19112 458
rect 19146 424 19180 458
rect 19214 424 19248 458
rect 19282 424 19316 458
rect 19350 424 19384 458
rect 19418 424 19452 458
rect 19486 424 19520 458
rect 19554 424 19588 458
rect 19622 424 19656 458
rect 19690 424 19724 458
rect 19758 424 19792 458
rect 19826 424 19860 458
rect 19894 424 19928 458
rect 19962 424 19996 458
rect 20030 424 20064 458
rect 20098 424 20132 458
rect 20166 424 20200 458
rect 20234 424 20268 458
rect 20302 424 20336 458
rect 20370 424 20404 458
rect 20438 424 20472 458
rect 20506 424 20540 458
rect 20574 424 20608 458
rect 20642 424 20676 458
rect 20710 424 20744 458
rect 20778 424 20812 458
rect 20846 424 20880 458
rect 20914 424 20948 458
rect 20982 424 21016 458
rect 21050 424 21084 458
rect 21118 424 21152 458
rect 21186 424 21220 458
rect 21254 424 21288 458
rect 21322 424 21356 458
rect 21390 424 21424 458
rect 21458 424 21492 458
rect 21526 424 21560 458
rect 21594 424 21628 458
rect 21662 424 21696 458
rect 21730 424 21764 458
rect 21798 424 21832 458
rect 21866 424 21900 458
rect 21934 424 21968 458
rect 22002 424 22036 458
rect 22070 424 22104 458
rect 22138 424 22172 458
rect 22206 424 22240 458
rect 22274 424 22308 458
rect 22342 424 22376 458
rect 22410 424 22444 458
rect 22478 424 22512 458
rect 22546 424 22580 458
rect 22614 424 22648 458
rect 22682 424 22716 458
rect 22750 424 22784 458
rect 22818 424 22852 458
rect 22886 424 22920 458
rect 22954 424 22988 458
rect 23022 424 23056 458
rect 23090 424 23124 458
rect 23158 424 23192 458
rect 23226 424 23260 458
rect 23294 424 23328 458
rect 23362 424 23396 458
rect 23430 424 23464 458
rect 23498 424 23532 458
rect 23566 424 23600 458
rect 23634 424 23668 458
rect 23702 424 23736 458
rect 23770 424 23804 458
rect 23838 424 23872 458
rect 23906 424 23940 458
rect 23974 424 24008 458
rect 24042 424 24076 458
rect 24110 424 24144 458
rect 24178 424 24212 458
rect 24246 424 24280 458
rect 24314 424 24348 458
rect 24382 424 24416 458
rect 24450 424 24484 458
rect 24518 424 24552 458
rect 24586 424 24620 458
rect 24654 424 24688 458
rect 24722 424 24756 458
rect 24790 424 24824 458
rect 24858 424 24892 458
rect 24926 424 24960 458
rect 24994 424 25028 458
rect 25062 424 25096 458
rect 25130 424 25164 458
rect 25198 424 25232 458
rect 25266 424 25300 458
rect 25334 424 25368 458
rect 25402 424 25436 458
rect 25470 424 25504 458
rect 25538 424 25572 458
rect 25606 424 25640 458
rect 25674 424 25708 458
rect 25742 424 25776 458
rect 25810 424 25844 458
rect 25878 424 25912 458
rect 25946 424 25980 458
rect 26014 424 26048 458
rect 26082 424 26116 458
rect 26150 424 26184 458
rect 26218 424 26252 458
rect 26286 424 26320 458
rect 26354 424 26388 458
rect 26422 424 26456 458
rect 26490 424 26524 458
rect 26558 424 26592 458
rect 26626 424 26660 458
rect 26694 424 26728 458
rect 26762 424 26796 458
rect 26830 424 26864 458
rect 26898 424 26932 458
rect 26966 424 27000 458
rect 27034 424 27068 458
rect 27102 424 27136 458
rect 27170 424 27204 458
rect 27238 424 27272 458
rect 27306 424 27340 458
rect 27374 424 27408 458
rect 27442 424 27476 458
rect 27510 424 27544 458
rect 27578 424 27612 458
rect 27646 424 27680 458
rect 27714 424 27748 458
rect 27782 424 27816 458
rect 27850 424 27884 458
rect 27918 424 27952 458
rect 27986 424 28020 458
rect 28054 424 28088 458
rect 28122 424 28156 458
rect 28190 424 28224 458
rect 28258 424 28292 458
rect 28326 424 28360 458
rect 28394 424 28428 458
rect 28462 424 28496 458
rect 28530 424 28564 458
rect 28598 424 28632 458
rect 28666 424 28700 458
rect 28734 424 28768 458
rect 28802 424 28836 458
rect 28870 424 28904 458
rect 28938 424 28972 458
rect 29006 424 29040 458
rect 29074 424 29108 458
rect 29142 424 29176 458
rect 29210 424 29244 458
rect 29278 424 29312 458
rect 29346 424 29380 458
rect 29414 424 29448 458
rect 29482 424 29516 458
rect 29550 424 29584 458
rect 29618 424 29652 458
rect 29686 424 29720 458
rect 29754 424 29788 458
rect 29822 424 29856 458
rect 29890 424 29924 458
rect 29958 424 29992 458
rect 30026 424 30060 458
rect 30094 424 30128 458
rect 30162 424 30196 458
rect 30230 424 30264 458
rect 30298 424 30332 458
rect 30366 424 30400 458
rect 30434 424 30468 458
rect 30502 424 30536 458
rect 30570 424 30604 458
rect 30638 424 30672 458
rect 30706 424 30740 458
rect 30774 424 30808 458
rect 30842 424 30876 458
rect 30910 424 30944 458
rect 30978 424 31012 458
rect 31046 424 31080 458
rect 31114 424 31148 458
rect 31182 424 31216 458
rect 31250 424 31284 458
rect 31318 424 31352 458
rect 31386 424 31420 458
rect 31454 424 31488 458
rect 31522 424 31556 458
rect 31590 424 31624 458
rect 31658 424 31692 458
rect 31726 424 31760 458
rect 31794 424 31828 458
rect 31862 424 31896 458
rect 31930 424 31964 458
rect 31998 424 32032 458
rect 32066 424 32100 458
rect 32134 424 32168 458
rect 32202 424 32236 458
rect 32270 424 32304 458
rect 32338 424 32372 458
rect 32406 424 32440 458
rect 32474 424 32508 458
rect 32542 424 32576 458
rect 32610 424 32644 458
rect 32678 424 32712 458
rect 32746 424 32780 458
rect 32814 424 32848 458
rect 32882 424 32916 458
rect 32950 424 32984 458
rect 33018 424 33052 458
rect 33086 424 33120 458
rect 33154 424 33188 458
rect 33222 424 33256 458
rect 33290 424 33324 458
rect 33358 424 33392 458
rect 33426 424 33460 458
rect 33494 424 33528 458
rect 33562 424 33596 458
rect 33630 424 33664 458
rect 33698 424 33732 458
rect 33766 424 33800 458
rect 33834 424 33868 458
rect 33902 424 33936 458
rect 33970 424 34004 458
rect 34038 424 34072 458
rect 34106 424 34140 458
rect 34174 424 34208 458
rect 34242 424 34276 458
rect 34310 424 34344 458
rect 34378 424 34412 458
rect 34446 424 34480 458
rect 34514 424 34548 458
rect 34582 424 34616 458
rect 34650 424 34684 458
rect 34718 424 34752 458
rect 34786 424 34820 458
rect 34854 424 34888 458
rect 34922 424 34956 458
rect 34990 424 35024 458
rect 35058 424 35092 458
rect 35126 424 35160 458
rect 35194 424 35228 458
rect 35262 424 35296 458
rect 35330 424 35364 458
rect 35398 424 35432 458
rect 35466 424 35500 458
rect 35534 424 35568 458
rect 35602 424 35636 458
rect 35670 424 35704 458
rect 35738 424 35772 458
rect 35806 424 35840 458
rect 35874 424 35908 458
rect 35942 424 35976 458
rect 36010 424 36044 458
rect 36078 424 36112 458
rect 36146 424 36180 458
rect 36214 424 36248 458
rect 36282 424 36316 458
rect 36350 424 36384 458
rect 36418 424 36452 458
rect 36486 424 36520 458
rect 36554 424 36588 458
rect 36622 424 36656 458
rect 36690 424 36724 458
rect 36758 424 36792 458
rect 36826 424 36860 458
rect 36894 424 36928 458
rect 36962 424 36996 458
rect 37030 424 37064 458
rect 37098 424 37132 458
rect 37166 424 37200 458
rect 37234 424 37268 458
rect 37302 424 37336 458
rect 37370 424 37404 458
rect 37438 424 37472 458
rect 37506 424 37540 458
rect 37574 424 37608 458
rect 37642 424 37676 458
rect 37710 424 37744 458
rect 37778 424 37812 458
rect 37846 424 37880 458
rect 37914 424 37948 458
rect 37982 424 38016 458
rect 38050 424 38084 458
rect 38118 424 38152 458
rect 38186 424 38220 458
rect 38254 424 38288 458
rect 38322 424 38356 458
rect 38390 424 38424 458
rect 38458 424 38492 458
rect 38526 424 38560 458
rect 38594 424 38628 458
rect 38662 424 38696 458
rect 38730 424 38764 458
rect 38798 424 38832 458
rect 38866 424 38900 458
rect 38934 424 38968 458
rect 39002 424 39036 458
rect 39070 424 39104 458
rect 39138 424 39172 458
rect 39206 424 39240 458
rect 39274 424 39308 458
rect 39342 424 39376 458
rect 39410 424 39444 458
rect 39478 424 39512 458
rect 39546 424 39580 458
rect 39614 424 39648 458
rect 39682 424 39716 458
rect 39750 424 39784 458
rect 39818 424 39852 458
rect 39886 424 39920 458
rect 39954 424 39988 458
rect 40022 424 40056 458
rect 40090 424 40124 458
rect 40158 424 40192 458
rect 40226 424 40260 458
rect 40294 424 40328 458
rect 40362 424 40396 458
rect 40430 424 40464 458
rect 40498 424 40532 458
rect 40566 424 40600 458
rect 40634 424 40668 458
rect 40702 424 40736 458
rect 40770 424 40804 458
rect 40838 424 40872 458
rect 40906 424 40940 458
rect 40974 424 41008 458
rect 41042 424 41076 458
rect 41110 424 41144 458
rect 41178 424 41212 458
rect 41246 424 41280 458
rect 41314 424 41348 458
rect 41382 424 41416 458
rect 41450 424 41484 458
rect 41518 424 41552 458
rect 41586 424 41620 458
rect 41654 424 41688 458
rect 41722 424 41756 458
rect 41790 424 41824 458
<< locali >>
rect 15694 15053 20241 15073
rect 15694 15019 15740 15053
rect 15774 15031 20241 15053
rect 15774 15019 15879 15031
rect 15694 14997 15879 15019
rect 15913 14997 15947 15031
rect 15981 14997 16015 15031
rect 16049 14997 16083 15031
rect 16117 14997 16151 15031
rect 16185 14997 16219 15031
rect 16253 14997 16287 15031
rect 16321 14997 16355 15031
rect 16389 14997 16423 15031
rect 16457 14997 16491 15031
rect 16525 14997 16559 15031
rect 16593 14997 16627 15031
rect 16661 14997 16695 15031
rect 16729 14997 16763 15031
rect 16797 14997 16831 15031
rect 16865 14997 16899 15031
rect 16933 14997 16967 15031
rect 17001 14997 17035 15031
rect 17069 14997 17103 15031
rect 17137 14997 17171 15031
rect 17205 14997 17239 15031
rect 17273 14997 17307 15031
rect 17341 14997 17375 15031
rect 17409 14997 17443 15031
rect 17477 14997 17511 15031
rect 17545 14997 17579 15031
rect 17613 14997 17647 15031
rect 17681 14997 17715 15031
rect 17749 14997 17783 15031
rect 17817 14997 17851 15031
rect 17885 14997 17919 15031
rect 17953 14997 17987 15031
rect 18021 14997 18055 15031
rect 18089 14997 18123 15031
rect 18157 14997 18191 15031
rect 18225 14997 18259 15031
rect 18293 14997 18327 15031
rect 18361 14997 18395 15031
rect 18429 14997 18463 15031
rect 18497 14997 18531 15031
rect 18565 14997 18599 15031
rect 18633 14997 18667 15031
rect 18701 14997 18735 15031
rect 18769 14997 18803 15031
rect 18837 14997 18871 15031
rect 18905 14997 18939 15031
rect 18973 14997 19007 15031
rect 19041 14997 19075 15031
rect 19109 14997 19143 15031
rect 19177 14997 19211 15031
rect 19245 14997 19279 15031
rect 19313 14997 19347 15031
rect 19381 14997 19415 15031
rect 19449 14997 19483 15031
rect 19517 14997 19551 15031
rect 19585 14997 19619 15031
rect 19653 14997 19687 15031
rect 19721 14997 19755 15031
rect 19789 14997 19823 15031
rect 19857 14997 19891 15031
rect 19925 14997 19959 15031
rect 19993 14997 20027 15031
rect 20061 15026 20241 15031
rect 20061 14997 20152 15026
rect 15694 14992 20152 14997
rect 20186 14992 20241 15026
rect 15694 14985 20241 14992
rect 15694 14951 15740 14985
rect 15774 14964 20241 14985
rect 15774 14951 15841 14964
rect 11930 14791 14414 14936
rect 11930 12377 12181 14791
rect 14187 12377 14414 14791
rect 15694 14917 15841 14951
rect 15694 14883 15740 14917
rect 15774 14883 15841 14917
rect 15694 14849 15841 14883
rect 15694 14815 15740 14849
rect 15774 14815 15841 14849
rect 15694 14781 15841 14815
rect 15694 14747 15740 14781
rect 15774 14747 15841 14781
rect 15694 14713 15841 14747
rect 15694 14679 15740 14713
rect 15774 14679 15841 14713
rect 15694 14645 15841 14679
rect 15694 14611 15740 14645
rect 15774 14611 15841 14645
rect 20095 14959 20241 14964
rect 20095 14954 20242 14959
rect 20095 14920 20152 14954
rect 20186 14920 20242 14954
rect 20095 14886 20242 14920
rect 20095 14852 20152 14886
rect 20186 14852 20242 14886
rect 20095 14818 20242 14852
rect 20095 14784 20152 14818
rect 20186 14784 20242 14818
rect 20095 14750 20242 14784
rect 20095 14716 20152 14750
rect 20186 14716 20242 14750
rect 20095 14682 20242 14716
rect 20095 14648 20152 14682
rect 20186 14648 20242 14682
rect 15694 14577 15841 14611
rect 15694 14543 15740 14577
rect 15774 14543 15841 14577
rect 15694 14509 15841 14543
rect 15694 14475 15740 14509
rect 15774 14475 15841 14509
rect 15694 14441 15841 14475
rect 15694 14407 15740 14441
rect 15774 14407 15841 14441
rect 15694 14373 15841 14407
rect 15694 14339 15740 14373
rect 15774 14339 15841 14373
rect 15694 14305 15841 14339
rect 15694 14271 15740 14305
rect 15774 14271 15841 14305
rect 15694 14237 15841 14271
rect 15694 14203 15740 14237
rect 15774 14203 15841 14237
rect 15694 14169 15841 14203
rect 15694 14135 15740 14169
rect 15774 14135 15841 14169
rect 15694 14101 15841 14135
rect 15694 14067 15740 14101
rect 15774 14067 15841 14101
rect 15694 14033 15841 14067
rect 15694 13999 15740 14033
rect 15774 13999 15841 14033
rect 15694 13965 15841 13999
rect 15694 13931 15740 13965
rect 15774 13931 15841 13965
rect 15694 13897 15841 13931
rect 15694 13863 15740 13897
rect 15774 13863 15841 13897
rect 15694 13829 15841 13863
rect 15694 13795 15740 13829
rect 15774 13795 15841 13829
rect 15694 13761 15841 13795
rect 15694 13727 15740 13761
rect 15774 13727 15841 13761
rect 15694 13693 15841 13727
rect 15694 13659 15740 13693
rect 15774 13659 15841 13693
rect 15694 13625 15841 13659
rect 15694 13591 15740 13625
rect 15774 13591 15841 13625
rect 15694 13557 15841 13591
rect 15694 13523 15740 13557
rect 15774 13523 15841 13557
rect 15694 13489 15841 13523
rect 15694 13455 15740 13489
rect 15774 13455 15841 13489
rect 15694 13421 15841 13455
rect 15694 13387 15740 13421
rect 15774 13387 15841 13421
rect 15694 13353 15841 13387
rect 15694 13319 15740 13353
rect 15774 13319 15841 13353
rect 15694 13285 15841 13319
rect 15694 13251 15740 13285
rect 15774 13251 15841 13285
rect 15694 13217 15841 13251
rect 15694 13183 15740 13217
rect 15774 13183 15841 13217
rect 15694 13149 15841 13183
rect 15694 13115 15740 13149
rect 15774 13115 15841 13149
rect 17468 14592 17615 14641
rect 17468 14558 17525 14592
rect 17559 14558 17615 14592
rect 17468 14524 17615 14558
rect 17468 14490 17525 14524
rect 17559 14490 17615 14524
rect 17468 14456 17615 14490
rect 17468 14422 17525 14456
rect 17559 14422 17615 14456
rect 17468 14388 17615 14422
rect 17468 14354 17525 14388
rect 17559 14354 17615 14388
rect 17468 14320 17615 14354
rect 17468 14286 17525 14320
rect 17559 14286 17615 14320
rect 17468 14166 17615 14286
rect 17468 14132 17525 14166
rect 17559 14132 17615 14166
rect 17468 14098 17615 14132
rect 17468 14064 17525 14098
rect 17559 14064 17615 14098
rect 17468 14030 17615 14064
rect 17468 13996 17525 14030
rect 17559 13996 17615 14030
rect 17468 13962 17615 13996
rect 17468 13928 17525 13962
rect 17559 13928 17615 13962
rect 17468 13894 17615 13928
rect 17468 13860 17525 13894
rect 17559 13860 17615 13894
rect 17468 13826 17615 13860
rect 17468 13792 17525 13826
rect 17559 13792 17615 13826
rect 17468 13758 17615 13792
rect 17468 13724 17525 13758
rect 17559 13724 17615 13758
rect 17468 13690 17615 13724
rect 17468 13656 17525 13690
rect 17559 13656 17615 13690
rect 17468 13622 17615 13656
rect 17468 13588 17525 13622
rect 17559 13588 17615 13622
rect 17468 13554 17615 13588
rect 17468 13520 17525 13554
rect 17559 13520 17615 13554
rect 17468 13486 17615 13520
rect 17468 13452 17525 13486
rect 17559 13452 17615 13486
rect 17468 13418 17615 13452
rect 17468 13384 17525 13418
rect 17559 13384 17615 13418
rect 17468 13350 17615 13384
rect 17468 13316 17525 13350
rect 17559 13316 17615 13350
rect 17468 13282 17615 13316
rect 17468 13248 17525 13282
rect 17559 13248 17615 13282
rect 17468 13214 17615 13248
rect 17468 13180 17525 13214
rect 17559 13180 17615 13214
rect 17468 13136 17615 13180
rect 19247 14579 19391 14635
rect 19247 14545 19304 14579
rect 19338 14545 19391 14579
rect 19247 14511 19391 14545
rect 19247 14477 19304 14511
rect 19338 14477 19391 14511
rect 19247 14443 19391 14477
rect 19247 14409 19304 14443
rect 19338 14409 19391 14443
rect 19247 14375 19391 14409
rect 19247 14341 19304 14375
rect 19338 14341 19391 14375
rect 19247 14307 19391 14341
rect 19247 14273 19304 14307
rect 19338 14273 19391 14307
rect 19247 14239 19391 14273
rect 19247 14205 19304 14239
rect 19338 14205 19391 14239
rect 19247 14171 19391 14205
rect 19247 14137 19304 14171
rect 19338 14137 19391 14171
rect 19247 14103 19391 14137
rect 19247 14069 19304 14103
rect 19338 14069 19391 14103
rect 19247 14035 19391 14069
rect 19247 14001 19304 14035
rect 19338 14001 19391 14035
rect 19247 13967 19391 14001
rect 19247 13933 19304 13967
rect 19338 13933 19391 13967
rect 19247 13899 19391 13933
rect 19247 13865 19304 13899
rect 19338 13865 19391 13899
rect 19247 13831 19391 13865
rect 19247 13797 19304 13831
rect 19338 13797 19391 13831
rect 19247 13763 19391 13797
rect 19247 13729 19304 13763
rect 19338 13729 19391 13763
rect 19247 13695 19391 13729
rect 19247 13661 19304 13695
rect 19338 13661 19391 13695
rect 19247 13627 19391 13661
rect 19247 13593 19304 13627
rect 19338 13593 19391 13627
rect 19247 13559 19391 13593
rect 19247 13525 19304 13559
rect 19338 13525 19391 13559
rect 19247 13491 19391 13525
rect 19247 13457 19304 13491
rect 19338 13457 19391 13491
rect 19247 13423 19391 13457
rect 19247 13389 19304 13423
rect 19338 13389 19391 13423
rect 19247 13355 19391 13389
rect 19247 13321 19304 13355
rect 19338 13321 19391 13355
rect 19247 13287 19391 13321
rect 19247 13253 19304 13287
rect 19338 13253 19391 13287
rect 19247 13219 19391 13253
rect 19247 13185 19304 13219
rect 19338 13185 19391 13219
rect 19247 13139 19391 13185
rect 20095 14614 20242 14648
rect 20095 14580 20152 14614
rect 20186 14580 20242 14614
rect 20095 14546 20242 14580
rect 20095 14512 20152 14546
rect 20186 14512 20242 14546
rect 20095 14478 20242 14512
rect 20095 14444 20152 14478
rect 20186 14444 20242 14478
rect 20095 14402 20242 14444
rect 20095 14341 20241 14402
rect 20095 14307 20152 14341
rect 20186 14307 20241 14341
rect 20095 14273 20241 14307
rect 20095 14239 20152 14273
rect 20186 14239 20241 14273
rect 20095 14205 20241 14239
rect 20095 14171 20152 14205
rect 20186 14171 20241 14205
rect 20095 14137 20241 14171
rect 20095 14103 20152 14137
rect 20186 14103 20241 14137
rect 20095 14069 20241 14103
rect 20095 14035 20152 14069
rect 20186 14035 20241 14069
rect 20095 14001 20241 14035
rect 20095 13967 20152 14001
rect 20186 13967 20241 14001
rect 20095 13933 20241 13967
rect 20095 13899 20152 13933
rect 20186 13899 20241 13933
rect 20095 13865 20241 13899
rect 20095 13831 20152 13865
rect 20186 13831 20241 13865
rect 20095 13797 20241 13831
rect 20095 13763 20152 13797
rect 20186 13763 20241 13797
rect 20095 13729 20241 13763
rect 20095 13695 20152 13729
rect 20186 13695 20241 13729
rect 20095 13661 20241 13695
rect 20095 13627 20152 13661
rect 20186 13627 20241 13661
rect 20095 13593 20241 13627
rect 20095 13559 20152 13593
rect 20186 13559 20241 13593
rect 20095 13525 20241 13559
rect 20095 13491 20152 13525
rect 20186 13491 20241 13525
rect 20095 13457 20241 13491
rect 20095 13423 20152 13457
rect 20186 13423 20241 13457
rect 20095 13389 20241 13423
rect 20095 13355 20152 13389
rect 20186 13355 20241 13389
rect 20095 13321 20241 13355
rect 20095 13287 20152 13321
rect 20186 13287 20241 13321
rect 20095 13253 20241 13287
rect 20095 13219 20152 13253
rect 20186 13219 20241 13253
rect 20095 13185 20241 13219
rect 20095 13151 20152 13185
rect 20186 13151 20241 13185
rect 15694 13081 15841 13115
rect 15694 13047 15740 13081
rect 15774 13047 15841 13081
rect 15694 13013 15841 13047
rect 15694 12979 15740 13013
rect 15774 12979 15841 13013
rect 15694 12973 15841 12979
rect 20095 13117 20241 13151
rect 20095 13083 20152 13117
rect 20186 13083 20241 13117
rect 20095 13049 20241 13083
rect 20095 13015 20152 13049
rect 20186 13015 20241 13049
rect 20095 12973 20241 13015
rect 15694 12945 20241 12973
rect 15694 12843 15740 12945
rect 20194 12843 20241 12945
rect 15694 12821 20241 12843
rect 11930 12218 14414 12377
rect 15700 11941 20246 11971
rect 15700 11907 15746 11941
rect 15780 11907 15814 11941
rect 15848 11907 15882 11941
rect 15916 11907 15950 11941
rect 15984 11907 16018 11941
rect 16052 11907 16086 11941
rect 16120 11907 16154 11941
rect 16188 11907 16222 11941
rect 16256 11907 16290 11941
rect 16324 11907 16358 11941
rect 16392 11907 16426 11941
rect 16460 11907 16494 11941
rect 16528 11907 16562 11941
rect 16596 11907 16630 11941
rect 16664 11907 16698 11941
rect 16732 11907 16766 11941
rect 16800 11907 16834 11941
rect 16868 11907 16902 11941
rect 16936 11907 16970 11941
rect 17004 11907 17038 11941
rect 17072 11907 17106 11941
rect 17140 11907 17174 11941
rect 17208 11907 17242 11941
rect 17276 11907 17310 11941
rect 17344 11907 17378 11941
rect 17412 11907 17446 11941
rect 17480 11907 17514 11941
rect 17548 11907 17582 11941
rect 17616 11907 17650 11941
rect 17684 11907 17718 11941
rect 17752 11907 17786 11941
rect 17820 11907 17854 11941
rect 17888 11907 17922 11941
rect 17956 11907 17990 11941
rect 18024 11907 18058 11941
rect 18092 11907 18126 11941
rect 18160 11907 18194 11941
rect 18228 11907 18262 11941
rect 18296 11907 18330 11941
rect 18364 11907 18398 11941
rect 18432 11907 18466 11941
rect 18500 11907 18534 11941
rect 18568 11907 18602 11941
rect 18636 11907 18670 11941
rect 18704 11907 18738 11941
rect 18772 11907 18806 11941
rect 18840 11907 18874 11941
rect 18908 11907 18942 11941
rect 18976 11907 19010 11941
rect 19044 11907 19078 11941
rect 19112 11907 19146 11941
rect 19180 11907 19214 11941
rect 19248 11907 19282 11941
rect 19316 11907 19350 11941
rect 19384 11907 19418 11941
rect 19452 11907 19486 11941
rect 19520 11907 19554 11941
rect 19588 11907 19622 11941
rect 19656 11907 19690 11941
rect 19724 11907 19758 11941
rect 19792 11907 19826 11941
rect 19860 11907 19894 11941
rect 19928 11907 19962 11941
rect 19996 11907 20030 11941
rect 20064 11907 20098 11941
rect 20132 11907 20166 11941
rect 20200 11907 20246 11941
rect 15700 11873 20246 11907
rect 15700 11839 15746 11873
rect 15780 11839 20166 11873
rect 20200 11839 20246 11873
rect 15700 11822 20246 11839
rect 15700 11805 15838 11822
rect 15700 11771 15746 11805
rect 15780 11771 15838 11805
rect 15700 11737 15838 11771
rect 15700 11703 15746 11737
rect 15780 11703 15838 11737
rect 15700 11669 15838 11703
rect 15700 11635 15746 11669
rect 15780 11635 15838 11669
rect 15700 11601 15838 11635
rect 15700 11567 15746 11601
rect 15780 11567 15838 11601
rect 15700 11533 15838 11567
rect 15700 11499 15746 11533
rect 15780 11499 15838 11533
rect 15700 11465 15838 11499
rect 15700 11431 15746 11465
rect 15780 11431 15838 11465
rect 15700 11397 15838 11431
rect 15700 11363 15746 11397
rect 15780 11363 15838 11397
rect 15700 11329 15838 11363
rect 15700 11295 15746 11329
rect 15780 11295 15838 11329
rect 15700 11261 15838 11295
rect 15700 11227 15746 11261
rect 15780 11227 15838 11261
rect 15700 11193 15838 11227
rect 10755 11151 11235 11172
rect 10755 11117 10789 11151
rect 10823 11117 10876 11151
rect 10910 11117 10944 11151
rect 10978 11117 11012 11151
rect 11046 11117 11080 11151
rect 11114 11117 11168 11151
rect 11202 11117 11235 11151
rect 10755 11096 11235 11117
rect 10755 11084 10856 11096
rect 10755 11042 10789 11084
rect 10823 11042 10856 11084
rect 10755 11012 10856 11042
rect 10755 10974 10789 11012
rect 10823 10974 10856 11012
rect 10755 10940 10856 10974
rect 10755 10906 10789 10940
rect 10823 10906 10856 10940
rect 10755 10872 10856 10906
rect 10755 10834 10789 10872
rect 10823 10834 10856 10872
rect 10755 10804 10856 10834
rect 10755 10762 10789 10804
rect 10823 10762 10856 10804
rect 10755 10750 10856 10762
rect 11134 11076 11235 11096
rect 11134 11042 11168 11076
rect 11202 11042 11235 11076
rect 11134 11008 11235 11042
rect 11134 10974 11168 11008
rect 11202 10974 11235 11008
rect 11134 10954 11235 10974
rect 15700 11159 15746 11193
rect 15780 11159 15838 11193
rect 15700 11125 15838 11159
rect 15700 11091 15746 11125
rect 15780 11091 15838 11125
rect 15700 11057 15838 11091
rect 15700 11023 15746 11057
rect 15780 11023 15838 11057
rect 15700 10989 15838 11023
rect 15700 10955 15746 10989
rect 15780 10955 15838 10989
rect 11134 10940 11236 10954
rect 11134 10906 11168 10940
rect 11202 10906 11236 10940
rect 11134 10874 11236 10906
rect 15700 10950 15838 10955
rect 20106 11805 20246 11822
rect 20106 11771 20166 11805
rect 20200 11771 20246 11805
rect 20106 11737 20246 11771
rect 20106 11703 20166 11737
rect 20200 11703 20246 11737
rect 20106 11669 20246 11703
rect 20106 11635 20166 11669
rect 20200 11635 20246 11669
rect 20106 11601 20246 11635
rect 20106 11567 20166 11601
rect 20200 11567 20246 11601
rect 20106 11533 20246 11567
rect 20106 11499 20166 11533
rect 20200 11499 20246 11533
rect 20106 11465 20246 11499
rect 20106 11431 20166 11465
rect 20200 11431 20246 11465
rect 20106 11397 20246 11431
rect 20106 11363 20166 11397
rect 20200 11363 20246 11397
rect 20106 11329 20246 11363
rect 20106 11295 20166 11329
rect 20200 11295 20246 11329
rect 20106 11261 20246 11295
rect 20106 11227 20166 11261
rect 20200 11227 20246 11261
rect 20106 11193 20246 11227
rect 20106 11159 20166 11193
rect 20200 11159 20246 11193
rect 20106 11125 20246 11159
rect 20106 11091 20166 11125
rect 20200 11091 20246 11125
rect 20106 11057 20246 11091
rect 20106 11023 20166 11057
rect 20200 11023 20246 11057
rect 20106 10989 20246 11023
rect 20106 10955 20166 10989
rect 20200 10955 20246 10989
rect 20106 10950 20246 10955
rect 15700 10921 20246 10950
rect 11134 10872 11235 10874
rect 11134 10838 11168 10872
rect 11202 10838 11235 10872
rect 11134 10804 11235 10838
rect 11134 10770 11168 10804
rect 11202 10770 11235 10804
rect 15700 10819 15746 10921
rect 20200 10819 20246 10921
rect 15700 10791 20246 10819
rect 11134 10750 11235 10770
rect 10755 10728 11235 10750
rect 10755 10694 10789 10728
rect 10823 10694 10876 10728
rect 10910 10694 10944 10728
rect 10978 10694 11012 10728
rect 11046 10694 11080 10728
rect 11114 10694 11168 10728
rect 11202 10694 11235 10728
rect 10755 10671 11235 10694
rect 5615 10619 10162 10639
rect 5615 10597 10082 10619
rect 5615 10592 5794 10597
rect 5615 10558 5670 10592
rect 5704 10563 5794 10592
rect 5828 10563 5862 10597
rect 5896 10563 5930 10597
rect 5964 10563 5998 10597
rect 6032 10563 6066 10597
rect 6100 10563 6134 10597
rect 6168 10563 6202 10597
rect 6236 10563 6270 10597
rect 6304 10563 6338 10597
rect 6372 10563 6406 10597
rect 6440 10563 6474 10597
rect 6508 10563 6542 10597
rect 6576 10563 6610 10597
rect 6644 10563 6678 10597
rect 6712 10563 6746 10597
rect 6780 10563 6814 10597
rect 6848 10563 6882 10597
rect 6916 10563 6950 10597
rect 6984 10563 7018 10597
rect 7052 10563 7086 10597
rect 7120 10563 7154 10597
rect 7188 10563 7222 10597
rect 7256 10563 7290 10597
rect 7324 10563 7358 10597
rect 7392 10563 7426 10597
rect 7460 10563 7494 10597
rect 7528 10563 7562 10597
rect 7596 10563 7630 10597
rect 7664 10563 7698 10597
rect 7732 10563 7766 10597
rect 7800 10563 7834 10597
rect 7868 10563 7902 10597
rect 7936 10563 7970 10597
rect 8004 10563 8038 10597
rect 8072 10563 8106 10597
rect 8140 10563 8174 10597
rect 8208 10563 8242 10597
rect 8276 10563 8310 10597
rect 8344 10563 8378 10597
rect 8412 10563 8446 10597
rect 8480 10563 8514 10597
rect 8548 10563 8582 10597
rect 8616 10563 8650 10597
rect 8684 10563 8718 10597
rect 8752 10563 8786 10597
rect 8820 10563 8854 10597
rect 8888 10563 8922 10597
rect 8956 10563 8990 10597
rect 9024 10563 9058 10597
rect 9092 10563 9126 10597
rect 9160 10563 9194 10597
rect 9228 10563 9262 10597
rect 9296 10563 9330 10597
rect 9364 10563 9398 10597
rect 9432 10563 9466 10597
rect 9500 10563 9534 10597
rect 9568 10563 9602 10597
rect 9636 10563 9670 10597
rect 9704 10563 9738 10597
rect 9772 10563 9806 10597
rect 9840 10563 9874 10597
rect 9908 10563 9942 10597
rect 9976 10585 10082 10597
rect 10116 10585 10162 10619
rect 9976 10563 10162 10585
rect 5704 10558 10162 10563
rect 5615 10551 10162 10558
rect 5615 10530 10082 10551
rect 5615 10525 5761 10530
rect 5614 10486 5761 10525
rect 5614 10452 5669 10486
rect 5703 10452 5761 10486
rect 5614 10418 5761 10452
rect 5614 10384 5669 10418
rect 5703 10384 5761 10418
rect 5614 10350 5761 10384
rect 5614 10316 5669 10350
rect 5703 10316 5761 10350
rect 5614 10282 5761 10316
rect 5614 10248 5669 10282
rect 5703 10248 5761 10282
rect 5614 10214 5761 10248
rect 5614 10180 5669 10214
rect 5703 10180 5761 10214
rect 10015 10517 10082 10530
rect 10116 10517 10162 10551
rect 10015 10483 10162 10517
rect 10015 10449 10082 10483
rect 10116 10449 10162 10483
rect 10741 10533 11253 10553
rect 10741 10499 10776 10533
rect 10810 10499 10879 10533
rect 10913 10499 10947 10533
rect 10981 10499 11015 10533
rect 11049 10499 11083 10533
rect 11117 10499 11187 10533
rect 11221 10499 11253 10533
rect 10741 10476 11253 10499
rect 10015 10415 10162 10449
rect 10015 10381 10082 10415
rect 10116 10381 10162 10415
rect 10015 10347 10162 10381
rect 10015 10313 10082 10347
rect 10116 10313 10162 10347
rect 10015 10279 10162 10313
rect 10015 10245 10082 10279
rect 10116 10245 10162 10279
rect 10015 10211 10162 10245
rect 5614 10146 5761 10180
rect 5614 10112 5669 10146
rect 5703 10112 5761 10146
rect 5614 10078 5761 10112
rect 5614 10044 5669 10078
rect 5703 10044 5761 10078
rect 5614 10010 5761 10044
rect 5614 9976 5669 10010
rect 5703 9976 5761 10010
rect 5614 9968 5761 9976
rect 5615 9907 5761 9968
rect 5615 9873 5670 9907
rect 5704 9873 5761 9907
rect 5615 9839 5761 9873
rect 5615 9805 5670 9839
rect 5704 9805 5761 9839
rect 5615 9771 5761 9805
rect 5615 9737 5670 9771
rect 5704 9737 5761 9771
rect 5615 9703 5761 9737
rect 5615 9669 5670 9703
rect 5704 9669 5761 9703
rect 5615 9635 5761 9669
rect 5615 9601 5670 9635
rect 5704 9601 5761 9635
rect 5615 9567 5761 9601
rect 5615 9533 5670 9567
rect 5704 9533 5761 9567
rect 5615 9499 5761 9533
rect 5615 9465 5670 9499
rect 5704 9465 5761 9499
rect 5615 9431 5761 9465
rect 5615 9397 5670 9431
rect 5704 9397 5761 9431
rect 5615 9363 5761 9397
rect 5615 9329 5670 9363
rect 5704 9329 5761 9363
rect 5615 9295 5761 9329
rect 5615 9261 5670 9295
rect 5704 9261 5761 9295
rect 5615 9227 5761 9261
rect 5615 9193 5670 9227
rect 5704 9193 5761 9227
rect 5615 9159 5761 9193
rect 5615 9125 5670 9159
rect 5704 9125 5761 9159
rect 5615 9091 5761 9125
rect 5615 9057 5670 9091
rect 5704 9057 5761 9091
rect 5615 9023 5761 9057
rect 5615 8989 5670 9023
rect 5704 8989 5761 9023
rect 5615 8955 5761 8989
rect 5615 8921 5670 8955
rect 5704 8921 5761 8955
rect 5615 8887 5761 8921
rect 5615 8853 5670 8887
rect 5704 8853 5761 8887
rect 5615 8819 5761 8853
rect 5615 8785 5670 8819
rect 5704 8785 5761 8819
rect 5615 8751 5761 8785
rect 5615 8717 5670 8751
rect 5704 8717 5761 8751
rect 5615 8683 5761 8717
rect 6465 10145 6609 10201
rect 6465 10111 6518 10145
rect 6552 10111 6609 10145
rect 6465 10077 6609 10111
rect 6465 10043 6518 10077
rect 6552 10043 6609 10077
rect 6465 10009 6609 10043
rect 6465 9975 6518 10009
rect 6552 9975 6609 10009
rect 6465 9941 6609 9975
rect 6465 9907 6518 9941
rect 6552 9907 6609 9941
rect 6465 9873 6609 9907
rect 6465 9839 6518 9873
rect 6552 9839 6609 9873
rect 6465 9805 6609 9839
rect 6465 9771 6518 9805
rect 6552 9771 6609 9805
rect 6465 9737 6609 9771
rect 6465 9703 6518 9737
rect 6552 9703 6609 9737
rect 6465 9669 6609 9703
rect 6465 9635 6518 9669
rect 6552 9635 6609 9669
rect 6465 9601 6609 9635
rect 6465 9567 6518 9601
rect 6552 9567 6609 9601
rect 6465 9533 6609 9567
rect 6465 9499 6518 9533
rect 6552 9499 6609 9533
rect 6465 9465 6609 9499
rect 6465 9431 6518 9465
rect 6552 9431 6609 9465
rect 6465 9397 6609 9431
rect 6465 9363 6518 9397
rect 6552 9363 6609 9397
rect 6465 9329 6609 9363
rect 6465 9295 6518 9329
rect 6552 9295 6609 9329
rect 6465 9261 6609 9295
rect 6465 9227 6518 9261
rect 6552 9227 6609 9261
rect 6465 9193 6609 9227
rect 6465 9159 6518 9193
rect 6552 9159 6609 9193
rect 6465 9125 6609 9159
rect 6465 9091 6518 9125
rect 6552 9091 6609 9125
rect 6465 9057 6609 9091
rect 6465 9023 6518 9057
rect 6552 9023 6609 9057
rect 6465 8989 6609 9023
rect 6465 8955 6518 8989
rect 6552 8955 6609 8989
rect 6465 8921 6609 8955
rect 6465 8887 6518 8921
rect 6552 8887 6609 8921
rect 6465 8853 6609 8887
rect 6465 8819 6518 8853
rect 6552 8819 6609 8853
rect 6465 8785 6609 8819
rect 6465 8751 6518 8785
rect 6552 8751 6609 8785
rect 6465 8705 6609 8751
rect 8241 10175 8388 10207
rect 8241 10141 8296 10175
rect 8330 10141 8388 10175
rect 8241 10107 8388 10141
rect 8241 10073 8296 10107
rect 8330 10073 8388 10107
rect 8241 10039 8388 10073
rect 8241 10005 8296 10039
rect 8330 10005 8388 10039
rect 8241 9971 8388 10005
rect 8241 9937 8296 9971
rect 8330 9937 8388 9971
rect 8241 9903 8388 9937
rect 8241 9869 8296 9903
rect 8330 9869 8388 9903
rect 8241 9835 8388 9869
rect 8241 9801 8296 9835
rect 8330 9801 8388 9835
rect 8241 9732 8388 9801
rect 8241 9698 8297 9732
rect 8331 9698 8388 9732
rect 8241 9664 8388 9698
rect 8241 9630 8297 9664
rect 8331 9630 8388 9664
rect 8241 9596 8388 9630
rect 8241 9562 8297 9596
rect 8331 9562 8388 9596
rect 8241 9528 8388 9562
rect 8241 9494 8297 9528
rect 8331 9494 8388 9528
rect 8241 9460 8388 9494
rect 8241 9426 8297 9460
rect 8331 9426 8388 9460
rect 8241 9392 8388 9426
rect 8241 9358 8297 9392
rect 8331 9358 8388 9392
rect 8241 9324 8388 9358
rect 8241 9290 8297 9324
rect 8331 9290 8388 9324
rect 8241 9256 8388 9290
rect 8241 9222 8297 9256
rect 8331 9222 8388 9256
rect 8241 9188 8388 9222
rect 8241 9154 8297 9188
rect 8331 9154 8388 9188
rect 8241 9120 8388 9154
rect 8241 9086 8297 9120
rect 8331 9086 8388 9120
rect 8241 9052 8388 9086
rect 8241 9018 8297 9052
rect 8331 9018 8388 9052
rect 8241 8984 8388 9018
rect 8241 8950 8297 8984
rect 8331 8950 8388 8984
rect 8241 8916 8388 8950
rect 8241 8882 8297 8916
rect 8331 8882 8388 8916
rect 8241 8848 8388 8882
rect 8241 8814 8297 8848
rect 8331 8814 8388 8848
rect 8241 8780 8388 8814
rect 8241 8746 8297 8780
rect 8331 8746 8388 8780
rect 8241 8702 8388 8746
rect 10015 10177 10082 10211
rect 10116 10177 10162 10211
rect 10015 10143 10162 10177
rect 10015 10109 10082 10143
rect 10116 10109 10162 10143
rect 10015 10075 10162 10109
rect 10015 10041 10082 10075
rect 10116 10041 10162 10075
rect 10015 10007 10162 10041
rect 10015 9973 10082 10007
rect 10116 9973 10162 10007
rect 10015 9939 10162 9973
rect 10015 9905 10082 9939
rect 10116 9905 10162 9939
rect 10015 9871 10162 9905
rect 10015 9837 10082 9871
rect 10116 9837 10162 9871
rect 10015 9803 10162 9837
rect 10015 9769 10082 9803
rect 10116 9769 10162 9803
rect 10015 9735 10162 9769
rect 10015 9701 10082 9735
rect 10116 9701 10162 9735
rect 10015 9667 10162 9701
rect 10015 9633 10082 9667
rect 10116 9633 10162 9667
rect 10015 9599 10162 9633
rect 10015 9565 10082 9599
rect 10116 9565 10162 9599
rect 10015 9531 10162 9565
rect 10015 9497 10082 9531
rect 10116 9497 10162 9531
rect 10015 9463 10162 9497
rect 10015 9429 10082 9463
rect 10116 9429 10162 9463
rect 10015 9395 10162 9429
rect 10015 9361 10082 9395
rect 10116 9361 10162 9395
rect 10015 9327 10162 9361
rect 10015 9293 10082 9327
rect 10116 9293 10162 9327
rect 10015 9259 10162 9293
rect 10015 9225 10082 9259
rect 10116 9225 10162 9259
rect 10015 9191 10162 9225
rect 10015 9157 10082 9191
rect 10116 9157 10162 9191
rect 10015 9123 10162 9157
rect 10015 9089 10082 9123
rect 10116 9089 10162 9123
rect 10015 9055 10162 9089
rect 10015 9021 10082 9055
rect 10116 9021 10162 9055
rect 10015 8987 10162 9021
rect 10015 8953 10082 8987
rect 10116 8953 10162 8987
rect 10015 8919 10162 8953
rect 10015 8885 10082 8919
rect 10116 8885 10162 8919
rect 10015 8851 10162 8885
rect 10015 8817 10082 8851
rect 10116 8817 10162 8851
rect 10015 8783 10162 8817
rect 10015 8749 10082 8783
rect 10116 8749 10162 8783
rect 10015 8715 10162 8749
rect 5615 8649 5670 8683
rect 5704 8649 5761 8683
rect 5615 8615 5761 8649
rect 5615 8581 5670 8615
rect 5704 8581 5761 8615
rect 5615 8542 5761 8581
rect 5615 8511 5664 8542
rect 5698 8539 5761 8542
rect 10015 8681 10082 8715
rect 10116 8681 10162 8715
rect 10015 8647 10162 8681
rect 10015 8613 10082 8647
rect 10116 8613 10162 8647
rect 10015 8579 10162 8613
rect 10015 8545 10082 8579
rect 10116 8545 10162 8579
rect 10747 10448 10833 10476
rect 10747 10414 10776 10448
rect 10810 10414 10833 10448
rect 10747 10380 10833 10414
rect 10747 10346 10776 10380
rect 10810 10346 10833 10380
rect 10747 10312 10833 10346
rect 10747 10278 10776 10312
rect 10810 10278 10833 10312
rect 10747 10244 10833 10278
rect 10747 10210 10776 10244
rect 10810 10210 10833 10244
rect 10747 10176 10833 10210
rect 10747 10142 10776 10176
rect 10810 10142 10833 10176
rect 10747 10108 10833 10142
rect 10747 10074 10776 10108
rect 10810 10074 10833 10108
rect 10747 10040 10833 10074
rect 10747 10006 10776 10040
rect 10810 10006 10833 10040
rect 10747 9972 10833 10006
rect 10747 9938 10776 9972
rect 10810 9938 10833 9972
rect 10747 9904 10833 9938
rect 10747 9870 10776 9904
rect 10810 9870 10833 9904
rect 10747 9836 10833 9870
rect 10747 9802 10776 9836
rect 10810 9802 10833 9836
rect 10747 9768 10833 9802
rect 10747 9734 10776 9768
rect 10810 9734 10833 9768
rect 10747 9700 10833 9734
rect 10747 9666 10776 9700
rect 10810 9666 10833 9700
rect 10747 9632 10833 9666
rect 10747 9598 10776 9632
rect 10810 9598 10833 9632
rect 10747 9564 10833 9598
rect 10747 9530 10776 9564
rect 10810 9530 10833 9564
rect 10747 9496 10833 9530
rect 10747 9462 10776 9496
rect 10810 9462 10833 9496
rect 10747 9428 10833 9462
rect 10747 9394 10776 9428
rect 10810 9394 10833 9428
rect 10747 9360 10833 9394
rect 10747 9326 10776 9360
rect 10810 9326 10833 9360
rect 10747 9292 10833 9326
rect 10747 9258 10776 9292
rect 10810 9258 10833 9292
rect 10747 9224 10833 9258
rect 10747 9190 10776 9224
rect 10810 9190 10833 9224
rect 10747 9156 10833 9190
rect 10747 9122 10776 9156
rect 10810 9122 10833 9156
rect 10747 9088 10833 9122
rect 10747 9054 10776 9088
rect 10810 9054 10833 9088
rect 10747 9020 10833 9054
rect 10747 8986 10776 9020
rect 10810 8986 10833 9020
rect 10747 8952 10833 8986
rect 10747 8918 10776 8952
rect 10810 8918 10833 8952
rect 10747 8884 10833 8918
rect 10747 8850 10776 8884
rect 10810 8850 10833 8884
rect 10747 8816 10833 8850
rect 10747 8782 10776 8816
rect 10810 8782 10833 8816
rect 10747 8748 10833 8782
rect 10747 8714 10776 8748
rect 10810 8714 10833 8748
rect 10747 8680 10833 8714
rect 10747 8646 10776 8680
rect 10810 8646 10833 8680
rect 10747 8616 10833 8646
rect 11158 10448 11253 10476
rect 11158 10414 11187 10448
rect 11221 10414 11253 10448
rect 11158 10380 11253 10414
rect 11158 10346 11187 10380
rect 11221 10346 11253 10380
rect 11158 10312 11253 10346
rect 11158 10278 11187 10312
rect 11221 10278 11253 10312
rect 11158 10244 11253 10278
rect 11158 10210 11187 10244
rect 11221 10210 11253 10244
rect 11158 10176 11253 10210
rect 11158 10142 11187 10176
rect 11221 10142 11253 10176
rect 11158 10108 11253 10142
rect 11158 10074 11187 10108
rect 11221 10074 11253 10108
rect 11158 10040 11253 10074
rect 11158 10006 11187 10040
rect 11221 10006 11253 10040
rect 11158 9972 11253 10006
rect 11158 9938 11187 9972
rect 11221 9938 11253 9972
rect 11158 9904 11253 9938
rect 11158 9870 11187 9904
rect 11221 9870 11253 9904
rect 11158 9836 11253 9870
rect 11158 9802 11187 9836
rect 11221 9802 11253 9836
rect 11158 9768 11253 9802
rect 11158 9734 11187 9768
rect 11221 9734 11253 9768
rect 11158 9700 11253 9734
rect 11158 9666 11187 9700
rect 11221 9666 11253 9700
rect 11158 9632 11253 9666
rect 11158 9598 11187 9632
rect 11221 9598 11253 9632
rect 11158 9564 11253 9598
rect 11158 9530 11187 9564
rect 11221 9530 11253 9564
rect 11158 9496 11253 9530
rect 11158 9462 11187 9496
rect 11221 9462 11253 9496
rect 11158 9428 11253 9462
rect 16361 9877 16965 9896
rect 16361 9843 16395 9877
rect 16429 9843 16509 9877
rect 16543 9843 16577 9877
rect 16611 9843 16645 9877
rect 16679 9843 16713 9877
rect 16747 9843 16781 9877
rect 16815 9843 16895 9877
rect 16929 9843 16965 9877
rect 16361 9830 16965 9843
rect 16361 9793 16465 9830
rect 16361 9759 16395 9793
rect 16429 9759 16465 9793
rect 16361 9725 16465 9759
rect 16361 9691 16395 9725
rect 16429 9691 16465 9725
rect 16361 9657 16465 9691
rect 16361 9623 16395 9657
rect 16429 9623 16465 9657
rect 16361 9589 16465 9623
rect 16361 9555 16395 9589
rect 16429 9555 16465 9589
rect 16361 9516 16465 9555
rect 16859 9793 16965 9830
rect 16859 9759 16895 9793
rect 16929 9759 16965 9793
rect 16859 9725 16965 9759
rect 16859 9676 16895 9725
rect 16929 9676 16965 9725
rect 16859 9657 16965 9676
rect 16859 9604 16895 9657
rect 16929 9604 16965 9657
rect 16859 9589 16965 9604
rect 16859 9555 16895 9589
rect 16929 9555 16965 9589
rect 16859 9516 16965 9555
rect 16361 9501 16965 9516
rect 16361 9467 16395 9501
rect 16429 9467 16509 9501
rect 16543 9467 16577 9501
rect 16611 9467 16645 9501
rect 16679 9467 16713 9501
rect 16747 9467 16781 9501
rect 16815 9467 16895 9501
rect 16929 9467 16965 9501
rect 16361 9449 16965 9467
rect 19828 9873 20432 9892
rect 19828 9839 19862 9873
rect 19896 9839 19976 9873
rect 20010 9839 20044 9873
rect 20078 9839 20112 9873
rect 20146 9839 20180 9873
rect 20214 9839 20248 9873
rect 20282 9839 20362 9873
rect 20396 9839 20432 9873
rect 19828 9826 20432 9839
rect 19828 9789 19932 9826
rect 19828 9755 19862 9789
rect 19896 9755 19932 9789
rect 19828 9721 19932 9755
rect 19828 9687 19862 9721
rect 19896 9687 19932 9721
rect 19828 9653 19932 9687
rect 19828 9619 19862 9653
rect 19896 9619 19932 9653
rect 19828 9585 19932 9619
rect 19828 9551 19862 9585
rect 19896 9551 19932 9585
rect 19828 9512 19932 9551
rect 20326 9789 20432 9826
rect 20326 9755 20362 9789
rect 20396 9755 20432 9789
rect 20326 9721 20432 9755
rect 20326 9687 20362 9721
rect 20396 9687 20432 9721
rect 20326 9653 20432 9687
rect 20326 9619 20362 9653
rect 20396 9652 20432 9653
rect 20326 9618 20367 9619
rect 20401 9618 20432 9652
rect 20326 9585 20432 9618
rect 20326 9551 20362 9585
rect 20396 9551 20432 9585
rect 20326 9512 20432 9551
rect 19828 9497 20432 9512
rect 19828 9463 19862 9497
rect 19896 9463 19976 9497
rect 20010 9463 20044 9497
rect 20078 9463 20112 9497
rect 20146 9463 20180 9497
rect 20214 9463 20248 9497
rect 20282 9463 20362 9497
rect 20396 9463 20432 9497
rect 19828 9445 20432 9463
rect 11158 9394 11187 9428
rect 11221 9394 11253 9428
rect 11158 9360 11253 9394
rect 17420 9407 18253 9423
rect 17420 9373 17443 9407
rect 17477 9373 17519 9407
rect 17553 9373 17587 9407
rect 17621 9373 17655 9407
rect 17689 9373 17723 9407
rect 17757 9373 17791 9407
rect 17825 9373 17859 9407
rect 17893 9373 17927 9407
rect 17961 9373 17995 9407
rect 18029 9373 18063 9407
rect 18097 9373 18131 9407
rect 18165 9373 18203 9407
rect 18237 9373 18253 9407
rect 11158 9326 11187 9360
rect 11221 9326 11253 9360
rect 11158 9292 11253 9326
rect 11158 9258 11187 9292
rect 11221 9258 11253 9292
rect 11158 9224 11253 9258
rect 11158 9190 11187 9224
rect 11221 9190 11253 9224
rect 11158 9156 11253 9190
rect 11158 9122 11187 9156
rect 11221 9122 11253 9156
rect 11158 9088 11253 9122
rect 11158 9054 11187 9088
rect 11221 9054 11253 9088
rect 11158 9020 11253 9054
rect 11158 8986 11187 9020
rect 11221 8986 11253 9020
rect 11158 8952 11253 8986
rect 11158 8918 11187 8952
rect 11221 8918 11253 8952
rect 11158 8884 11253 8918
rect 11158 8850 11187 8884
rect 11221 8850 11253 8884
rect 11158 8816 11253 8850
rect 11158 8782 11187 8816
rect 11221 8782 11253 8816
rect 11158 8748 11253 8782
rect 16452 9357 16966 9371
rect 16452 9344 16490 9357
rect 16452 9310 16489 9344
rect 16524 9323 16588 9357
rect 16622 9323 16656 9357
rect 16690 9323 16724 9357
rect 16758 9323 16792 9357
rect 16826 9323 16890 9357
rect 16924 9323 16966 9357
rect 16523 9312 16966 9323
rect 16523 9310 16563 9312
rect 16452 9285 16563 9310
rect 16452 9272 16490 9285
rect 16452 9238 16489 9272
rect 16524 9251 16563 9285
rect 16523 9238 16563 9251
rect 16452 9217 16563 9238
rect 16452 9183 16490 9217
rect 16524 9183 16563 9217
rect 16452 9149 16563 9183
rect 16452 9115 16490 9149
rect 16524 9115 16563 9149
rect 16452 9081 16563 9115
rect 16452 9047 16490 9081
rect 16524 9047 16563 9081
rect 16452 9013 16563 9047
rect 16452 8979 16490 9013
rect 16524 8979 16563 9013
rect 16452 8945 16563 8979
rect 16452 8911 16490 8945
rect 16524 8911 16563 8945
rect 16452 8877 16563 8911
rect 16452 8843 16490 8877
rect 16524 8843 16563 8877
rect 16452 8818 16563 8843
rect 16846 9285 16966 9312
rect 16846 9251 16890 9285
rect 16924 9251 16966 9285
rect 16846 9217 16966 9251
rect 16846 9183 16890 9217
rect 16924 9183 16966 9217
rect 16846 9149 16966 9183
rect 16846 9115 16890 9149
rect 16924 9115 16966 9149
rect 16846 9081 16966 9115
rect 16846 9047 16890 9081
rect 16924 9047 16966 9081
rect 16846 9013 16966 9047
rect 16846 8979 16890 9013
rect 16924 8979 16966 9013
rect 16846 8945 16966 8979
rect 16846 8911 16890 8945
rect 16924 8911 16966 8945
rect 16846 8877 16966 8911
rect 16846 8843 16890 8877
rect 16924 8843 16966 8877
rect 16846 8818 16966 8843
rect 16452 8805 16966 8818
rect 16452 8771 16490 8805
rect 16524 8771 16588 8805
rect 16622 8771 16656 8805
rect 16690 8771 16724 8805
rect 16758 8771 16792 8805
rect 16826 8771 16890 8805
rect 16924 8771 16966 8805
rect 16452 8755 16966 8771
rect 17420 9366 18253 9373
rect 17420 9312 17498 9366
rect 17420 9278 17443 9312
rect 17477 9278 17498 9312
rect 17420 9244 17498 9278
rect 17420 9210 17443 9244
rect 17477 9210 17498 9244
rect 17420 9176 17498 9210
rect 17420 9142 17443 9176
rect 17477 9142 17498 9176
rect 17420 9108 17498 9142
rect 17420 9074 17443 9108
rect 17477 9074 17498 9108
rect 17420 9040 17498 9074
rect 17420 9006 17443 9040
rect 17477 9006 17498 9040
rect 17420 8972 17498 9006
rect 17420 8938 17443 8972
rect 17477 8938 17498 8972
rect 18189 9312 18253 9366
rect 18189 9278 18203 9312
rect 18237 9278 18253 9312
rect 18189 9244 18253 9278
rect 18189 9210 18203 9244
rect 18237 9210 18253 9244
rect 18189 9176 18253 9210
rect 18189 9142 18203 9176
rect 18237 9142 18253 9176
rect 18189 9108 18253 9142
rect 18189 9074 18203 9108
rect 18237 9074 18253 9108
rect 18189 9040 18253 9074
rect 18189 9006 18203 9040
rect 18237 9006 18253 9040
rect 18189 8972 18253 9006
rect 17420 8904 17498 8938
rect 17420 8870 17443 8904
rect 17477 8870 17498 8904
rect 17570 8938 18075 8954
rect 17570 8904 17602 8938
rect 17636 8904 17670 8938
rect 17704 8904 17738 8938
rect 17772 8904 17806 8938
rect 17840 8904 17874 8938
rect 17908 8904 17942 8938
rect 17976 8904 18010 8938
rect 18044 8904 18075 8938
rect 17570 8888 18075 8904
rect 18189 8938 18203 8972
rect 18237 8938 18253 8972
rect 18189 8904 18253 8938
rect 17420 8836 17498 8870
rect 17420 8802 17443 8836
rect 17477 8802 17498 8836
rect 17420 8768 17498 8802
rect 11158 8714 11187 8748
rect 11221 8714 11253 8748
rect 11158 8680 11253 8714
rect 11158 8665 11187 8680
rect 11158 8631 11185 8665
rect 11221 8646 11253 8680
rect 11219 8631 11253 8646
rect 11158 8616 11253 8631
rect 10747 8604 11253 8616
rect 10747 8570 10776 8604
rect 10810 8570 10879 8604
rect 10913 8570 10947 8604
rect 10981 8570 11015 8604
rect 11049 8570 11083 8604
rect 11117 8570 11187 8604
rect 11221 8570 11253 8604
rect 10747 8553 11253 8570
rect 17420 8734 17443 8768
rect 17477 8734 17498 8768
rect 17420 8700 17498 8734
rect 17420 8666 17443 8700
rect 17477 8666 17498 8700
rect 17420 8632 17498 8666
rect 17420 8598 17443 8632
rect 17477 8598 17498 8632
rect 17420 8564 17498 8598
rect 10015 8539 10162 8545
rect 5698 8511 10162 8539
rect 5615 8409 5662 8511
rect 10116 8409 10162 8511
rect 17420 8530 17443 8564
rect 17477 8530 17498 8564
rect 5615 8387 10162 8409
rect 16357 8482 16961 8501
rect 16357 8448 16391 8482
rect 16425 8448 16505 8482
rect 16539 8448 16573 8482
rect 16607 8448 16641 8482
rect 16675 8448 16709 8482
rect 16743 8448 16777 8482
rect 16811 8474 16891 8482
rect 16811 8448 16889 8474
rect 16925 8448 16961 8482
rect 16357 8440 16889 8448
rect 16923 8440 16961 8448
rect 16357 8435 16961 8440
rect 16357 8398 16461 8435
rect 16357 8364 16391 8398
rect 16425 8364 16461 8398
rect 16357 8330 16461 8364
rect 16357 8296 16391 8330
rect 16425 8296 16461 8330
rect 16357 8262 16461 8296
rect 16357 8228 16391 8262
rect 16425 8228 16461 8262
rect 16357 8194 16461 8228
rect 10757 8154 11237 8175
rect 10757 8120 10791 8154
rect 10825 8120 10878 8154
rect 10912 8120 10946 8154
rect 10980 8120 11014 8154
rect 11048 8120 11082 8154
rect 11116 8120 11170 8154
rect 11204 8120 11237 8154
rect 10757 8099 11237 8120
rect 10757 8079 10858 8099
rect 10757 8045 10791 8079
rect 10825 8045 10858 8079
rect 10757 8011 10858 8045
rect 10757 7977 10791 8011
rect 10825 7977 10858 8011
rect 10757 7963 10858 7977
rect 10757 7929 10790 7963
rect 10824 7943 10858 7963
rect 10757 7909 10791 7929
rect 10825 7909 10858 7943
rect 10757 7891 10858 7909
rect 10757 7857 10790 7891
rect 10824 7875 10858 7891
rect 10757 7841 10791 7857
rect 10825 7841 10858 7875
rect 10757 7807 10858 7841
rect 10757 7773 10791 7807
rect 10825 7773 10858 7807
rect 10757 7753 10858 7773
rect 11136 8079 11237 8099
rect 11136 8045 11170 8079
rect 11204 8045 11237 8079
rect 16357 8160 16391 8194
rect 16425 8160 16461 8194
rect 16357 8121 16461 8160
rect 16855 8402 16961 8435
rect 16855 8368 16889 8402
rect 16923 8398 16961 8402
rect 16855 8364 16891 8368
rect 16925 8364 16961 8398
rect 16855 8330 16961 8364
rect 16855 8296 16891 8330
rect 16925 8296 16961 8330
rect 16855 8262 16961 8296
rect 16855 8228 16891 8262
rect 16925 8228 16961 8262
rect 16855 8194 16961 8228
rect 16855 8160 16891 8194
rect 16925 8160 16961 8194
rect 16855 8121 16961 8160
rect 16357 8106 16961 8121
rect 16357 8072 16391 8106
rect 16425 8072 16505 8106
rect 16539 8072 16573 8106
rect 16607 8072 16641 8106
rect 16675 8072 16709 8106
rect 16743 8072 16777 8106
rect 16811 8072 16891 8106
rect 16925 8072 16961 8106
rect 16357 8054 16961 8072
rect 17420 8496 17498 8530
rect 17420 8462 17443 8496
rect 17477 8462 17498 8496
rect 17420 8428 17498 8462
rect 17420 8394 17443 8428
rect 17477 8394 17498 8428
rect 17420 8360 17498 8394
rect 17420 8326 17443 8360
rect 17477 8326 17498 8360
rect 17420 8292 17498 8326
rect 17420 8258 17443 8292
rect 17477 8258 17498 8292
rect 17420 8224 17498 8258
rect 17420 8190 17443 8224
rect 17477 8190 17498 8224
rect 17420 8156 17498 8190
rect 17420 8122 17443 8156
rect 17477 8122 17498 8156
rect 17420 8088 17498 8122
rect 17420 8054 17443 8088
rect 17477 8054 17498 8088
rect 11136 8011 11237 8045
rect 11136 7977 11170 8011
rect 11204 7977 11237 8011
rect 11136 7957 11237 7977
rect 17420 8020 17498 8054
rect 17420 7986 17443 8020
rect 17477 7986 17498 8020
rect 16446 7961 16960 7975
rect 11136 7943 11238 7957
rect 11136 7909 11170 7943
rect 11204 7909 11238 7943
rect 11136 7877 11238 7909
rect 16446 7928 16484 7961
rect 16446 7894 16479 7928
rect 16518 7927 16582 7961
rect 16616 7927 16650 7961
rect 16684 7927 16718 7961
rect 16752 7927 16786 7961
rect 16820 7927 16884 7961
rect 16918 7927 16960 7961
rect 16513 7916 16960 7927
rect 16513 7894 16557 7916
rect 16446 7889 16557 7894
rect 11136 7875 11237 7877
rect 11136 7841 11170 7875
rect 11204 7841 11237 7875
rect 11136 7807 11237 7841
rect 11136 7773 11170 7807
rect 11204 7773 11237 7807
rect 11136 7753 11237 7773
rect 10757 7731 11237 7753
rect 10757 7697 10791 7731
rect 10825 7697 10878 7731
rect 10912 7697 10946 7731
rect 10980 7697 11014 7731
rect 11048 7697 11082 7731
rect 11116 7697 11170 7731
rect 11204 7697 11237 7731
rect 10757 7674 11237 7697
rect 16446 7856 16484 7889
rect 16446 7822 16479 7856
rect 16518 7855 16557 7889
rect 16513 7822 16557 7855
rect 16446 7821 16557 7822
rect 16446 7787 16484 7821
rect 16518 7787 16557 7821
rect 16446 7753 16557 7787
rect 16446 7719 16484 7753
rect 16518 7719 16557 7753
rect 16446 7685 16557 7719
rect 16446 7651 16484 7685
rect 16518 7651 16557 7685
rect 16446 7617 16557 7651
rect 16446 7583 16484 7617
rect 16518 7583 16557 7617
rect 10748 7540 11260 7560
rect 5613 7507 10159 7537
rect 5613 7473 5659 7507
rect 5693 7473 5727 7507
rect 5761 7473 5795 7507
rect 5829 7473 5863 7507
rect 5897 7473 5931 7507
rect 5965 7473 5999 7507
rect 6033 7473 6067 7507
rect 6101 7473 6135 7507
rect 6169 7473 6203 7507
rect 6237 7473 6271 7507
rect 6305 7473 6339 7507
rect 6373 7473 6407 7507
rect 6441 7473 6475 7507
rect 6509 7473 6543 7507
rect 6577 7473 6611 7507
rect 6645 7473 6679 7507
rect 6713 7473 6747 7507
rect 6781 7473 6815 7507
rect 6849 7473 6883 7507
rect 6917 7473 6951 7507
rect 6985 7473 7019 7507
rect 7053 7473 7087 7507
rect 7121 7473 7155 7507
rect 7189 7473 7223 7507
rect 7257 7473 7291 7507
rect 7325 7473 7359 7507
rect 7393 7473 7427 7507
rect 7461 7473 7495 7507
rect 7529 7473 7563 7507
rect 7597 7473 7631 7507
rect 7665 7473 7699 7507
rect 7733 7473 7767 7507
rect 7801 7473 7835 7507
rect 7869 7473 7903 7507
rect 7937 7473 7971 7507
rect 8005 7473 8039 7507
rect 8073 7473 8107 7507
rect 8141 7473 8175 7507
rect 8209 7473 8243 7507
rect 8277 7473 8311 7507
rect 8345 7473 8379 7507
rect 8413 7473 8447 7507
rect 8481 7473 8515 7507
rect 8549 7473 8583 7507
rect 8617 7473 8651 7507
rect 8685 7473 8719 7507
rect 8753 7473 8787 7507
rect 8821 7473 8855 7507
rect 8889 7473 8923 7507
rect 8957 7473 8991 7507
rect 9025 7473 9059 7507
rect 9093 7473 9127 7507
rect 9161 7473 9195 7507
rect 9229 7473 9263 7507
rect 9297 7473 9331 7507
rect 9365 7473 9399 7507
rect 9433 7473 9467 7507
rect 9501 7473 9535 7507
rect 9569 7473 9603 7507
rect 9637 7473 9671 7507
rect 9705 7473 9739 7507
rect 9773 7473 9807 7507
rect 9841 7473 9875 7507
rect 9909 7473 9943 7507
rect 9977 7473 10011 7507
rect 10045 7473 10079 7507
rect 10113 7473 10159 7507
rect 10748 7506 10783 7540
rect 10817 7506 10886 7540
rect 10920 7506 10954 7540
rect 10988 7506 11022 7540
rect 11056 7506 11090 7540
rect 11124 7506 11194 7540
rect 11228 7506 11260 7540
rect 10748 7483 11260 7506
rect 5613 7439 10159 7473
rect 5613 7405 5659 7439
rect 5693 7405 10079 7439
rect 10113 7405 10159 7439
rect 5613 7388 10159 7405
rect 5613 7371 5753 7388
rect 5613 7337 5659 7371
rect 5693 7337 5753 7371
rect 5613 7303 5753 7337
rect 5613 7269 5659 7303
rect 5693 7269 5753 7303
rect 5613 7235 5753 7269
rect 5613 7201 5659 7235
rect 5693 7201 5753 7235
rect 5613 7167 5753 7201
rect 5613 7133 5659 7167
rect 5693 7133 5753 7167
rect 5613 7099 5753 7133
rect 5613 7065 5659 7099
rect 5693 7065 5753 7099
rect 5613 7031 5753 7065
rect 5613 6997 5659 7031
rect 5693 6997 5753 7031
rect 5613 6963 5753 6997
rect 5613 6929 5659 6963
rect 5693 6929 5753 6963
rect 5613 6895 5753 6929
rect 5613 6861 5659 6895
rect 5693 6861 5753 6895
rect 5613 6827 5753 6861
rect 5613 6793 5659 6827
rect 5693 6793 5753 6827
rect 5613 6759 5753 6793
rect 5613 6725 5659 6759
rect 5693 6725 5753 6759
rect 5613 6691 5753 6725
rect 5613 6657 5659 6691
rect 5693 6657 5753 6691
rect 5613 6623 5753 6657
rect 5613 6589 5659 6623
rect 5693 6589 5753 6623
rect 5613 6555 5753 6589
rect 5613 6521 5659 6555
rect 5693 6521 5753 6555
rect 5613 6516 5753 6521
rect 10021 7371 10159 7388
rect 10021 7337 10079 7371
rect 10113 7337 10159 7371
rect 10021 7303 10159 7337
rect 10021 7269 10079 7303
rect 10113 7269 10159 7303
rect 10021 7235 10159 7269
rect 10021 7201 10079 7235
rect 10113 7201 10159 7235
rect 10021 7167 10159 7201
rect 10021 7133 10079 7167
rect 10113 7133 10159 7167
rect 10021 7099 10159 7133
rect 10021 7065 10079 7099
rect 10113 7065 10159 7099
rect 10021 7031 10159 7065
rect 10021 6997 10079 7031
rect 10113 6997 10159 7031
rect 10021 6963 10159 6997
rect 10021 6929 10079 6963
rect 10113 6929 10159 6963
rect 10021 6895 10159 6929
rect 10021 6861 10079 6895
rect 10113 6861 10159 6895
rect 10021 6827 10159 6861
rect 10021 6793 10079 6827
rect 10113 6793 10159 6827
rect 10021 6759 10159 6793
rect 10021 6725 10079 6759
rect 10113 6725 10159 6759
rect 10021 6691 10159 6725
rect 10021 6657 10079 6691
rect 10113 6657 10159 6691
rect 10021 6623 10159 6657
rect 10021 6589 10079 6623
rect 10113 6589 10159 6623
rect 10021 6555 10159 6589
rect 10021 6521 10079 6555
rect 10113 6521 10159 6555
rect 10021 6516 10159 6521
rect 5613 6487 10159 6516
rect 5613 6385 5659 6487
rect 10113 6385 10159 6487
rect 5613 6357 10159 6385
rect 10754 7455 10840 7483
rect 10754 7421 10783 7455
rect 10817 7421 10840 7455
rect 10754 7387 10840 7421
rect 10754 7353 10783 7387
rect 10817 7353 10840 7387
rect 10754 7319 10840 7353
rect 10754 7285 10783 7319
rect 10817 7285 10840 7319
rect 10754 7251 10840 7285
rect 10754 7217 10783 7251
rect 10817 7217 10840 7251
rect 10754 7183 10840 7217
rect 10754 7149 10783 7183
rect 10817 7149 10840 7183
rect 10754 7115 10840 7149
rect 10754 7081 10783 7115
rect 10817 7081 10840 7115
rect 10754 7047 10840 7081
rect 10754 7013 10783 7047
rect 10817 7013 10840 7047
rect 10754 6979 10840 7013
rect 10754 6945 10783 6979
rect 10817 6945 10840 6979
rect 10754 6911 10840 6945
rect 10754 6877 10783 6911
rect 10817 6877 10840 6911
rect 10754 6843 10840 6877
rect 10754 6809 10783 6843
rect 10817 6809 10840 6843
rect 10754 6775 10840 6809
rect 10754 6741 10783 6775
rect 10817 6741 10840 6775
rect 10754 6707 10840 6741
rect 10754 6673 10783 6707
rect 10817 6673 10840 6707
rect 10754 6639 10840 6673
rect 10754 6605 10783 6639
rect 10817 6605 10840 6639
rect 10754 6571 10840 6605
rect 10754 6537 10783 6571
rect 10817 6537 10840 6571
rect 10754 6503 10840 6537
rect 10754 6469 10783 6503
rect 10817 6469 10840 6503
rect 10754 6435 10840 6469
rect 10754 6401 10783 6435
rect 10817 6401 10840 6435
rect 10754 6367 10840 6401
rect 10754 6333 10783 6367
rect 10817 6333 10840 6367
rect 10754 6299 10840 6333
rect 10754 6265 10783 6299
rect 10817 6265 10840 6299
rect 10754 6231 10840 6265
rect 10754 6197 10783 6231
rect 10817 6197 10840 6231
rect 10754 6163 10840 6197
rect 10754 6129 10783 6163
rect 10817 6129 10840 6163
rect 10754 6095 10840 6129
rect 10754 6061 10783 6095
rect 10817 6061 10840 6095
rect 10754 6027 10840 6061
rect 10754 5993 10783 6027
rect 10817 5993 10840 6027
rect 10754 5959 10840 5993
rect 10754 5925 10783 5959
rect 10817 5925 10840 5959
rect 10754 5891 10840 5925
rect 10754 5857 10783 5891
rect 10817 5857 10840 5891
rect 10754 5823 10840 5857
rect 10754 5789 10783 5823
rect 10817 5789 10840 5823
rect 10754 5755 10840 5789
rect 10754 5721 10783 5755
rect 10817 5721 10840 5755
rect 10754 5687 10840 5721
rect 10754 5653 10783 5687
rect 10817 5653 10840 5687
rect 10754 5623 10840 5653
rect 11165 7455 11260 7483
rect 11165 7421 11194 7455
rect 11228 7421 11260 7455
rect 11165 7387 11260 7421
rect 11165 7353 11194 7387
rect 11228 7353 11260 7387
rect 16446 7549 16557 7583
rect 16446 7515 16484 7549
rect 16518 7515 16557 7549
rect 16446 7481 16557 7515
rect 16446 7447 16484 7481
rect 16518 7447 16557 7481
rect 16446 7422 16557 7447
rect 16840 7889 16960 7916
rect 16840 7855 16884 7889
rect 16918 7855 16960 7889
rect 17420 7944 17498 7986
rect 18189 8870 18203 8904
rect 18237 8870 18253 8904
rect 18189 8836 18253 8870
rect 18189 8802 18203 8836
rect 18237 8802 18253 8836
rect 18189 8768 18253 8802
rect 18189 8734 18203 8768
rect 18237 8734 18253 8768
rect 18189 8700 18253 8734
rect 18189 8666 18203 8700
rect 18237 8666 18253 8700
rect 18189 8632 18253 8666
rect 18189 8598 18203 8632
rect 18237 8598 18253 8632
rect 18189 8564 18253 8598
rect 18189 8530 18203 8564
rect 18237 8530 18253 8564
rect 18189 8496 18253 8530
rect 18189 8462 18203 8496
rect 18237 8462 18253 8496
rect 18189 8428 18253 8462
rect 18189 8394 18203 8428
rect 18237 8394 18253 8428
rect 18189 8360 18253 8394
rect 18189 8326 18203 8360
rect 18237 8326 18253 8360
rect 18189 8292 18253 8326
rect 18189 8258 18203 8292
rect 18237 8258 18253 8292
rect 18189 8224 18253 8258
rect 18189 8190 18203 8224
rect 18237 8190 18253 8224
rect 18189 8156 18253 8190
rect 18189 8122 18203 8156
rect 18237 8122 18253 8156
rect 18189 8088 18253 8122
rect 18189 8054 18203 8088
rect 18237 8054 18253 8088
rect 18189 8020 18253 8054
rect 18189 7986 18203 8020
rect 18237 7986 18253 8020
rect 18189 7944 18253 7986
rect 18539 9396 19429 9424
rect 18539 9392 19284 9396
rect 19318 9392 19356 9396
rect 19390 9392 19429 9396
rect 18539 9358 18554 9392
rect 18588 9358 18627 9392
rect 18661 9358 18695 9392
rect 18729 9358 18763 9392
rect 18797 9358 18831 9392
rect 18865 9358 18899 9392
rect 18933 9358 18967 9392
rect 19001 9358 19035 9392
rect 19069 9358 19103 9392
rect 19137 9358 19171 9392
rect 19205 9358 19239 9392
rect 19273 9362 19284 9392
rect 19341 9362 19356 9392
rect 19273 9358 19307 9362
rect 19341 9358 19380 9362
rect 19414 9358 19429 9392
rect 18539 9330 19429 9358
rect 18539 9303 18603 9330
rect 18539 9269 18554 9303
rect 18588 9269 18603 9303
rect 18539 9235 18603 9269
rect 18539 9201 18554 9235
rect 18588 9201 18603 9235
rect 18539 9167 18603 9201
rect 18539 9133 18554 9167
rect 18588 9133 18603 9167
rect 18539 9099 18603 9133
rect 18539 9065 18554 9099
rect 18588 9065 18603 9099
rect 18539 9031 18603 9065
rect 18539 8997 18554 9031
rect 18588 8997 18603 9031
rect 18539 8963 18603 8997
rect 18539 8929 18554 8963
rect 18588 8929 18603 8963
rect 18539 8895 18603 8929
rect 18539 8861 18554 8895
rect 18588 8861 18603 8895
rect 18539 8827 18603 8861
rect 18539 8793 18554 8827
rect 18588 8793 18603 8827
rect 18539 8759 18603 8793
rect 18539 8725 18554 8759
rect 18588 8725 18603 8759
rect 18539 8691 18603 8725
rect 18539 8657 18554 8691
rect 18588 8657 18603 8691
rect 18539 8623 18603 8657
rect 18539 8589 18554 8623
rect 18588 8589 18603 8623
rect 18539 8555 18603 8589
rect 18539 8521 18554 8555
rect 18588 8521 18603 8555
rect 18539 8487 18603 8521
rect 18539 8453 18554 8487
rect 18588 8453 18603 8487
rect 18539 8419 18603 8453
rect 18539 8385 18554 8419
rect 18588 8385 18603 8419
rect 18539 8351 18603 8385
rect 18539 8317 18554 8351
rect 18588 8317 18603 8351
rect 18539 8283 18603 8317
rect 18539 8249 18554 8283
rect 18588 8249 18603 8283
rect 18539 8215 18603 8249
rect 18539 8181 18554 8215
rect 18588 8181 18603 8215
rect 18539 8147 18603 8181
rect 18539 8113 18554 8147
rect 18588 8113 18603 8147
rect 18539 8079 18603 8113
rect 18539 8045 18554 8079
rect 18588 8045 18603 8079
rect 18539 8011 18603 8045
rect 18539 7977 18554 8011
rect 18588 7977 18603 8011
rect 18539 7951 18603 7977
rect 19365 9303 19429 9330
rect 19365 9269 19380 9303
rect 19414 9269 19429 9303
rect 19365 9235 19429 9269
rect 19365 9201 19380 9235
rect 19414 9201 19429 9235
rect 19365 9167 19429 9201
rect 19365 9133 19380 9167
rect 19414 9133 19429 9167
rect 19365 9099 19429 9133
rect 19365 9065 19380 9099
rect 19414 9065 19429 9099
rect 19365 9031 19429 9065
rect 19365 8997 19380 9031
rect 19414 8997 19429 9031
rect 19365 8963 19429 8997
rect 19365 8929 19380 8963
rect 19414 8929 19429 8963
rect 19365 8895 19429 8929
rect 19365 8861 19380 8895
rect 19414 8861 19429 8895
rect 19365 8827 19429 8861
rect 19365 8793 19380 8827
rect 19414 8793 19429 8827
rect 19365 8759 19429 8793
rect 19365 8725 19380 8759
rect 19414 8725 19429 8759
rect 19919 9352 20433 9366
rect 19919 9318 19957 9352
rect 19991 9318 20055 9352
rect 20089 9318 20123 9352
rect 20157 9318 20191 9352
rect 20225 9318 20259 9352
rect 20293 9318 20357 9352
rect 20391 9318 20433 9352
rect 19919 9307 20433 9318
rect 19919 9280 20030 9307
rect 19919 9246 19957 9280
rect 19991 9246 20030 9280
rect 19919 9212 20030 9246
rect 19919 9178 19957 9212
rect 19991 9178 20030 9212
rect 19919 9144 20030 9178
rect 19919 9110 19957 9144
rect 19991 9110 20030 9144
rect 19919 9076 20030 9110
rect 19919 9042 19957 9076
rect 19991 9042 20030 9076
rect 19919 9016 20030 9042
rect 19919 9008 19959 9016
rect 19919 8974 19957 9008
rect 19993 8982 20030 9016
rect 19991 8974 20030 8982
rect 19919 8940 20030 8974
rect 19919 8906 19957 8940
rect 19991 8906 20030 8940
rect 19919 8872 20030 8906
rect 19919 8838 19957 8872
rect 19991 8838 20030 8872
rect 19919 8813 20030 8838
rect 20313 9280 20433 9307
rect 20313 9246 20357 9280
rect 20391 9246 20433 9280
rect 20313 9212 20433 9246
rect 20313 9178 20357 9212
rect 20391 9178 20433 9212
rect 20313 9144 20433 9178
rect 20313 9110 20357 9144
rect 20391 9110 20433 9144
rect 20313 9076 20433 9110
rect 20313 9042 20357 9076
rect 20391 9042 20433 9076
rect 20313 9008 20433 9042
rect 20313 8974 20357 9008
rect 20391 8974 20433 9008
rect 20313 8940 20433 8974
rect 20313 8906 20357 8940
rect 20391 8906 20433 8940
rect 20313 8872 20433 8906
rect 20313 8838 20357 8872
rect 20391 8838 20433 8872
rect 20313 8813 20433 8838
rect 19919 8800 20433 8813
rect 19919 8766 19957 8800
rect 19991 8766 20055 8800
rect 20089 8766 20123 8800
rect 20157 8766 20191 8800
rect 20225 8766 20259 8800
rect 20293 8766 20357 8800
rect 20391 8766 20433 8800
rect 19919 8750 20433 8766
rect 19365 8691 19429 8725
rect 19365 8657 19380 8691
rect 19414 8657 19429 8691
rect 19365 8623 19429 8657
rect 19365 8589 19380 8623
rect 19414 8589 19429 8623
rect 19365 8555 19429 8589
rect 19365 8521 19380 8555
rect 19414 8521 19429 8555
rect 19365 8487 19429 8521
rect 19365 8453 19380 8487
rect 19414 8453 19429 8487
rect 19365 8419 19429 8453
rect 19365 8385 19380 8419
rect 19414 8385 19429 8419
rect 19365 8351 19429 8385
rect 19365 8317 19380 8351
rect 19414 8317 19429 8351
rect 19365 8283 19429 8317
rect 19365 8249 19380 8283
rect 19414 8249 19429 8283
rect 19365 8215 19429 8249
rect 19365 8181 19380 8215
rect 19414 8181 19429 8215
rect 19365 8147 19429 8181
rect 19365 8113 19380 8147
rect 19414 8113 19429 8147
rect 19825 8542 20429 8561
rect 19825 8508 19859 8542
rect 19893 8508 19973 8542
rect 20007 8508 20041 8542
rect 20075 8508 20109 8542
rect 20143 8508 20177 8542
rect 20211 8508 20245 8542
rect 20279 8508 20359 8542
rect 20393 8508 20429 8542
rect 19825 8495 20429 8508
rect 19825 8458 19929 8495
rect 19825 8424 19859 8458
rect 19893 8424 19929 8458
rect 19825 8390 19929 8424
rect 19825 8356 19859 8390
rect 19893 8356 19929 8390
rect 19825 8322 19929 8356
rect 19825 8288 19859 8322
rect 19893 8288 19929 8322
rect 19825 8254 19929 8288
rect 19825 8220 19859 8254
rect 19893 8220 19929 8254
rect 19825 8181 19929 8220
rect 20323 8458 20429 8495
rect 20323 8424 20359 8458
rect 20393 8424 20429 8458
rect 20323 8390 20429 8424
rect 20323 8356 20359 8390
rect 20393 8356 20429 8390
rect 20323 8322 20429 8356
rect 20323 8288 20359 8322
rect 20393 8300 20429 8322
rect 20323 8266 20363 8288
rect 20397 8266 20429 8300
rect 20323 8254 20429 8266
rect 20323 8220 20359 8254
rect 20393 8220 20429 8254
rect 20323 8181 20429 8220
rect 19825 8166 20429 8181
rect 19825 8132 19859 8166
rect 19893 8132 19973 8166
rect 20007 8132 20041 8166
rect 20075 8132 20109 8166
rect 20143 8132 20177 8166
rect 20211 8132 20245 8166
rect 20279 8132 20359 8166
rect 20393 8132 20429 8166
rect 19825 8114 20429 8132
rect 19365 8079 19429 8113
rect 19365 8045 19380 8079
rect 19414 8045 19429 8079
rect 19365 8011 19429 8045
rect 19365 7977 19380 8011
rect 19414 7977 19429 8011
rect 19365 7951 19429 7977
rect 17420 7919 18253 7944
rect 17420 7885 17443 7919
rect 17478 7885 17516 7919
rect 17553 7885 17587 7919
rect 17622 7885 17655 7919
rect 17694 7885 17723 7919
rect 17766 7885 17791 7919
rect 17825 7885 17859 7919
rect 17893 7885 17927 7919
rect 17961 7885 17995 7919
rect 18029 7885 18063 7919
rect 18097 7885 18131 7919
rect 18165 7885 18203 7919
rect 18237 7885 18253 7919
rect 17420 7858 18253 7885
rect 18537 7950 19429 7951
rect 19915 8021 20429 8035
rect 19915 7987 19953 8021
rect 19987 7987 20051 8021
rect 20085 7987 20119 8021
rect 20153 7987 20187 8021
rect 20221 7987 20255 8021
rect 20289 7987 20353 8021
rect 20387 7987 20429 8021
rect 19915 7976 20429 7987
rect 18537 7921 19435 7950
rect 18537 7887 18554 7921
rect 18588 7887 18627 7921
rect 18661 7887 18695 7921
rect 18729 7887 18763 7921
rect 18797 7887 18831 7921
rect 18865 7887 18899 7921
rect 18933 7887 18967 7921
rect 19001 7887 19035 7921
rect 19069 7887 19103 7921
rect 19137 7887 19171 7921
rect 19205 7887 19239 7921
rect 19273 7887 19307 7921
rect 19341 7887 19380 7921
rect 19414 7887 19435 7921
rect 18537 7858 19435 7887
rect 19915 7949 20026 7976
rect 19915 7910 19953 7949
rect 19987 7910 20026 7949
rect 19915 7881 20026 7910
rect 18537 7857 19429 7858
rect 16840 7821 16960 7855
rect 16840 7787 16884 7821
rect 16918 7787 16960 7821
rect 16840 7753 16960 7787
rect 16840 7719 16884 7753
rect 16918 7719 16960 7753
rect 16840 7685 16960 7719
rect 16840 7651 16884 7685
rect 16918 7651 16960 7685
rect 16840 7617 16960 7651
rect 16840 7583 16884 7617
rect 16918 7583 16960 7617
rect 16840 7549 16960 7583
rect 16840 7515 16884 7549
rect 16918 7515 16960 7549
rect 16840 7481 16960 7515
rect 16840 7447 16884 7481
rect 16918 7447 16960 7481
rect 16840 7422 16960 7447
rect 16446 7409 16960 7422
rect 19915 7847 19953 7881
rect 19987 7847 20026 7881
rect 19915 7813 20026 7847
rect 19915 7779 19953 7813
rect 19987 7779 20026 7813
rect 19915 7745 20026 7779
rect 19915 7711 19953 7745
rect 19987 7711 20026 7745
rect 19915 7677 20026 7711
rect 19915 7643 19953 7677
rect 19987 7643 20026 7677
rect 19915 7609 20026 7643
rect 19915 7575 19953 7609
rect 19987 7575 20026 7609
rect 19915 7541 20026 7575
rect 19915 7507 19953 7541
rect 19987 7507 20026 7541
rect 19915 7482 20026 7507
rect 20309 7949 20429 7976
rect 20309 7915 20353 7949
rect 20387 7915 20429 7949
rect 20309 7881 20429 7915
rect 20309 7847 20353 7881
rect 20387 7847 20429 7881
rect 20309 7813 20429 7847
rect 20309 7779 20353 7813
rect 20387 7779 20429 7813
rect 20309 7745 20429 7779
rect 20309 7711 20353 7745
rect 20387 7711 20429 7745
rect 20309 7677 20429 7711
rect 20309 7643 20353 7677
rect 20387 7643 20429 7677
rect 20309 7609 20429 7643
rect 20309 7575 20353 7609
rect 20387 7575 20429 7609
rect 20309 7541 20429 7575
rect 20309 7507 20353 7541
rect 20387 7507 20429 7541
rect 20309 7482 20429 7507
rect 19915 7469 20429 7482
rect 19915 7435 19953 7469
rect 19987 7435 20051 7469
rect 20085 7435 20119 7469
rect 20153 7435 20187 7469
rect 20221 7435 20255 7469
rect 20289 7435 20353 7469
rect 20387 7435 20429 7469
rect 19915 7419 20429 7435
rect 16446 7375 16484 7409
rect 16518 7375 16582 7409
rect 16616 7375 16650 7409
rect 16684 7375 16718 7409
rect 16752 7375 16786 7409
rect 16820 7375 16884 7409
rect 16918 7375 16960 7409
rect 16446 7359 16960 7375
rect 11165 7319 11260 7353
rect 11165 7285 11194 7319
rect 11228 7285 11260 7319
rect 11165 7251 11260 7285
rect 11165 7217 11194 7251
rect 11228 7217 11260 7251
rect 11165 7183 11260 7217
rect 11165 7149 11194 7183
rect 11228 7149 11260 7183
rect 11165 7115 11260 7149
rect 11165 7081 11194 7115
rect 11228 7081 11260 7115
rect 11165 7047 11260 7081
rect 11165 7013 11194 7047
rect 11228 7013 11260 7047
rect 11165 6979 11260 7013
rect 11165 6945 11194 6979
rect 11228 6945 11260 6979
rect 11165 6911 11260 6945
rect 11165 6877 11194 6911
rect 11228 6877 11260 6911
rect 11165 6843 11260 6877
rect 19839 7300 20443 7319
rect 19839 7266 19873 7300
rect 19907 7266 19987 7300
rect 20021 7266 20055 7300
rect 20089 7266 20123 7300
rect 20157 7266 20191 7300
rect 20225 7266 20259 7300
rect 20293 7266 20373 7300
rect 20407 7266 20443 7300
rect 19839 7253 20443 7266
rect 19839 7216 19943 7253
rect 19839 7182 19873 7216
rect 19907 7182 19943 7216
rect 19839 7148 19943 7182
rect 19839 7114 19873 7148
rect 19907 7114 19943 7148
rect 19839 7080 19943 7114
rect 19839 7046 19873 7080
rect 19907 7046 19943 7080
rect 19839 7012 19943 7046
rect 19839 6978 19873 7012
rect 19907 6978 19943 7012
rect 19839 6939 19943 6978
rect 20337 7216 20443 7253
rect 20337 7182 20373 7216
rect 20407 7182 20443 7216
rect 20337 7148 20443 7182
rect 20337 7114 20373 7148
rect 20407 7114 20443 7148
rect 20337 7085 20443 7114
rect 20337 7046 20373 7085
rect 20407 7046 20443 7085
rect 20337 7012 20443 7046
rect 20337 6978 20373 7012
rect 20407 6978 20443 7012
rect 20337 6939 20443 6978
rect 19839 6924 20443 6939
rect 19839 6890 19873 6924
rect 19907 6890 19987 6924
rect 20021 6890 20055 6924
rect 20089 6890 20123 6924
rect 20157 6890 20191 6924
rect 20225 6890 20259 6924
rect 20293 6890 20373 6924
rect 20407 6890 20443 6924
rect 19839 6872 20443 6890
rect 11165 6809 11194 6843
rect 11228 6809 11260 6843
rect 11165 6775 11260 6809
rect 11165 6741 11194 6775
rect 11228 6741 11260 6775
rect 11165 6707 11260 6741
rect 11165 6673 11194 6707
rect 11228 6673 11260 6707
rect 11165 6639 11260 6673
rect 11165 6605 11194 6639
rect 11228 6605 11260 6639
rect 11165 6571 11260 6605
rect 11165 6537 11194 6571
rect 11228 6537 11260 6571
rect 11165 6503 11260 6537
rect 11165 6469 11194 6503
rect 11228 6469 11260 6503
rect 11165 6435 11260 6469
rect 11165 6401 11194 6435
rect 11228 6401 11260 6435
rect 11165 6367 11260 6401
rect 11165 6333 11194 6367
rect 11228 6333 11260 6367
rect 11165 6299 11260 6333
rect 11165 6265 11194 6299
rect 11228 6265 11260 6299
rect 11165 6231 11260 6265
rect 11165 6197 11194 6231
rect 11228 6197 11260 6231
rect 11165 6163 11260 6197
rect 19933 6779 20447 6793
rect 19933 6745 19971 6779
rect 20005 6745 20069 6779
rect 20103 6745 20137 6779
rect 20171 6745 20205 6779
rect 20239 6745 20273 6779
rect 20307 6745 20371 6779
rect 20405 6745 20447 6779
rect 19933 6734 20447 6745
rect 19933 6707 20044 6734
rect 19933 6673 19971 6707
rect 20005 6673 20044 6707
rect 19933 6639 20044 6673
rect 19933 6605 19971 6639
rect 20005 6605 20044 6639
rect 19933 6571 20044 6605
rect 19933 6537 19971 6571
rect 20005 6537 20044 6571
rect 19933 6503 20044 6537
rect 19933 6469 19971 6503
rect 20005 6469 20044 6503
rect 19933 6435 20044 6469
rect 19933 6401 19971 6435
rect 20005 6401 20044 6435
rect 19933 6367 20044 6401
rect 19933 6333 19971 6367
rect 20005 6333 20044 6367
rect 19933 6299 20044 6333
rect 19933 6265 19971 6299
rect 20005 6265 20044 6299
rect 19933 6258 20044 6265
rect 19933 6224 19959 6258
rect 19993 6240 20044 6258
rect 20327 6707 20447 6734
rect 20327 6673 20371 6707
rect 20405 6673 20447 6707
rect 20327 6639 20447 6673
rect 20327 6605 20371 6639
rect 20405 6605 20447 6639
rect 20327 6571 20447 6605
rect 20327 6537 20371 6571
rect 20405 6537 20447 6571
rect 20327 6503 20447 6537
rect 20327 6469 20371 6503
rect 20405 6469 20447 6503
rect 20327 6435 20447 6469
rect 20327 6401 20371 6435
rect 20405 6401 20447 6435
rect 20327 6367 20447 6401
rect 20327 6333 20371 6367
rect 20405 6333 20447 6367
rect 20327 6299 20447 6333
rect 20327 6265 20371 6299
rect 20405 6265 20447 6299
rect 20327 6240 20447 6265
rect 19993 6227 20447 6240
rect 19933 6193 19971 6224
rect 20005 6193 20069 6227
rect 20103 6193 20137 6227
rect 20171 6193 20205 6227
rect 20239 6193 20273 6227
rect 20307 6193 20371 6227
rect 20405 6193 20447 6227
rect 19933 6177 20447 6193
rect 11165 6129 11194 6163
rect 11228 6129 11260 6163
rect 11165 6095 11260 6129
rect 11165 6061 11194 6095
rect 11228 6061 11260 6095
rect 11165 6027 11260 6061
rect 11165 5993 11194 6027
rect 11228 5993 11260 6027
rect 11165 5959 11260 5993
rect 11165 5925 11194 5959
rect 11228 5925 11260 5959
rect 12603 5940 12683 5941
rect 11165 5891 11260 5925
rect 11165 5857 11194 5891
rect 11228 5857 11260 5891
rect 11165 5823 11260 5857
rect 11165 5789 11194 5823
rect 11228 5789 11260 5823
rect 11165 5755 11260 5789
rect 11165 5721 11194 5755
rect 11228 5721 11260 5755
rect 11165 5687 11260 5721
rect 11165 5653 11194 5687
rect 11228 5665 11260 5687
rect 11165 5631 11197 5653
rect 11231 5631 11260 5665
rect 11165 5623 11260 5631
rect 10754 5611 11260 5623
rect 10754 5577 10783 5611
rect 10817 5577 10886 5611
rect 10920 5577 10954 5611
rect 10988 5577 11022 5611
rect 11056 5577 11090 5611
rect 11124 5577 11194 5611
rect 11228 5577 11260 5611
rect 10754 5560 11260 5577
rect 12385 5907 12886 5940
rect 12385 5873 12405 5907
rect 12439 5873 12481 5907
rect 12515 5873 12549 5907
rect 12583 5873 12617 5907
rect 12651 5873 12685 5907
rect 12719 5873 12753 5907
rect 12787 5873 12828 5907
rect 12862 5873 12886 5907
rect 12385 5839 12886 5873
rect 12385 5819 12461 5839
rect 12385 5785 12405 5819
rect 12439 5785 12461 5819
rect 12385 5751 12461 5785
rect 12385 5717 12405 5751
rect 12439 5717 12461 5751
rect 12385 5683 12461 5717
rect 12385 5649 12405 5683
rect 12439 5649 12461 5683
rect 12385 5615 12461 5649
rect 12385 5581 12405 5615
rect 12439 5581 12461 5615
rect 12385 5561 12461 5581
rect 12807 5819 12886 5839
rect 12807 5785 12828 5819
rect 12862 5785 12886 5819
rect 12807 5751 12886 5785
rect 12807 5717 12828 5751
rect 12862 5717 12886 5751
rect 12807 5683 12886 5717
rect 12807 5649 12828 5683
rect 12862 5649 12886 5683
rect 12807 5615 12886 5649
rect 12807 5581 12828 5615
rect 12862 5581 12886 5615
rect 12807 5561 12886 5581
rect 12385 5528 12886 5561
rect 12385 5494 12405 5528
rect 12439 5494 12449 5528
rect 12515 5494 12521 5528
rect 12583 5494 12593 5528
rect 12651 5494 12685 5528
rect 12719 5494 12753 5528
rect 12787 5494 12828 5528
rect 12862 5494 12886 5528
rect 12385 5460 12886 5494
rect 13000 5913 15000 5945
rect 13000 5879 13020 5913
rect 13054 5879 13105 5913
rect 13139 5879 13173 5913
rect 13207 5879 13241 5913
rect 13275 5879 13309 5913
rect 13343 5879 13377 5913
rect 13411 5879 13445 5913
rect 13479 5879 13513 5913
rect 13547 5879 13581 5913
rect 13615 5879 13649 5913
rect 13683 5879 13717 5913
rect 13751 5879 13785 5913
rect 13819 5879 13853 5913
rect 13887 5879 13921 5913
rect 13955 5879 13989 5913
rect 14023 5879 14057 5913
rect 14091 5879 14125 5913
rect 14159 5879 14193 5913
rect 14227 5879 14261 5913
rect 14295 5879 14329 5913
rect 14363 5879 14397 5913
rect 14431 5879 14465 5913
rect 14499 5879 14533 5913
rect 14567 5879 14601 5913
rect 14635 5879 14669 5913
rect 14703 5879 14737 5913
rect 14771 5879 14805 5913
rect 14839 5879 14873 5913
rect 14907 5879 14949 5913
rect 14983 5879 15000 5913
rect 13000 5850 15000 5879
rect 13000 5809 13077 5850
rect 13000 5775 13020 5809
rect 13054 5775 13077 5809
rect 13000 5741 13077 5775
rect 13000 5707 13020 5741
rect 13054 5707 13077 5741
rect 13000 5673 13077 5707
rect 13000 5639 13020 5673
rect 13054 5639 13077 5673
rect 13000 5605 13077 5639
rect 13000 5571 13020 5605
rect 13054 5571 13077 5605
rect 13000 5525 13077 5571
rect 14937 5809 15000 5850
rect 14937 5775 14949 5809
rect 14983 5775 15000 5809
rect 14937 5741 15000 5775
rect 14937 5707 14949 5741
rect 14983 5707 15000 5741
rect 14937 5673 15000 5707
rect 14937 5639 14949 5673
rect 14983 5639 15000 5673
rect 14937 5605 15000 5639
rect 14937 5571 14949 5605
rect 14983 5571 15000 5605
rect 14937 5525 15000 5571
rect 13000 5521 15000 5525
rect 13000 5487 13017 5521
rect 13051 5502 15000 5521
rect 13051 5500 13105 5502
rect 13000 5466 13020 5487
rect 13054 5468 13105 5500
rect 13139 5468 13173 5502
rect 13207 5468 13241 5502
rect 13275 5468 13309 5502
rect 13343 5468 13377 5502
rect 13411 5468 13445 5502
rect 13479 5468 13513 5502
rect 13547 5468 13581 5502
rect 13615 5468 13649 5502
rect 13683 5468 13717 5502
rect 13751 5468 13785 5502
rect 13819 5468 13853 5502
rect 13887 5468 13921 5502
rect 13955 5468 13989 5502
rect 14023 5468 14057 5502
rect 14091 5468 14125 5502
rect 14159 5468 14193 5502
rect 14227 5468 14261 5502
rect 14295 5468 14329 5502
rect 14363 5468 14397 5502
rect 14431 5468 14465 5502
rect 14499 5468 14533 5502
rect 14567 5468 14601 5502
rect 14635 5468 14669 5502
rect 14703 5468 14737 5502
rect 14771 5468 14805 5502
rect 14839 5468 14873 5502
rect 14907 5468 14949 5502
rect 14983 5468 15000 5502
rect 13054 5466 15000 5468
rect 13000 5439 15000 5466
rect 13000 5433 13077 5439
rect 5440 2572 5546 2606
rect 5580 2572 5614 2606
rect 5648 2572 5682 2606
rect 5716 2572 5750 2606
rect 5784 2572 5818 2606
rect 5852 2572 5886 2606
rect 5920 2572 5954 2606
rect 5988 2572 6022 2606
rect 6056 2572 6090 2606
rect 6124 2572 6158 2606
rect 6192 2572 6226 2606
rect 6260 2572 6294 2606
rect 6328 2572 6362 2606
rect 6396 2572 6430 2606
rect 6464 2572 6498 2606
rect 6532 2572 6566 2606
rect 6600 2572 6634 2606
rect 6668 2572 6702 2606
rect 6736 2572 6770 2606
rect 6804 2572 6838 2606
rect 6872 2572 6906 2606
rect 6940 2572 6974 2606
rect 7008 2572 7042 2606
rect 7076 2572 7110 2606
rect 7144 2572 7178 2606
rect 7212 2572 7246 2606
rect 7280 2572 7314 2606
rect 7348 2572 7382 2606
rect 7416 2572 7450 2606
rect 7484 2572 7518 2606
rect 7552 2572 7586 2606
rect 7620 2572 7654 2606
rect 7688 2572 7722 2606
rect 7756 2572 7790 2606
rect 7824 2572 7858 2606
rect 7892 2572 7926 2606
rect 7960 2572 7994 2606
rect 8028 2572 8062 2606
rect 8096 2572 8130 2606
rect 8164 2572 8198 2606
rect 8232 2572 8266 2606
rect 8300 2572 8334 2606
rect 8368 2572 8402 2606
rect 8436 2572 8470 2606
rect 8504 2572 8538 2606
rect 8572 2572 8606 2606
rect 8640 2572 8674 2606
rect 8708 2572 8742 2606
rect 8776 2572 8810 2606
rect 8844 2572 8878 2606
rect 8912 2572 8946 2606
rect 8980 2572 9014 2606
rect 9048 2572 9082 2606
rect 9116 2572 9150 2606
rect 9184 2572 9218 2606
rect 9252 2572 9286 2606
rect 9320 2572 9354 2606
rect 9388 2572 9422 2606
rect 9456 2572 9490 2606
rect 9524 2572 9558 2606
rect 9592 2572 9626 2606
rect 9660 2572 9694 2606
rect 9728 2572 9762 2606
rect 9796 2572 9830 2606
rect 9864 2572 9898 2606
rect 9932 2572 9966 2606
rect 10000 2572 10034 2606
rect 10068 2572 10102 2606
rect 10136 2572 10170 2606
rect 10204 2572 10238 2606
rect 10272 2572 10306 2606
rect 10340 2572 10374 2606
rect 10408 2572 10442 2606
rect 10476 2572 10510 2606
rect 10544 2572 10578 2606
rect 10612 2572 10646 2606
rect 10680 2572 10714 2606
rect 10748 2572 10782 2606
rect 10816 2572 10850 2606
rect 10884 2572 10918 2606
rect 10952 2572 10986 2606
rect 11020 2572 11054 2606
rect 11088 2572 11122 2606
rect 11156 2572 11190 2606
rect 11224 2572 11258 2606
rect 11292 2572 11326 2606
rect 11360 2572 11394 2606
rect 11428 2572 11462 2606
rect 11496 2572 11530 2606
rect 11564 2572 11598 2606
rect 11632 2572 11666 2606
rect 11700 2572 11734 2606
rect 11768 2572 11802 2606
rect 11836 2572 11870 2606
rect 11904 2572 11938 2606
rect 11972 2572 12006 2606
rect 12040 2572 12074 2606
rect 12108 2572 12142 2606
rect 12176 2572 12210 2606
rect 12244 2572 12278 2606
rect 12312 2572 12346 2606
rect 12380 2572 12414 2606
rect 12448 2572 12482 2606
rect 12516 2572 12550 2606
rect 12584 2572 12618 2606
rect 12652 2572 12686 2606
rect 12720 2572 12754 2606
rect 12788 2572 12822 2606
rect 12856 2572 12890 2606
rect 12924 2572 12958 2606
rect 12992 2572 13026 2606
rect 13060 2572 13094 2606
rect 13128 2572 13162 2606
rect 13196 2572 13230 2606
rect 13264 2572 13298 2606
rect 13332 2572 13366 2606
rect 13400 2572 13434 2606
rect 13468 2572 13502 2606
rect 13536 2572 13570 2606
rect 13604 2572 13638 2606
rect 13672 2572 13706 2606
rect 13740 2572 13774 2606
rect 13808 2572 13842 2606
rect 13876 2572 13910 2606
rect 13944 2572 13978 2606
rect 14012 2572 14046 2606
rect 14080 2572 14114 2606
rect 14148 2572 14182 2606
rect 14216 2572 14250 2606
rect 14284 2572 14318 2606
rect 14352 2572 14386 2606
rect 14420 2572 14454 2606
rect 14488 2572 14522 2606
rect 14556 2572 14590 2606
rect 14624 2572 14658 2606
rect 14692 2572 14726 2606
rect 14760 2572 14794 2606
rect 14828 2572 14862 2606
rect 14896 2572 14930 2606
rect 14964 2572 14998 2606
rect 15032 2572 15066 2606
rect 15100 2572 15134 2606
rect 15168 2572 15202 2606
rect 15236 2572 15270 2606
rect 15304 2572 15338 2606
rect 15372 2572 15406 2606
rect 15440 2572 15474 2606
rect 15508 2572 15542 2606
rect 15576 2572 15610 2606
rect 15644 2572 15678 2606
rect 15712 2572 15746 2606
rect 15780 2572 15814 2606
rect 15848 2572 15882 2606
rect 15916 2572 15950 2606
rect 15984 2572 16018 2606
rect 16052 2572 16086 2606
rect 16120 2572 16154 2606
rect 16188 2572 16222 2606
rect 16256 2572 16290 2606
rect 16324 2572 16358 2606
rect 16392 2572 16426 2606
rect 16460 2572 16494 2606
rect 16528 2572 16562 2606
rect 16596 2572 16630 2606
rect 16664 2572 16698 2606
rect 16732 2572 16766 2606
rect 16800 2572 16834 2606
rect 16868 2572 16902 2606
rect 16936 2572 16970 2606
rect 17004 2572 17038 2606
rect 17072 2572 17106 2606
rect 17140 2572 17174 2606
rect 17208 2572 17242 2606
rect 17276 2572 17310 2606
rect 17344 2572 17378 2606
rect 17412 2572 17446 2606
rect 17480 2572 17514 2606
rect 17548 2572 17582 2606
rect 17616 2572 17650 2606
rect 17684 2572 17718 2606
rect 17752 2572 17786 2606
rect 17820 2572 17854 2606
rect 17888 2572 17922 2606
rect 17956 2572 17990 2606
rect 18024 2572 18058 2606
rect 18092 2572 18126 2606
rect 18160 2572 18194 2606
rect 18228 2572 18262 2606
rect 18296 2572 18330 2606
rect 18364 2572 18398 2606
rect 18432 2572 18466 2606
rect 18500 2572 18534 2606
rect 18568 2572 18602 2606
rect 18636 2572 18670 2606
rect 18704 2572 18738 2606
rect 18772 2572 18806 2606
rect 18840 2572 18874 2606
rect 18908 2572 18942 2606
rect 18976 2572 19010 2606
rect 19044 2572 19078 2606
rect 19112 2572 19146 2606
rect 19180 2572 19214 2606
rect 19248 2572 19282 2606
rect 19316 2572 19350 2606
rect 19384 2572 19418 2606
rect 19452 2572 19486 2606
rect 19520 2572 19554 2606
rect 19588 2572 19622 2606
rect 19656 2572 19690 2606
rect 19724 2572 19758 2606
rect 19792 2572 19826 2606
rect 19860 2572 19894 2606
rect 19928 2572 19962 2606
rect 19996 2572 20030 2606
rect 20064 2572 20098 2606
rect 20132 2572 20166 2606
rect 20200 2572 20234 2606
rect 20268 2572 20302 2606
rect 20336 2572 20370 2606
rect 20404 2572 20438 2606
rect 20472 2572 20506 2606
rect 20540 2572 20574 2606
rect 20608 2572 20642 2606
rect 20676 2572 20710 2606
rect 20744 2572 20778 2606
rect 20812 2572 20846 2606
rect 20880 2572 20914 2606
rect 20948 2572 20982 2606
rect 21016 2572 21050 2606
rect 21084 2572 21118 2606
rect 21152 2572 21186 2606
rect 21220 2572 21254 2606
rect 21288 2572 21322 2606
rect 21356 2572 21390 2606
rect 21424 2572 21458 2606
rect 21492 2572 21526 2606
rect 21560 2572 21594 2606
rect 21628 2572 21662 2606
rect 21696 2572 21730 2606
rect 21764 2572 21798 2606
rect 21832 2572 21866 2606
rect 21900 2572 21934 2606
rect 21968 2572 22002 2606
rect 22036 2572 22070 2606
rect 22104 2572 22138 2606
rect 22172 2572 22206 2606
rect 22240 2572 22274 2606
rect 22308 2572 22342 2606
rect 22376 2572 22410 2606
rect 22444 2572 22478 2606
rect 22512 2572 22546 2606
rect 22580 2572 22614 2606
rect 22648 2572 22682 2606
rect 22716 2572 22750 2606
rect 22784 2572 22818 2606
rect 22852 2572 22886 2606
rect 22920 2572 22954 2606
rect 22988 2572 23022 2606
rect 23056 2572 23090 2606
rect 23124 2572 23158 2606
rect 23192 2572 23226 2606
rect 23260 2572 23294 2606
rect 23328 2572 23362 2606
rect 23396 2572 23430 2606
rect 23464 2572 23498 2606
rect 23532 2572 23566 2606
rect 23600 2572 23634 2606
rect 23668 2572 23702 2606
rect 23736 2572 23770 2606
rect 23804 2572 23838 2606
rect 23872 2572 23906 2606
rect 23940 2572 23974 2606
rect 24008 2572 24042 2606
rect 24076 2572 24110 2606
rect 24144 2572 24178 2606
rect 24212 2572 24246 2606
rect 24280 2572 24314 2606
rect 24348 2572 24382 2606
rect 24416 2572 24450 2606
rect 24484 2572 24518 2606
rect 24552 2572 24586 2606
rect 24620 2572 24654 2606
rect 24688 2572 24722 2606
rect 24756 2572 24790 2606
rect 24824 2572 24858 2606
rect 24892 2572 24926 2606
rect 24960 2572 24994 2606
rect 25028 2572 25062 2606
rect 25096 2572 25130 2606
rect 25164 2572 25198 2606
rect 25232 2572 25266 2606
rect 25300 2572 25334 2606
rect 25368 2572 25402 2606
rect 25436 2572 25470 2606
rect 25504 2572 25538 2606
rect 25572 2572 25606 2606
rect 25640 2572 25674 2606
rect 25708 2572 25742 2606
rect 25776 2572 25810 2606
rect 25844 2572 25878 2606
rect 25912 2572 25946 2606
rect 25980 2572 26014 2606
rect 26048 2572 26082 2606
rect 26116 2572 26150 2606
rect 26184 2572 26218 2606
rect 26252 2572 26286 2606
rect 26320 2572 26354 2606
rect 26388 2572 26422 2606
rect 26456 2572 26490 2606
rect 26524 2572 26558 2606
rect 26592 2572 26626 2606
rect 26660 2572 26694 2606
rect 26728 2572 26762 2606
rect 26796 2572 26830 2606
rect 26864 2572 26898 2606
rect 26932 2572 26966 2606
rect 27000 2572 27034 2606
rect 27068 2572 27102 2606
rect 27136 2572 27170 2606
rect 27204 2572 27238 2606
rect 27272 2572 27306 2606
rect 27340 2572 27374 2606
rect 27408 2572 27442 2606
rect 27476 2572 27510 2606
rect 27544 2572 27578 2606
rect 27612 2572 27646 2606
rect 27680 2572 27714 2606
rect 27748 2572 27782 2606
rect 27816 2572 27850 2606
rect 27884 2572 27918 2606
rect 27952 2572 27986 2606
rect 28020 2572 28054 2606
rect 28088 2572 28122 2606
rect 28156 2572 28190 2606
rect 28224 2572 28258 2606
rect 28292 2572 28326 2606
rect 28360 2572 28394 2606
rect 28428 2572 28462 2606
rect 28496 2572 28530 2606
rect 28564 2572 28598 2606
rect 28632 2572 28666 2606
rect 28700 2572 28734 2606
rect 28768 2572 28802 2606
rect 28836 2572 28870 2606
rect 28904 2572 28938 2606
rect 28972 2572 29006 2606
rect 29040 2572 29074 2606
rect 29108 2572 29142 2606
rect 29176 2572 29210 2606
rect 29244 2572 29278 2606
rect 29312 2572 29346 2606
rect 29380 2572 29414 2606
rect 29448 2572 29482 2606
rect 29516 2572 29550 2606
rect 29584 2572 29618 2606
rect 29652 2572 29686 2606
rect 29720 2572 29754 2606
rect 29788 2572 29822 2606
rect 29856 2572 29890 2606
rect 29924 2572 29958 2606
rect 29992 2572 30026 2606
rect 30060 2572 30094 2606
rect 30128 2572 30162 2606
rect 30196 2572 30230 2606
rect 30264 2572 30298 2606
rect 30332 2572 30366 2606
rect 30400 2572 30434 2606
rect 30468 2572 30502 2606
rect 30536 2572 30570 2606
rect 30604 2572 30638 2606
rect 30672 2572 30706 2606
rect 30740 2572 30774 2606
rect 30808 2572 30842 2606
rect 30876 2572 30910 2606
rect 30944 2572 30978 2606
rect 31012 2572 31046 2606
rect 31080 2572 31114 2606
rect 31148 2572 31182 2606
rect 31216 2572 31250 2606
rect 31284 2572 31318 2606
rect 31352 2572 31386 2606
rect 31420 2572 31454 2606
rect 31488 2572 31522 2606
rect 31556 2572 31590 2606
rect 31624 2572 31658 2606
rect 31692 2572 31726 2606
rect 31760 2572 31794 2606
rect 31828 2572 31862 2606
rect 31896 2572 31930 2606
rect 31964 2572 31998 2606
rect 32032 2572 32066 2606
rect 32100 2572 32134 2606
rect 32168 2572 32202 2606
rect 32236 2572 32270 2606
rect 32304 2572 32338 2606
rect 32372 2572 32406 2606
rect 32440 2572 32474 2606
rect 32508 2572 32542 2606
rect 32576 2572 32610 2606
rect 32644 2572 32678 2606
rect 32712 2572 32746 2606
rect 32780 2572 32814 2606
rect 32848 2572 32882 2606
rect 32916 2572 32950 2606
rect 32984 2572 33018 2606
rect 33052 2572 33086 2606
rect 33120 2572 33154 2606
rect 33188 2572 33222 2606
rect 33256 2572 33290 2606
rect 33324 2572 33358 2606
rect 33392 2572 33426 2606
rect 33460 2572 33494 2606
rect 33528 2572 33562 2606
rect 33596 2572 33630 2606
rect 33664 2572 33698 2606
rect 33732 2572 33766 2606
rect 33800 2572 33834 2606
rect 33868 2572 33902 2606
rect 33936 2572 33970 2606
rect 34004 2572 34038 2606
rect 34072 2572 34106 2606
rect 34140 2572 34174 2606
rect 34208 2572 34242 2606
rect 34276 2572 34310 2606
rect 34344 2572 34378 2606
rect 34412 2572 34446 2606
rect 34480 2572 34514 2606
rect 34548 2572 34582 2606
rect 34616 2572 34650 2606
rect 34684 2572 34718 2606
rect 34752 2572 34786 2606
rect 34820 2572 34854 2606
rect 34888 2572 34922 2606
rect 34956 2572 34990 2606
rect 35024 2572 35058 2606
rect 35092 2572 35126 2606
rect 35160 2572 35194 2606
rect 35228 2572 35262 2606
rect 35296 2572 35330 2606
rect 35364 2572 35398 2606
rect 35432 2572 35466 2606
rect 35500 2572 35534 2606
rect 35568 2572 35602 2606
rect 35636 2572 35670 2606
rect 35704 2572 35738 2606
rect 35772 2572 35806 2606
rect 35840 2572 35874 2606
rect 35908 2572 35942 2606
rect 35976 2572 36010 2606
rect 36044 2572 36078 2606
rect 36112 2572 36146 2606
rect 36180 2572 36214 2606
rect 36248 2572 36282 2606
rect 36316 2572 36350 2606
rect 36384 2572 36418 2606
rect 36452 2572 36486 2606
rect 36520 2572 36554 2606
rect 36588 2572 36622 2606
rect 36656 2572 36690 2606
rect 36724 2572 36758 2606
rect 36792 2572 36826 2606
rect 36860 2572 36894 2606
rect 36928 2572 36962 2606
rect 36996 2572 37030 2606
rect 37064 2572 37098 2606
rect 37132 2572 37166 2606
rect 37200 2572 37234 2606
rect 37268 2572 37302 2606
rect 37336 2572 37370 2606
rect 37404 2572 37438 2606
rect 37472 2572 37506 2606
rect 37540 2572 37574 2606
rect 37608 2572 37642 2606
rect 37676 2572 37710 2606
rect 37744 2572 37778 2606
rect 37812 2572 37846 2606
rect 37880 2572 37914 2606
rect 37948 2572 37982 2606
rect 38016 2572 38050 2606
rect 38084 2572 38118 2606
rect 38152 2572 38186 2606
rect 38220 2572 38254 2606
rect 38288 2572 38322 2606
rect 38356 2572 38390 2606
rect 38424 2572 38458 2606
rect 38492 2572 38526 2606
rect 38560 2572 38594 2606
rect 38628 2572 38662 2606
rect 38696 2572 38730 2606
rect 38764 2572 38798 2606
rect 38832 2572 38866 2606
rect 38900 2572 38934 2606
rect 38968 2572 39002 2606
rect 39036 2572 39070 2606
rect 39104 2572 39138 2606
rect 39172 2572 39206 2606
rect 39240 2572 39274 2606
rect 39308 2572 39342 2606
rect 39376 2572 39410 2606
rect 39444 2572 39478 2606
rect 39512 2572 39546 2606
rect 39580 2572 39614 2606
rect 39648 2572 39682 2606
rect 39716 2572 39750 2606
rect 39784 2572 39818 2606
rect 39852 2572 39886 2606
rect 39920 2572 39954 2606
rect 39988 2572 40022 2606
rect 40056 2572 40090 2606
rect 40124 2572 40158 2606
rect 40192 2572 40226 2606
rect 40260 2572 40294 2606
rect 40328 2572 40362 2606
rect 40396 2572 40430 2606
rect 40464 2572 40498 2606
rect 40532 2572 40566 2606
rect 40600 2572 40634 2606
rect 40668 2572 40702 2606
rect 40736 2572 40770 2606
rect 40804 2572 40838 2606
rect 40872 2572 40906 2606
rect 40940 2572 40974 2606
rect 41008 2572 41042 2606
rect 41076 2572 41110 2606
rect 41144 2572 41178 2606
rect 41212 2572 41246 2606
rect 41280 2572 41314 2606
rect 41348 2572 41382 2606
rect 41416 2572 41450 2606
rect 41484 2572 41518 2606
rect 41552 2572 41586 2606
rect 41620 2572 41654 2606
rect 41688 2572 41722 2606
rect 41756 2572 41790 2606
rect 41824 2572 41896 2606
rect 5440 2484 5474 2572
rect 5440 2416 5474 2450
rect 5440 2348 5474 2382
rect 5440 2280 5474 2314
rect 5440 2212 5474 2246
rect 5440 2144 5474 2178
rect 5440 2076 5474 2110
rect 5440 2008 5474 2042
rect 5440 1940 5474 1974
rect 5440 1872 5474 1906
rect 5440 1804 5474 1838
rect 5440 1736 5474 1770
rect 5440 1668 5474 1702
rect 5440 1600 5474 1634
rect 5440 1532 5474 1566
rect 5440 1464 5474 1498
rect 5440 1396 5474 1430
rect 5440 1328 5474 1362
rect 5440 1260 5474 1294
rect 5440 1192 5474 1226
rect 5440 1124 5474 1158
rect 5440 1056 5474 1090
rect 5440 988 5474 1022
rect 5440 920 5474 954
rect 5440 852 5474 886
rect 5440 784 5474 818
rect 5440 716 5474 750
rect 5440 648 5474 682
rect 5440 580 5474 614
rect 5440 458 5474 546
rect 22324 465 23410 470
rect 11401 458 12487 463
rect 15028 458 16114 461
rect 18681 458 19767 460
rect 22324 458 22346 465
rect 22380 458 22418 465
rect 22452 458 22490 465
rect 22524 458 22562 465
rect 22596 458 22634 465
rect 22668 458 22706 465
rect 22740 458 22778 465
rect 22812 458 22850 465
rect 22884 458 22922 465
rect 22956 458 22994 465
rect 23028 458 23066 465
rect 23100 458 23138 465
rect 23172 458 23210 465
rect 23244 458 23282 465
rect 23316 458 23354 465
rect 23388 458 23410 465
rect 25949 460 27035 465
rect 33227 460 34313 465
rect 25949 458 25971 460
rect 26005 458 26043 460
rect 26077 458 26115 460
rect 26149 458 26187 460
rect 26221 458 26259 460
rect 26293 458 26331 460
rect 26365 458 26403 460
rect 26437 458 26475 460
rect 26509 458 26547 460
rect 26581 458 26619 460
rect 26653 458 26691 460
rect 26725 458 26763 460
rect 26797 458 26835 460
rect 26869 458 26907 460
rect 26941 458 26979 460
rect 27013 458 27035 460
rect 29580 458 30666 460
rect 33227 458 33249 460
rect 33283 458 33321 460
rect 33355 458 33393 460
rect 33427 458 33465 460
rect 33499 458 33537 460
rect 33571 458 33609 460
rect 33643 458 33681 460
rect 33715 458 33753 460
rect 33787 458 33825 460
rect 33859 458 33897 460
rect 33931 458 33969 460
rect 34003 458 34041 460
rect 34075 458 34113 460
rect 34147 458 34185 460
rect 34219 458 34257 460
rect 34291 458 34313 460
rect 36856 462 37942 467
rect 36856 458 36878 462
rect 36912 458 36950 462
rect 36984 458 37022 462
rect 37056 458 37094 462
rect 37128 458 37166 462
rect 37200 458 37238 462
rect 37272 458 37310 462
rect 37344 458 37382 462
rect 37416 458 37454 462
rect 37488 458 37526 462
rect 37560 458 37598 462
rect 37632 458 37670 462
rect 37704 458 37742 462
rect 37776 458 37814 462
rect 37848 458 37886 462
rect 37920 458 37942 462
rect 40551 458 41637 461
rect 5440 424 5546 458
rect 5580 424 5614 458
rect 5648 424 5682 458
rect 5716 424 5750 458
rect 5784 424 5818 458
rect 5852 424 5886 458
rect 5920 424 5954 458
rect 5988 424 6022 458
rect 6056 424 6090 458
rect 6124 424 6158 458
rect 6192 424 6226 458
rect 6260 424 6294 458
rect 6328 424 6362 458
rect 6396 424 6430 458
rect 6464 424 6498 458
rect 6532 424 6566 458
rect 6600 424 6634 458
rect 6668 424 6702 458
rect 6736 424 6770 458
rect 6804 424 6838 458
rect 6872 424 6906 458
rect 6940 424 6974 458
rect 7008 424 7042 458
rect 7076 424 7110 458
rect 7144 424 7178 458
rect 7212 424 7246 458
rect 7280 424 7314 458
rect 7348 424 7382 458
rect 7416 424 7450 458
rect 7484 424 7518 458
rect 7552 424 7586 458
rect 7620 424 7654 458
rect 7688 424 7722 458
rect 7756 453 7790 458
rect 7824 453 7858 458
rect 7892 453 7926 458
rect 7960 453 7994 458
rect 8028 453 8062 458
rect 7756 424 7772 453
rect 7824 424 7844 453
rect 7892 424 7916 453
rect 7960 424 7988 453
rect 8028 424 8060 453
rect 8096 424 8130 458
rect 8164 453 8198 458
rect 8232 453 8266 458
rect 8300 453 8334 458
rect 8368 453 8402 458
rect 8436 453 8470 458
rect 8504 453 8538 458
rect 8572 453 8606 458
rect 8640 453 8674 458
rect 8166 424 8198 453
rect 8238 424 8266 453
rect 8310 424 8334 453
rect 8382 424 8402 453
rect 8454 424 8470 453
rect 8526 424 8538 453
rect 8598 424 8606 453
rect 8670 424 8674 453
rect 8708 453 8742 458
rect 7750 419 7772 424
rect 7806 419 7844 424
rect 7878 419 7916 424
rect 7950 419 7988 424
rect 8022 419 8060 424
rect 8094 419 8132 424
rect 8166 419 8204 424
rect 8238 419 8276 424
rect 8310 419 8348 424
rect 8382 419 8420 424
rect 8454 419 8492 424
rect 8526 419 8564 424
rect 8598 419 8636 424
rect 8670 419 8708 424
rect 8776 453 8810 458
rect 8776 424 8780 453
rect 8844 424 8878 458
rect 8912 424 8946 458
rect 8980 424 9014 458
rect 9048 424 9082 458
rect 9116 424 9150 458
rect 9184 424 9218 458
rect 9252 424 9286 458
rect 9320 424 9354 458
rect 9388 424 9422 458
rect 9456 424 9490 458
rect 9524 424 9558 458
rect 9592 424 9626 458
rect 9660 424 9694 458
rect 9728 424 9762 458
rect 9796 424 9830 458
rect 9864 424 9898 458
rect 9932 424 9966 458
rect 10000 424 10034 458
rect 10068 424 10102 458
rect 10136 424 10170 458
rect 10204 424 10238 458
rect 10272 424 10306 458
rect 10340 424 10374 458
rect 10408 424 10442 458
rect 10476 424 10510 458
rect 10544 424 10578 458
rect 10612 424 10646 458
rect 10680 424 10714 458
rect 10748 424 10782 458
rect 10816 424 10850 458
rect 10884 424 10918 458
rect 10952 424 10986 458
rect 11020 424 11054 458
rect 11088 424 11122 458
rect 11156 424 11190 458
rect 11224 424 11258 458
rect 11292 424 11326 458
rect 11360 424 11394 458
rect 11457 424 11462 458
rect 11529 424 11530 458
rect 11564 424 11567 458
rect 11632 424 11639 458
rect 11700 424 11711 458
rect 11768 424 11783 458
rect 11836 424 11855 458
rect 11904 424 11927 458
rect 11972 424 11999 458
rect 12040 424 12071 458
rect 12108 424 12142 458
rect 12177 424 12210 458
rect 12249 424 12278 458
rect 12321 424 12346 458
rect 12393 424 12414 458
rect 12465 424 12482 458
rect 12516 424 12550 458
rect 12584 424 12618 458
rect 12652 424 12686 458
rect 12720 424 12754 458
rect 12788 424 12822 458
rect 12856 424 12890 458
rect 12924 424 12958 458
rect 12992 424 13026 458
rect 13060 424 13094 458
rect 13128 424 13162 458
rect 13196 424 13230 458
rect 13264 424 13298 458
rect 13332 424 13366 458
rect 13400 424 13434 458
rect 13468 424 13502 458
rect 13536 424 13570 458
rect 13604 424 13638 458
rect 13672 424 13706 458
rect 13740 424 13774 458
rect 13808 424 13842 458
rect 13876 424 13910 458
rect 13944 424 13978 458
rect 14012 424 14046 458
rect 14080 424 14114 458
rect 14148 424 14182 458
rect 14216 424 14250 458
rect 14284 424 14318 458
rect 14352 424 14386 458
rect 14420 424 14454 458
rect 14488 424 14522 458
rect 14556 424 14590 458
rect 14624 424 14658 458
rect 14692 424 14726 458
rect 14760 424 14794 458
rect 14828 424 14862 458
rect 14896 424 14930 458
rect 14964 424 14998 458
rect 15032 456 15066 458
rect 15100 456 15134 458
rect 15168 456 15202 458
rect 15236 456 15270 458
rect 15032 424 15050 456
rect 15100 424 15122 456
rect 15168 424 15194 456
rect 15236 424 15266 456
rect 15304 424 15338 458
rect 15372 424 15406 458
rect 15440 456 15474 458
rect 15508 456 15542 458
rect 15576 456 15610 458
rect 15644 456 15678 458
rect 15712 456 15746 458
rect 15780 456 15814 458
rect 15848 456 15882 458
rect 15916 456 15950 458
rect 15444 424 15474 456
rect 15516 424 15542 456
rect 15588 424 15610 456
rect 15660 424 15678 456
rect 15732 424 15746 456
rect 15804 424 15814 456
rect 15876 424 15882 456
rect 15948 424 15950 456
rect 15984 456 16018 458
rect 16052 456 16086 458
rect 15984 424 15986 456
rect 16052 424 16058 456
rect 16120 424 16154 458
rect 16188 424 16222 458
rect 16256 424 16290 458
rect 16324 424 16358 458
rect 16392 424 16426 458
rect 16460 424 16494 458
rect 16528 424 16562 458
rect 16596 424 16630 458
rect 16664 424 16698 458
rect 16732 424 16766 458
rect 16800 424 16834 458
rect 16868 424 16902 458
rect 16936 424 16970 458
rect 17004 424 17038 458
rect 17072 424 17106 458
rect 17140 424 17174 458
rect 17208 424 17242 458
rect 17276 424 17310 458
rect 17344 424 17378 458
rect 17412 424 17446 458
rect 17480 424 17514 458
rect 17548 424 17582 458
rect 17616 424 17650 458
rect 17684 424 17718 458
rect 17752 424 17786 458
rect 17820 424 17854 458
rect 17888 424 17922 458
rect 17956 424 17990 458
rect 18024 424 18058 458
rect 18092 424 18126 458
rect 18160 424 18194 458
rect 18228 424 18262 458
rect 18296 424 18330 458
rect 18364 424 18398 458
rect 18432 424 18466 458
rect 18500 424 18534 458
rect 18568 424 18602 458
rect 18636 424 18670 458
rect 18704 455 18738 458
rect 18737 424 18738 455
rect 18772 455 18806 458
rect 18840 455 18874 458
rect 18908 455 18942 458
rect 18976 455 19010 458
rect 19044 455 19078 458
rect 19112 455 19146 458
rect 19180 455 19214 458
rect 19248 455 19282 458
rect 18772 424 18775 455
rect 18840 424 18847 455
rect 18908 424 18919 455
rect 18976 424 18991 455
rect 19044 424 19063 455
rect 19112 424 19135 455
rect 19180 424 19207 455
rect 19248 424 19279 455
rect 19316 424 19350 458
rect 19384 455 19418 458
rect 19452 455 19486 458
rect 19520 455 19554 458
rect 19588 455 19622 458
rect 19656 455 19690 458
rect 19724 455 19758 458
rect 19385 424 19418 455
rect 19457 424 19486 455
rect 19529 424 19554 455
rect 19601 424 19622 455
rect 19673 424 19690 455
rect 19745 424 19758 455
rect 19792 424 19826 458
rect 19860 424 19894 458
rect 19928 424 19962 458
rect 19996 424 20030 458
rect 20064 424 20098 458
rect 20132 424 20166 458
rect 20200 424 20234 458
rect 20268 424 20302 458
rect 20336 424 20370 458
rect 20404 424 20438 458
rect 20472 424 20506 458
rect 20540 424 20574 458
rect 20608 424 20642 458
rect 20676 424 20710 458
rect 20744 424 20778 458
rect 20812 424 20846 458
rect 20880 424 20914 458
rect 20948 424 20982 458
rect 21016 424 21050 458
rect 21084 424 21118 458
rect 21152 424 21186 458
rect 21220 424 21254 458
rect 21288 424 21322 458
rect 21356 424 21390 458
rect 21424 424 21458 458
rect 21492 424 21526 458
rect 21560 424 21594 458
rect 21628 424 21662 458
rect 21696 424 21730 458
rect 21764 424 21798 458
rect 21832 424 21866 458
rect 21900 424 21934 458
rect 21968 424 22002 458
rect 22036 424 22070 458
rect 22104 424 22138 458
rect 22172 424 22206 458
rect 22240 424 22274 458
rect 22308 424 22342 458
rect 22380 431 22410 458
rect 22452 431 22478 458
rect 22524 431 22546 458
rect 22596 431 22614 458
rect 22668 431 22682 458
rect 22740 431 22750 458
rect 22812 431 22818 458
rect 22884 431 22886 458
rect 22376 424 22410 431
rect 22444 424 22478 431
rect 22512 424 22546 431
rect 22580 424 22614 431
rect 22648 424 22682 431
rect 22716 424 22750 431
rect 22784 424 22818 431
rect 22852 424 22886 431
rect 22920 431 22922 458
rect 22988 431 22994 458
rect 23056 431 23066 458
rect 23124 431 23138 458
rect 23192 431 23210 458
rect 23260 431 23282 458
rect 23328 431 23354 458
rect 22920 424 22954 431
rect 22988 424 23022 431
rect 23056 424 23090 431
rect 23124 424 23158 431
rect 23192 424 23226 431
rect 23260 424 23294 431
rect 23328 424 23362 431
rect 23396 424 23430 458
rect 23464 424 23498 458
rect 23532 424 23566 458
rect 23600 424 23634 458
rect 23668 424 23702 458
rect 23736 424 23770 458
rect 23804 424 23838 458
rect 23872 424 23906 458
rect 23940 424 23974 458
rect 24008 424 24042 458
rect 24076 424 24110 458
rect 24144 424 24178 458
rect 24212 424 24246 458
rect 24280 424 24314 458
rect 24348 424 24382 458
rect 24416 424 24450 458
rect 24484 424 24518 458
rect 24552 424 24586 458
rect 24620 424 24654 458
rect 24688 424 24722 458
rect 24756 424 24790 458
rect 24824 424 24858 458
rect 24892 424 24926 458
rect 24960 424 24994 458
rect 25028 424 25062 458
rect 25096 424 25130 458
rect 25164 424 25198 458
rect 25232 424 25266 458
rect 25300 424 25334 458
rect 25368 424 25402 458
rect 25436 424 25470 458
rect 25504 424 25538 458
rect 25572 424 25606 458
rect 25640 424 25674 458
rect 25708 424 25742 458
rect 25776 424 25810 458
rect 25844 424 25878 458
rect 25912 424 25946 458
rect 26005 426 26014 458
rect 26077 426 26082 458
rect 26149 426 26150 458
rect 25980 424 26014 426
rect 26048 424 26082 426
rect 26116 424 26150 426
rect 26184 426 26187 458
rect 26252 426 26259 458
rect 26320 426 26331 458
rect 26388 426 26403 458
rect 26456 426 26475 458
rect 26524 426 26547 458
rect 26592 426 26619 458
rect 26660 426 26691 458
rect 26184 424 26218 426
rect 26252 424 26286 426
rect 26320 424 26354 426
rect 26388 424 26422 426
rect 26456 424 26490 426
rect 26524 424 26558 426
rect 26592 424 26626 426
rect 26660 424 26694 426
rect 26728 424 26762 458
rect 26797 426 26830 458
rect 26869 426 26898 458
rect 26941 426 26966 458
rect 27013 426 27034 458
rect 26796 424 26830 426
rect 26864 424 26898 426
rect 26932 424 26966 426
rect 27000 424 27034 426
rect 27068 424 27102 458
rect 27136 424 27170 458
rect 27204 424 27238 458
rect 27272 424 27306 458
rect 27340 424 27374 458
rect 27408 424 27442 458
rect 27476 424 27510 458
rect 27544 424 27578 458
rect 27612 424 27646 458
rect 27680 424 27714 458
rect 27748 424 27782 458
rect 27816 424 27850 458
rect 27884 424 27918 458
rect 27952 424 27986 458
rect 28020 424 28054 458
rect 28088 424 28122 458
rect 28156 424 28190 458
rect 28224 424 28258 458
rect 28292 424 28326 458
rect 28360 424 28394 458
rect 28428 424 28462 458
rect 28496 424 28530 458
rect 28564 424 28598 458
rect 28632 424 28666 458
rect 28700 424 28734 458
rect 28768 424 28802 458
rect 28836 424 28870 458
rect 28904 424 28938 458
rect 28972 424 29006 458
rect 29040 424 29074 458
rect 29108 424 29142 458
rect 29176 424 29210 458
rect 29244 424 29278 458
rect 29312 424 29346 458
rect 29380 424 29414 458
rect 29448 424 29482 458
rect 29516 424 29550 458
rect 29584 455 29618 458
rect 29652 455 29686 458
rect 29720 455 29754 458
rect 29788 455 29822 458
rect 29584 424 29602 455
rect 29652 424 29674 455
rect 29720 424 29746 455
rect 29788 424 29818 455
rect 29856 424 29890 458
rect 29924 424 29958 458
rect 29992 455 30026 458
rect 30060 455 30094 458
rect 30128 455 30162 458
rect 30196 455 30230 458
rect 30264 455 30298 458
rect 30332 455 30366 458
rect 30400 455 30434 458
rect 30468 455 30502 458
rect 29996 424 30026 455
rect 30068 424 30094 455
rect 30140 424 30162 455
rect 30212 424 30230 455
rect 30284 424 30298 455
rect 30356 424 30366 455
rect 30428 424 30434 455
rect 30500 424 30502 455
rect 30536 455 30570 458
rect 30604 455 30638 458
rect 30536 424 30538 455
rect 30604 424 30610 455
rect 30672 424 30706 458
rect 30740 424 30774 458
rect 30808 424 30842 458
rect 30876 424 30910 458
rect 30944 424 30978 458
rect 31012 424 31046 458
rect 31080 424 31114 458
rect 31148 424 31182 458
rect 31216 424 31250 458
rect 31284 424 31318 458
rect 31352 424 31386 458
rect 31420 424 31454 458
rect 31488 424 31522 458
rect 31556 424 31590 458
rect 31624 424 31658 458
rect 31692 424 31726 458
rect 31760 424 31794 458
rect 31828 424 31862 458
rect 31896 424 31930 458
rect 31964 424 31998 458
rect 32032 424 32066 458
rect 32100 424 32134 458
rect 32168 424 32202 458
rect 32236 424 32270 458
rect 32304 424 32338 458
rect 32372 424 32406 458
rect 32440 424 32474 458
rect 32508 424 32542 458
rect 32576 424 32610 458
rect 32644 424 32678 458
rect 32712 424 32746 458
rect 32780 424 32814 458
rect 32848 424 32882 458
rect 32916 424 32950 458
rect 32984 424 33018 458
rect 33052 424 33086 458
rect 33120 424 33154 458
rect 33188 424 33222 458
rect 33283 426 33290 458
rect 33355 426 33358 458
rect 33256 424 33290 426
rect 33324 424 33358 426
rect 33392 426 33393 458
rect 33460 426 33465 458
rect 33528 426 33537 458
rect 33596 426 33609 458
rect 33664 426 33681 458
rect 33732 426 33753 458
rect 33800 426 33825 458
rect 33868 426 33897 458
rect 33936 426 33969 458
rect 33392 424 33426 426
rect 33460 424 33494 426
rect 33528 424 33562 426
rect 33596 424 33630 426
rect 33664 424 33698 426
rect 33732 424 33766 426
rect 33800 424 33834 426
rect 33868 424 33902 426
rect 33936 424 33970 426
rect 34004 424 34038 458
rect 34075 426 34106 458
rect 34147 426 34174 458
rect 34219 426 34242 458
rect 34291 426 34310 458
rect 34072 424 34106 426
rect 34140 424 34174 426
rect 34208 424 34242 426
rect 34276 424 34310 426
rect 34344 424 34378 458
rect 34412 424 34446 458
rect 34480 424 34514 458
rect 34548 424 34582 458
rect 34616 424 34650 458
rect 34684 424 34718 458
rect 34752 424 34786 458
rect 34820 424 34854 458
rect 34888 424 34922 458
rect 34956 424 34990 458
rect 35024 424 35058 458
rect 35092 424 35126 458
rect 35160 424 35194 458
rect 35228 424 35262 458
rect 35296 424 35330 458
rect 35364 424 35398 458
rect 35432 424 35466 458
rect 35500 424 35534 458
rect 35568 424 35602 458
rect 35636 424 35670 458
rect 35704 424 35738 458
rect 35772 424 35806 458
rect 35840 424 35874 458
rect 35908 424 35942 458
rect 35976 424 36010 458
rect 36044 424 36078 458
rect 36112 424 36146 458
rect 36180 424 36214 458
rect 36248 424 36282 458
rect 36316 424 36350 458
rect 36384 424 36418 458
rect 36452 424 36486 458
rect 36520 424 36554 458
rect 36588 424 36622 458
rect 36656 424 36690 458
rect 36724 424 36758 458
rect 36792 424 36826 458
rect 36860 428 36878 458
rect 36928 428 36950 458
rect 36996 428 37022 458
rect 37064 428 37094 458
rect 36860 424 36894 428
rect 36928 424 36962 428
rect 36996 424 37030 428
rect 37064 424 37098 428
rect 37132 424 37166 458
rect 37200 424 37234 458
rect 37272 428 37302 458
rect 37344 428 37370 458
rect 37416 428 37438 458
rect 37488 428 37506 458
rect 37560 428 37574 458
rect 37632 428 37642 458
rect 37704 428 37710 458
rect 37776 428 37778 458
rect 37268 424 37302 428
rect 37336 424 37370 428
rect 37404 424 37438 428
rect 37472 424 37506 428
rect 37540 424 37574 428
rect 37608 424 37642 428
rect 37676 424 37710 428
rect 37744 424 37778 428
rect 37812 428 37814 458
rect 37880 428 37886 458
rect 37812 424 37846 428
rect 37880 424 37914 428
rect 37948 424 37982 458
rect 38016 424 38050 458
rect 38084 424 38118 458
rect 38152 424 38186 458
rect 38220 424 38254 458
rect 38288 424 38322 458
rect 38356 424 38390 458
rect 38424 424 38458 458
rect 38492 424 38526 458
rect 38560 424 38594 458
rect 38628 424 38662 458
rect 38696 424 38730 458
rect 38764 424 38798 458
rect 38832 424 38866 458
rect 38900 424 38934 458
rect 38968 424 39002 458
rect 39036 424 39070 458
rect 39104 424 39138 458
rect 39172 424 39206 458
rect 39240 424 39274 458
rect 39308 424 39342 458
rect 39376 424 39410 458
rect 39444 424 39478 458
rect 39512 424 39546 458
rect 39580 424 39614 458
rect 39648 424 39682 458
rect 39716 424 39750 458
rect 39784 424 39818 458
rect 39852 424 39886 458
rect 39920 424 39954 458
rect 39988 424 40022 458
rect 40056 424 40090 458
rect 40124 424 40158 458
rect 40192 424 40226 458
rect 40260 424 40294 458
rect 40328 424 40362 458
rect 40396 424 40430 458
rect 40464 424 40498 458
rect 40532 424 40566 458
rect 40600 456 40634 458
rect 40668 456 40702 458
rect 40736 456 40770 458
rect 40804 456 40838 458
rect 40872 456 40906 458
rect 40940 456 40974 458
rect 41008 456 41042 458
rect 40607 424 40634 456
rect 40679 424 40702 456
rect 40751 424 40770 456
rect 40823 424 40838 456
rect 40895 424 40906 456
rect 40967 424 40974 456
rect 41039 424 41042 456
rect 41076 456 41110 458
rect 41144 456 41178 458
rect 41212 456 41246 458
rect 41280 456 41314 458
rect 41348 456 41382 458
rect 41416 456 41450 458
rect 41484 456 41518 458
rect 41552 456 41586 458
rect 41076 424 41077 456
rect 41144 424 41149 456
rect 41212 424 41221 456
rect 41280 424 41293 456
rect 41348 424 41365 456
rect 41416 424 41437 456
rect 41484 424 41509 456
rect 41552 424 41581 456
rect 41620 424 41654 458
rect 41688 424 41722 458
rect 41756 424 41790 458
rect 41824 424 41896 458
rect 8742 419 8780 424
rect 8814 419 8836 424
rect 11401 420 12487 424
rect 15028 422 15050 424
rect 15084 422 15122 424
rect 15156 422 15194 424
rect 15228 422 15266 424
rect 15300 422 15338 424
rect 15372 422 15410 424
rect 15444 422 15482 424
rect 15516 422 15554 424
rect 15588 422 15626 424
rect 15660 422 15698 424
rect 15732 422 15770 424
rect 15804 422 15842 424
rect 15876 422 15914 424
rect 15948 422 15986 424
rect 16020 422 16058 424
rect 16092 422 16114 424
rect 7750 415 8836 419
rect 15028 418 16114 422
rect 18681 421 18703 424
rect 18737 421 18775 424
rect 18809 421 18847 424
rect 18881 421 18919 424
rect 18953 421 18991 424
rect 19025 421 19063 424
rect 19097 421 19135 424
rect 19169 421 19207 424
rect 19241 421 19279 424
rect 19313 421 19351 424
rect 19385 421 19423 424
rect 19457 421 19495 424
rect 19529 421 19567 424
rect 19601 421 19639 424
rect 19673 421 19711 424
rect 19745 421 19767 424
rect 25949 422 27035 424
rect 18681 417 19767 421
rect 29580 421 29602 424
rect 29636 421 29674 424
rect 29708 421 29746 424
rect 29780 421 29818 424
rect 29852 421 29890 424
rect 29924 421 29962 424
rect 29996 421 30034 424
rect 30068 421 30106 424
rect 30140 421 30178 424
rect 30212 421 30250 424
rect 30284 421 30322 424
rect 30356 421 30394 424
rect 30428 421 30466 424
rect 30500 421 30538 424
rect 30572 421 30610 424
rect 30644 421 30666 424
rect 33227 422 34313 424
rect 40551 422 40573 424
rect 40607 422 40645 424
rect 40679 422 40717 424
rect 40751 422 40789 424
rect 40823 422 40861 424
rect 40895 422 40933 424
rect 40967 422 41005 424
rect 41039 422 41077 424
rect 41111 422 41149 424
rect 41183 422 41221 424
rect 41255 422 41293 424
rect 41327 422 41365 424
rect 41399 422 41437 424
rect 41471 422 41509 424
rect 41543 422 41581 424
rect 41615 422 41637 424
rect 29580 417 30666 421
rect 40551 418 41637 422
<< viali >>
rect 12406 12503 14024 12753
rect 15858 12867 15892 12901
rect 15930 12867 15964 12901
rect 10789 11076 10823 11084
rect 10789 11050 10823 11076
rect 10789 11008 10823 11012
rect 10789 10978 10823 11008
rect 10789 10906 10823 10940
rect 10789 10838 10823 10868
rect 10789 10834 10823 10838
rect 10789 10770 10823 10796
rect 10789 10762 10823 10770
rect 15758 10856 15792 10890
rect 15830 10856 15864 10890
rect 15902 10856 15936 10890
rect 15974 10856 16008 10890
rect 16046 10856 16080 10890
rect 16118 10856 16152 10890
rect 5664 8511 5698 8542
rect 16895 9691 16929 9710
rect 16895 9676 16929 9691
rect 16895 9623 16929 9638
rect 16895 9604 16929 9623
rect 20367 9619 20396 9652
rect 20396 9619 20401 9652
rect 20367 9618 20401 9619
rect 16489 9323 16490 9344
rect 16490 9323 16523 9344
rect 16489 9310 16523 9323
rect 16489 9251 16490 9272
rect 16490 9251 16523 9272
rect 16489 9238 16523 9251
rect 11185 8646 11187 8665
rect 11187 8646 11219 8665
rect 11185 8631 11219 8646
rect 5664 8508 5698 8511
rect 5664 8436 5698 8470
rect 16889 8448 16891 8474
rect 16891 8448 16923 8474
rect 16889 8440 16923 8448
rect 10790 7943 10824 7963
rect 10790 7929 10791 7943
rect 10791 7929 10824 7943
rect 10790 7875 10824 7891
rect 10790 7857 10791 7875
rect 10791 7857 10824 7875
rect 16889 8398 16923 8402
rect 16889 8368 16891 8398
rect 16891 8368 16923 8398
rect 16479 7927 16484 7928
rect 16484 7927 16513 7928
rect 16479 7894 16513 7927
rect 16479 7855 16484 7856
rect 16484 7855 16513 7856
rect 16479 7822 16513 7855
rect 9719 6423 9753 6457
rect 9791 6423 9825 6457
rect 9863 6423 9897 6457
rect 9935 6423 9969 6457
rect 10007 6423 10041 6457
rect 10079 6423 10113 6457
rect 19284 9392 19318 9396
rect 19356 9392 19390 9396
rect 19284 9362 19307 9392
rect 19307 9362 19318 9392
rect 19356 9362 19380 9392
rect 19380 9362 19390 9392
rect 19959 9008 19993 9016
rect 19959 8982 19991 9008
rect 19991 8982 19993 9008
rect 20363 8288 20393 8300
rect 20393 8288 20397 8300
rect 20363 8266 20397 8288
rect 17444 7885 17477 7919
rect 17477 7885 17478 7919
rect 17516 7885 17519 7919
rect 17519 7885 17550 7919
rect 17588 7885 17621 7919
rect 17621 7885 17622 7919
rect 17660 7885 17689 7919
rect 17689 7885 17694 7919
rect 17732 7885 17757 7919
rect 17757 7885 17766 7919
rect 19953 7915 19987 7944
rect 19953 7910 19987 7915
rect 20373 7080 20407 7085
rect 20373 7051 20407 7080
rect 19959 6227 19993 6258
rect 19959 6224 19971 6227
rect 19971 6224 19993 6227
rect 11197 5653 11228 5665
rect 11228 5653 11231 5665
rect 11197 5631 11231 5653
rect 12449 5494 12481 5528
rect 12481 5494 12483 5528
rect 12521 5494 12549 5528
rect 12549 5494 12555 5528
rect 12593 5494 12617 5528
rect 12617 5494 12627 5528
rect 13017 5500 13051 5521
rect 13017 5487 13020 5500
rect 13020 5487 13051 5500
rect 22346 458 22380 465
rect 22418 458 22452 465
rect 22490 458 22524 465
rect 22562 458 22596 465
rect 22634 458 22668 465
rect 22706 458 22740 465
rect 22778 458 22812 465
rect 22850 458 22884 465
rect 22922 458 22956 465
rect 22994 458 23028 465
rect 23066 458 23100 465
rect 23138 458 23172 465
rect 23210 458 23244 465
rect 23282 458 23316 465
rect 23354 458 23388 465
rect 25971 458 26005 460
rect 26043 458 26077 460
rect 26115 458 26149 460
rect 26187 458 26221 460
rect 26259 458 26293 460
rect 26331 458 26365 460
rect 26403 458 26437 460
rect 26475 458 26509 460
rect 26547 458 26581 460
rect 26619 458 26653 460
rect 26691 458 26725 460
rect 26763 458 26797 460
rect 26835 458 26869 460
rect 26907 458 26941 460
rect 26979 458 27013 460
rect 33249 458 33283 460
rect 33321 458 33355 460
rect 33393 458 33427 460
rect 33465 458 33499 460
rect 33537 458 33571 460
rect 33609 458 33643 460
rect 33681 458 33715 460
rect 33753 458 33787 460
rect 33825 458 33859 460
rect 33897 458 33931 460
rect 33969 458 34003 460
rect 34041 458 34075 460
rect 34113 458 34147 460
rect 34185 458 34219 460
rect 34257 458 34291 460
rect 36878 458 36912 462
rect 36950 458 36984 462
rect 37022 458 37056 462
rect 37094 458 37128 462
rect 37166 458 37200 462
rect 37238 458 37272 462
rect 37310 458 37344 462
rect 37382 458 37416 462
rect 37454 458 37488 462
rect 37526 458 37560 462
rect 37598 458 37632 462
rect 37670 458 37704 462
rect 37742 458 37776 462
rect 37814 458 37848 462
rect 37886 458 37920 462
rect 7772 424 7790 453
rect 7790 424 7806 453
rect 7844 424 7858 453
rect 7858 424 7878 453
rect 7916 424 7926 453
rect 7926 424 7950 453
rect 7988 424 7994 453
rect 7994 424 8022 453
rect 8060 424 8062 453
rect 8062 424 8094 453
rect 8132 424 8164 453
rect 8164 424 8166 453
rect 8204 424 8232 453
rect 8232 424 8238 453
rect 8276 424 8300 453
rect 8300 424 8310 453
rect 8348 424 8368 453
rect 8368 424 8382 453
rect 8420 424 8436 453
rect 8436 424 8454 453
rect 8492 424 8504 453
rect 8504 424 8526 453
rect 8564 424 8572 453
rect 8572 424 8598 453
rect 8636 424 8640 453
rect 8640 424 8670 453
rect 7772 419 7806 424
rect 7844 419 7878 424
rect 7916 419 7950 424
rect 7988 419 8022 424
rect 8060 419 8094 424
rect 8132 419 8166 424
rect 8204 419 8238 424
rect 8276 419 8310 424
rect 8348 419 8382 424
rect 8420 419 8454 424
rect 8492 419 8526 424
rect 8564 419 8598 424
rect 8636 419 8670 424
rect 8708 419 8742 453
rect 8780 424 8810 453
rect 8810 424 8814 453
rect 11423 424 11428 458
rect 11428 424 11457 458
rect 11495 424 11496 458
rect 11496 424 11529 458
rect 11567 424 11598 458
rect 11598 424 11601 458
rect 11639 424 11666 458
rect 11666 424 11673 458
rect 11711 424 11734 458
rect 11734 424 11745 458
rect 11783 424 11802 458
rect 11802 424 11817 458
rect 11855 424 11870 458
rect 11870 424 11889 458
rect 11927 424 11938 458
rect 11938 424 11961 458
rect 11999 424 12006 458
rect 12006 424 12033 458
rect 12071 424 12074 458
rect 12074 424 12105 458
rect 12143 424 12176 458
rect 12176 424 12177 458
rect 12215 424 12244 458
rect 12244 424 12249 458
rect 12287 424 12312 458
rect 12312 424 12321 458
rect 12359 424 12380 458
rect 12380 424 12393 458
rect 12431 424 12448 458
rect 12448 424 12465 458
rect 15050 424 15066 456
rect 15066 424 15084 456
rect 15122 424 15134 456
rect 15134 424 15156 456
rect 15194 424 15202 456
rect 15202 424 15228 456
rect 15266 424 15270 456
rect 15270 424 15300 456
rect 15338 424 15372 456
rect 15410 424 15440 456
rect 15440 424 15444 456
rect 15482 424 15508 456
rect 15508 424 15516 456
rect 15554 424 15576 456
rect 15576 424 15588 456
rect 15626 424 15644 456
rect 15644 424 15660 456
rect 15698 424 15712 456
rect 15712 424 15732 456
rect 15770 424 15780 456
rect 15780 424 15804 456
rect 15842 424 15848 456
rect 15848 424 15876 456
rect 15914 424 15916 456
rect 15916 424 15948 456
rect 15986 424 16018 456
rect 16018 424 16020 456
rect 16058 424 16086 456
rect 16086 424 16092 456
rect 18703 424 18704 455
rect 18704 424 18737 455
rect 18775 424 18806 455
rect 18806 424 18809 455
rect 18847 424 18874 455
rect 18874 424 18881 455
rect 18919 424 18942 455
rect 18942 424 18953 455
rect 18991 424 19010 455
rect 19010 424 19025 455
rect 19063 424 19078 455
rect 19078 424 19097 455
rect 19135 424 19146 455
rect 19146 424 19169 455
rect 19207 424 19214 455
rect 19214 424 19241 455
rect 19279 424 19282 455
rect 19282 424 19313 455
rect 19351 424 19384 455
rect 19384 424 19385 455
rect 19423 424 19452 455
rect 19452 424 19457 455
rect 19495 424 19520 455
rect 19520 424 19529 455
rect 19567 424 19588 455
rect 19588 424 19601 455
rect 19639 424 19656 455
rect 19656 424 19673 455
rect 19711 424 19724 455
rect 19724 424 19745 455
rect 22346 431 22376 458
rect 22376 431 22380 458
rect 22418 431 22444 458
rect 22444 431 22452 458
rect 22490 431 22512 458
rect 22512 431 22524 458
rect 22562 431 22580 458
rect 22580 431 22596 458
rect 22634 431 22648 458
rect 22648 431 22668 458
rect 22706 431 22716 458
rect 22716 431 22740 458
rect 22778 431 22784 458
rect 22784 431 22812 458
rect 22850 431 22852 458
rect 22852 431 22884 458
rect 22922 431 22954 458
rect 22954 431 22956 458
rect 22994 431 23022 458
rect 23022 431 23028 458
rect 23066 431 23090 458
rect 23090 431 23100 458
rect 23138 431 23158 458
rect 23158 431 23172 458
rect 23210 431 23226 458
rect 23226 431 23244 458
rect 23282 431 23294 458
rect 23294 431 23316 458
rect 23354 431 23362 458
rect 23362 431 23388 458
rect 25971 426 25980 458
rect 25980 426 26005 458
rect 26043 426 26048 458
rect 26048 426 26077 458
rect 26115 426 26116 458
rect 26116 426 26149 458
rect 26187 426 26218 458
rect 26218 426 26221 458
rect 26259 426 26286 458
rect 26286 426 26293 458
rect 26331 426 26354 458
rect 26354 426 26365 458
rect 26403 426 26422 458
rect 26422 426 26437 458
rect 26475 426 26490 458
rect 26490 426 26509 458
rect 26547 426 26558 458
rect 26558 426 26581 458
rect 26619 426 26626 458
rect 26626 426 26653 458
rect 26691 426 26694 458
rect 26694 426 26725 458
rect 26763 426 26796 458
rect 26796 426 26797 458
rect 26835 426 26864 458
rect 26864 426 26869 458
rect 26907 426 26932 458
rect 26932 426 26941 458
rect 26979 426 27000 458
rect 27000 426 27013 458
rect 29602 424 29618 455
rect 29618 424 29636 455
rect 29674 424 29686 455
rect 29686 424 29708 455
rect 29746 424 29754 455
rect 29754 424 29780 455
rect 29818 424 29822 455
rect 29822 424 29852 455
rect 29890 424 29924 455
rect 29962 424 29992 455
rect 29992 424 29996 455
rect 30034 424 30060 455
rect 30060 424 30068 455
rect 30106 424 30128 455
rect 30128 424 30140 455
rect 30178 424 30196 455
rect 30196 424 30212 455
rect 30250 424 30264 455
rect 30264 424 30284 455
rect 30322 424 30332 455
rect 30332 424 30356 455
rect 30394 424 30400 455
rect 30400 424 30428 455
rect 30466 424 30468 455
rect 30468 424 30500 455
rect 30538 424 30570 455
rect 30570 424 30572 455
rect 30610 424 30638 455
rect 30638 424 30644 455
rect 33249 426 33256 458
rect 33256 426 33283 458
rect 33321 426 33324 458
rect 33324 426 33355 458
rect 33393 426 33426 458
rect 33426 426 33427 458
rect 33465 426 33494 458
rect 33494 426 33499 458
rect 33537 426 33562 458
rect 33562 426 33571 458
rect 33609 426 33630 458
rect 33630 426 33643 458
rect 33681 426 33698 458
rect 33698 426 33715 458
rect 33753 426 33766 458
rect 33766 426 33787 458
rect 33825 426 33834 458
rect 33834 426 33859 458
rect 33897 426 33902 458
rect 33902 426 33931 458
rect 33969 426 33970 458
rect 33970 426 34003 458
rect 34041 426 34072 458
rect 34072 426 34075 458
rect 34113 426 34140 458
rect 34140 426 34147 458
rect 34185 426 34208 458
rect 34208 426 34219 458
rect 34257 426 34276 458
rect 34276 426 34291 458
rect 36878 428 36894 458
rect 36894 428 36912 458
rect 36950 428 36962 458
rect 36962 428 36984 458
rect 37022 428 37030 458
rect 37030 428 37056 458
rect 37094 428 37098 458
rect 37098 428 37128 458
rect 37166 428 37200 458
rect 37238 428 37268 458
rect 37268 428 37272 458
rect 37310 428 37336 458
rect 37336 428 37344 458
rect 37382 428 37404 458
rect 37404 428 37416 458
rect 37454 428 37472 458
rect 37472 428 37488 458
rect 37526 428 37540 458
rect 37540 428 37560 458
rect 37598 428 37608 458
rect 37608 428 37632 458
rect 37670 428 37676 458
rect 37676 428 37704 458
rect 37742 428 37744 458
rect 37744 428 37776 458
rect 37814 428 37846 458
rect 37846 428 37848 458
rect 37886 428 37914 458
rect 37914 428 37920 458
rect 40573 424 40600 456
rect 40600 424 40607 456
rect 40645 424 40668 456
rect 40668 424 40679 456
rect 40717 424 40736 456
rect 40736 424 40751 456
rect 40789 424 40804 456
rect 40804 424 40823 456
rect 40861 424 40872 456
rect 40872 424 40895 456
rect 40933 424 40940 456
rect 40940 424 40967 456
rect 41005 424 41008 456
rect 41008 424 41039 456
rect 41077 424 41110 456
rect 41110 424 41111 456
rect 41149 424 41178 456
rect 41178 424 41183 456
rect 41221 424 41246 456
rect 41246 424 41255 456
rect 41293 424 41314 456
rect 41314 424 41327 456
rect 41365 424 41382 456
rect 41382 424 41399 456
rect 41437 424 41450 456
rect 41450 424 41471 456
rect 41509 424 41518 456
rect 41518 424 41543 456
rect 41581 424 41586 456
rect 41586 424 41615 456
rect 8780 419 8814 424
rect 15050 422 15084 424
rect 15122 422 15156 424
rect 15194 422 15228 424
rect 15266 422 15300 424
rect 15338 422 15372 424
rect 15410 422 15444 424
rect 15482 422 15516 424
rect 15554 422 15588 424
rect 15626 422 15660 424
rect 15698 422 15732 424
rect 15770 422 15804 424
rect 15842 422 15876 424
rect 15914 422 15948 424
rect 15986 422 16020 424
rect 16058 422 16092 424
rect 18703 421 18737 424
rect 18775 421 18809 424
rect 18847 421 18881 424
rect 18919 421 18953 424
rect 18991 421 19025 424
rect 19063 421 19097 424
rect 19135 421 19169 424
rect 19207 421 19241 424
rect 19279 421 19313 424
rect 19351 421 19385 424
rect 19423 421 19457 424
rect 19495 421 19529 424
rect 19567 421 19601 424
rect 19639 421 19673 424
rect 19711 421 19745 424
rect 29602 421 29636 424
rect 29674 421 29708 424
rect 29746 421 29780 424
rect 29818 421 29852 424
rect 29890 421 29924 424
rect 29962 421 29996 424
rect 30034 421 30068 424
rect 30106 421 30140 424
rect 30178 421 30212 424
rect 30250 421 30284 424
rect 30322 421 30356 424
rect 30394 421 30428 424
rect 30466 421 30500 424
rect 30538 421 30572 424
rect 30610 421 30644 424
rect 40573 422 40607 424
rect 40645 422 40679 424
rect 40717 422 40751 424
rect 40789 422 40823 424
rect 40861 422 40895 424
rect 40933 422 40967 424
rect 41005 422 41039 424
rect 41077 422 41111 424
rect 41149 422 41183 424
rect 41221 422 41255 424
rect 41293 422 41327 424
rect 41365 422 41399 424
rect 41437 422 41471 424
rect 41509 422 41543 424
rect 41581 422 41615 424
<< metal1 >>
rect 15842 12921 15994 12960
rect 10425 12902 12152 12906
rect 10425 12753 14210 12902
rect 15842 12867 15858 12921
rect 15910 12869 15922 12921
rect 15974 12869 15994 12921
rect 15892 12867 15930 12869
rect 15964 12867 15994 12869
rect 15842 12826 15994 12867
rect 10425 12503 12406 12753
rect 14024 12503 14210 12753
rect 10425 12380 14210 12503
rect 10425 11478 10595 12380
rect 12156 12370 14210 12380
rect 19709 12278 19810 12363
rect 15398 11478 15573 11482
rect 10425 11255 15576 11478
rect 10425 10964 10595 11255
rect 10774 11084 10838 11110
rect 10774 11050 10789 11084
rect 10823 11050 10838 11084
rect 10774 11012 10838 11050
rect 10774 10978 10789 11012
rect 10823 10978 10838 11012
rect 10774 10964 10838 10978
rect 10983 11024 11086 11034
rect 10983 10972 11009 11024
rect 11061 10972 11086 11024
rect 10983 10967 11086 10972
rect 10425 10940 10838 10964
rect 10425 10906 10789 10940
rect 10823 10906 10838 10940
rect 10425 10868 10838 10906
rect 10425 10834 10789 10868
rect 10823 10834 10838 10868
rect 10425 10810 10838 10834
rect 15398 10937 15573 11255
rect 15398 10890 16519 10937
rect 15398 10856 15758 10890
rect 15792 10856 15830 10890
rect 15864 10856 15902 10890
rect 15936 10856 15974 10890
rect 16008 10856 16046 10890
rect 16080 10856 16118 10890
rect 16152 10856 16519 10890
rect 15398 10817 16519 10856
rect 15398 10815 15573 10817
rect 4417 8586 5486 8587
rect 4417 8542 5746 8586
rect 4417 8508 5664 8542
rect 5698 8508 5746 8542
rect 4417 8470 5746 8508
rect 4417 8436 5664 8470
rect 5698 8436 5746 8470
rect 4417 8398 5746 8436
rect 4417 5140 5153 8398
rect 10425 7987 10595 10810
rect 10774 10796 10838 10810
rect 10774 10762 10789 10796
rect 10823 10762 10838 10796
rect 10774 10736 10838 10762
rect 16333 10111 16519 10817
rect 16333 10109 17650 10111
rect 16333 10107 18381 10109
rect 16333 10103 19462 10107
rect 16333 9985 20702 10103
rect 16339 9983 20702 9985
rect 17070 9981 20702 9983
rect 16671 9797 16761 9813
rect 16671 9745 16689 9797
rect 16741 9745 16761 9797
rect 16671 9732 16761 9745
rect 16882 9710 16944 9724
rect 16882 9676 16895 9710
rect 16929 9676 16944 9710
rect 16882 9647 16944 9676
rect 17078 9647 17179 9981
rect 18151 9979 20702 9981
rect 19255 9976 20702 9979
rect 16880 9638 17179 9647
rect 16880 9604 16895 9638
rect 16929 9604 17179 9638
rect 16880 9591 17179 9604
rect 17078 9572 17179 9591
rect 16442 9345 16554 9360
rect 16442 9293 16480 9345
rect 16532 9293 16554 9345
rect 16442 9281 16554 9293
rect 16442 9229 16480 9281
rect 16532 9229 16554 9281
rect 16442 9216 16554 9229
rect 16648 8904 16758 8914
rect 16648 8852 16676 8904
rect 16728 8852 16758 8904
rect 16648 8842 16758 8852
rect 10966 8749 11073 8760
rect 10966 8697 10983 8749
rect 11035 8697 11073 8749
rect 10966 8688 11073 8697
rect 11160 8665 11634 8710
rect 11160 8631 11185 8665
rect 11219 8631 11634 8665
rect 11160 8584 11634 8631
rect 10967 8025 11073 8033
rect 10425 7963 10842 7987
rect 10967 7973 10993 8025
rect 11045 7973 11073 8025
rect 10967 7967 11073 7973
rect 6050 7863 6163 7937
rect 10425 7929 10790 7963
rect 10824 7929 10842 7963
rect 10425 7891 10842 7929
rect 10425 7857 10790 7891
rect 10824 7857 10842 7891
rect 10425 7833 10842 7857
rect 10425 6861 10595 7833
rect 10425 6860 10592 6861
rect 10422 6678 10592 6860
rect 10422 6677 10587 6678
rect 10420 6503 10587 6677
rect 9679 6457 10587 6503
rect 9679 6423 9719 6457
rect 9753 6423 9791 6457
rect 9825 6423 9863 6457
rect 9897 6423 9935 6457
rect 9969 6423 10007 6457
rect 10041 6423 10079 6457
rect 10113 6423 10587 6457
rect 9679 6374 10587 6423
rect 10420 5330 10587 6374
rect 10943 5758 11058 5768
rect 10943 5706 10975 5758
rect 11027 5706 11058 5758
rect 11508 5717 11634 8584
rect 17081 8491 17177 9572
rect 19256 9410 19387 9976
rect 20589 9974 20702 9976
rect 20589 9904 20703 9974
rect 20139 9798 20221 9813
rect 20139 9746 20154 9798
rect 20206 9746 20221 9798
rect 20139 9732 20221 9746
rect 20589 9683 20704 9904
rect 20343 9652 20704 9683
rect 20343 9618 20367 9652
rect 20401 9618 20704 9652
rect 20343 9587 20704 9618
rect 17438 9372 18239 9408
rect 17438 9130 17482 9372
rect 17595 9298 17731 9313
rect 17595 9246 17636 9298
rect 17688 9246 17731 9298
rect 17595 9232 17731 9246
rect 17759 9298 17837 9301
rect 17759 9246 17771 9298
rect 17823 9246 17837 9298
rect 17759 9240 17837 9246
rect 17759 9212 17821 9240
rect 17759 9068 17820 9212
rect 18202 8948 18239 9372
rect 19256 9396 19414 9410
rect 19256 9362 19284 9396
rect 19318 9362 19356 9396
rect 19390 9362 19414 9396
rect 19256 9345 19414 9362
rect 18942 9286 19099 9312
rect 18942 9234 18960 9286
rect 19012 9234 19024 9286
rect 19076 9234 19099 9286
rect 18942 9212 19099 9234
rect 17591 8905 18239 8948
rect 19377 8943 19414 9345
rect 19590 9016 20033 9064
rect 19590 8982 19959 9016
rect 19993 8982 20033 9016
rect 17591 8904 18061 8905
rect 16874 8474 17177 8491
rect 16874 8440 16889 8474
rect 16923 8440 17177 8474
rect 16874 8428 17177 8440
rect 16641 8408 16737 8425
rect 16641 8356 16664 8408
rect 16716 8356 16737 8408
rect 16641 8340 16737 8356
rect 16874 8402 16940 8428
rect 17081 8427 17177 8428
rect 17538 8718 17686 8720
rect 17538 8697 17689 8718
rect 17538 8645 17590 8697
rect 17642 8645 17689 8697
rect 17538 8633 17689 8645
rect 17538 8581 17590 8633
rect 17642 8581 17689 8633
rect 17538 8569 17689 8581
rect 17538 8517 17590 8569
rect 17642 8517 17689 8569
rect 17538 8505 17689 8517
rect 17538 8453 17590 8505
rect 17642 8453 17689 8505
rect 17538 8441 17689 8453
rect 16874 8368 16889 8402
rect 16923 8368 16940 8402
rect 16874 8344 16940 8368
rect 17538 8389 17590 8441
rect 17642 8389 17689 8441
rect 17538 8365 17689 8389
rect 17538 8359 17686 8365
rect 16446 7940 16548 7964
rect 16446 7888 16471 7940
rect 16523 7888 16548 7940
rect 16446 7876 16548 7888
rect 16446 7824 16471 7876
rect 16523 7824 16548 7876
rect 16446 7822 16479 7824
rect 16513 7822 16548 7824
rect 16446 7798 16548 7822
rect 17399 7929 17623 7942
rect 18202 7929 18238 8905
rect 18995 8903 19416 8943
rect 19590 8921 20033 8982
rect 19590 8847 19782 8921
rect 20133 8902 20217 8914
rect 20133 8850 20151 8902
rect 20203 8850 20217 8902
rect 19591 8001 19781 8847
rect 20133 8839 20217 8850
rect 20137 8454 20214 8466
rect 20137 8402 20149 8454
rect 20201 8402 20214 8454
rect 20137 8395 20214 8402
rect 20589 8334 20704 9587
rect 20339 8300 20704 8334
rect 20339 8266 20363 8300
rect 20397 8266 20704 8300
rect 20339 8238 20704 8266
rect 19591 7944 20033 8001
rect 17399 7919 18241 7929
rect 17399 7885 17444 7919
rect 17478 7885 17516 7919
rect 17550 7885 17588 7919
rect 17622 7885 17660 7919
rect 17694 7885 17732 7919
rect 17766 7885 18241 7919
rect 17399 7879 18241 7885
rect 19591 7910 19953 7944
rect 19987 7910 20033 7944
rect 17399 7870 18240 7879
rect 16636 7502 16766 7520
rect 16636 7450 16673 7502
rect 16725 7450 16766 7502
rect 16636 7435 16766 7450
rect 12514 5769 12591 5770
rect 12507 5758 12591 5769
rect 10943 5697 11058 5706
rect 11174 5665 11636 5717
rect 12507 5706 12529 5758
rect 12581 5706 12591 5758
rect 12507 5697 12591 5706
rect 14797 5722 14882 5738
rect 11174 5631 11197 5665
rect 11231 5631 11636 5665
rect 14797 5670 14803 5722
rect 14855 5670 14882 5722
rect 14797 5656 14882 5670
rect 11174 5591 11636 5631
rect 10420 5278 10478 5330
rect 10530 5278 10587 5330
rect 10420 5246 10587 5278
rect 11508 5140 11634 5591
rect 12416 5544 12512 5546
rect 12414 5532 12666 5544
rect 12414 5480 12436 5532
rect 12488 5528 12666 5532
rect 12488 5494 12521 5528
rect 12555 5494 12593 5528
rect 12627 5494 12666 5528
rect 12488 5480 12666 5494
rect 12985 5521 13088 5566
rect 12985 5487 13017 5521
rect 13051 5487 13088 5521
rect 12416 5479 12512 5480
rect 4412 5138 11676 5140
rect 12985 5139 13088 5487
rect 17399 5163 17623 7870
rect 19591 7858 20033 7910
rect 19591 6304 19781 7858
rect 20132 7559 20222 7577
rect 20132 7507 20150 7559
rect 20202 7507 20222 7559
rect 20132 7487 20222 7507
rect 20152 7213 20231 7223
rect 20152 7161 20165 7213
rect 20217 7161 20231 7213
rect 20152 7152 20231 7161
rect 20354 7120 20426 7122
rect 20589 7120 20704 8238
rect 20351 7085 20704 7120
rect 20351 7051 20373 7085
rect 20407 7051 20704 7085
rect 20351 7042 20704 7051
rect 20351 7041 20692 7042
rect 20354 7010 20426 7041
rect 20146 6315 20231 6331
rect 19591 6258 20025 6304
rect 19591 6224 19959 6258
rect 19993 6224 20025 6258
rect 20146 6263 20163 6315
rect 20215 6263 20231 6315
rect 20146 6248 20231 6263
rect 19591 6161 20025 6224
rect 19591 5163 19781 6161
rect 27240 5376 27403 5404
rect 22419 5317 22547 5350
rect 22419 5265 22456 5317
rect 22508 5265 22547 5317
rect 23408 5313 23517 5337
rect 22846 5266 23087 5311
rect 22419 5233 22547 5265
rect 23408 5261 23437 5313
rect 23489 5261 23517 5313
rect 23408 5235 23517 5261
rect 27240 5260 27262 5376
rect 27378 5260 27403 5376
rect 15841 5142 15999 5147
rect 17399 5142 19781 5163
rect 15841 5140 19781 5142
rect 14520 5139 19781 5140
rect 12985 5138 19781 5139
rect 4412 5100 19781 5138
rect 4412 5048 15862 5100
rect 15914 5048 15926 5100
rect 15978 5048 19781 5100
rect 27240 5093 27403 5260
rect 4412 5013 19781 5048
rect 4412 5008 19743 5013
rect 4417 -474 5153 5008
rect 11508 5006 19743 5008
rect 11508 5004 17457 5006
rect 11508 5002 15999 5004
rect 11508 5001 14552 5002
rect 11594 5000 13088 5001
rect 15841 4998 15999 5002
rect 27239 569 27403 5093
rect 22324 465 23410 470
rect 11401 458 12487 463
rect 7750 453 8836 458
rect 7750 419 7772 453
rect 7806 419 7844 453
rect 7878 419 7916 453
rect 7950 419 7988 453
rect 8022 419 8060 453
rect 8094 419 8132 453
rect 8166 419 8204 453
rect 8238 419 8276 453
rect 8310 419 8348 453
rect 8382 419 8420 453
rect 8454 419 8492 453
rect 8526 419 8564 453
rect 8598 419 8636 453
rect 8670 419 8708 453
rect 8742 419 8780 453
rect 8814 419 8836 453
rect 11401 424 11423 458
rect 11457 424 11495 458
rect 11529 424 11567 458
rect 11601 424 11639 458
rect 11673 424 11711 458
rect 11745 424 11783 458
rect 11817 424 11855 458
rect 11889 424 11927 458
rect 11961 424 11999 458
rect 12033 424 12071 458
rect 12105 424 12143 458
rect 12177 424 12215 458
rect 12249 424 12287 458
rect 12321 424 12359 458
rect 12393 424 12431 458
rect 12465 424 12487 458
rect 11401 420 12487 424
rect 15028 456 16114 461
rect 15028 422 15050 456
rect 15084 422 15122 456
rect 15156 422 15194 456
rect 15228 422 15266 456
rect 15300 422 15338 456
rect 15372 422 15410 456
rect 15444 422 15482 456
rect 15516 422 15554 456
rect 15588 422 15626 456
rect 15660 422 15698 456
rect 15732 422 15770 456
rect 15804 422 15842 456
rect 15876 422 15914 456
rect 15948 422 15986 456
rect 16020 422 16058 456
rect 16092 422 16114 456
rect 7750 415 8836 419
rect 15028 418 16114 422
rect 18681 455 19767 460
rect 18681 421 18703 455
rect 18737 421 18775 455
rect 18809 421 18847 455
rect 18881 421 18919 455
rect 18953 421 18991 455
rect 19025 421 19063 455
rect 19097 421 19135 455
rect 19169 421 19207 455
rect 19241 421 19279 455
rect 19313 421 19351 455
rect 19385 421 19423 455
rect 19457 421 19495 455
rect 19529 421 19567 455
rect 19601 421 19639 455
rect 19673 421 19711 455
rect 19745 421 19767 455
rect 22324 431 22346 465
rect 22380 431 22418 465
rect 22452 431 22490 465
rect 22524 431 22562 465
rect 22596 431 22634 465
rect 22668 431 22706 465
rect 22740 431 22778 465
rect 22812 431 22850 465
rect 22884 431 22922 465
rect 22956 431 22994 465
rect 23028 431 23066 465
rect 23100 431 23138 465
rect 23172 431 23210 465
rect 23244 431 23282 465
rect 23316 431 23354 465
rect 23388 431 23410 465
rect 22324 427 23410 431
rect 25949 460 27035 465
rect 33227 460 34313 465
rect 25949 426 25971 460
rect 26005 426 26043 460
rect 26077 426 26115 460
rect 26149 426 26187 460
rect 26221 426 26259 460
rect 26293 426 26331 460
rect 26365 426 26403 460
rect 26437 426 26475 460
rect 26509 426 26547 460
rect 26581 426 26619 460
rect 26653 426 26691 460
rect 26725 426 26763 460
rect 26797 426 26835 460
rect 26869 426 26907 460
rect 26941 426 26979 460
rect 27013 426 27035 460
rect 25949 422 27035 426
rect 29580 455 30666 460
rect 18681 417 19767 421
rect 29580 421 29602 455
rect 29636 421 29674 455
rect 29708 421 29746 455
rect 29780 421 29818 455
rect 29852 421 29890 455
rect 29924 421 29962 455
rect 29996 421 30034 455
rect 30068 421 30106 455
rect 30140 421 30178 455
rect 30212 421 30250 455
rect 30284 421 30322 455
rect 30356 421 30394 455
rect 30428 421 30466 455
rect 30500 421 30538 455
rect 30572 421 30610 455
rect 30644 421 30666 455
rect 33227 426 33249 460
rect 33283 426 33321 460
rect 33355 426 33393 460
rect 33427 426 33465 460
rect 33499 426 33537 460
rect 33571 426 33609 460
rect 33643 426 33681 460
rect 33715 426 33753 460
rect 33787 426 33825 460
rect 33859 426 33897 460
rect 33931 426 33969 460
rect 34003 426 34041 460
rect 34075 426 34113 460
rect 34147 426 34185 460
rect 34219 426 34257 460
rect 34291 426 34313 460
rect 33227 422 34313 426
rect 36856 462 37942 467
rect 36856 428 36878 462
rect 36912 428 36950 462
rect 36984 428 37022 462
rect 37056 428 37094 462
rect 37128 428 37166 462
rect 37200 428 37238 462
rect 37272 428 37310 462
rect 37344 428 37382 462
rect 37416 428 37454 462
rect 37488 428 37526 462
rect 37560 428 37598 462
rect 37632 428 37670 462
rect 37704 428 37742 462
rect 37776 428 37814 462
rect 37848 428 37886 462
rect 37920 428 37942 462
rect 36856 424 37942 428
rect 40551 456 41637 461
rect 40551 422 40573 456
rect 40607 422 40645 456
rect 40679 422 40717 456
rect 40751 422 40789 456
rect 40823 422 40861 456
rect 40895 422 40933 456
rect 40967 422 41005 456
rect 41039 422 41077 456
rect 41111 422 41149 456
rect 41183 422 41221 456
rect 41255 422 41293 456
rect 41327 422 41365 456
rect 41399 422 41437 456
rect 41471 422 41509 456
rect 41543 422 41581 456
rect 41615 422 41637 456
rect 29580 417 30666 421
rect 40551 418 41637 422
rect 4417 -543 5171 -474
rect 4417 -1107 4514 -543
rect 5078 -1107 5171 -543
rect 4417 -1169 5171 -1107
<< via1 >>
rect 15858 12901 15910 12921
rect 15858 12869 15892 12901
rect 15892 12869 15910 12901
rect 15922 12901 15974 12921
rect 15922 12869 15930 12901
rect 15930 12869 15964 12901
rect 15964 12869 15974 12901
rect 11009 10972 11061 11024
rect 16689 9745 16741 9797
rect 16480 9344 16532 9345
rect 16480 9310 16489 9344
rect 16489 9310 16523 9344
rect 16523 9310 16532 9344
rect 16480 9293 16532 9310
rect 16480 9272 16532 9281
rect 16480 9238 16489 9272
rect 16489 9238 16523 9272
rect 16523 9238 16532 9272
rect 16480 9229 16532 9238
rect 16676 8852 16728 8904
rect 10983 8697 11035 8749
rect 10993 7973 11045 8025
rect 10975 5706 11027 5758
rect 20154 9746 20206 9798
rect 17636 9246 17688 9298
rect 17771 9246 17823 9298
rect 18960 9234 19012 9286
rect 19024 9234 19076 9286
rect 16664 8356 16716 8408
rect 17590 8645 17642 8697
rect 17590 8581 17642 8633
rect 17590 8517 17642 8569
rect 17590 8453 17642 8505
rect 17590 8389 17642 8441
rect 16471 7928 16523 7940
rect 16471 7894 16479 7928
rect 16479 7894 16513 7928
rect 16513 7894 16523 7928
rect 16471 7888 16523 7894
rect 16471 7856 16523 7876
rect 16471 7824 16479 7856
rect 16479 7824 16513 7856
rect 16513 7824 16523 7856
rect 20151 8850 20203 8902
rect 20149 8402 20201 8454
rect 16673 7450 16725 7502
rect 12529 5706 12581 5758
rect 14803 5670 14855 5722
rect 10478 5278 10530 5330
rect 12436 5528 12488 5532
rect 12436 5494 12449 5528
rect 12449 5494 12483 5528
rect 12483 5494 12488 5528
rect 12436 5480 12488 5494
rect 20150 7507 20202 7559
rect 20165 7161 20217 7213
rect 20163 6263 20215 6315
rect 22456 5265 22508 5317
rect 23437 5261 23489 5313
rect 27262 5260 27378 5376
rect 15862 5048 15914 5100
rect 15926 5048 15978 5100
rect 4514 -1107 5078 -543
<< metal2 >>
rect 15842 12921 15994 12960
rect 15842 12869 15858 12921
rect 15910 12869 15922 12921
rect 15974 12869 15994 12921
rect 10983 11028 11086 11034
rect 10983 10972 11007 11028
rect 11063 10972 11086 11028
rect 10983 10967 11086 10972
rect 11033 10359 11114 10400
rect 11033 10303 11034 10359
rect 11090 10303 11114 10359
rect 11033 10279 11114 10303
rect 11033 10223 11034 10279
rect 11090 10223 11114 10279
rect 11033 10199 11114 10223
rect 11033 10143 11034 10199
rect 11090 10143 11114 10199
rect 11033 10119 11114 10143
rect 11033 10063 11034 10119
rect 11090 10063 11114 10119
rect 11033 10039 11114 10063
rect 11033 9983 11034 10039
rect 11090 9983 11114 10039
rect 11033 9959 11114 9983
rect 11033 9903 11034 9959
rect 11090 9903 11114 9959
rect 11033 9879 11114 9903
rect 11033 9823 11034 9879
rect 11090 9823 11114 9879
rect 11033 9799 11114 9823
rect 11033 9743 11034 9799
rect 11090 9743 11114 9799
rect 11033 9719 11114 9743
rect 11033 9663 11034 9719
rect 11090 9663 11114 9719
rect 11033 9639 11114 9663
rect 11033 9583 11034 9639
rect 11090 9583 11114 9639
rect 11033 9559 11114 9583
rect 11033 9503 11034 9559
rect 11090 9503 11114 9559
rect 11033 9479 11114 9503
rect 11033 9423 11034 9479
rect 11090 9423 11114 9479
rect 11033 9399 11114 9423
rect 11033 9343 11034 9399
rect 11090 9343 11114 9399
rect 11033 9319 11114 9343
rect 11033 9263 11034 9319
rect 11090 9263 11114 9319
rect 11033 9239 11114 9263
rect 10918 9168 10966 9228
rect 11033 9183 11034 9239
rect 11090 9183 11114 9239
rect 15842 9360 15994 12869
rect 16192 11613 16327 11643
rect 16192 11557 16230 11613
rect 16286 11557 16327 11613
rect 16192 11531 16327 11557
rect 16801 11591 16904 11637
rect 16801 11535 16826 11591
rect 16882 11535 16904 11591
rect 16801 11487 16904 11535
rect 18943 10553 19099 10591
rect 18943 10497 18991 10553
rect 19047 10497 19099 10553
rect 16671 9799 16761 9813
rect 16671 9743 16687 9799
rect 16743 9743 16761 9799
rect 16671 9732 16761 9743
rect 17759 9799 17837 9813
rect 17759 9743 17769 9799
rect 17825 9743 17837 9799
rect 15842 9345 16554 9360
rect 15842 9293 16480 9345
rect 16532 9293 16554 9345
rect 15842 9281 16554 9293
rect 15842 9229 16480 9281
rect 16532 9229 16554 9281
rect 17595 9300 17731 9313
rect 17595 9244 17634 9300
rect 17690 9244 17731 9300
rect 17595 9232 17731 9244
rect 17759 9298 17837 9743
rect 18943 9313 19099 10497
rect 20139 9800 20221 9813
rect 20139 9744 20152 9800
rect 20208 9744 20221 9800
rect 20139 9732 20221 9744
rect 19626 9314 19703 9315
rect 19543 9313 19704 9314
rect 17759 9246 17771 9298
rect 17823 9246 17837 9298
rect 17759 9240 17837 9246
rect 18941 9286 19704 9313
rect 18941 9234 18960 9286
rect 19012 9234 19024 9286
rect 19076 9234 19704 9286
rect 15842 9216 16554 9229
rect 11033 9159 11114 9183
rect 11033 9103 11034 9159
rect 11090 9103 11114 9159
rect 11033 9079 11114 9103
rect 11033 9023 11034 9079
rect 11090 9023 11114 9079
rect 11033 8999 11114 9023
rect 11033 8943 11034 8999
rect 11090 8943 11114 8999
rect 11033 8919 11114 8943
rect 11033 8863 11034 8919
rect 11090 8863 11114 8919
rect 11033 8842 11114 8863
rect 11076 8799 11114 8842
rect 10966 8749 11073 8760
rect 10966 8697 10983 8749
rect 11035 8747 11073 8749
rect 10966 8691 10990 8697
rect 11046 8691 11073 8747
rect 10966 8679 11073 8691
rect 10967 8037 11073 8051
rect 15844 8047 16002 9216
rect 18941 9214 19704 9234
rect 18941 9213 19548 9214
rect 18943 9212 19099 9213
rect 16609 9113 16692 9147
rect 16609 9057 16626 9113
rect 16682 9057 16692 9113
rect 16609 9033 16692 9057
rect 16609 8977 16626 9033
rect 16682 8977 16692 9033
rect 16609 8946 16692 8977
rect 16726 9115 16826 9149
rect 16726 9059 16759 9115
rect 16815 9059 16826 9115
rect 16726 9035 16826 9059
rect 16726 8979 16759 9035
rect 16815 8979 16826 9035
rect 16726 8946 16826 8979
rect 17631 9022 17713 9033
rect 17631 8966 17644 9022
rect 17700 8966 17713 9022
rect 17631 8956 17713 8966
rect 19626 8914 19703 9214
rect 20076 9131 20095 9140
rect 20076 9096 20150 9131
rect 20076 9040 20091 9096
rect 20147 9040 20150 9096
rect 20076 9006 20150 9040
rect 20196 9128 20326 9162
rect 20196 9072 20245 9128
rect 20301 9072 20326 9128
rect 20196 9048 20326 9072
rect 20076 8997 20095 9006
rect 20196 8992 20245 9048
rect 20301 8992 20326 9048
rect 20196 8962 20326 8992
rect 16648 8904 16758 8914
rect 16648 8852 16676 8904
rect 16728 8852 16758 8904
rect 19626 8902 20217 8914
rect 16648 8815 16758 8852
rect 16648 8759 16673 8815
rect 16729 8759 16758 8815
rect 17974 8847 18099 8876
rect 17974 8791 18006 8847
rect 18062 8791 18099 8847
rect 17974 8763 18099 8791
rect 18770 8837 18887 8864
rect 19626 8850 20151 8902
rect 20203 8850 20217 8902
rect 18770 8781 18798 8837
rect 18854 8781 18887 8837
rect 16648 8734 16758 8759
rect 18770 8758 18887 8781
rect 19136 8827 19244 8846
rect 19136 8771 19160 8827
rect 19216 8771 19244 8827
rect 19136 8753 19244 8771
rect 19626 8839 20217 8850
rect 17538 8718 17686 8720
rect 17538 8697 17689 8718
rect 17538 8691 17590 8697
rect 17642 8691 17689 8697
rect 17538 8635 17588 8691
rect 17644 8635 17689 8691
rect 17538 8633 17689 8635
rect 17538 8611 17590 8633
rect 17642 8611 17689 8633
rect 17538 8555 17588 8611
rect 17644 8555 17689 8611
rect 17538 8531 17590 8555
rect 17642 8531 17689 8555
rect 18354 8553 18395 8597
rect 17538 8475 17588 8531
rect 17644 8475 17689 8531
rect 17538 8453 17590 8475
rect 17642 8453 17689 8475
rect 17538 8451 17689 8453
rect 16641 8410 16737 8425
rect 16641 8354 16660 8410
rect 16716 8354 16737 8410
rect 17538 8395 17588 8451
rect 17644 8395 17689 8451
rect 17538 8389 17590 8395
rect 17642 8389 17689 8395
rect 17538 8365 17689 8389
rect 17538 8359 17686 8365
rect 16641 8340 16737 8354
rect 10967 7981 10991 8037
rect 11047 7981 11073 8037
rect 10967 7973 10993 7981
rect 11045 7973 11073 7981
rect 10967 7967 11073 7973
rect 15843 7964 16002 8047
rect 15843 7940 16548 7964
rect 15843 7888 16471 7940
rect 16523 7888 16548 7940
rect 15843 7876 16548 7888
rect 15843 7824 16471 7876
rect 16523 7824 16548 7876
rect 15843 7798 16548 7824
rect 10909 7360 10986 7396
rect 10909 7304 10919 7360
rect 10975 7304 10986 7360
rect 10909 7280 10986 7304
rect 10909 7224 10919 7280
rect 10975 7224 10986 7280
rect 8973 7191 9030 7202
rect 10909 7200 10986 7224
rect 9029 7135 9030 7191
rect 8973 7124 9030 7135
rect 9555 7184 9633 7191
rect 9555 7128 9566 7184
rect 9622 7128 9633 7184
rect 9555 7121 9633 7128
rect 10909 7144 10919 7200
rect 10975 7144 10986 7200
rect 10909 7120 10986 7144
rect 10909 7064 10919 7120
rect 10975 7064 10986 7120
rect 10909 7040 10986 7064
rect 10909 6984 10919 7040
rect 10975 6984 10986 7040
rect 10909 6960 10986 6984
rect 10909 6904 10919 6960
rect 10975 6904 10986 6960
rect 10909 6880 10986 6904
rect 10909 6824 10919 6880
rect 10975 6824 10986 6880
rect 10909 6800 10986 6824
rect 10909 6744 10919 6800
rect 10975 6744 10986 6800
rect 10909 6720 10986 6744
rect 10909 6664 10919 6720
rect 10975 6664 10986 6720
rect 10909 6640 10986 6664
rect 10909 6584 10919 6640
rect 10975 6584 10986 6640
rect 10909 6560 10986 6584
rect 10909 6504 10919 6560
rect 10975 6504 10986 6560
rect 10909 6480 10986 6504
rect 10909 6424 10919 6480
rect 10975 6424 10986 6480
rect 10909 6400 10986 6424
rect 10909 6344 10919 6400
rect 10975 6344 10986 6400
rect 10909 6320 10986 6344
rect 10909 6264 10919 6320
rect 10975 6264 10986 6320
rect 10909 6240 10986 6264
rect 10909 6184 10919 6240
rect 10975 6184 10986 6240
rect 10909 6160 10986 6184
rect 10909 6104 10919 6160
rect 10975 6104 10986 6160
rect 10909 6080 10986 6104
rect 10909 6024 10919 6080
rect 10975 6024 10986 6080
rect 10909 6000 10986 6024
rect 10909 5944 10919 6000
rect 10975 5944 10986 6000
rect 10909 5920 10986 5944
rect 10909 5864 10919 5920
rect 10975 5864 10986 5920
rect 10909 5829 10986 5864
rect 11049 6469 11140 6491
rect 11049 6413 11065 6469
rect 11121 6413 11140 6469
rect 11049 6389 11140 6413
rect 11049 6333 11065 6389
rect 11121 6333 11140 6389
rect 11049 6309 11140 6333
rect 11049 6253 11065 6309
rect 11121 6253 11140 6309
rect 11049 6229 11140 6253
rect 11049 6173 11065 6229
rect 11121 6173 11140 6229
rect 11049 6149 11140 6173
rect 11049 6093 11065 6149
rect 11121 6093 11140 6149
rect 11049 6069 11140 6093
rect 11049 6013 11065 6069
rect 11121 6013 11140 6069
rect 11049 5989 11140 6013
rect 11049 5933 11065 5989
rect 11121 5933 11140 5989
rect 11049 5909 11140 5933
rect 11049 5853 11065 5909
rect 11121 5853 11140 5909
rect 11049 5837 11140 5853
rect 10943 5760 11058 5768
rect 10943 5704 10972 5760
rect 11028 5704 11058 5760
rect 10943 5697 11058 5704
rect 12507 5761 12591 5770
rect 12507 5705 12520 5761
rect 12576 5758 12591 5761
rect 12581 5706 12591 5758
rect 13169 5719 13199 5775
rect 13255 5719 13279 5775
rect 13335 5719 13359 5775
rect 13415 5719 13439 5775
rect 13495 5719 13519 5775
rect 13575 5719 13599 5775
rect 13655 5719 13679 5775
rect 13735 5719 13759 5775
rect 13815 5719 13839 5775
rect 13895 5719 13919 5775
rect 13975 5719 13999 5775
rect 14055 5719 14079 5775
rect 14135 5719 14159 5775
rect 14215 5719 14239 5775
rect 14295 5719 14319 5775
rect 14375 5719 14399 5775
rect 14455 5719 14479 5775
rect 14535 5719 14559 5775
rect 14615 5719 14639 5775
rect 14695 5719 14726 5775
rect 14797 5722 14882 5738
rect 12576 5705 12591 5706
rect 12507 5697 12591 5705
rect 14797 5670 14803 5722
rect 14855 5720 14882 5722
rect 14797 5664 14807 5670
rect 14863 5664 14882 5720
rect 14797 5656 14882 5664
rect 13159 5548 14759 5618
rect 12415 5532 12512 5545
rect 12415 5480 12436 5532
rect 12488 5480 12512 5532
rect 12415 5366 12512 5480
rect 13159 5492 13211 5548
rect 13267 5492 13291 5548
rect 13347 5492 13371 5548
rect 13427 5492 13451 5548
rect 13507 5492 13531 5548
rect 13587 5492 13611 5548
rect 13667 5492 13691 5548
rect 13747 5492 13771 5548
rect 13827 5492 13851 5548
rect 13907 5492 13931 5548
rect 13987 5492 14011 5548
rect 14067 5492 14091 5548
rect 14147 5492 14171 5548
rect 14227 5492 14251 5548
rect 14307 5492 14331 5548
rect 14387 5492 14411 5548
rect 14467 5492 14491 5548
rect 14547 5492 14571 5548
rect 14627 5492 14651 5548
rect 14707 5492 14759 5548
rect 13159 5467 14759 5492
rect 10428 5330 12512 5366
rect 10428 5278 10478 5330
rect 10530 5278 12512 5330
rect 10428 5246 12512 5278
rect 15843 5147 16000 7798
rect 16612 7719 16686 7752
rect 16612 7663 16622 7719
rect 16678 7663 16686 7719
rect 16612 7639 16686 7663
rect 16612 7583 16622 7639
rect 16678 7583 16686 7639
rect 16612 7550 16686 7583
rect 16722 7720 16825 7754
rect 16722 7664 16757 7720
rect 16813 7664 16825 7720
rect 16722 7640 16825 7664
rect 16722 7584 16757 7640
rect 16813 7584 16825 7640
rect 16722 7551 16825 7584
rect 19626 7577 19702 8839
rect 20137 8458 20214 8466
rect 20137 8402 20147 8458
rect 20203 8402 20214 8458
rect 20137 8395 20214 8402
rect 20028 7771 20146 7800
rect 20028 7715 20060 7771
rect 20116 7715 20146 7771
rect 20028 7691 20146 7715
rect 20028 7635 20060 7691
rect 20116 7635 20146 7691
rect 20196 7668 20228 7698
rect 20028 7606 20146 7635
rect 19626 7559 20222 7577
rect 16636 7502 16766 7520
rect 16636 7450 16673 7502
rect 16725 7450 16766 7502
rect 16636 7418 16766 7450
rect 16636 7362 16672 7418
rect 16728 7362 16766 7418
rect 16636 7343 16766 7362
rect 19626 7507 20150 7559
rect 20202 7507 20222 7559
rect 19626 7467 20222 7507
rect 19626 6331 19702 7467
rect 20152 7219 20231 7231
rect 20152 7163 20163 7219
rect 20219 7163 20231 7219
rect 20152 7161 20165 7163
rect 20217 7161 20231 7163
rect 20152 7154 20231 7161
rect 20056 6535 20162 6566
rect 20056 6479 20082 6535
rect 20138 6479 20162 6535
rect 20056 6455 20162 6479
rect 20218 6472 20234 6490
rect 20056 6399 20082 6455
rect 20138 6399 20162 6455
rect 20056 6369 20162 6399
rect 19626 6315 20231 6331
rect 19626 6263 20163 6315
rect 20215 6263 20231 6315
rect 19626 6244 20231 6263
rect 27240 5386 27403 5405
rect 22419 5319 22547 5350
rect 22419 5263 22454 5319
rect 22510 5263 22547 5319
rect 22419 5233 22547 5263
rect 23408 5315 23517 5337
rect 23408 5259 23435 5315
rect 23491 5259 23517 5315
rect 23408 5235 23517 5259
rect 27240 5250 27252 5386
rect 27388 5250 27403 5386
rect 27240 5229 27403 5250
rect 15841 5100 16000 5147
rect 15841 5048 15862 5100
rect 15914 5048 15926 5100
rect 15978 5048 16000 5100
rect 15841 5023 16000 5048
rect 15841 4998 15999 5023
rect 4417 -543 5171 -474
rect 4417 -557 4514 -543
rect 5078 -557 5171 -543
rect 4417 -1093 4488 -557
rect 5104 -1093 5171 -557
rect 4417 -1107 4514 -1093
rect 5078 -1107 5171 -1093
rect 4417 -1169 5171 -1107
<< via2 >>
rect 11007 11024 11063 11028
rect 11007 10972 11009 11024
rect 11009 10972 11061 11024
rect 11061 10972 11063 11024
rect 11034 10303 11090 10359
rect 11034 10223 11090 10279
rect 11034 10143 11090 10199
rect 11034 10063 11090 10119
rect 11034 9983 11090 10039
rect 11034 9903 11090 9959
rect 11034 9823 11090 9879
rect 11034 9743 11090 9799
rect 11034 9663 11090 9719
rect 11034 9583 11090 9639
rect 11034 9503 11090 9559
rect 11034 9423 11090 9479
rect 11034 9343 11090 9399
rect 11034 9263 11090 9319
rect 11034 9183 11090 9239
rect 16230 11557 16286 11613
rect 16826 11535 16882 11591
rect 18991 10497 19047 10553
rect 16687 9797 16743 9799
rect 16687 9745 16689 9797
rect 16689 9745 16741 9797
rect 16741 9745 16743 9797
rect 16687 9743 16743 9745
rect 17769 9743 17825 9799
rect 17634 9298 17690 9300
rect 17634 9246 17636 9298
rect 17636 9246 17688 9298
rect 17688 9246 17690 9298
rect 17634 9244 17690 9246
rect 20152 9798 20208 9800
rect 20152 9746 20154 9798
rect 20154 9746 20206 9798
rect 20206 9746 20208 9798
rect 20152 9744 20208 9746
rect 11034 9103 11090 9159
rect 11034 9023 11090 9079
rect 11034 8943 11090 8999
rect 11034 8863 11090 8919
rect 10990 8697 11035 8747
rect 11035 8697 11046 8747
rect 10990 8691 11046 8697
rect 16626 9057 16682 9113
rect 16626 8977 16682 9033
rect 16759 9059 16815 9115
rect 16759 8979 16815 9035
rect 17644 8966 17700 9022
rect 20091 9040 20147 9096
rect 20245 9072 20301 9128
rect 20245 8992 20301 9048
rect 16673 8759 16729 8815
rect 18006 8791 18062 8847
rect 18798 8781 18854 8837
rect 19160 8771 19216 8827
rect 17588 8645 17590 8691
rect 17590 8645 17642 8691
rect 17642 8645 17644 8691
rect 17588 8635 17644 8645
rect 17588 8581 17590 8611
rect 17590 8581 17642 8611
rect 17642 8581 17644 8611
rect 17588 8569 17644 8581
rect 17588 8555 17590 8569
rect 17590 8555 17642 8569
rect 17642 8555 17644 8569
rect 17588 8517 17590 8531
rect 17590 8517 17642 8531
rect 17642 8517 17644 8531
rect 17588 8505 17644 8517
rect 17588 8475 17590 8505
rect 17590 8475 17642 8505
rect 17642 8475 17644 8505
rect 16660 8408 16716 8410
rect 16660 8356 16664 8408
rect 16664 8356 16716 8408
rect 16660 8354 16716 8356
rect 17588 8441 17644 8451
rect 17588 8395 17590 8441
rect 17590 8395 17642 8441
rect 17642 8395 17644 8441
rect 10991 8025 11047 8037
rect 10991 7981 10993 8025
rect 10993 7981 11045 8025
rect 11045 7981 11047 8025
rect 10919 7304 10975 7360
rect 10919 7224 10975 7280
rect 8973 7135 9029 7191
rect 9566 7128 9622 7184
rect 10919 7144 10975 7200
rect 10919 7064 10975 7120
rect 10919 6984 10975 7040
rect 10919 6904 10975 6960
rect 10919 6824 10975 6880
rect 10919 6744 10975 6800
rect 10919 6664 10975 6720
rect 10919 6584 10975 6640
rect 10919 6504 10975 6560
rect 10919 6424 10975 6480
rect 10919 6344 10975 6400
rect 10919 6264 10975 6320
rect 10919 6184 10975 6240
rect 10919 6104 10975 6160
rect 10919 6024 10975 6080
rect 10919 5944 10975 6000
rect 10919 5864 10975 5920
rect 11065 6413 11121 6469
rect 11065 6333 11121 6389
rect 11065 6253 11121 6309
rect 11065 6173 11121 6229
rect 11065 6093 11121 6149
rect 11065 6013 11121 6069
rect 11065 5933 11121 5989
rect 11065 5853 11121 5909
rect 10972 5758 11028 5760
rect 10972 5706 10975 5758
rect 10975 5706 11027 5758
rect 11027 5706 11028 5758
rect 10972 5704 11028 5706
rect 12520 5758 12576 5761
rect 12520 5706 12529 5758
rect 12529 5706 12576 5758
rect 13199 5719 13255 5775
rect 13279 5719 13335 5775
rect 13359 5719 13415 5775
rect 13439 5719 13495 5775
rect 13519 5719 13575 5775
rect 13599 5719 13655 5775
rect 13679 5719 13735 5775
rect 13759 5719 13815 5775
rect 13839 5719 13895 5775
rect 13919 5719 13975 5775
rect 13999 5719 14055 5775
rect 14079 5719 14135 5775
rect 14159 5719 14215 5775
rect 14239 5719 14295 5775
rect 14319 5719 14375 5775
rect 14399 5719 14455 5775
rect 14479 5719 14535 5775
rect 14559 5719 14615 5775
rect 14639 5719 14695 5775
rect 12520 5705 12576 5706
rect 14807 5670 14855 5720
rect 14855 5670 14863 5720
rect 14807 5664 14863 5670
rect 13211 5492 13267 5548
rect 13291 5492 13347 5548
rect 13371 5492 13427 5548
rect 13451 5492 13507 5548
rect 13531 5492 13587 5548
rect 13611 5492 13667 5548
rect 13691 5492 13747 5548
rect 13771 5492 13827 5548
rect 13851 5492 13907 5548
rect 13931 5492 13987 5548
rect 14011 5492 14067 5548
rect 14091 5492 14147 5548
rect 14171 5492 14227 5548
rect 14251 5492 14307 5548
rect 14331 5492 14387 5548
rect 14411 5492 14467 5548
rect 14491 5492 14547 5548
rect 14571 5492 14627 5548
rect 14651 5492 14707 5548
rect 16622 7663 16678 7719
rect 16622 7583 16678 7639
rect 16757 7664 16813 7720
rect 16757 7584 16813 7640
rect 20147 8454 20203 8458
rect 20147 8402 20149 8454
rect 20149 8402 20201 8454
rect 20201 8402 20203 8454
rect 20060 7715 20116 7771
rect 20060 7635 20116 7691
rect 16672 7362 16728 7418
rect 20163 7213 20219 7219
rect 20163 7163 20165 7213
rect 20165 7163 20217 7213
rect 20217 7163 20219 7213
rect 20082 6479 20138 6535
rect 20082 6399 20138 6455
rect 22454 5317 22510 5319
rect 22454 5265 22456 5317
rect 22456 5265 22508 5317
rect 22508 5265 22510 5317
rect 22454 5263 22510 5265
rect 23435 5313 23491 5315
rect 23435 5261 23437 5313
rect 23437 5261 23489 5313
rect 23489 5261 23491 5313
rect 23435 5259 23491 5261
rect 27252 5376 27388 5386
rect 27252 5260 27262 5376
rect 27262 5260 27378 5376
rect 27378 5260 27388 5376
rect 27252 5250 27388 5260
rect 4488 -1093 4514 -557
rect 4514 -1093 5078 -557
rect 5078 -1093 5104 -557
<< metal3 >>
rect 16192 11613 16327 11643
rect 16192 11557 16230 11613
rect 16286 11557 16327 11613
rect 10738 11028 11086 11034
rect 10738 10972 11007 11028
rect 11063 10972 11086 11028
rect 10738 10957 11086 10972
rect 10738 10862 10843 10957
rect 8944 7198 9069 7215
rect 10737 7208 10843 10862
rect 16192 10662 16327 11557
rect 16801 11595 16904 11637
rect 16801 11531 16822 11595
rect 16886 11531 16904 11595
rect 16801 11487 16904 11531
rect 16191 10553 16327 10662
rect 18943 10557 19098 10594
rect 11028 10362 11099 10388
rect 11028 10298 11033 10362
rect 11097 10298 11099 10362
rect 16191 10345 16326 10553
rect 18943 10493 18987 10557
rect 19051 10493 19098 10557
rect 18943 10460 19098 10493
rect 11028 10282 11099 10298
rect 11028 10218 11033 10282
rect 11097 10218 11099 10282
rect 11028 10202 11099 10218
rect 11028 10138 11033 10202
rect 11097 10138 11099 10202
rect 11028 10122 11099 10138
rect 11028 10058 11033 10122
rect 11097 10058 11099 10122
rect 11028 10042 11099 10058
rect 11028 9978 11033 10042
rect 11097 9978 11099 10042
rect 11028 9962 11099 9978
rect 11028 9898 11033 9962
rect 11097 9898 11099 9962
rect 11028 9882 11099 9898
rect 11028 9818 11033 9882
rect 11097 9818 11099 9882
rect 11028 9802 11099 9818
rect 11028 9738 11033 9802
rect 11097 9738 11099 9802
rect 11028 9722 11099 9738
rect 11028 9658 11033 9722
rect 11097 9658 11099 9722
rect 11028 9642 11099 9658
rect 11028 9578 11033 9642
rect 11097 9578 11099 9642
rect 11028 9562 11099 9578
rect 11028 9498 11033 9562
rect 11097 9498 11099 9562
rect 11028 9482 11099 9498
rect 11028 9418 11033 9482
rect 11097 9418 11099 9482
rect 11028 9402 11099 9418
rect 11028 9338 11033 9402
rect 11097 9338 11099 9402
rect 11028 9322 11099 9338
rect 11028 9258 11033 9322
rect 11097 9258 11099 9322
rect 11028 9242 11099 9258
rect 11028 9178 11033 9242
rect 11097 9178 11099 9242
rect 11028 9162 11099 9178
rect 11028 9098 11033 9162
rect 11097 9098 11099 9162
rect 11028 9082 11099 9098
rect 11028 9018 11033 9082
rect 11097 9018 11099 9082
rect 16190 10145 16326 10345
rect 16190 9813 16325 10145
rect 16190 9800 20529 9813
rect 16190 9799 20152 9800
rect 16190 9743 16687 9799
rect 16743 9743 17769 9799
rect 17825 9744 20152 9799
rect 20208 9744 20529 9800
rect 17825 9743 20529 9744
rect 16190 9732 20529 9743
rect 16190 9051 16325 9732
rect 17594 9410 20326 9498
rect 17594 9300 17731 9410
rect 17594 9244 17634 9300
rect 17690 9244 17731 9300
rect 17594 9232 17731 9244
rect 11028 9002 11099 9018
rect 11028 8938 11033 9002
rect 11097 8938 11099 9002
rect 11028 8922 11099 8938
rect 11028 8858 11033 8922
rect 11097 8858 11099 8922
rect 11028 8835 11099 8858
rect 10967 8747 11073 8769
rect 10967 8691 10990 8747
rect 11046 8691 11073 8747
rect 10967 8387 11073 8691
rect 16189 8579 16325 9051
rect 16609 9119 16692 9147
rect 16609 9055 16618 9119
rect 16682 9055 16692 9119
rect 16609 9039 16692 9055
rect 16609 8975 16618 9039
rect 16682 8975 16692 9039
rect 16609 8946 16692 8975
rect 16752 9115 16850 9150
rect 16752 9059 16759 9115
rect 16815 9059 16850 9115
rect 16752 9048 16850 9059
rect 18596 9096 20158 9140
rect 16752 9035 17725 9048
rect 16752 8979 16759 9035
rect 16815 9022 17725 9035
rect 16815 8979 17644 9022
rect 16752 8966 17644 8979
rect 17700 8966 17725 9022
rect 16752 8946 17725 8966
rect 18596 9040 20091 9096
rect 20147 9040 20158 9096
rect 18596 8997 20158 9040
rect 20224 9132 20326 9410
rect 20224 9068 20241 9132
rect 20305 9068 20326 9132
rect 20224 9052 20326 9068
rect 20224 9027 20241 9052
rect 17974 8851 18099 8876
rect 16648 8819 16758 8842
rect 16648 8755 16669 8819
rect 16733 8755 16758 8819
rect 17974 8787 18002 8851
rect 18066 8787 18099 8851
rect 17974 8763 18099 8787
rect 16648 8734 16758 8755
rect 17538 8718 17686 8720
rect 17538 8695 17689 8718
rect 18596 8714 18703 8997
rect 20225 8988 20241 9027
rect 20305 8988 20326 9052
rect 20225 8962 20326 8988
rect 18770 8841 18887 8864
rect 18770 8777 18794 8841
rect 18858 8777 18887 8841
rect 18770 8758 18887 8777
rect 19136 8827 19277 8846
rect 19136 8771 19160 8827
rect 19216 8771 19277 8827
rect 19136 8753 19277 8771
rect 17538 8631 17584 8695
rect 17648 8631 17689 8695
rect 17538 8615 17689 8631
rect 16189 8425 16324 8579
rect 17538 8551 17584 8615
rect 17648 8551 17689 8615
rect 17538 8535 17689 8551
rect 17538 8471 17584 8535
rect 17648 8471 17689 8535
rect 17538 8455 17689 8471
rect 16189 8410 16737 8425
rect 10967 8354 11349 8387
rect 10967 8290 10986 8354
rect 11050 8290 11349 8354
rect 16189 8354 16660 8410
rect 16716 8354 16737 8410
rect 17538 8391 17584 8455
rect 17648 8391 17689 8455
rect 18594 8397 18703 8714
rect 17538 8365 17689 8391
rect 17538 8359 17686 8365
rect 16189 8339 16737 8354
rect 10967 8261 11349 8290
rect 10967 8037 11073 8261
rect 10967 7981 10991 8037
rect 11047 7981 11073 8037
rect 10967 7957 11073 7981
rect 10909 7364 10986 7396
rect 10909 7300 10915 7364
rect 10979 7300 10986 7364
rect 10909 7284 10986 7300
rect 10909 7220 10915 7284
rect 10979 7220 10986 7284
rect 8944 7191 8976 7198
rect 8944 7135 8973 7191
rect 8944 7134 8976 7135
rect 9040 7134 9069 7198
rect 8944 7114 9069 7134
rect 9547 7184 10842 7208
rect 9547 7128 9566 7184
rect 9622 7128 10842 7184
rect 9547 7108 10842 7128
rect 10736 5769 10842 7108
rect 10909 7204 10986 7220
rect 10909 7140 10915 7204
rect 10979 7140 10986 7204
rect 10909 7124 10986 7140
rect 10909 7060 10915 7124
rect 10979 7060 10986 7124
rect 10909 7044 10986 7060
rect 10909 6980 10915 7044
rect 10979 6980 10986 7044
rect 10909 6964 10986 6980
rect 10909 6900 10915 6964
rect 10979 6900 10986 6964
rect 10909 6884 10986 6900
rect 10909 6820 10915 6884
rect 10979 6820 10986 6884
rect 10909 6804 10986 6820
rect 10909 6740 10915 6804
rect 10979 6740 10986 6804
rect 10909 6724 10986 6740
rect 10909 6660 10915 6724
rect 10979 6660 10986 6724
rect 10909 6644 10986 6660
rect 10909 6580 10915 6644
rect 10979 6580 10986 6644
rect 10909 6564 10986 6580
rect 10909 6500 10915 6564
rect 10979 6500 10986 6564
rect 10909 6484 10986 6500
rect 10909 6420 10915 6484
rect 10979 6420 10986 6484
rect 10909 6404 10986 6420
rect 10909 6340 10915 6404
rect 10979 6340 10986 6404
rect 10909 6324 10986 6340
rect 10909 6260 10915 6324
rect 10979 6260 10986 6324
rect 10909 6244 10986 6260
rect 10909 6180 10915 6244
rect 10979 6180 10986 6244
rect 10909 6164 10986 6180
rect 10909 6100 10915 6164
rect 10979 6100 10986 6164
rect 10909 6084 10986 6100
rect 10909 6020 10915 6084
rect 10979 6020 10986 6084
rect 10909 6004 10986 6020
rect 10909 5940 10915 6004
rect 10979 5940 10986 6004
rect 10909 5924 10986 5940
rect 10909 5860 10915 5924
rect 10979 5860 10986 5924
rect 10909 5829 10986 5860
rect 11049 6469 11140 6491
rect 11049 6434 11065 6469
rect 11121 6434 11140 6469
rect 11049 6370 11064 6434
rect 11128 6370 11140 6434
rect 11049 6354 11065 6370
rect 11121 6354 11140 6370
rect 11049 6290 11064 6354
rect 11128 6290 11140 6354
rect 11049 6274 11065 6290
rect 11121 6274 11140 6290
rect 11049 6210 11064 6274
rect 11128 6210 11140 6274
rect 11049 6194 11065 6210
rect 11121 6194 11140 6210
rect 11049 6130 11064 6194
rect 11128 6130 11140 6194
rect 11049 6114 11065 6130
rect 11121 6114 11140 6130
rect 11049 6050 11064 6114
rect 11128 6050 11140 6114
rect 11049 6034 11065 6050
rect 11121 6034 11140 6050
rect 11049 5970 11064 6034
rect 11128 5970 11140 6034
rect 11049 5954 11065 5970
rect 11121 5954 11140 5970
rect 11049 5890 11064 5954
rect 11128 5890 11140 5954
rect 11049 5853 11065 5890
rect 11121 5853 11140 5890
rect 11248 5980 11349 8261
rect 19165 7757 19277 8753
rect 20137 8462 20214 8466
rect 20460 8462 20529 9732
rect 20137 8458 20529 8462
rect 20137 8402 20147 8458
rect 20203 8402 20529 8458
rect 20137 8392 20529 8402
rect 20460 8168 20529 8392
rect 20459 7930 20529 8168
rect 18528 7756 19277 7757
rect 17963 7755 19277 7756
rect 17401 7754 19277 7755
rect 16599 7722 16686 7753
rect 16599 7658 16612 7722
rect 16676 7719 16686 7722
rect 16678 7663 16686 7719
rect 16676 7658 16686 7663
rect 16599 7642 16686 7658
rect 16599 7578 16612 7642
rect 16676 7639 16686 7642
rect 16678 7583 16686 7639
rect 16676 7578 16686 7583
rect 16599 7550 16686 7578
rect 16748 7720 19277 7754
rect 16748 7664 16757 7720
rect 16813 7664 19277 7720
rect 16748 7640 19277 7664
rect 16748 7584 16757 7640
rect 16813 7584 19277 7640
rect 20028 7775 20146 7800
rect 20028 7711 20056 7775
rect 20120 7711 20146 7775
rect 20028 7695 20146 7711
rect 20028 7631 20056 7695
rect 20120 7631 20146 7695
rect 20028 7606 20146 7631
rect 16748 7554 19277 7584
rect 16748 7553 18556 7554
rect 19081 7553 19244 7554
rect 16748 7552 17994 7553
rect 16748 7551 17417 7552
rect 16636 7422 16766 7435
rect 16636 7358 16668 7422
rect 16732 7358 16766 7422
rect 16636 7343 16766 7358
rect 20459 7227 20528 7930
rect 20152 7219 20528 7227
rect 20152 7163 20163 7219
rect 20219 7163 20528 7219
rect 20152 7152 20528 7163
rect 20056 6539 20162 6566
rect 20056 6475 20078 6539
rect 20142 6475 20162 6539
rect 20056 6459 20162 6475
rect 20056 6395 20078 6459
rect 20142 6395 20162 6459
rect 20056 6369 20162 6395
rect 11248 5867 14882 5980
rect 11049 5837 11140 5853
rect 13158 5786 14735 5799
rect 10736 5761 12599 5769
rect 10736 5760 12520 5761
rect 10736 5704 10972 5760
rect 11028 5705 12520 5760
rect 12576 5705 12599 5761
rect 13158 5722 13196 5786
rect 13260 5722 13276 5786
rect 13340 5722 13356 5786
rect 13420 5722 13436 5786
rect 13500 5722 13516 5786
rect 13580 5722 13596 5786
rect 13660 5722 13676 5786
rect 13740 5722 13756 5786
rect 13820 5722 13836 5786
rect 13900 5722 13916 5786
rect 13980 5722 13996 5786
rect 14060 5722 14076 5786
rect 14140 5722 14156 5786
rect 14220 5722 14236 5786
rect 14300 5722 14316 5786
rect 14380 5722 14396 5786
rect 14460 5722 14476 5786
rect 14540 5722 14556 5786
rect 14620 5722 14636 5786
rect 14700 5776 14735 5786
rect 14700 5722 14736 5776
rect 13158 5719 13199 5722
rect 13255 5719 13279 5722
rect 13335 5719 13359 5722
rect 13415 5719 13439 5722
rect 13495 5719 13519 5722
rect 13575 5719 13599 5722
rect 13655 5719 13679 5722
rect 13735 5719 13759 5722
rect 13815 5719 13839 5722
rect 13895 5719 13919 5722
rect 13975 5719 13999 5722
rect 14055 5719 14079 5722
rect 14135 5719 14159 5722
rect 14215 5719 14239 5722
rect 14295 5719 14319 5722
rect 14375 5719 14399 5722
rect 14455 5719 14479 5722
rect 14535 5719 14559 5722
rect 14615 5719 14639 5722
rect 14695 5719 14736 5722
rect 13158 5710 14736 5719
rect 14797 5720 14882 5867
rect 13158 5709 14735 5710
rect 11028 5704 12599 5705
rect 10736 5697 12599 5704
rect 14797 5664 14807 5720
rect 14863 5664 14882 5720
rect 14797 5656 14882 5664
rect 13159 5552 14759 5578
rect 13159 5488 13207 5552
rect 13271 5488 13287 5552
rect 13351 5488 13367 5552
rect 13431 5488 13447 5552
rect 13511 5488 13527 5552
rect 13591 5488 13607 5552
rect 13671 5488 13687 5552
rect 13751 5488 13767 5552
rect 13831 5488 13847 5552
rect 13911 5488 13927 5552
rect 13991 5488 14007 5552
rect 14071 5488 14087 5552
rect 14151 5488 14167 5552
rect 14231 5488 14247 5552
rect 14311 5488 14327 5552
rect 14391 5488 14407 5552
rect 14471 5488 14487 5552
rect 14551 5488 14567 5552
rect 14631 5488 14647 5552
rect 14711 5488 14759 5552
rect 13159 5467 14759 5488
rect 27240 5390 27403 5405
rect 27240 5386 27288 5390
rect 27352 5386 27403 5390
rect 22419 5323 22547 5350
rect 22419 5259 22450 5323
rect 22514 5259 22547 5323
rect 22419 5233 22547 5259
rect 23402 5318 23525 5343
rect 23402 5254 23431 5318
rect 23495 5254 23525 5318
rect 23402 5230 23525 5254
rect 27240 5250 27252 5386
rect 27388 5250 27403 5386
rect 27240 5246 27288 5250
rect 27352 5246 27403 5250
rect 27240 5229 27403 5246
rect 4417 -476 5171 -474
rect 4417 -557 6104 -476
rect 4417 -1093 4488 -557
rect 5104 -1093 6104 -557
rect 4417 -1169 6104 -1093
rect 5136 -1170 6104 -1169
<< via3 >>
rect 16822 11591 16886 11595
rect 16822 11535 16826 11591
rect 16826 11535 16882 11591
rect 16882 11535 16886 11591
rect 16822 11531 16886 11535
rect 11033 10359 11097 10362
rect 11033 10303 11034 10359
rect 11034 10303 11090 10359
rect 11090 10303 11097 10359
rect 11033 10298 11097 10303
rect 18987 10553 19051 10557
rect 18987 10497 18991 10553
rect 18991 10497 19047 10553
rect 19047 10497 19051 10553
rect 18987 10493 19051 10497
rect 11033 10279 11097 10282
rect 11033 10223 11034 10279
rect 11034 10223 11090 10279
rect 11090 10223 11097 10279
rect 11033 10218 11097 10223
rect 11033 10199 11097 10202
rect 11033 10143 11034 10199
rect 11034 10143 11090 10199
rect 11090 10143 11097 10199
rect 11033 10138 11097 10143
rect 11033 10119 11097 10122
rect 11033 10063 11034 10119
rect 11034 10063 11090 10119
rect 11090 10063 11097 10119
rect 11033 10058 11097 10063
rect 11033 10039 11097 10042
rect 11033 9983 11034 10039
rect 11034 9983 11090 10039
rect 11090 9983 11097 10039
rect 11033 9978 11097 9983
rect 11033 9959 11097 9962
rect 11033 9903 11034 9959
rect 11034 9903 11090 9959
rect 11090 9903 11097 9959
rect 11033 9898 11097 9903
rect 11033 9879 11097 9882
rect 11033 9823 11034 9879
rect 11034 9823 11090 9879
rect 11090 9823 11097 9879
rect 11033 9818 11097 9823
rect 11033 9799 11097 9802
rect 11033 9743 11034 9799
rect 11034 9743 11090 9799
rect 11090 9743 11097 9799
rect 11033 9738 11097 9743
rect 11033 9719 11097 9722
rect 11033 9663 11034 9719
rect 11034 9663 11090 9719
rect 11090 9663 11097 9719
rect 11033 9658 11097 9663
rect 11033 9639 11097 9642
rect 11033 9583 11034 9639
rect 11034 9583 11090 9639
rect 11090 9583 11097 9639
rect 11033 9578 11097 9583
rect 11033 9559 11097 9562
rect 11033 9503 11034 9559
rect 11034 9503 11090 9559
rect 11090 9503 11097 9559
rect 11033 9498 11097 9503
rect 11033 9479 11097 9482
rect 11033 9423 11034 9479
rect 11034 9423 11090 9479
rect 11090 9423 11097 9479
rect 11033 9418 11097 9423
rect 11033 9399 11097 9402
rect 11033 9343 11034 9399
rect 11034 9343 11090 9399
rect 11090 9343 11097 9399
rect 11033 9338 11097 9343
rect 11033 9319 11097 9322
rect 11033 9263 11034 9319
rect 11034 9263 11090 9319
rect 11090 9263 11097 9319
rect 11033 9258 11097 9263
rect 11033 9239 11097 9242
rect 11033 9183 11034 9239
rect 11034 9183 11090 9239
rect 11090 9183 11097 9239
rect 11033 9178 11097 9183
rect 11033 9159 11097 9162
rect 11033 9103 11034 9159
rect 11034 9103 11090 9159
rect 11090 9103 11097 9159
rect 11033 9098 11097 9103
rect 11033 9079 11097 9082
rect 11033 9023 11034 9079
rect 11034 9023 11090 9079
rect 11090 9023 11097 9079
rect 11033 9018 11097 9023
rect 11033 8999 11097 9002
rect 11033 8943 11034 8999
rect 11034 8943 11090 8999
rect 11090 8943 11097 8999
rect 11033 8938 11097 8943
rect 11033 8919 11097 8922
rect 11033 8863 11034 8919
rect 11034 8863 11090 8919
rect 11090 8863 11097 8919
rect 11033 8858 11097 8863
rect 16618 9113 16682 9119
rect 16618 9057 16626 9113
rect 16626 9057 16682 9113
rect 16618 9055 16682 9057
rect 16618 9033 16682 9039
rect 16618 8977 16626 9033
rect 16626 8977 16682 9033
rect 16618 8975 16682 8977
rect 20241 9128 20305 9132
rect 20241 9072 20245 9128
rect 20245 9072 20301 9128
rect 20301 9072 20305 9128
rect 20241 9068 20305 9072
rect 20241 9048 20305 9052
rect 16669 8815 16733 8819
rect 16669 8759 16673 8815
rect 16673 8759 16729 8815
rect 16729 8759 16733 8815
rect 16669 8755 16733 8759
rect 18002 8847 18066 8851
rect 18002 8791 18006 8847
rect 18006 8791 18062 8847
rect 18062 8791 18066 8847
rect 18002 8787 18066 8791
rect 20241 8992 20245 9048
rect 20245 8992 20301 9048
rect 20301 8992 20305 9048
rect 20241 8988 20305 8992
rect 18794 8837 18858 8841
rect 18794 8781 18798 8837
rect 18798 8781 18854 8837
rect 18854 8781 18858 8837
rect 18794 8777 18858 8781
rect 17584 8691 17648 8695
rect 17584 8635 17588 8691
rect 17588 8635 17644 8691
rect 17644 8635 17648 8691
rect 17584 8631 17648 8635
rect 17584 8611 17648 8615
rect 17584 8555 17588 8611
rect 17588 8555 17644 8611
rect 17644 8555 17648 8611
rect 17584 8551 17648 8555
rect 17584 8531 17648 8535
rect 17584 8475 17588 8531
rect 17588 8475 17644 8531
rect 17644 8475 17648 8531
rect 17584 8471 17648 8475
rect 10986 8290 11050 8354
rect 17584 8451 17648 8455
rect 17584 8395 17588 8451
rect 17588 8395 17644 8451
rect 17644 8395 17648 8451
rect 17584 8391 17648 8395
rect 10915 7360 10979 7364
rect 10915 7304 10919 7360
rect 10919 7304 10975 7360
rect 10975 7304 10979 7360
rect 10915 7300 10979 7304
rect 10915 7280 10979 7284
rect 10915 7224 10919 7280
rect 10919 7224 10975 7280
rect 10975 7224 10979 7280
rect 10915 7220 10979 7224
rect 8976 7191 9040 7198
rect 8976 7135 9029 7191
rect 9029 7135 9040 7191
rect 8976 7134 9040 7135
rect 10915 7200 10979 7204
rect 10915 7144 10919 7200
rect 10919 7144 10975 7200
rect 10975 7144 10979 7200
rect 10915 7140 10979 7144
rect 10915 7120 10979 7124
rect 10915 7064 10919 7120
rect 10919 7064 10975 7120
rect 10975 7064 10979 7120
rect 10915 7060 10979 7064
rect 10915 7040 10979 7044
rect 10915 6984 10919 7040
rect 10919 6984 10975 7040
rect 10975 6984 10979 7040
rect 10915 6980 10979 6984
rect 10915 6960 10979 6964
rect 10915 6904 10919 6960
rect 10919 6904 10975 6960
rect 10975 6904 10979 6960
rect 10915 6900 10979 6904
rect 10915 6880 10979 6884
rect 10915 6824 10919 6880
rect 10919 6824 10975 6880
rect 10975 6824 10979 6880
rect 10915 6820 10979 6824
rect 10915 6800 10979 6804
rect 10915 6744 10919 6800
rect 10919 6744 10975 6800
rect 10975 6744 10979 6800
rect 10915 6740 10979 6744
rect 10915 6720 10979 6724
rect 10915 6664 10919 6720
rect 10919 6664 10975 6720
rect 10975 6664 10979 6720
rect 10915 6660 10979 6664
rect 10915 6640 10979 6644
rect 10915 6584 10919 6640
rect 10919 6584 10975 6640
rect 10975 6584 10979 6640
rect 10915 6580 10979 6584
rect 10915 6560 10979 6564
rect 10915 6504 10919 6560
rect 10919 6504 10975 6560
rect 10975 6504 10979 6560
rect 10915 6500 10979 6504
rect 10915 6480 10979 6484
rect 10915 6424 10919 6480
rect 10919 6424 10975 6480
rect 10975 6424 10979 6480
rect 10915 6420 10979 6424
rect 10915 6400 10979 6404
rect 10915 6344 10919 6400
rect 10919 6344 10975 6400
rect 10975 6344 10979 6400
rect 10915 6340 10979 6344
rect 10915 6320 10979 6324
rect 10915 6264 10919 6320
rect 10919 6264 10975 6320
rect 10975 6264 10979 6320
rect 10915 6260 10979 6264
rect 10915 6240 10979 6244
rect 10915 6184 10919 6240
rect 10919 6184 10975 6240
rect 10975 6184 10979 6240
rect 10915 6180 10979 6184
rect 10915 6160 10979 6164
rect 10915 6104 10919 6160
rect 10919 6104 10975 6160
rect 10975 6104 10979 6160
rect 10915 6100 10979 6104
rect 10915 6080 10979 6084
rect 10915 6024 10919 6080
rect 10919 6024 10975 6080
rect 10975 6024 10979 6080
rect 10915 6020 10979 6024
rect 10915 6000 10979 6004
rect 10915 5944 10919 6000
rect 10919 5944 10975 6000
rect 10975 5944 10979 6000
rect 10915 5940 10979 5944
rect 10915 5920 10979 5924
rect 10915 5864 10919 5920
rect 10919 5864 10975 5920
rect 10975 5864 10979 5920
rect 10915 5860 10979 5864
rect 11064 6413 11065 6434
rect 11065 6413 11121 6434
rect 11121 6413 11128 6434
rect 11064 6389 11128 6413
rect 11064 6370 11065 6389
rect 11065 6370 11121 6389
rect 11121 6370 11128 6389
rect 11064 6333 11065 6354
rect 11065 6333 11121 6354
rect 11121 6333 11128 6354
rect 11064 6309 11128 6333
rect 11064 6290 11065 6309
rect 11065 6290 11121 6309
rect 11121 6290 11128 6309
rect 11064 6253 11065 6274
rect 11065 6253 11121 6274
rect 11121 6253 11128 6274
rect 11064 6229 11128 6253
rect 11064 6210 11065 6229
rect 11065 6210 11121 6229
rect 11121 6210 11128 6229
rect 11064 6173 11065 6194
rect 11065 6173 11121 6194
rect 11121 6173 11128 6194
rect 11064 6149 11128 6173
rect 11064 6130 11065 6149
rect 11065 6130 11121 6149
rect 11121 6130 11128 6149
rect 11064 6093 11065 6114
rect 11065 6093 11121 6114
rect 11121 6093 11128 6114
rect 11064 6069 11128 6093
rect 11064 6050 11065 6069
rect 11065 6050 11121 6069
rect 11121 6050 11128 6069
rect 11064 6013 11065 6034
rect 11065 6013 11121 6034
rect 11121 6013 11128 6034
rect 11064 5989 11128 6013
rect 11064 5970 11065 5989
rect 11065 5970 11121 5989
rect 11121 5970 11128 5989
rect 11064 5933 11065 5954
rect 11065 5933 11121 5954
rect 11121 5933 11128 5954
rect 11064 5909 11128 5933
rect 11064 5890 11065 5909
rect 11065 5890 11121 5909
rect 11121 5890 11128 5909
rect 16612 7719 16676 7722
rect 16612 7663 16622 7719
rect 16622 7663 16676 7719
rect 16612 7658 16676 7663
rect 16612 7639 16676 7642
rect 16612 7583 16622 7639
rect 16622 7583 16676 7639
rect 16612 7578 16676 7583
rect 20056 7771 20120 7775
rect 20056 7715 20060 7771
rect 20060 7715 20116 7771
rect 20116 7715 20120 7771
rect 20056 7711 20120 7715
rect 20056 7691 20120 7695
rect 20056 7635 20060 7691
rect 20060 7635 20116 7691
rect 20116 7635 20120 7691
rect 20056 7631 20120 7635
rect 16668 7418 16732 7422
rect 16668 7362 16672 7418
rect 16672 7362 16728 7418
rect 16728 7362 16732 7418
rect 16668 7358 16732 7362
rect 20078 6535 20142 6539
rect 20078 6479 20082 6535
rect 20082 6479 20138 6535
rect 20138 6479 20142 6535
rect 20078 6475 20142 6479
rect 20078 6455 20142 6459
rect 20078 6399 20082 6455
rect 20082 6399 20138 6455
rect 20138 6399 20142 6455
rect 20078 6395 20142 6399
rect 13196 5775 13260 5786
rect 13196 5722 13199 5775
rect 13199 5722 13255 5775
rect 13255 5722 13260 5775
rect 13276 5775 13340 5786
rect 13276 5722 13279 5775
rect 13279 5722 13335 5775
rect 13335 5722 13340 5775
rect 13356 5775 13420 5786
rect 13356 5722 13359 5775
rect 13359 5722 13415 5775
rect 13415 5722 13420 5775
rect 13436 5775 13500 5786
rect 13436 5722 13439 5775
rect 13439 5722 13495 5775
rect 13495 5722 13500 5775
rect 13516 5775 13580 5786
rect 13516 5722 13519 5775
rect 13519 5722 13575 5775
rect 13575 5722 13580 5775
rect 13596 5775 13660 5786
rect 13596 5722 13599 5775
rect 13599 5722 13655 5775
rect 13655 5722 13660 5775
rect 13676 5775 13740 5786
rect 13676 5722 13679 5775
rect 13679 5722 13735 5775
rect 13735 5722 13740 5775
rect 13756 5775 13820 5786
rect 13756 5722 13759 5775
rect 13759 5722 13815 5775
rect 13815 5722 13820 5775
rect 13836 5775 13900 5786
rect 13836 5722 13839 5775
rect 13839 5722 13895 5775
rect 13895 5722 13900 5775
rect 13916 5775 13980 5786
rect 13916 5722 13919 5775
rect 13919 5722 13975 5775
rect 13975 5722 13980 5775
rect 13996 5775 14060 5786
rect 13996 5722 13999 5775
rect 13999 5722 14055 5775
rect 14055 5722 14060 5775
rect 14076 5775 14140 5786
rect 14076 5722 14079 5775
rect 14079 5722 14135 5775
rect 14135 5722 14140 5775
rect 14156 5775 14220 5786
rect 14156 5722 14159 5775
rect 14159 5722 14215 5775
rect 14215 5722 14220 5775
rect 14236 5775 14300 5786
rect 14236 5722 14239 5775
rect 14239 5722 14295 5775
rect 14295 5722 14300 5775
rect 14316 5775 14380 5786
rect 14316 5722 14319 5775
rect 14319 5722 14375 5775
rect 14375 5722 14380 5775
rect 14396 5775 14460 5786
rect 14396 5722 14399 5775
rect 14399 5722 14455 5775
rect 14455 5722 14460 5775
rect 14476 5775 14540 5786
rect 14476 5722 14479 5775
rect 14479 5722 14535 5775
rect 14535 5722 14540 5775
rect 14556 5775 14620 5786
rect 14556 5722 14559 5775
rect 14559 5722 14615 5775
rect 14615 5722 14620 5775
rect 14636 5775 14700 5786
rect 14636 5722 14639 5775
rect 14639 5722 14695 5775
rect 14695 5722 14700 5775
rect 13207 5548 13271 5552
rect 13207 5492 13211 5548
rect 13211 5492 13267 5548
rect 13267 5492 13271 5548
rect 13207 5488 13271 5492
rect 13287 5548 13351 5552
rect 13287 5492 13291 5548
rect 13291 5492 13347 5548
rect 13347 5492 13351 5548
rect 13287 5488 13351 5492
rect 13367 5548 13431 5552
rect 13367 5492 13371 5548
rect 13371 5492 13427 5548
rect 13427 5492 13431 5548
rect 13367 5488 13431 5492
rect 13447 5548 13511 5552
rect 13447 5492 13451 5548
rect 13451 5492 13507 5548
rect 13507 5492 13511 5548
rect 13447 5488 13511 5492
rect 13527 5548 13591 5552
rect 13527 5492 13531 5548
rect 13531 5492 13587 5548
rect 13587 5492 13591 5548
rect 13527 5488 13591 5492
rect 13607 5548 13671 5552
rect 13607 5492 13611 5548
rect 13611 5492 13667 5548
rect 13667 5492 13671 5548
rect 13607 5488 13671 5492
rect 13687 5548 13751 5552
rect 13687 5492 13691 5548
rect 13691 5492 13747 5548
rect 13747 5492 13751 5548
rect 13687 5488 13751 5492
rect 13767 5548 13831 5552
rect 13767 5492 13771 5548
rect 13771 5492 13827 5548
rect 13827 5492 13831 5548
rect 13767 5488 13831 5492
rect 13847 5548 13911 5552
rect 13847 5492 13851 5548
rect 13851 5492 13907 5548
rect 13907 5492 13911 5548
rect 13847 5488 13911 5492
rect 13927 5548 13991 5552
rect 13927 5492 13931 5548
rect 13931 5492 13987 5548
rect 13987 5492 13991 5548
rect 13927 5488 13991 5492
rect 14007 5548 14071 5552
rect 14007 5492 14011 5548
rect 14011 5492 14067 5548
rect 14067 5492 14071 5548
rect 14007 5488 14071 5492
rect 14087 5548 14151 5552
rect 14087 5492 14091 5548
rect 14091 5492 14147 5548
rect 14147 5492 14151 5548
rect 14087 5488 14151 5492
rect 14167 5548 14231 5552
rect 14167 5492 14171 5548
rect 14171 5492 14227 5548
rect 14227 5492 14231 5548
rect 14167 5488 14231 5492
rect 14247 5548 14311 5552
rect 14247 5492 14251 5548
rect 14251 5492 14307 5548
rect 14307 5492 14311 5548
rect 14247 5488 14311 5492
rect 14327 5548 14391 5552
rect 14327 5492 14331 5548
rect 14331 5492 14387 5548
rect 14387 5492 14391 5548
rect 14327 5488 14391 5492
rect 14407 5548 14471 5552
rect 14407 5492 14411 5548
rect 14411 5492 14467 5548
rect 14467 5492 14471 5548
rect 14407 5488 14471 5492
rect 14487 5548 14551 5552
rect 14487 5492 14491 5548
rect 14491 5492 14547 5548
rect 14547 5492 14551 5548
rect 14487 5488 14551 5492
rect 14567 5548 14631 5552
rect 14567 5492 14571 5548
rect 14571 5492 14627 5548
rect 14627 5492 14631 5548
rect 14567 5488 14631 5492
rect 14647 5548 14711 5552
rect 14647 5492 14651 5548
rect 14651 5492 14707 5548
rect 14707 5492 14711 5548
rect 14647 5488 14711 5492
rect 27288 5386 27352 5390
rect 22450 5319 22514 5323
rect 22450 5263 22454 5319
rect 22454 5263 22510 5319
rect 22510 5263 22514 5319
rect 22450 5259 22514 5263
rect 23431 5315 23495 5318
rect 23431 5259 23435 5315
rect 23435 5259 23491 5315
rect 23491 5259 23495 5315
rect 23431 5254 23495 5259
rect 27288 5326 27352 5386
rect 27288 5250 27352 5310
rect 27288 5246 27352 5250
<< metal4 >>
rect 16801 11595 16904 11637
rect 16801 11531 16822 11595
rect 16886 11531 16904 11595
rect 16801 11487 16904 11531
rect 16802 10592 16881 11487
rect 17581 10592 19099 10593
rect 16802 10557 19099 10592
rect 16802 10493 18987 10557
rect 19051 10493 19099 10557
rect 16802 10460 19099 10493
rect 16802 10459 17623 10460
rect 11028 10362 12098 10388
rect 11028 10298 11033 10362
rect 11097 10298 12098 10362
rect 11028 10282 12098 10298
rect 11028 10218 11033 10282
rect 11097 10218 12098 10282
rect 11028 10202 12098 10218
rect 11028 10138 11033 10202
rect 11097 10138 12098 10202
rect 11028 10122 12098 10138
rect 11028 10058 11033 10122
rect 11097 10058 12098 10122
rect 11028 10042 12098 10058
rect 11028 9978 11033 10042
rect 11097 9978 12098 10042
rect 11028 9962 12098 9978
rect 11028 9898 11033 9962
rect 11097 9898 12098 9962
rect 11028 9882 12098 9898
rect 11028 9818 11033 9882
rect 11097 9818 12098 9882
rect 11028 9802 12098 9818
rect 11028 9738 11033 9802
rect 11097 9738 12098 9802
rect 11028 9722 12098 9738
rect 11028 9658 11033 9722
rect 11097 9658 12098 9722
rect 11028 9642 12098 9658
rect 11028 9578 11033 9642
rect 11097 9578 12098 9642
rect 11028 9562 12098 9578
rect 11028 9498 11033 9562
rect 11097 9498 12098 9562
rect 11028 9482 12098 9498
rect 11028 9418 11033 9482
rect 11097 9418 12098 9482
rect 11028 9402 12098 9418
rect 11028 9338 11033 9402
rect 11097 9338 12098 9402
rect 11028 9322 12098 9338
rect 11028 9258 11033 9322
rect 11097 9258 12098 9322
rect 11028 9242 12098 9258
rect 11028 9178 11033 9242
rect 11097 9178 12098 9242
rect 11028 9162 12098 9178
rect 11028 9098 11033 9162
rect 11097 9098 12098 9162
rect 11028 9082 12098 9098
rect 11028 9018 11033 9082
rect 11097 9018 12098 9082
rect 11028 9002 12098 9018
rect 11028 8938 11033 9002
rect 11097 8938 12098 9002
rect 16211 9119 16692 9147
rect 16211 9055 16618 9119
rect 16682 9055 16692 9119
rect 16211 9039 16692 9055
rect 16211 8975 16618 9039
rect 16682 8975 16692 9039
rect 16211 8947 16692 8975
rect 11028 8922 12098 8938
rect 11028 8858 11033 8922
rect 11097 8858 12098 8922
rect 11028 8811 12098 8858
rect 10534 8354 11098 8386
rect 10534 8290 10986 8354
rect 11050 8290 11098 8354
rect 10534 8262 11098 8290
rect 10534 7342 10653 8262
rect 16212 7753 16329 8947
rect 16803 8842 16882 10459
rect 20225 9132 21793 9170
rect 20225 9068 20241 9132
rect 20305 9068 21793 9132
rect 20225 9052 21793 9068
rect 20225 8988 20241 9052
rect 20305 8988 21793 9052
rect 20225 8962 21793 8988
rect 16648 8819 16882 8842
rect 16648 8755 16669 8819
rect 16733 8755 16882 8819
rect 16648 8734 16882 8755
rect 16212 7722 16687 7753
rect 16212 7658 16612 7722
rect 16676 7658 16687 7722
rect 16212 7642 16687 7658
rect 16212 7578 16612 7642
rect 16676 7578 16687 7642
rect 16212 7550 16687 7578
rect 8959 7253 10653 7342
rect 10909 7390 10986 7396
rect 10909 7364 12051 7390
rect 10909 7300 10915 7364
rect 10979 7300 12051 7364
rect 10909 7284 12051 7300
rect 8959 7198 9049 7253
rect 8959 7134 8976 7198
rect 9040 7134 9049 7198
rect 8959 7114 9049 7134
rect 10909 7220 10915 7284
rect 10979 7220 12051 7284
rect 10909 7204 12051 7220
rect 10909 7140 10915 7204
rect 10979 7140 12051 7204
rect 10909 7124 12051 7140
rect 10909 7060 10915 7124
rect 10979 7060 12051 7124
rect 10909 7044 12051 7060
rect 10909 6980 10915 7044
rect 10979 6980 12051 7044
rect 10909 6964 12051 6980
rect 10909 6900 10915 6964
rect 10979 6900 12051 6964
rect 10909 6884 12051 6900
rect 10909 6820 10915 6884
rect 10979 6820 12051 6884
rect 10909 6804 12051 6820
rect 10909 6740 10915 6804
rect 10979 6740 12051 6804
rect 10909 6724 12051 6740
rect 10909 6660 10915 6724
rect 10979 6660 12051 6724
rect 10909 6644 12051 6660
rect 10909 6580 10915 6644
rect 10979 6580 12051 6644
rect 10909 6572 12051 6580
rect 10909 6564 10986 6572
rect 10909 6500 10915 6564
rect 10979 6500 10986 6564
rect 10909 6484 10986 6500
rect 10909 6420 10915 6484
rect 10979 6420 10986 6484
rect 10909 6404 10986 6420
rect 10909 6340 10915 6404
rect 10979 6340 10986 6404
rect 10909 6324 10986 6340
rect 10909 6260 10915 6324
rect 10979 6260 10986 6324
rect 10909 6244 10986 6260
rect 10909 6180 10915 6244
rect 10979 6180 10986 6244
rect 10909 6164 10986 6180
rect 10909 6100 10915 6164
rect 10979 6100 10986 6164
rect 10909 6084 10986 6100
rect 10909 6020 10915 6084
rect 10979 6020 10986 6084
rect 10909 6004 10986 6020
rect 10909 5940 10915 6004
rect 10979 5940 10986 6004
rect 10909 5924 10986 5940
rect 10909 5860 10915 5924
rect 10979 5860 10986 5924
rect 10909 5829 10986 5860
rect 11049 6434 11140 6491
rect 11049 6370 11064 6434
rect 11128 6370 11140 6434
rect 16212 6423 16329 7550
rect 16803 7435 16882 8734
rect 17969 8851 18102 8880
rect 18881 8864 18979 8865
rect 17969 8787 18002 8851
rect 18066 8787 18102 8851
rect 16636 7422 16882 7435
rect 16636 7358 16668 7422
rect 16732 7358 16882 7422
rect 16636 7343 16882 7358
rect 17538 8718 17686 8720
rect 17538 8695 17689 8718
rect 17538 8631 17584 8695
rect 17648 8631 17689 8695
rect 17538 8615 17689 8631
rect 17538 8551 17584 8615
rect 17648 8551 17689 8615
rect 17538 8535 17689 8551
rect 17538 8471 17584 8535
rect 17648 8471 17689 8535
rect 17538 8455 17689 8471
rect 17538 8391 17584 8455
rect 17648 8391 17689 8455
rect 11049 6354 11140 6370
rect 11049 6290 11064 6354
rect 11128 6290 11140 6354
rect 11049 6274 11140 6290
rect 11049 6210 11064 6274
rect 11128 6210 11140 6274
rect 11049 6194 11140 6210
rect 11049 6130 11064 6194
rect 11128 6130 11140 6194
rect 11049 6114 11140 6130
rect 11049 6050 11064 6114
rect 11128 6050 11140 6114
rect 11049 6034 11140 6050
rect 11049 5970 11064 6034
rect 11128 5970 11140 6034
rect 11049 5954 11140 5970
rect 11049 5890 11064 5954
rect 11128 5890 11140 5954
rect 11049 5752 11140 5890
rect 11048 5349 11140 5752
rect 13158 5786 14757 6418
rect 15785 6327 16329 6423
rect 15785 6326 16323 6327
rect 13158 5722 13196 5786
rect 13260 5722 13276 5786
rect 13340 5722 13356 5786
rect 13420 5722 13436 5786
rect 13500 5722 13516 5786
rect 13580 5722 13596 5786
rect 13660 5722 13676 5786
rect 13740 5722 13756 5786
rect 13820 5722 13836 5786
rect 13900 5722 13916 5786
rect 13980 5722 13996 5786
rect 14060 5722 14076 5786
rect 14140 5722 14156 5786
rect 14220 5722 14236 5786
rect 14300 5722 14316 5786
rect 14380 5722 14396 5786
rect 14460 5722 14476 5786
rect 14540 5722 14556 5786
rect 14620 5722 14636 5786
rect 14700 5722 14757 5786
rect 13158 5710 14757 5722
rect 17538 5579 17689 8391
rect 17969 8185 18102 8787
rect 18770 8841 18979 8864
rect 18770 8777 18794 8841
rect 18858 8777 18979 8841
rect 18770 8758 18979 8777
rect 18881 8600 18979 8758
rect 17968 7170 18102 8185
rect 18880 7909 18979 8600
rect 18880 7800 18978 7909
rect 18880 7775 20147 7800
rect 18880 7711 20056 7775
rect 20120 7711 20147 7775
rect 18880 7695 20147 7711
rect 18880 7631 20056 7695
rect 20120 7631 20147 7695
rect 18880 7596 20147 7631
rect 17968 6566 18101 7170
rect 17968 6539 20162 6566
rect 17968 6475 20078 6539
rect 20142 6475 20162 6539
rect 17968 6459 20162 6475
rect 17968 6395 20078 6459
rect 20142 6395 20162 6459
rect 17968 6369 20162 6395
rect 26109 6157 27403 6368
rect 13159 5552 17689 5579
rect 13159 5488 13207 5552
rect 13271 5488 13287 5552
rect 13351 5488 13367 5552
rect 13431 5488 13447 5552
rect 13511 5488 13527 5552
rect 13591 5488 13607 5552
rect 13671 5488 13687 5552
rect 13751 5488 13767 5552
rect 13831 5488 13847 5552
rect 13911 5488 13927 5552
rect 13991 5488 14007 5552
rect 14071 5488 14087 5552
rect 14151 5488 14167 5552
rect 14231 5488 14247 5552
rect 14311 5488 14327 5552
rect 14391 5488 14407 5552
rect 14471 5488 14487 5552
rect 14551 5488 14567 5552
rect 14631 5488 14647 5552
rect 14711 5488 17689 5552
rect 13159 5467 17689 5488
rect 11048 5323 22547 5349
rect 11048 5259 22450 5323
rect 22514 5259 22547 5323
rect 11048 5234 22547 5259
rect 11048 5233 13123 5234
rect 13309 5233 22547 5234
rect 23402 5318 23527 5718
rect 23402 5254 23431 5318
rect 23495 5254 23527 5318
rect 19120 4266 20674 5233
rect 23402 5230 23527 5254
rect 27240 5390 27403 6157
rect 27240 5326 27288 5390
rect 27352 5326 27403 5390
rect 27240 5310 27403 5326
rect 27240 5246 27288 5310
rect 27352 5246 27403 5310
rect 27240 5229 27403 5246
use pseudolayout  CLKgenerator
timestamp 1669522153
transform 1 0 5266 0 1 6298
box 356 74 4887 4325
use pseudolayout  ENgenerator
timestamp 1669522153
transform -1 0 20592 0 1 10732
box 356 74 4887 4325
use Liza_Tgate  amplify
timestamp 1669522153
transform 0 -1 15126 1 0 5215
box 173 68 787 2594
use Liza_Tgate  autozero
timestamp 1669522153
transform 1 0 10524 0 1 5429
box 173 68 787 2594
use Liza_enable  bottomleft_enable
timestamp 1669522153
transform 1 0 16070 0 1 7094
box 434 356 744 1300
use Liza_enable  n_enable
timestamp 1669522153
transform 1 0 19540 0 1 7153
box 434 356 744 1300
use Liza_enable  p_enable
timestamp 1669522153
transform 1 0 19556 0 1 5912
box 434 356 744 1300
use sky130_fd_pr__pfet_01v8_J2H2S6  pass
timestamp 1669522153
transform 0 1 23685 1 0 1515
box -3371 -18281 3401 18341
use rldo  rldo_0
timestamp 1669522153
transform 1 0 12335 0 1 4667
box 5103 3281 6955 4741
use Liza_Tgate  sample
timestamp 1669522153
transform 1 0 10523 0 1 8432
box 173 68 787 2594
use sky130_fd_pr__cap_mim_m3_1_3RKQ3N  sky130_fd_pr__cap_mim_m3_1_3RKQ3N_0
timestamp 1669522153
transform 0 1 23906 -1 0 7783
box -2150 -2600 2149 2600
use sky130_fd_pr__cap_mim_m3_1_BSSJ5K  sky130_fd_pr__cap_mim_m3_1_BSSJ5K_0
timestamp 1669522153
transform 0 1 13844 -1 0 8471
box -2150 -2100 2149 2100
use sky130_fd_pr__res_generic_po_B4RDC6  sky130_fd_pr__res_generic_po_B4RDC6_0
timestamp 1669522153
transform 0 -1 22968 1 0 5288
box -33 -528 33 528
use Liza_enable  topleft_enable
timestamp 1669522153
transform 1 0 16074 0 1 8490
box 434 356 744 1300
use Liza_enable  topright_enable
timestamp 1669522153
transform 1 0 19544 0 1 8486
box 434 356 744 1300
<< labels >>
rlabel locali s 13041 5889 13041 5889 4 Vin
port 1 nsew
rlabel locali s 11204 7519 11204 7519 4 Vin
port 1 nsew
rlabel locali s 16887 9284 16921 9357 4 Vin
port 1 nsew
rlabel locali s 11197 10512 11197 10512 4 Vin
port 1 nsew
rlabel metal1 s 19753 12322 19753 12322 4 ENPin
port 2 nsew
rlabel metal1 s 10510 11916 10510 11916 4 GND
port 3 nsew
rlabel metal1 s 6105 7900 6105 7900 4 CLKin
port 4 nsew
rlabel metal1 s 4811 0 4811 0 4 Vin
port 1 nsew
rlabel metal2 s 20212 7682 20212 7682 4 NMOS_DZ
port 5 nsew
rlabel metal2 s 20224 6482 20224 6482 4 PMOS_DZ
port 6 nsew
rlabel metal2 s 10940 9192 10940 9192 4 Vref
port 7 nsew
rlabel metal2 s 18373 8572 18373 8572 4 net3
port 8 nsew
rlabel metal4 s 22086 5298 22086 5298 4 Vout
port 9 nsew
rlabel metal4 s 20644 9030 20644 9030 4 net4
port 10 nsew
rlabel metal4 s 15660 5518 15660 5518 4 net1
port 11 nsew
rlabel metal4 s 16168 6370 16168 6370 4 net6
port 12 nsew
rlabel metal4 s 11552 9167 11552 9167 4 net5
port 13 nsew
rlabel metal4 s 16826 11045 16826 11045 4 ENinverted
port 14 nsew
rlabel metal4 s 9689 7306 9689 7306 4 CLKinverted
port 15 nsew
rlabel metal3 s 17238 7620 17238 7620 4 net8
port 16 nsew
rlabel metal3 s 18662 8786 18662 8786 4 net2
port 17 nsew
rlabel metal3 s 16261 10599 16262 10600 4 EN
port 18 nsew
rlabel metal3 s 17190 8974 17190 8974 4 net7
port 19 nsew
rlabel metal3 s 9688 7158 9688 7158 4 CLK
port 20 nsew
<< end >>
