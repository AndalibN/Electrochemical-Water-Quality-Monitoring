magic
tech sky130A
magscale 1 2
timestamp 1666966674
<< nwell >>
rect 2297 6567 2685 8167
rect 5298 6567 5686 8167
use sky130_fd_pr__cap_mim_m3_1_WYFAV5  XC1
timestamp 1666963525
transform 1 0 1590 0 1 5920
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_WYFAV5  XC2
timestamp 1666963525
transform 1 0 6319 0 1 5968
box -350 -300 349 300
use sky130_fd_pr__nfet_01v8_69TA9T  XM2
timestamp 1666965885
transform 1 0 663 0 1 4243
box -287 -788 287 788
use sky130_fd_pr__nfet_01v8_HVQB9X  XM3
timestamp 1666966019
transform 1 0 1437 0 1 4243
box -545 -788 545 788
use sky130_fd_pr__pfet_01v8_4398VV  XM4
timestamp 1666965119
transform 1 0 3346 0 1 7367
box -523 -800 523 800
use sky130_fd_pr__pfet_01v8_TQ88FE  XM5
timestamp 1666963525
transform 1 0 4262 0 1 7367
box -523 -800 523 800
use sky130_fd_pr__pfet_01v8_7AWYVM  XM6
timestamp 1666965350
transform 1 0 2630 0 1 7367
box -323 -800 323 800
use sky130_fd_pr__nfet_01v8_XWWVCW  XM8
timestamp 1666966402
transform 1 0 2785 0 1 4289
box -487 -1088 487 1088
use sky130_fd_pr__nfet_01v8_XWWVCW  XM9
timestamp 1666966402
transform 1 0 3701 0 1 4289
box -487 -1088 487 1088
use sky130_fd_pr__nfet_01v8_XWWVCW  XM10
timestamp 1666966402
transform 1 0 4617 0 1 4289
box -487 -1088 487 1088
use sky130_fd_pr__pfet_01v8_3H7JSM  XM13
timestamp 1666966402
transform 1 0 5555 0 1 7367
box -194 -800 194 800
use sky130_fd_pr__nfet_01v8_HVQB9X  XMNB
timestamp 1666966019
transform 1 0 7120 0 1 4352
box -545 -788 545 788
use sky130_fd_pr__nfet_01v8_69TA9T  sky130_fd_pr__nfet_01v8_69TA9T_0
timestamp 1666965885
transform 1 0 147 0 1 4243
box -287 -788 287 788
use sky130_fd_pr__nfet_01v8_HVQB9X  sky130_fd_pr__nfet_01v8_HVQB9X_0
timestamp 1666966019
transform 1 0 8152 0 1 4352
box -545 -788 545 788
use sky130_fd_pr__nfet_01v8_XWWVCW  sky130_fd_pr__nfet_01v8_XWWVCW_0
timestamp 1666966402
transform 1 0 5533 0 1 4289
box -487 -1088 487 1088
use sky130_fd_pr__pfet_01v8_3H7JSM  sky130_fd_pr__pfet_01v8_3H7JSM_0
timestamp 1666966402
transform 1 0 2104 0 1 7367
box -194 -800 194 800
use sky130_fd_pr__pfet_01v8_7AWYVM  sky130_fd_pr__pfet_01v8_7AWYVM_0
timestamp 1666965350
transform 1 0 4978 0 1 7367
box -323 -800 323 800
<< end >>
