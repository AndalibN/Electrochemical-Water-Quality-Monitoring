magic
tech sky130A
timestamp 1668130419
<< nmos >>
rect -15 -165 15 134
<< ndiff >>
rect -44 128 -15 134
rect -44 -159 -38 128
rect -21 -159 -15 128
rect -44 -165 -15 -159
rect 15 128 44 134
rect 15 -159 21 128
rect 38 -159 44 128
rect 15 -165 44 -159
<< ndiffc >>
rect -38 -159 -21 128
rect 21 -159 38 128
<< poly >>
rect -16 170 16 178
rect -16 153 -8 170
rect 8 153 16 170
rect -16 145 16 153
rect -15 134 15 145
rect -15 -178 15 -165
<< polycont >>
rect -8 153 8 170
<< locali >>
rect -16 153 -8 170
rect 8 153 16 170
rect -38 128 -21 136
rect -38 -167 -21 -159
rect 21 128 38 136
rect 21 -167 38 -159
<< viali >>
rect -8 153 8 170
rect -38 -159 -21 128
rect 21 -159 38 128
<< metal1 >>
rect -14 170 14 173
rect -14 153 -8 170
rect 8 153 14 170
rect -14 150 14 153
rect -41 128 -18 134
rect -41 -159 -38 128
rect -21 -159 -18 128
rect -41 -165 -18 -159
rect 18 128 41 134
rect 18 -159 21 128
rect 38 -159 41 128
rect 18 -165 41 -159
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
