magic
tech sky130A
magscale 1 2
timestamp 1669744940
<< metal4 >>
rect 3400 -5532 4400 1099
rect 3400 -5768 3532 -5532
rect 3768 -5768 3932 -5532
rect 4168 -5768 4400 -5532
rect 3400 -5932 4400 -5768
rect 3400 -6168 3632 -5932
rect 3868 -6168 4032 -5932
rect 4268 -6168 4400 -5932
rect 3400 -6400 4400 -6168
<< via4 >>
rect 3532 -5768 3768 -5532
rect 3932 -5768 4168 -5532
rect 3632 -6168 3868 -5932
rect 4032 -6168 4268 -5932
<< metal5 >>
rect 1200 -3200 11600 -2200
rect 1800 -4800 10000 -3800
rect 1800 -11000 2800 -4800
rect 3400 -5532 4400 -5400
rect 3400 -5768 3532 -5532
rect 3768 -5768 3932 -5532
rect 4168 -5768 4400 -5532
rect 3400 -5932 4400 -5768
rect 3400 -6168 3632 -5932
rect 3868 -6168 4032 -5932
rect 4268 -6168 4400 -5932
rect 3400 -9200 4400 -6168
rect 9000 -9200 10000 -4800
rect 3400 -10400 10000 -9200
rect 10600 -11000 11600 -3200
rect 1800 -12000 11600 -11000
<< end >>
