magic
tech sky130A
magscale 1 2
timestamp 1666815934
<< metal3 >>
rect -3065 2987 3064 3015
rect -3065 -2987 2980 2987
rect 3044 -2987 3064 2987
rect -3065 -3015 3064 -2987
<< via3 >>
rect 2980 -2987 3044 2987
<< mimcap >>
rect -2965 2875 2865 2915
rect -2965 -2875 -2925 2875
rect 2825 -2875 2865 2875
rect -2965 -2915 2865 -2875
<< mimcapcontact >>
rect -2925 -2875 2825 2875
<< metal4 >>
rect 2964 2987 3060 3003
rect -2926 2875 2826 2876
rect -2926 -2875 -2925 2875
rect 2825 -2875 2826 2875
rect -2926 -2876 2826 -2875
rect 2964 -2987 2980 2987
rect 3044 -2987 3060 2987
rect 2964 -3003 3060 -2987
<< properties >>
string FIXED_BBOX -3065 -3015 2965 3015
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 29.15 l 29.15 val 1.721k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
