magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -23 509 23 524
rect -23 475 -17 509
rect -23 460 23 475
rect -23 105 23 120
rect -23 71 -17 105
rect -23 56 23 71
rect -23 -71 23 -56
rect -23 -105 -17 -71
rect -23 -120 23 -105
rect -23 -475 23 -460
rect -23 -509 -17 -475
rect -23 -524 23 -509
<< poly >>
rect -33 512 33 528
rect -33 478 -17 512
rect 17 478 33 512
rect -33 455 33 478
rect -33 102 33 125
rect -33 68 -17 102
rect 17 68 33 102
rect -33 52 33 68
rect -33 -68 33 -52
rect -33 -102 -17 -68
rect 17 -102 33 -68
rect -33 -125 33 -102
rect -33 -478 33 -455
rect -33 -512 -17 -478
rect 17 -512 33 -478
rect -33 -528 33 -512
<< polycont >>
rect -17 478 17 512
rect -17 68 17 102
rect -17 -102 17 -68
rect -17 -512 17 -478
<< npolyres >>
rect -33 125 33 455
rect -33 -455 33 -125
<< locali >>
rect -33 478 -17 512
rect 17 478 33 512
rect -17 472 17 475
rect -17 105 17 108
rect -33 68 -17 102
rect 17 68 33 102
rect -33 -102 -17 -68
rect 17 -102 33 -68
rect -17 -108 17 -105
rect -17 -475 17 -472
rect -33 -512 -17 -478
rect 17 -512 33 -478
<< viali >>
rect -17 478 17 509
rect -17 475 17 478
rect -17 102 17 105
rect -17 71 17 102
rect -17 -102 17 -71
rect -17 -105 17 -102
rect -17 -478 17 -475
rect -17 -509 17 -478
<< metal1 >>
rect -23 509 23 524
rect -23 475 -17 509
rect 17 475 23 509
rect -23 460 23 475
rect -23 105 23 120
rect -23 71 -17 105
rect 17 71 23 105
rect -23 56 23 71
rect -23 -71 23 -56
rect -23 -105 -17 -71
rect 17 -105 23 -71
rect -23 -120 23 -105
rect -23 -475 23 -460
rect -23 -509 -17 -475
rect 17 -509 23 -475
rect -23 -524 23 -509
<< end >>
