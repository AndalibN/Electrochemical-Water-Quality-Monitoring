magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -213 -1057 213 995
<< nmos >>
rect -129 -1031 -29 969
rect 29 -1031 129 969
<< ndiff >>
rect -187 938 -129 969
rect -187 904 -175 938
rect -141 904 -129 938
rect -187 870 -129 904
rect -187 836 -175 870
rect -141 836 -129 870
rect -187 802 -129 836
rect -187 768 -175 802
rect -141 768 -129 802
rect -187 734 -129 768
rect -187 700 -175 734
rect -141 700 -129 734
rect -187 666 -129 700
rect -187 632 -175 666
rect -141 632 -129 666
rect -187 598 -129 632
rect -187 564 -175 598
rect -141 564 -129 598
rect -187 530 -129 564
rect -187 496 -175 530
rect -141 496 -129 530
rect -187 462 -129 496
rect -187 428 -175 462
rect -141 428 -129 462
rect -187 394 -129 428
rect -187 360 -175 394
rect -141 360 -129 394
rect -187 326 -129 360
rect -187 292 -175 326
rect -141 292 -129 326
rect -187 258 -129 292
rect -187 224 -175 258
rect -141 224 -129 258
rect -187 190 -129 224
rect -187 156 -175 190
rect -141 156 -129 190
rect -187 122 -129 156
rect -187 88 -175 122
rect -141 88 -129 122
rect -187 54 -129 88
rect -187 20 -175 54
rect -141 20 -129 54
rect -187 -14 -129 20
rect -187 -48 -175 -14
rect -141 -48 -129 -14
rect -187 -82 -129 -48
rect -187 -116 -175 -82
rect -141 -116 -129 -82
rect -187 -150 -129 -116
rect -187 -184 -175 -150
rect -141 -184 -129 -150
rect -187 -218 -129 -184
rect -187 -252 -175 -218
rect -141 -252 -129 -218
rect -187 -286 -129 -252
rect -187 -320 -175 -286
rect -141 -320 -129 -286
rect -187 -354 -129 -320
rect -187 -388 -175 -354
rect -141 -388 -129 -354
rect -187 -422 -129 -388
rect -187 -456 -175 -422
rect -141 -456 -129 -422
rect -187 -490 -129 -456
rect -187 -524 -175 -490
rect -141 -524 -129 -490
rect -187 -558 -129 -524
rect -187 -592 -175 -558
rect -141 -592 -129 -558
rect -187 -626 -129 -592
rect -187 -660 -175 -626
rect -141 -660 -129 -626
rect -187 -694 -129 -660
rect -187 -728 -175 -694
rect -141 -728 -129 -694
rect -187 -762 -129 -728
rect -187 -796 -175 -762
rect -141 -796 -129 -762
rect -187 -830 -129 -796
rect -187 -864 -175 -830
rect -141 -864 -129 -830
rect -187 -898 -129 -864
rect -187 -932 -175 -898
rect -141 -932 -129 -898
rect -187 -966 -129 -932
rect -187 -1000 -175 -966
rect -141 -1000 -129 -966
rect -187 -1031 -129 -1000
rect -29 938 29 969
rect -29 904 -17 938
rect 17 904 29 938
rect -29 870 29 904
rect -29 836 -17 870
rect 17 836 29 870
rect -29 802 29 836
rect -29 768 -17 802
rect 17 768 29 802
rect -29 734 29 768
rect -29 700 -17 734
rect 17 700 29 734
rect -29 666 29 700
rect -29 632 -17 666
rect 17 632 29 666
rect -29 598 29 632
rect -29 564 -17 598
rect 17 564 29 598
rect -29 530 29 564
rect -29 496 -17 530
rect 17 496 29 530
rect -29 462 29 496
rect -29 428 -17 462
rect 17 428 29 462
rect -29 394 29 428
rect -29 360 -17 394
rect 17 360 29 394
rect -29 326 29 360
rect -29 292 -17 326
rect 17 292 29 326
rect -29 258 29 292
rect -29 224 -17 258
rect 17 224 29 258
rect -29 190 29 224
rect -29 156 -17 190
rect 17 156 29 190
rect -29 122 29 156
rect -29 88 -17 122
rect 17 88 29 122
rect -29 54 29 88
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -150 29 -116
rect -29 -184 -17 -150
rect 17 -184 29 -150
rect -29 -218 29 -184
rect -29 -252 -17 -218
rect 17 -252 29 -218
rect -29 -286 29 -252
rect -29 -320 -17 -286
rect 17 -320 29 -286
rect -29 -354 29 -320
rect -29 -388 -17 -354
rect 17 -388 29 -354
rect -29 -422 29 -388
rect -29 -456 -17 -422
rect 17 -456 29 -422
rect -29 -490 29 -456
rect -29 -524 -17 -490
rect 17 -524 29 -490
rect -29 -558 29 -524
rect -29 -592 -17 -558
rect 17 -592 29 -558
rect -29 -626 29 -592
rect -29 -660 -17 -626
rect 17 -660 29 -626
rect -29 -694 29 -660
rect -29 -728 -17 -694
rect 17 -728 29 -694
rect -29 -762 29 -728
rect -29 -796 -17 -762
rect 17 -796 29 -762
rect -29 -830 29 -796
rect -29 -864 -17 -830
rect 17 -864 29 -830
rect -29 -898 29 -864
rect -29 -932 -17 -898
rect 17 -932 29 -898
rect -29 -966 29 -932
rect -29 -1000 -17 -966
rect 17 -1000 29 -966
rect -29 -1031 29 -1000
rect 129 938 187 969
rect 129 904 141 938
rect 175 904 187 938
rect 129 870 187 904
rect 129 836 141 870
rect 175 836 187 870
rect 129 802 187 836
rect 129 768 141 802
rect 175 768 187 802
rect 129 734 187 768
rect 129 700 141 734
rect 175 700 187 734
rect 129 666 187 700
rect 129 632 141 666
rect 175 632 187 666
rect 129 598 187 632
rect 129 564 141 598
rect 175 564 187 598
rect 129 530 187 564
rect 129 496 141 530
rect 175 496 187 530
rect 129 462 187 496
rect 129 428 141 462
rect 175 428 187 462
rect 129 394 187 428
rect 129 360 141 394
rect 175 360 187 394
rect 129 326 187 360
rect 129 292 141 326
rect 175 292 187 326
rect 129 258 187 292
rect 129 224 141 258
rect 175 224 187 258
rect 129 190 187 224
rect 129 156 141 190
rect 175 156 187 190
rect 129 122 187 156
rect 129 88 141 122
rect 175 88 187 122
rect 129 54 187 88
rect 129 20 141 54
rect 175 20 187 54
rect 129 -14 187 20
rect 129 -48 141 -14
rect 175 -48 187 -14
rect 129 -82 187 -48
rect 129 -116 141 -82
rect 175 -116 187 -82
rect 129 -150 187 -116
rect 129 -184 141 -150
rect 175 -184 187 -150
rect 129 -218 187 -184
rect 129 -252 141 -218
rect 175 -252 187 -218
rect 129 -286 187 -252
rect 129 -320 141 -286
rect 175 -320 187 -286
rect 129 -354 187 -320
rect 129 -388 141 -354
rect 175 -388 187 -354
rect 129 -422 187 -388
rect 129 -456 141 -422
rect 175 -456 187 -422
rect 129 -490 187 -456
rect 129 -524 141 -490
rect 175 -524 187 -490
rect 129 -558 187 -524
rect 129 -592 141 -558
rect 175 -592 187 -558
rect 129 -626 187 -592
rect 129 -660 141 -626
rect 175 -660 187 -626
rect 129 -694 187 -660
rect 129 -728 141 -694
rect 175 -728 187 -694
rect 129 -762 187 -728
rect 129 -796 141 -762
rect 175 -796 187 -762
rect 129 -830 187 -796
rect 129 -864 141 -830
rect 175 -864 187 -830
rect 129 -898 187 -864
rect 129 -932 141 -898
rect 175 -932 187 -898
rect 129 -966 187 -932
rect 129 -1000 141 -966
rect 175 -1000 187 -966
rect 129 -1031 187 -1000
<< ndiffc >>
rect -175 904 -141 938
rect -175 836 -141 870
rect -175 768 -141 802
rect -175 700 -141 734
rect -175 632 -141 666
rect -175 564 -141 598
rect -175 496 -141 530
rect -175 428 -141 462
rect -175 360 -141 394
rect -175 292 -141 326
rect -175 224 -141 258
rect -175 156 -141 190
rect -175 88 -141 122
rect -175 20 -141 54
rect -175 -48 -141 -14
rect -175 -116 -141 -82
rect -175 -184 -141 -150
rect -175 -252 -141 -218
rect -175 -320 -141 -286
rect -175 -388 -141 -354
rect -175 -456 -141 -422
rect -175 -524 -141 -490
rect -175 -592 -141 -558
rect -175 -660 -141 -626
rect -175 -728 -141 -694
rect -175 -796 -141 -762
rect -175 -864 -141 -830
rect -175 -932 -141 -898
rect -175 -1000 -141 -966
rect -17 904 17 938
rect -17 836 17 870
rect -17 768 17 802
rect -17 700 17 734
rect -17 632 17 666
rect -17 564 17 598
rect -17 496 17 530
rect -17 428 17 462
rect -17 360 17 394
rect -17 292 17 326
rect -17 224 17 258
rect -17 156 17 190
rect -17 88 17 122
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect -17 -184 17 -150
rect -17 -252 17 -218
rect -17 -320 17 -286
rect -17 -388 17 -354
rect -17 -456 17 -422
rect -17 -524 17 -490
rect -17 -592 17 -558
rect -17 -660 17 -626
rect -17 -728 17 -694
rect -17 -796 17 -762
rect -17 -864 17 -830
rect -17 -932 17 -898
rect -17 -1000 17 -966
rect 141 904 175 938
rect 141 836 175 870
rect 141 768 175 802
rect 141 700 175 734
rect 141 632 175 666
rect 141 564 175 598
rect 141 496 175 530
rect 141 428 175 462
rect 141 360 175 394
rect 141 292 175 326
rect 141 224 175 258
rect 141 156 175 190
rect 141 88 175 122
rect 141 20 175 54
rect 141 -48 175 -14
rect 141 -116 175 -82
rect 141 -184 175 -150
rect 141 -252 175 -218
rect 141 -320 175 -286
rect 141 -388 175 -354
rect 141 -456 175 -422
rect 141 -524 175 -490
rect 141 -592 175 -558
rect 141 -660 175 -626
rect 141 -728 175 -694
rect 141 -796 175 -762
rect 141 -864 175 -830
rect 141 -932 175 -898
rect 141 -1000 175 -966
<< poly >>
rect -129 1041 -29 1057
rect -129 1007 -96 1041
rect -62 1007 -29 1041
rect -129 969 -29 1007
rect 29 1041 129 1057
rect 29 1007 62 1041
rect 96 1007 129 1041
rect 29 969 129 1007
rect -129 -1057 -29 -1031
rect 29 -1057 129 -1031
<< polycont >>
rect -96 1007 -62 1041
rect 62 1007 96 1041
<< locali >>
rect -129 1007 -96 1041
rect -62 1007 -29 1041
rect 29 1007 62 1041
rect 96 1007 129 1041
rect -175 938 -141 973
rect -175 870 -141 888
rect -175 802 -141 816
rect -175 734 -141 744
rect -175 666 -141 672
rect -175 598 -141 600
rect -175 562 -141 564
rect -175 490 -141 496
rect -175 418 -141 428
rect -175 346 -141 360
rect -175 274 -141 292
rect -175 202 -141 224
rect -175 130 -141 156
rect -175 58 -141 88
rect -175 -14 -141 20
rect -175 -82 -141 -48
rect -175 -150 -141 -120
rect -175 -218 -141 -192
rect -175 -286 -141 -264
rect -175 -354 -141 -336
rect -175 -422 -141 -408
rect -175 -490 -141 -480
rect -175 -558 -141 -552
rect -175 -626 -141 -624
rect -175 -662 -141 -660
rect -175 -734 -141 -728
rect -175 -806 -141 -796
rect -175 -878 -141 -864
rect -175 -950 -141 -932
rect -175 -1035 -141 -1000
rect -17 938 17 973
rect -17 870 17 888
rect -17 802 17 816
rect -17 734 17 744
rect -17 666 17 672
rect -17 598 17 600
rect -17 562 17 564
rect -17 490 17 496
rect -17 418 17 428
rect -17 346 17 360
rect -17 274 17 292
rect -17 202 17 224
rect -17 130 17 156
rect -17 58 17 88
rect -17 -14 17 20
rect -17 -82 17 -48
rect -17 -150 17 -120
rect -17 -218 17 -192
rect -17 -286 17 -264
rect -17 -354 17 -336
rect -17 -422 17 -408
rect -17 -490 17 -480
rect -17 -558 17 -552
rect -17 -626 17 -624
rect -17 -662 17 -660
rect -17 -734 17 -728
rect -17 -806 17 -796
rect -17 -878 17 -864
rect -17 -950 17 -932
rect -17 -1035 17 -1000
rect 141 938 175 973
rect 141 870 175 888
rect 141 802 175 816
rect 141 734 175 744
rect 141 666 175 672
rect 141 598 175 600
rect 141 562 175 564
rect 141 490 175 496
rect 141 418 175 428
rect 141 346 175 360
rect 141 274 175 292
rect 141 202 175 224
rect 141 130 175 156
rect 141 58 175 88
rect 141 -14 175 20
rect 141 -82 175 -48
rect 141 -150 175 -120
rect 141 -218 175 -192
rect 141 -286 175 -264
rect 141 -354 175 -336
rect 141 -422 175 -408
rect 141 -490 175 -480
rect 141 -558 175 -552
rect 141 -626 175 -624
rect 141 -662 175 -660
rect 141 -734 175 -728
rect 141 -806 175 -796
rect 141 -878 175 -864
rect 141 -950 175 -932
rect 141 -1035 175 -1000
<< viali >>
rect -96 1007 -62 1041
rect 62 1007 96 1041
rect -175 904 -141 922
rect -175 888 -141 904
rect -175 836 -141 850
rect -175 816 -141 836
rect -175 768 -141 778
rect -175 744 -141 768
rect -175 700 -141 706
rect -175 672 -141 700
rect -175 632 -141 634
rect -175 600 -141 632
rect -175 530 -141 562
rect -175 528 -141 530
rect -175 462 -141 490
rect -175 456 -141 462
rect -175 394 -141 418
rect -175 384 -141 394
rect -175 326 -141 346
rect -175 312 -141 326
rect -175 258 -141 274
rect -175 240 -141 258
rect -175 190 -141 202
rect -175 168 -141 190
rect -175 122 -141 130
rect -175 96 -141 122
rect -175 54 -141 58
rect -175 24 -141 54
rect -175 -48 -141 -14
rect -175 -116 -141 -86
rect -175 -120 -141 -116
rect -175 -184 -141 -158
rect -175 -192 -141 -184
rect -175 -252 -141 -230
rect -175 -264 -141 -252
rect -175 -320 -141 -302
rect -175 -336 -141 -320
rect -175 -388 -141 -374
rect -175 -408 -141 -388
rect -175 -456 -141 -446
rect -175 -480 -141 -456
rect -175 -524 -141 -518
rect -175 -552 -141 -524
rect -175 -592 -141 -590
rect -175 -624 -141 -592
rect -175 -694 -141 -662
rect -175 -696 -141 -694
rect -175 -762 -141 -734
rect -175 -768 -141 -762
rect -175 -830 -141 -806
rect -175 -840 -141 -830
rect -175 -898 -141 -878
rect -175 -912 -141 -898
rect -175 -966 -141 -950
rect -175 -984 -141 -966
rect -17 904 17 922
rect -17 888 17 904
rect -17 836 17 850
rect -17 816 17 836
rect -17 768 17 778
rect -17 744 17 768
rect -17 700 17 706
rect -17 672 17 700
rect -17 632 17 634
rect -17 600 17 632
rect -17 530 17 562
rect -17 528 17 530
rect -17 462 17 490
rect -17 456 17 462
rect -17 394 17 418
rect -17 384 17 394
rect -17 326 17 346
rect -17 312 17 326
rect -17 258 17 274
rect -17 240 17 258
rect -17 190 17 202
rect -17 168 17 190
rect -17 122 17 130
rect -17 96 17 122
rect -17 54 17 58
rect -17 24 17 54
rect -17 -48 17 -14
rect -17 -116 17 -86
rect -17 -120 17 -116
rect -17 -184 17 -158
rect -17 -192 17 -184
rect -17 -252 17 -230
rect -17 -264 17 -252
rect -17 -320 17 -302
rect -17 -336 17 -320
rect -17 -388 17 -374
rect -17 -408 17 -388
rect -17 -456 17 -446
rect -17 -480 17 -456
rect -17 -524 17 -518
rect -17 -552 17 -524
rect -17 -592 17 -590
rect -17 -624 17 -592
rect -17 -694 17 -662
rect -17 -696 17 -694
rect -17 -762 17 -734
rect -17 -768 17 -762
rect -17 -830 17 -806
rect -17 -840 17 -830
rect -17 -898 17 -878
rect -17 -912 17 -898
rect -17 -966 17 -950
rect -17 -984 17 -966
rect 141 904 175 922
rect 141 888 175 904
rect 141 836 175 850
rect 141 816 175 836
rect 141 768 175 778
rect 141 744 175 768
rect 141 700 175 706
rect 141 672 175 700
rect 141 632 175 634
rect 141 600 175 632
rect 141 530 175 562
rect 141 528 175 530
rect 141 462 175 490
rect 141 456 175 462
rect 141 394 175 418
rect 141 384 175 394
rect 141 326 175 346
rect 141 312 175 326
rect 141 258 175 274
rect 141 240 175 258
rect 141 190 175 202
rect 141 168 175 190
rect 141 122 175 130
rect 141 96 175 122
rect 141 54 175 58
rect 141 24 175 54
rect 141 -48 175 -14
rect 141 -116 175 -86
rect 141 -120 175 -116
rect 141 -184 175 -158
rect 141 -192 175 -184
rect 141 -252 175 -230
rect 141 -264 175 -252
rect 141 -320 175 -302
rect 141 -336 175 -320
rect 141 -388 175 -374
rect 141 -408 175 -388
rect 141 -456 175 -446
rect 141 -480 175 -456
rect 141 -524 175 -518
rect 141 -552 175 -524
rect 141 -592 175 -590
rect 141 -624 175 -592
rect 141 -694 175 -662
rect 141 -696 175 -694
rect 141 -762 175 -734
rect 141 -768 175 -762
rect 141 -830 175 -806
rect 141 -840 175 -830
rect 141 -898 175 -878
rect 141 -912 175 -898
rect 141 -966 175 -950
rect 141 -984 175 -966
<< metal1 >>
rect -125 1041 -33 1047
rect -125 1007 -96 1041
rect -62 1007 -33 1041
rect -125 1001 -33 1007
rect 33 1041 125 1047
rect 33 1007 62 1041
rect 96 1007 125 1041
rect 33 1001 125 1007
rect -181 922 -135 969
rect -181 888 -175 922
rect -141 888 -135 922
rect -181 850 -135 888
rect -181 816 -175 850
rect -141 816 -135 850
rect -181 778 -135 816
rect -181 744 -175 778
rect -141 744 -135 778
rect -181 706 -135 744
rect -181 672 -175 706
rect -141 672 -135 706
rect -181 634 -135 672
rect -181 600 -175 634
rect -141 600 -135 634
rect -181 562 -135 600
rect -181 528 -175 562
rect -141 528 -135 562
rect -181 490 -135 528
rect -181 456 -175 490
rect -141 456 -135 490
rect -181 418 -135 456
rect -181 384 -175 418
rect -141 384 -135 418
rect -181 346 -135 384
rect -181 312 -175 346
rect -141 312 -135 346
rect -181 274 -135 312
rect -181 240 -175 274
rect -141 240 -135 274
rect -181 202 -135 240
rect -181 168 -175 202
rect -141 168 -135 202
rect -181 130 -135 168
rect -181 96 -175 130
rect -141 96 -135 130
rect -181 58 -135 96
rect -181 24 -175 58
rect -141 24 -135 58
rect -181 -14 -135 24
rect -181 -48 -175 -14
rect -141 -48 -135 -14
rect -181 -86 -135 -48
rect -181 -120 -175 -86
rect -141 -120 -135 -86
rect -181 -158 -135 -120
rect -181 -192 -175 -158
rect -141 -192 -135 -158
rect -181 -230 -135 -192
rect -181 -264 -175 -230
rect -141 -264 -135 -230
rect -181 -302 -135 -264
rect -181 -336 -175 -302
rect -141 -336 -135 -302
rect -181 -374 -135 -336
rect -181 -408 -175 -374
rect -141 -408 -135 -374
rect -181 -446 -135 -408
rect -181 -480 -175 -446
rect -141 -480 -135 -446
rect -181 -518 -135 -480
rect -181 -552 -175 -518
rect -141 -552 -135 -518
rect -181 -590 -135 -552
rect -181 -624 -175 -590
rect -141 -624 -135 -590
rect -181 -662 -135 -624
rect -181 -696 -175 -662
rect -141 -696 -135 -662
rect -181 -734 -135 -696
rect -181 -768 -175 -734
rect -141 -768 -135 -734
rect -181 -806 -135 -768
rect -181 -840 -175 -806
rect -141 -840 -135 -806
rect -181 -878 -135 -840
rect -181 -912 -175 -878
rect -141 -912 -135 -878
rect -181 -950 -135 -912
rect -181 -984 -175 -950
rect -141 -984 -135 -950
rect -181 -1031 -135 -984
rect -23 922 23 969
rect -23 888 -17 922
rect 17 888 23 922
rect -23 850 23 888
rect -23 816 -17 850
rect 17 816 23 850
rect -23 778 23 816
rect -23 744 -17 778
rect 17 744 23 778
rect -23 706 23 744
rect -23 672 -17 706
rect 17 672 23 706
rect -23 634 23 672
rect -23 600 -17 634
rect 17 600 23 634
rect -23 562 23 600
rect -23 528 -17 562
rect 17 528 23 562
rect -23 490 23 528
rect -23 456 -17 490
rect 17 456 23 490
rect -23 418 23 456
rect -23 384 -17 418
rect 17 384 23 418
rect -23 346 23 384
rect -23 312 -17 346
rect 17 312 23 346
rect -23 274 23 312
rect -23 240 -17 274
rect 17 240 23 274
rect -23 202 23 240
rect -23 168 -17 202
rect 17 168 23 202
rect -23 130 23 168
rect -23 96 -17 130
rect 17 96 23 130
rect -23 58 23 96
rect -23 24 -17 58
rect 17 24 23 58
rect -23 -14 23 24
rect -23 -48 -17 -14
rect 17 -48 23 -14
rect -23 -86 23 -48
rect -23 -120 -17 -86
rect 17 -120 23 -86
rect -23 -158 23 -120
rect -23 -192 -17 -158
rect 17 -192 23 -158
rect -23 -230 23 -192
rect -23 -264 -17 -230
rect 17 -264 23 -230
rect -23 -302 23 -264
rect -23 -336 -17 -302
rect 17 -336 23 -302
rect -23 -374 23 -336
rect -23 -408 -17 -374
rect 17 -408 23 -374
rect -23 -446 23 -408
rect -23 -480 -17 -446
rect 17 -480 23 -446
rect -23 -518 23 -480
rect -23 -552 -17 -518
rect 17 -552 23 -518
rect -23 -590 23 -552
rect -23 -624 -17 -590
rect 17 -624 23 -590
rect -23 -662 23 -624
rect -23 -696 -17 -662
rect 17 -696 23 -662
rect -23 -734 23 -696
rect -23 -768 -17 -734
rect 17 -768 23 -734
rect -23 -806 23 -768
rect -23 -840 -17 -806
rect 17 -840 23 -806
rect -23 -878 23 -840
rect -23 -912 -17 -878
rect 17 -912 23 -878
rect -23 -950 23 -912
rect -23 -984 -17 -950
rect 17 -984 23 -950
rect -23 -1031 23 -984
rect 135 922 181 969
rect 135 888 141 922
rect 175 888 181 922
rect 135 850 181 888
rect 135 816 141 850
rect 175 816 181 850
rect 135 778 181 816
rect 135 744 141 778
rect 175 744 181 778
rect 135 706 181 744
rect 135 672 141 706
rect 175 672 181 706
rect 135 634 181 672
rect 135 600 141 634
rect 175 600 181 634
rect 135 562 181 600
rect 135 528 141 562
rect 175 528 181 562
rect 135 490 181 528
rect 135 456 141 490
rect 175 456 181 490
rect 135 418 181 456
rect 135 384 141 418
rect 175 384 181 418
rect 135 346 181 384
rect 135 312 141 346
rect 175 312 181 346
rect 135 274 181 312
rect 135 240 141 274
rect 175 240 181 274
rect 135 202 181 240
rect 135 168 141 202
rect 175 168 181 202
rect 135 130 181 168
rect 135 96 141 130
rect 175 96 181 130
rect 135 58 181 96
rect 135 24 141 58
rect 175 24 181 58
rect 135 -14 181 24
rect 135 -48 141 -14
rect 175 -48 181 -14
rect 135 -86 181 -48
rect 135 -120 141 -86
rect 175 -120 181 -86
rect 135 -158 181 -120
rect 135 -192 141 -158
rect 175 -192 181 -158
rect 135 -230 181 -192
rect 135 -264 141 -230
rect 175 -264 181 -230
rect 135 -302 181 -264
rect 135 -336 141 -302
rect 175 -336 181 -302
rect 135 -374 181 -336
rect 135 -408 141 -374
rect 175 -408 181 -374
rect 135 -446 181 -408
rect 135 -480 141 -446
rect 175 -480 181 -446
rect 135 -518 181 -480
rect 135 -552 141 -518
rect 175 -552 181 -518
rect 135 -590 181 -552
rect 135 -624 141 -590
rect 175 -624 181 -590
rect 135 -662 181 -624
rect 135 -696 141 -662
rect 175 -696 181 -662
rect 135 -734 181 -696
rect 135 -768 141 -734
rect 175 -768 181 -734
rect 135 -806 181 -768
rect 135 -840 141 -806
rect 175 -840 181 -806
rect 135 -878 181 -840
rect 135 -912 141 -878
rect 175 -912 181 -878
rect 135 -950 181 -912
rect 135 -984 141 -950
rect 175 -984 181 -950
rect 135 -1031 181 -984
<< end >>
