magic
tech sky130A
magscale 1 2
timestamp 1667788396
<< xpolycontact >>
rect -35 2000 35 2432
rect -35 -2432 35 -2000
<< ppolyres >>
rect -35 -2000 35 2000
<< viali >>
rect -19 2017 19 2414
rect -19 -2414 19 -2017
<< metal1 >>
rect -25 2414 25 2426
rect -25 2017 -19 2414
rect 19 2017 25 2414
rect -25 2005 25 2017
rect -25 -2017 25 -2005
rect -25 -2414 -19 -2017
rect 19 -2414 25 -2017
rect -25 -2426 25 -2414
<< res0p35 >>
rect -37 -2002 37 2002
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 20 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 19.387k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
