magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -8394 8272 -4048 9318
rect -8394 8242 -7276 8272
rect -7226 8242 -4048 8272
rect -8394 8095 -4048 8242
rect -8394 8094 -8379 8095
rect -6384 8094 -4048 8095
rect -8394 6800 -4048 8094
rect -8394 6624 -8370 6800
rect -8192 6624 -4048 6800
rect -8394 6598 -4048 6624
rect -8394 6586 -5768 6598
rect -4118 6586 -4048 6598
<< pwell >>
rect -9048 8112 -8850 8258
rect -6404 4070 -6012 4220
rect -8304 3432 -4010 3838
<< psubdiff >>
rect -9022 8202 -8876 8232
rect -9022 8168 -8966 8202
rect -8932 8168 -8876 8202
rect -9022 8138 -8876 8168
rect -6378 4162 -6038 4194
rect -6378 4128 -6327 4162
rect -6293 4128 -6259 4162
rect -6225 4128 -6191 4162
rect -6157 4128 -6123 4162
rect -6089 4128 -6038 4162
rect -6378 4096 -6038 4128
rect -8278 3754 -4036 3812
rect -8278 3516 -8214 3754
rect -4100 3516 -4036 3754
rect -8278 3458 -4036 3516
<< nsubdiff >>
rect -8334 9202 -4092 9260
rect -8334 8964 -8270 9202
rect -4156 8964 -4092 9202
rect -8334 8906 -4092 8964
<< psubdiffcont >>
rect -8966 8168 -8932 8202
rect -6327 4128 -6293 4162
rect -6259 4128 -6225 4162
rect -6191 4128 -6157 4162
rect -6123 4128 -6089 4162
rect -8214 3516 -4100 3754
<< nsubdiffcont >>
rect -8270 8964 -4156 9202
<< poly >>
rect -5834 8724 -5672 8796
rect -5832 6600 -5574 6642
<< locali >>
rect -8318 9208 -4108 9244
rect -8318 8958 -8282 9208
rect -4144 8958 -4108 9208
rect -8318 8922 -4108 8958
rect -9014 8202 -8884 8224
rect -9014 8168 -9002 8202
rect -8968 8168 -8966 8202
rect -8932 8168 -8930 8202
rect -8896 8168 -8884 8202
rect -9014 8146 -8884 8168
rect -8352 8051 -8208 8070
rect -8352 7945 -8333 8051
rect -8227 7945 -8208 8051
rect -8352 7926 -8208 7945
rect -6370 4162 -6046 4186
rect -6370 4128 -6333 4162
rect -6293 4128 -6261 4162
rect -6225 4128 -6191 4162
rect -6155 4128 -6123 4162
rect -6083 4128 -6046 4162
rect -6370 4104 -6046 4128
rect -8262 3760 -4052 3796
rect -8262 3510 -8226 3760
rect -4088 3510 -4052 3760
rect -8262 3474 -4052 3510
<< viali >>
rect -8282 9202 -4144 9208
rect -8282 8964 -8270 9202
rect -8270 8964 -4156 9202
rect -4156 8964 -4144 9202
rect -8282 8958 -4144 8964
rect -9002 8168 -8968 8202
rect -8930 8168 -8896 8202
rect -8333 7945 -8227 8051
rect -6333 4128 -6327 4162
rect -6327 4128 -6299 4162
rect -6261 4128 -6259 4162
rect -6259 4128 -6227 4162
rect -6189 4128 -6157 4162
rect -6157 4128 -6155 4162
rect -6117 4128 -6089 4162
rect -6089 4128 -6083 4162
rect -8226 3754 -4088 3760
rect -8226 3516 -8214 3754
rect -8214 3516 -4100 3754
rect -4100 3516 -4088 3754
rect -8226 3510 -4088 3516
<< metal1 >>
rect -8318 9208 -4108 9244
rect -8318 8958 -8282 9208
rect -4144 8958 -4108 9208
rect -8318 8922 -4108 8958
rect -5726 8830 -4152 8922
rect -8330 8740 -8244 8788
rect -7284 8740 -7218 8788
rect -8330 8688 -8288 8740
rect -8326 8684 -8288 8688
rect -7280 8686 -7222 8706
rect -9186 8572 -9008 8638
rect -7280 8634 -7277 8686
rect -7225 8634 -7222 8686
rect -7280 8622 -7222 8634
rect -9186 8540 -8880 8572
rect -7280 8570 -7277 8622
rect -7225 8570 -7222 8622
rect -7280 8558 -7222 8570
rect -9186 8462 -9008 8540
rect -7280 8506 -7277 8558
rect -7225 8506 -7222 8558
rect -7280 8494 -7222 8506
rect -8972 8224 -8926 8432
rect -8508 8312 -8292 8488
rect -7280 8442 -7277 8494
rect -7225 8442 -7222 8494
rect -7280 8430 -7222 8442
rect -7280 8378 -7277 8430
rect -7225 8378 -7222 8430
rect -7280 8366 -7222 8378
rect -7280 8314 -7277 8366
rect -7225 8314 -7222 8366
rect -7280 8294 -7222 8314
rect -9014 8202 -8884 8224
rect -9014 8168 -9002 8202
rect -8968 8168 -8930 8202
rect -8896 8168 -8884 8202
rect -9014 8146 -8884 8168
rect -6216 8132 -6170 8302
rect -6582 8098 -6170 8132
rect -8370 8051 -8192 8086
rect -8370 7945 -8333 8051
rect -8227 7945 -8192 8051
rect -8370 7910 -8192 7945
rect -8370 6624 -8192 6800
rect -5884 6658 -5838 6714
rect -6202 6606 -6102 6612
rect -6202 6554 -6178 6606
rect -6126 6554 -6102 6606
rect -5884 6610 -5732 6658
rect -5884 6600 -5782 6610
rect -6630 6484 -6596 6488
rect -6614 6278 -6580 6484
rect -6202 6356 -6102 6554
rect -6472 6310 -5944 6356
rect -6614 6246 -6478 6278
rect -6254 6262 -6208 6310
rect -5832 6278 -5782 6600
rect -3874 6580 -3540 6700
rect -5726 6534 -5568 6580
rect -4258 6538 -3540 6580
rect -4258 6534 -3718 6538
rect -5726 6486 -3718 6534
rect -3666 6486 -3540 6538
rect -5726 6484 -3540 6486
rect -4110 6438 -3540 6484
rect -3874 6320 -3540 6438
rect -5932 6234 -5782 6278
rect -6524 4020 -6478 4290
rect -6366 4182 -6318 4284
rect -6096 4182 -6050 4288
rect -6366 4171 -6050 4182
rect -6366 4162 -6329 4171
rect -6366 4128 -6333 4162
rect -6366 4119 -6329 4128
rect -6277 4119 -6265 4171
rect -6213 4119 -6201 4171
rect -6149 4119 -6137 4171
rect -6085 4162 -6050 4171
rect -6083 4128 -6050 4162
rect -6085 4119 -6050 4128
rect -6366 4108 -6050 4119
rect -5702 4268 -5596 4324
rect -5702 4020 -5624 4268
rect -6524 3986 -5624 4020
rect -6524 3934 -6448 3986
rect -6396 3934 -5624 3986
rect -6524 3900 -5624 3934
rect -5568 3796 -4258 4234
rect -8262 3760 -4052 3796
rect -8262 3510 -8226 3760
rect -4088 3510 -4052 3760
rect -8262 3474 -4052 3510
<< via1 >>
rect -7277 9033 -7225 9085
rect -7277 8969 -7225 9021
rect -7277 8634 -7225 8686
rect -7277 8570 -7225 8622
rect -7277 8506 -7225 8558
rect -7277 8442 -7225 8494
rect -7277 8378 -7225 8430
rect -7277 8314 -7225 8366
rect -6178 6554 -6126 6606
rect -3718 6486 -3666 6538
rect -6329 4162 -6277 4171
rect -6329 4128 -6299 4162
rect -6299 4128 -6277 4162
rect -6329 4119 -6277 4128
rect -6265 4162 -6213 4171
rect -6265 4128 -6261 4162
rect -6261 4128 -6227 4162
rect -6227 4128 -6213 4162
rect -6265 4119 -6213 4128
rect -6201 4162 -6149 4171
rect -6201 4128 -6189 4162
rect -6189 4128 -6155 4162
rect -6155 4128 -6149 4162
rect -6201 4119 -6149 4128
rect -6137 4162 -6085 4171
rect -6137 4128 -6117 4162
rect -6117 4128 -6085 4162
rect -6137 4119 -6085 4128
rect -6448 3934 -6396 3986
rect -6236 3646 -6184 3698
<< metal2 >>
rect -7280 9085 -7222 9114
rect -7280 9033 -7277 9085
rect -7225 9033 -7222 9085
rect -7280 9021 -7222 9033
rect -7280 8969 -7277 9021
rect -7225 8969 -7222 9021
rect -7280 8686 -7222 8969
rect -7280 8634 -7277 8686
rect -7225 8634 -7222 8686
rect -7280 8622 -7222 8634
rect -7280 8570 -7277 8622
rect -7225 8570 -7222 8622
rect -7280 8558 -7222 8570
rect -7280 8506 -7277 8558
rect -7225 8506 -7222 8558
rect -7280 8494 -7222 8506
rect -7280 8442 -7277 8494
rect -7225 8442 -7222 8494
rect -7280 8430 -7222 8442
rect -7280 8378 -7277 8430
rect -7225 8378 -7222 8430
rect -7280 8366 -7222 8378
rect -7280 8314 -7277 8366
rect -7225 8314 -7222 8366
rect -7280 8294 -7222 8314
rect -6648 6606 -6102 6612
rect -6648 6554 -6178 6606
rect -6126 6554 -6102 6606
rect -6648 6548 -6102 6554
rect -3728 6540 -3656 6566
rect -3728 6484 -3720 6540
rect -3664 6484 -3656 6540
rect -3728 6458 -3656 6484
rect -6366 4171 -6050 4182
rect -6366 4119 -6329 4171
rect -6277 4119 -6265 4171
rect -6213 4119 -6201 4171
rect -6149 4119 -6137 4171
rect -6085 4119 -6050 4171
rect -6366 4108 -6050 4119
rect -6458 3988 -6386 4014
rect -6458 3932 -6450 3988
rect -6394 3932 -6386 3988
rect -6458 3906 -6386 3932
rect -6228 3704 -6194 4108
rect -6260 3698 -6160 3704
rect -6260 3646 -6236 3698
rect -6184 3646 -6160 3698
rect -6260 3640 -6160 3646
<< via2 >>
rect -3720 6538 -3664 6540
rect -3720 6486 -3718 6538
rect -3718 6486 -3666 6538
rect -3666 6486 -3664 6538
rect -3720 6484 -3664 6486
rect -6450 3986 -6394 3988
rect -6450 3934 -6448 3986
rect -6448 3934 -6396 3986
rect -6396 3934 -6394 3986
rect -6450 3932 -6394 3934
<< metal3 >>
rect -3734 6544 -3634 6572
rect -3734 6480 -3724 6544
rect -3660 6480 -3634 6544
rect -3734 6452 -3634 6480
rect -6464 3992 -6380 4020
rect -6464 3928 -6454 3992
rect -6390 3928 -6380 3992
rect -6464 3900 -6380 3928
<< via3 >>
rect -3724 6540 -3660 6544
rect -3724 6484 -3720 6540
rect -3720 6484 -3664 6540
rect -3664 6484 -3660 6540
rect -3724 6480 -3660 6484
rect -6454 3988 -6390 3992
rect -6454 3932 -6450 3988
rect -6450 3932 -6394 3988
rect -6394 3932 -6390 3988
rect -6454 3928 -6390 3932
<< metal4 >>
rect -3872 6544 -2242 6730
rect -3872 6480 -3724 6544
rect -3660 6480 -2242 6544
rect -9003 3264 -8351 4396
rect -6748 4020 -6634 4204
rect -6748 3992 -6380 4020
rect -6748 3928 -6454 3992
rect -6390 3928 -6380 3992
rect -6748 3900 -6380 3928
rect -3872 3264 -2242 6480
rect -9003 2577 -2242 3264
rect -8989 2573 -2242 2577
rect -8989 2572 -3337 2573
use sky130_fd_pr__nfet_01v8_JSTS37  XM4
timestamp 1669522153
transform 1 0 -6073 0 1 5309
box -213 -1057 213 1057
use sky130_fd_pr__pfet_01v8_G3EKZ5  XM6
timestamp 1669522153
transform 1 0 -5782 0 1 7662
box -144 -1064 144 1098
use sky130_fd_pr__pfet_01v8_GCY946  XM7
timestamp 1669522153
transform 1 0 -4916 0 1 7698
box -852 -1174 858 1174
use sky130_fd_pr__nfet_01v8_U894CR  XM8
timestamp 1669522153
transform 1 0 -4914 0 1 5324
box -844 -1136 846 1186
use sky130_fd_pr__pfet_01v8_MV88VP  XM9
timestamp 1669522153
transform 1 0 -7251 0 1 8536
box -1123 -298 1123 264
use sky130_fd_pr__nfet_01v8_N3YEAS  XM10
timestamp 1669522153
transform 1 0 -8720 0 1 8432
box -284 -157 284 157
use sky130_fd_pr__cap_mim_m3_1_A5GGR2  sky130_fd_pr__cap_mim_m3_1_A5GGR2_0
timestamp 1669522153
transform 1 0 -7893 0 1 5219
box -1249 -1199 1248 1199
use sky130_fd_pr__nfet_01v8_QAUSEG  sky130_fd_pr__nfet_01v8_QAUSEG_0
timestamp 1669522153
transform 1 0 -6422 0 1 5309
box -134 -1057 134 1057
use sky130_fd_pr__pfet_01v8_NDY9L5  sky130_fd_pr__pfet_01v8_NDY9L5_0
timestamp 1669522153
transform 1 0 -5037 0 1 7675
box -3343 -1193 -1297 457
<< labels >>
rlabel metal1 s -8352 7926 -8208 8070 4 nVin
port 1 nsew
rlabel metal1 s -8352 6640 -8208 6784 4 pVin
port 2 nsew
rlabel metal1 s -3874 6320 -3540 6700 4 Vout
port 3 nsew
rlabel metal1 s -9186 8462 -9008 8638 4 VBias
port 4 nsew
rlabel metal1 s -8302 8938 -4124 9228 4 VDD
port 5 nsew
rlabel metal1 s -8246 3490 -4068 3780 4 AGND
port 6 nsew
<< end >>
