magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 332 35 764
rect -35 -764 35 -332
<< xpolyres >>
rect -35 -332 35 332
<< viali >>
rect -17 710 17 744
rect -17 638 17 672
rect -17 566 17 600
rect -17 494 17 528
rect -17 422 17 456
rect -17 350 17 384
rect -17 -385 17 -351
rect -17 -457 17 -423
rect -17 -529 17 -495
rect -17 -601 17 -567
rect -17 -673 17 -639
rect -17 -745 17 -711
<< metal1 >>
rect -25 744 25 758
rect -25 710 -17 744
rect 17 710 25 744
rect -25 672 25 710
rect -25 638 -17 672
rect 17 638 25 672
rect -25 600 25 638
rect -25 566 -17 600
rect 17 566 25 600
rect -25 528 25 566
rect -25 494 -17 528
rect 17 494 25 528
rect -25 456 25 494
rect -25 422 -17 456
rect 17 422 25 456
rect -25 384 25 422
rect -25 350 -17 384
rect 17 350 25 384
rect -25 337 25 350
rect -25 -351 25 -337
rect -25 -385 -17 -351
rect 17 -385 25 -351
rect -25 -423 25 -385
rect -25 -457 -17 -423
rect 17 -457 25 -423
rect -25 -495 25 -457
rect -25 -529 -17 -495
rect 17 -529 25 -495
rect -25 -567 25 -529
rect -25 -601 -17 -567
rect 17 -601 25 -567
rect -25 -639 25 -601
rect -25 -673 -17 -639
rect 17 -673 25 -639
rect -25 -711 25 -673
rect -25 -745 -17 -711
rect 17 -745 25 -711
rect -25 -758 25 -745
<< end >>
