magic
tech sky130A
magscale 1 2
timestamp 1668369161
<< error_p >>
rect -2813 9672 -2755 9678
rect -2581 9672 -2523 9678
rect -2349 9672 -2291 9678
rect -2117 9672 -2059 9678
rect -1885 9672 -1827 9678
rect -1653 9672 -1595 9678
rect -1421 9672 -1363 9678
rect -1189 9672 -1131 9678
rect -957 9672 -899 9678
rect -725 9672 -667 9678
rect -493 9672 -435 9678
rect -261 9672 -203 9678
rect -29 9672 29 9678
rect 203 9672 261 9678
rect 435 9672 493 9678
rect 667 9672 725 9678
rect 899 9672 957 9678
rect 1131 9672 1189 9678
rect 1363 9672 1421 9678
rect 1595 9672 1653 9678
rect 1827 9672 1885 9678
rect 2059 9672 2117 9678
rect 2291 9672 2349 9678
rect 2523 9672 2581 9678
rect 2755 9672 2813 9678
rect -2813 9638 -2801 9672
rect -2581 9638 -2569 9672
rect -2349 9638 -2337 9672
rect -2117 9638 -2105 9672
rect -1885 9638 -1873 9672
rect -1653 9638 -1641 9672
rect -1421 9638 -1409 9672
rect -1189 9638 -1177 9672
rect -957 9638 -945 9672
rect -725 9638 -713 9672
rect -493 9638 -481 9672
rect -261 9638 -249 9672
rect -29 9638 -17 9672
rect 203 9638 215 9672
rect 435 9638 447 9672
rect 667 9638 679 9672
rect 899 9638 911 9672
rect 1131 9638 1143 9672
rect 1363 9638 1375 9672
rect 1595 9638 1607 9672
rect 1827 9638 1839 9672
rect 2059 9638 2071 9672
rect 2291 9638 2303 9672
rect 2523 9638 2535 9672
rect 2755 9638 2767 9672
rect -2813 9632 -2755 9638
rect -2581 9632 -2523 9638
rect -2349 9632 -2291 9638
rect -2117 9632 -2059 9638
rect -1885 9632 -1827 9638
rect -1653 9632 -1595 9638
rect -1421 9632 -1363 9638
rect -1189 9632 -1131 9638
rect -957 9632 -899 9638
rect -725 9632 -667 9638
rect -493 9632 -435 9638
rect -261 9632 -203 9638
rect -29 9632 29 9638
rect 203 9632 261 9638
rect 435 9632 493 9638
rect 667 9632 725 9638
rect 899 9632 957 9638
rect 1131 9632 1189 9638
rect 1363 9632 1421 9638
rect 1595 9632 1653 9638
rect 1827 9632 1885 9638
rect 2059 9632 2117 9638
rect 2291 9632 2349 9638
rect 2523 9632 2581 9638
rect 2755 9632 2813 9638
rect -2813 -9638 -2755 -9632
rect -2581 -9638 -2523 -9632
rect -2349 -9638 -2291 -9632
rect -2117 -9638 -2059 -9632
rect -1885 -9638 -1827 -9632
rect -1653 -9638 -1595 -9632
rect -1421 -9638 -1363 -9632
rect -1189 -9638 -1131 -9632
rect -957 -9638 -899 -9632
rect -725 -9638 -667 -9632
rect -493 -9638 -435 -9632
rect -261 -9638 -203 -9632
rect -29 -9638 29 -9632
rect 203 -9638 261 -9632
rect 435 -9638 493 -9632
rect 667 -9638 725 -9632
rect 899 -9638 957 -9632
rect 1131 -9638 1189 -9632
rect 1363 -9638 1421 -9632
rect 1595 -9638 1653 -9632
rect 1827 -9638 1885 -9632
rect 2059 -9638 2117 -9632
rect 2291 -9638 2349 -9632
rect 2523 -9638 2581 -9632
rect 2755 -9638 2813 -9632
rect -2813 -9672 -2801 -9638
rect -2581 -9672 -2569 -9638
rect -2349 -9672 -2337 -9638
rect -2117 -9672 -2105 -9638
rect -1885 -9672 -1873 -9638
rect -1653 -9672 -1641 -9638
rect -1421 -9672 -1409 -9638
rect -1189 -9672 -1177 -9638
rect -957 -9672 -945 -9638
rect -725 -9672 -713 -9638
rect -493 -9672 -481 -9638
rect -261 -9672 -249 -9638
rect -29 -9672 -17 -9638
rect 203 -9672 215 -9638
rect 435 -9672 447 -9638
rect 667 -9672 679 -9638
rect 899 -9672 911 -9638
rect 1131 -9672 1143 -9638
rect 1363 -9672 1375 -9638
rect 1595 -9672 1607 -9638
rect 1827 -9672 1839 -9638
rect 2059 -9672 2071 -9638
rect 2291 -9672 2303 -9638
rect 2523 -9672 2535 -9638
rect 2755 -9672 2767 -9638
rect -2813 -9678 -2755 -9672
rect -2581 -9678 -2523 -9672
rect -2349 -9678 -2291 -9672
rect -2117 -9678 -2059 -9672
rect -1885 -9678 -1827 -9672
rect -1653 -9678 -1595 -9672
rect -1421 -9678 -1363 -9672
rect -1189 -9678 -1131 -9672
rect -957 -9678 -899 -9672
rect -725 -9678 -667 -9672
rect -493 -9678 -435 -9672
rect -261 -9678 -203 -9672
rect -29 -9678 29 -9672
rect 203 -9678 261 -9672
rect 435 -9678 493 -9672
rect 667 -9678 725 -9672
rect 899 -9678 957 -9672
rect 1131 -9678 1189 -9672
rect 1363 -9678 1421 -9672
rect 1595 -9678 1653 -9672
rect 1827 -9678 1885 -9672
rect 2059 -9678 2117 -9672
rect 2291 -9678 2349 -9672
rect 2523 -9678 2581 -9672
rect 2755 -9678 2813 -9672
<< nmos >>
rect -2814 -9600 -2754 9600
rect -2582 -9600 -2522 9600
rect -2350 -9600 -2290 9600
rect -2118 -9600 -2058 9600
rect -1886 -9600 -1826 9600
rect -1654 -9600 -1594 9600
rect -1422 -9600 -1362 9600
rect -1190 -9600 -1130 9600
rect -958 -9600 -898 9600
rect -726 -9600 -666 9600
rect -494 -9600 -434 9600
rect -262 -9600 -202 9600
rect -30 -9600 30 9600
rect 202 -9600 262 9600
rect 434 -9600 494 9600
rect 666 -9600 726 9600
rect 898 -9600 958 9600
rect 1130 -9600 1190 9600
rect 1362 -9600 1422 9600
rect 1594 -9600 1654 9600
rect 1826 -9600 1886 9600
rect 2058 -9600 2118 9600
rect 2290 -9600 2350 9600
rect 2522 -9600 2582 9600
rect 2754 -9600 2814 9600
<< ndiff >>
rect -2872 9588 -2814 9600
rect -2872 -9588 -2860 9588
rect -2826 -9588 -2814 9588
rect -2872 -9600 -2814 -9588
rect -2754 9588 -2696 9600
rect -2754 -9588 -2742 9588
rect -2708 -9588 -2696 9588
rect -2754 -9600 -2696 -9588
rect -2640 9588 -2582 9600
rect -2640 -9588 -2628 9588
rect -2594 -9588 -2582 9588
rect -2640 -9600 -2582 -9588
rect -2522 9588 -2464 9600
rect -2522 -9588 -2510 9588
rect -2476 -9588 -2464 9588
rect -2522 -9600 -2464 -9588
rect -2408 9588 -2350 9600
rect -2408 -9588 -2396 9588
rect -2362 -9588 -2350 9588
rect -2408 -9600 -2350 -9588
rect -2290 9588 -2232 9600
rect -2290 -9588 -2278 9588
rect -2244 -9588 -2232 9588
rect -2290 -9600 -2232 -9588
rect -2176 9588 -2118 9600
rect -2176 -9588 -2164 9588
rect -2130 -9588 -2118 9588
rect -2176 -9600 -2118 -9588
rect -2058 9588 -2000 9600
rect -2058 -9588 -2046 9588
rect -2012 -9588 -2000 9588
rect -2058 -9600 -2000 -9588
rect -1944 9588 -1886 9600
rect -1944 -9588 -1932 9588
rect -1898 -9588 -1886 9588
rect -1944 -9600 -1886 -9588
rect -1826 9588 -1768 9600
rect -1826 -9588 -1814 9588
rect -1780 -9588 -1768 9588
rect -1826 -9600 -1768 -9588
rect -1712 9588 -1654 9600
rect -1712 -9588 -1700 9588
rect -1666 -9588 -1654 9588
rect -1712 -9600 -1654 -9588
rect -1594 9588 -1536 9600
rect -1594 -9588 -1582 9588
rect -1548 -9588 -1536 9588
rect -1594 -9600 -1536 -9588
rect -1480 9588 -1422 9600
rect -1480 -9588 -1468 9588
rect -1434 -9588 -1422 9588
rect -1480 -9600 -1422 -9588
rect -1362 9588 -1304 9600
rect -1362 -9588 -1350 9588
rect -1316 -9588 -1304 9588
rect -1362 -9600 -1304 -9588
rect -1248 9588 -1190 9600
rect -1248 -9588 -1236 9588
rect -1202 -9588 -1190 9588
rect -1248 -9600 -1190 -9588
rect -1130 9588 -1072 9600
rect -1130 -9588 -1118 9588
rect -1084 -9588 -1072 9588
rect -1130 -9600 -1072 -9588
rect -1016 9588 -958 9600
rect -1016 -9588 -1004 9588
rect -970 -9588 -958 9588
rect -1016 -9600 -958 -9588
rect -898 9588 -840 9600
rect -898 -9588 -886 9588
rect -852 -9588 -840 9588
rect -898 -9600 -840 -9588
rect -784 9588 -726 9600
rect -784 -9588 -772 9588
rect -738 -9588 -726 9588
rect -784 -9600 -726 -9588
rect -666 9588 -608 9600
rect -666 -9588 -654 9588
rect -620 -9588 -608 9588
rect -666 -9600 -608 -9588
rect -552 9588 -494 9600
rect -552 -9588 -540 9588
rect -506 -9588 -494 9588
rect -552 -9600 -494 -9588
rect -434 9588 -376 9600
rect -434 -9588 -422 9588
rect -388 -9588 -376 9588
rect -434 -9600 -376 -9588
rect -320 9588 -262 9600
rect -320 -9588 -308 9588
rect -274 -9588 -262 9588
rect -320 -9600 -262 -9588
rect -202 9588 -144 9600
rect -202 -9588 -190 9588
rect -156 -9588 -144 9588
rect -202 -9600 -144 -9588
rect -88 9588 -30 9600
rect -88 -9588 -76 9588
rect -42 -9588 -30 9588
rect -88 -9600 -30 -9588
rect 30 9588 88 9600
rect 30 -9588 42 9588
rect 76 -9588 88 9588
rect 30 -9600 88 -9588
rect 144 9588 202 9600
rect 144 -9588 156 9588
rect 190 -9588 202 9588
rect 144 -9600 202 -9588
rect 262 9588 320 9600
rect 262 -9588 274 9588
rect 308 -9588 320 9588
rect 262 -9600 320 -9588
rect 376 9588 434 9600
rect 376 -9588 388 9588
rect 422 -9588 434 9588
rect 376 -9600 434 -9588
rect 494 9588 552 9600
rect 494 -9588 506 9588
rect 540 -9588 552 9588
rect 494 -9600 552 -9588
rect 608 9588 666 9600
rect 608 -9588 620 9588
rect 654 -9588 666 9588
rect 608 -9600 666 -9588
rect 726 9588 784 9600
rect 726 -9588 738 9588
rect 772 -9588 784 9588
rect 726 -9600 784 -9588
rect 840 9588 898 9600
rect 840 -9588 852 9588
rect 886 -9588 898 9588
rect 840 -9600 898 -9588
rect 958 9588 1016 9600
rect 958 -9588 970 9588
rect 1004 -9588 1016 9588
rect 958 -9600 1016 -9588
rect 1072 9588 1130 9600
rect 1072 -9588 1084 9588
rect 1118 -9588 1130 9588
rect 1072 -9600 1130 -9588
rect 1190 9588 1248 9600
rect 1190 -9588 1202 9588
rect 1236 -9588 1248 9588
rect 1190 -9600 1248 -9588
rect 1304 9588 1362 9600
rect 1304 -9588 1316 9588
rect 1350 -9588 1362 9588
rect 1304 -9600 1362 -9588
rect 1422 9588 1480 9600
rect 1422 -9588 1434 9588
rect 1468 -9588 1480 9588
rect 1422 -9600 1480 -9588
rect 1536 9588 1594 9600
rect 1536 -9588 1548 9588
rect 1582 -9588 1594 9588
rect 1536 -9600 1594 -9588
rect 1654 9588 1712 9600
rect 1654 -9588 1666 9588
rect 1700 -9588 1712 9588
rect 1654 -9600 1712 -9588
rect 1768 9588 1826 9600
rect 1768 -9588 1780 9588
rect 1814 -9588 1826 9588
rect 1768 -9600 1826 -9588
rect 1886 9588 1944 9600
rect 1886 -9588 1898 9588
rect 1932 -9588 1944 9588
rect 1886 -9600 1944 -9588
rect 2000 9588 2058 9600
rect 2000 -9588 2012 9588
rect 2046 -9588 2058 9588
rect 2000 -9600 2058 -9588
rect 2118 9588 2176 9600
rect 2118 -9588 2130 9588
rect 2164 -9588 2176 9588
rect 2118 -9600 2176 -9588
rect 2232 9588 2290 9600
rect 2232 -9588 2244 9588
rect 2278 -9588 2290 9588
rect 2232 -9600 2290 -9588
rect 2350 9588 2408 9600
rect 2350 -9588 2362 9588
rect 2396 -9588 2408 9588
rect 2350 -9600 2408 -9588
rect 2464 9588 2522 9600
rect 2464 -9588 2476 9588
rect 2510 -9588 2522 9588
rect 2464 -9600 2522 -9588
rect 2582 9588 2640 9600
rect 2582 -9588 2594 9588
rect 2628 -9588 2640 9588
rect 2582 -9600 2640 -9588
rect 2696 9588 2754 9600
rect 2696 -9588 2708 9588
rect 2742 -9588 2754 9588
rect 2696 -9600 2754 -9588
rect 2814 9588 2872 9600
rect 2814 -9588 2826 9588
rect 2860 -9588 2872 9588
rect 2814 -9600 2872 -9588
<< ndiffc >>
rect -2860 -9588 -2826 9588
rect -2742 -9588 -2708 9588
rect -2628 -9588 -2594 9588
rect -2510 -9588 -2476 9588
rect -2396 -9588 -2362 9588
rect -2278 -9588 -2244 9588
rect -2164 -9588 -2130 9588
rect -2046 -9588 -2012 9588
rect -1932 -9588 -1898 9588
rect -1814 -9588 -1780 9588
rect -1700 -9588 -1666 9588
rect -1582 -9588 -1548 9588
rect -1468 -9588 -1434 9588
rect -1350 -9588 -1316 9588
rect -1236 -9588 -1202 9588
rect -1118 -9588 -1084 9588
rect -1004 -9588 -970 9588
rect -886 -9588 -852 9588
rect -772 -9588 -738 9588
rect -654 -9588 -620 9588
rect -540 -9588 -506 9588
rect -422 -9588 -388 9588
rect -308 -9588 -274 9588
rect -190 -9588 -156 9588
rect -76 -9588 -42 9588
rect 42 -9588 76 9588
rect 156 -9588 190 9588
rect 274 -9588 308 9588
rect 388 -9588 422 9588
rect 506 -9588 540 9588
rect 620 -9588 654 9588
rect 738 -9588 772 9588
rect 852 -9588 886 9588
rect 970 -9588 1004 9588
rect 1084 -9588 1118 9588
rect 1202 -9588 1236 9588
rect 1316 -9588 1350 9588
rect 1434 -9588 1468 9588
rect 1548 -9588 1582 9588
rect 1666 -9588 1700 9588
rect 1780 -9588 1814 9588
rect 1898 -9588 1932 9588
rect 2012 -9588 2046 9588
rect 2130 -9588 2164 9588
rect 2244 -9588 2278 9588
rect 2362 -9588 2396 9588
rect 2476 -9588 2510 9588
rect 2594 -9588 2628 9588
rect 2708 -9588 2742 9588
rect 2826 -9588 2860 9588
<< poly >>
rect -2817 9672 -2751 9688
rect -2817 9638 -2801 9672
rect -2767 9638 -2751 9672
rect -2817 9622 -2751 9638
rect -2585 9672 -2519 9688
rect -2585 9638 -2569 9672
rect -2535 9638 -2519 9672
rect -2585 9622 -2519 9638
rect -2353 9672 -2287 9688
rect -2353 9638 -2337 9672
rect -2303 9638 -2287 9672
rect -2353 9622 -2287 9638
rect -2121 9672 -2055 9688
rect -2121 9638 -2105 9672
rect -2071 9638 -2055 9672
rect -2121 9622 -2055 9638
rect -1889 9672 -1823 9688
rect -1889 9638 -1873 9672
rect -1839 9638 -1823 9672
rect -1889 9622 -1823 9638
rect -1657 9672 -1591 9688
rect -1657 9638 -1641 9672
rect -1607 9638 -1591 9672
rect -1657 9622 -1591 9638
rect -1425 9672 -1359 9688
rect -1425 9638 -1409 9672
rect -1375 9638 -1359 9672
rect -1425 9622 -1359 9638
rect -1193 9672 -1127 9688
rect -1193 9638 -1177 9672
rect -1143 9638 -1127 9672
rect -1193 9622 -1127 9638
rect -961 9672 -895 9688
rect -961 9638 -945 9672
rect -911 9638 -895 9672
rect -961 9622 -895 9638
rect -729 9672 -663 9688
rect -729 9638 -713 9672
rect -679 9638 -663 9672
rect -729 9622 -663 9638
rect -497 9672 -431 9688
rect -497 9638 -481 9672
rect -447 9638 -431 9672
rect -497 9622 -431 9638
rect -265 9672 -199 9688
rect -265 9638 -249 9672
rect -215 9638 -199 9672
rect -265 9622 -199 9638
rect -33 9672 33 9688
rect -33 9638 -17 9672
rect 17 9638 33 9672
rect -33 9622 33 9638
rect 199 9672 265 9688
rect 199 9638 215 9672
rect 249 9638 265 9672
rect 199 9622 265 9638
rect 431 9672 497 9688
rect 431 9638 447 9672
rect 481 9638 497 9672
rect 431 9622 497 9638
rect 663 9672 729 9688
rect 663 9638 679 9672
rect 713 9638 729 9672
rect 663 9622 729 9638
rect 895 9672 961 9688
rect 895 9638 911 9672
rect 945 9638 961 9672
rect 895 9622 961 9638
rect 1127 9672 1193 9688
rect 1127 9638 1143 9672
rect 1177 9638 1193 9672
rect 1127 9622 1193 9638
rect 1359 9672 1425 9688
rect 1359 9638 1375 9672
rect 1409 9638 1425 9672
rect 1359 9622 1425 9638
rect 1591 9672 1657 9688
rect 1591 9638 1607 9672
rect 1641 9638 1657 9672
rect 1591 9622 1657 9638
rect 1823 9672 1889 9688
rect 1823 9638 1839 9672
rect 1873 9638 1889 9672
rect 1823 9622 1889 9638
rect 2055 9672 2121 9688
rect 2055 9638 2071 9672
rect 2105 9638 2121 9672
rect 2055 9622 2121 9638
rect 2287 9672 2353 9688
rect 2287 9638 2303 9672
rect 2337 9638 2353 9672
rect 2287 9622 2353 9638
rect 2519 9672 2585 9688
rect 2519 9638 2535 9672
rect 2569 9638 2585 9672
rect 2519 9622 2585 9638
rect 2751 9672 2817 9688
rect 2751 9638 2767 9672
rect 2801 9638 2817 9672
rect 2751 9622 2817 9638
rect -2814 9600 -2754 9622
rect -2582 9600 -2522 9622
rect -2350 9600 -2290 9622
rect -2118 9600 -2058 9622
rect -1886 9600 -1826 9622
rect -1654 9600 -1594 9622
rect -1422 9600 -1362 9622
rect -1190 9600 -1130 9622
rect -958 9600 -898 9622
rect -726 9600 -666 9622
rect -494 9600 -434 9622
rect -262 9600 -202 9622
rect -30 9600 30 9622
rect 202 9600 262 9622
rect 434 9600 494 9622
rect 666 9600 726 9622
rect 898 9600 958 9622
rect 1130 9600 1190 9622
rect 1362 9600 1422 9622
rect 1594 9600 1654 9622
rect 1826 9600 1886 9622
rect 2058 9600 2118 9622
rect 2290 9600 2350 9622
rect 2522 9600 2582 9622
rect 2754 9600 2814 9622
rect -2814 -9622 -2754 -9600
rect -2582 -9622 -2522 -9600
rect -2350 -9622 -2290 -9600
rect -2118 -9622 -2058 -9600
rect -1886 -9622 -1826 -9600
rect -1654 -9622 -1594 -9600
rect -1422 -9622 -1362 -9600
rect -1190 -9622 -1130 -9600
rect -958 -9622 -898 -9600
rect -726 -9622 -666 -9600
rect -494 -9622 -434 -9600
rect -262 -9622 -202 -9600
rect -30 -9622 30 -9600
rect 202 -9622 262 -9600
rect 434 -9622 494 -9600
rect 666 -9622 726 -9600
rect 898 -9622 958 -9600
rect 1130 -9622 1190 -9600
rect 1362 -9622 1422 -9600
rect 1594 -9622 1654 -9600
rect 1826 -9622 1886 -9600
rect 2058 -9622 2118 -9600
rect 2290 -9622 2350 -9600
rect 2522 -9622 2582 -9600
rect 2754 -9622 2814 -9600
rect -2817 -9638 -2751 -9622
rect -2817 -9672 -2801 -9638
rect -2767 -9672 -2751 -9638
rect -2817 -9688 -2751 -9672
rect -2585 -9638 -2519 -9622
rect -2585 -9672 -2569 -9638
rect -2535 -9672 -2519 -9638
rect -2585 -9688 -2519 -9672
rect -2353 -9638 -2287 -9622
rect -2353 -9672 -2337 -9638
rect -2303 -9672 -2287 -9638
rect -2353 -9688 -2287 -9672
rect -2121 -9638 -2055 -9622
rect -2121 -9672 -2105 -9638
rect -2071 -9672 -2055 -9638
rect -2121 -9688 -2055 -9672
rect -1889 -9638 -1823 -9622
rect -1889 -9672 -1873 -9638
rect -1839 -9672 -1823 -9638
rect -1889 -9688 -1823 -9672
rect -1657 -9638 -1591 -9622
rect -1657 -9672 -1641 -9638
rect -1607 -9672 -1591 -9638
rect -1657 -9688 -1591 -9672
rect -1425 -9638 -1359 -9622
rect -1425 -9672 -1409 -9638
rect -1375 -9672 -1359 -9638
rect -1425 -9688 -1359 -9672
rect -1193 -9638 -1127 -9622
rect -1193 -9672 -1177 -9638
rect -1143 -9672 -1127 -9638
rect -1193 -9688 -1127 -9672
rect -961 -9638 -895 -9622
rect -961 -9672 -945 -9638
rect -911 -9672 -895 -9638
rect -961 -9688 -895 -9672
rect -729 -9638 -663 -9622
rect -729 -9672 -713 -9638
rect -679 -9672 -663 -9638
rect -729 -9688 -663 -9672
rect -497 -9638 -431 -9622
rect -497 -9672 -481 -9638
rect -447 -9672 -431 -9638
rect -497 -9688 -431 -9672
rect -265 -9638 -199 -9622
rect -265 -9672 -249 -9638
rect -215 -9672 -199 -9638
rect -265 -9688 -199 -9672
rect -33 -9638 33 -9622
rect -33 -9672 -17 -9638
rect 17 -9672 33 -9638
rect -33 -9688 33 -9672
rect 199 -9638 265 -9622
rect 199 -9672 215 -9638
rect 249 -9672 265 -9638
rect 199 -9688 265 -9672
rect 431 -9638 497 -9622
rect 431 -9672 447 -9638
rect 481 -9672 497 -9638
rect 431 -9688 497 -9672
rect 663 -9638 729 -9622
rect 663 -9672 679 -9638
rect 713 -9672 729 -9638
rect 663 -9688 729 -9672
rect 895 -9638 961 -9622
rect 895 -9672 911 -9638
rect 945 -9672 961 -9638
rect 895 -9688 961 -9672
rect 1127 -9638 1193 -9622
rect 1127 -9672 1143 -9638
rect 1177 -9672 1193 -9638
rect 1127 -9688 1193 -9672
rect 1359 -9638 1425 -9622
rect 1359 -9672 1375 -9638
rect 1409 -9672 1425 -9638
rect 1359 -9688 1425 -9672
rect 1591 -9638 1657 -9622
rect 1591 -9672 1607 -9638
rect 1641 -9672 1657 -9638
rect 1591 -9688 1657 -9672
rect 1823 -9638 1889 -9622
rect 1823 -9672 1839 -9638
rect 1873 -9672 1889 -9638
rect 1823 -9688 1889 -9672
rect 2055 -9638 2121 -9622
rect 2055 -9672 2071 -9638
rect 2105 -9672 2121 -9638
rect 2055 -9688 2121 -9672
rect 2287 -9638 2353 -9622
rect 2287 -9672 2303 -9638
rect 2337 -9672 2353 -9638
rect 2287 -9688 2353 -9672
rect 2519 -9638 2585 -9622
rect 2519 -9672 2535 -9638
rect 2569 -9672 2585 -9638
rect 2519 -9688 2585 -9672
rect 2751 -9638 2817 -9622
rect 2751 -9672 2767 -9638
rect 2801 -9672 2817 -9638
rect 2751 -9688 2817 -9672
<< polycont >>
rect -2801 9638 -2767 9672
rect -2569 9638 -2535 9672
rect -2337 9638 -2303 9672
rect -2105 9638 -2071 9672
rect -1873 9638 -1839 9672
rect -1641 9638 -1607 9672
rect -1409 9638 -1375 9672
rect -1177 9638 -1143 9672
rect -945 9638 -911 9672
rect -713 9638 -679 9672
rect -481 9638 -447 9672
rect -249 9638 -215 9672
rect -17 9638 17 9672
rect 215 9638 249 9672
rect 447 9638 481 9672
rect 679 9638 713 9672
rect 911 9638 945 9672
rect 1143 9638 1177 9672
rect 1375 9638 1409 9672
rect 1607 9638 1641 9672
rect 1839 9638 1873 9672
rect 2071 9638 2105 9672
rect 2303 9638 2337 9672
rect 2535 9638 2569 9672
rect 2767 9638 2801 9672
rect -2801 -9672 -2767 -9638
rect -2569 -9672 -2535 -9638
rect -2337 -9672 -2303 -9638
rect -2105 -9672 -2071 -9638
rect -1873 -9672 -1839 -9638
rect -1641 -9672 -1607 -9638
rect -1409 -9672 -1375 -9638
rect -1177 -9672 -1143 -9638
rect -945 -9672 -911 -9638
rect -713 -9672 -679 -9638
rect -481 -9672 -447 -9638
rect -249 -9672 -215 -9638
rect -17 -9672 17 -9638
rect 215 -9672 249 -9638
rect 447 -9672 481 -9638
rect 679 -9672 713 -9638
rect 911 -9672 945 -9638
rect 1143 -9672 1177 -9638
rect 1375 -9672 1409 -9638
rect 1607 -9672 1641 -9638
rect 1839 -9672 1873 -9638
rect 2071 -9672 2105 -9638
rect 2303 -9672 2337 -9638
rect 2535 -9672 2569 -9638
rect 2767 -9672 2801 -9638
<< locali >>
rect -2817 9638 -2801 9672
rect -2767 9638 -2751 9672
rect -2585 9638 -2569 9672
rect -2535 9638 -2519 9672
rect -2353 9638 -2337 9672
rect -2303 9638 -2287 9672
rect -2121 9638 -2105 9672
rect -2071 9638 -2055 9672
rect -1889 9638 -1873 9672
rect -1839 9638 -1823 9672
rect -1657 9638 -1641 9672
rect -1607 9638 -1591 9672
rect -1425 9638 -1409 9672
rect -1375 9638 -1359 9672
rect -1193 9638 -1177 9672
rect -1143 9638 -1127 9672
rect -961 9638 -945 9672
rect -911 9638 -895 9672
rect -729 9638 -713 9672
rect -679 9638 -663 9672
rect -497 9638 -481 9672
rect -447 9638 -431 9672
rect -265 9638 -249 9672
rect -215 9638 -199 9672
rect -33 9638 -17 9672
rect 17 9638 33 9672
rect 199 9638 215 9672
rect 249 9638 265 9672
rect 431 9638 447 9672
rect 481 9638 497 9672
rect 663 9638 679 9672
rect 713 9638 729 9672
rect 895 9638 911 9672
rect 945 9638 961 9672
rect 1127 9638 1143 9672
rect 1177 9638 1193 9672
rect 1359 9638 1375 9672
rect 1409 9638 1425 9672
rect 1591 9638 1607 9672
rect 1641 9638 1657 9672
rect 1823 9638 1839 9672
rect 1873 9638 1889 9672
rect 2055 9638 2071 9672
rect 2105 9638 2121 9672
rect 2287 9638 2303 9672
rect 2337 9638 2353 9672
rect 2519 9638 2535 9672
rect 2569 9638 2585 9672
rect 2751 9638 2767 9672
rect 2801 9638 2817 9672
rect -2860 9588 -2826 9604
rect -2860 -9604 -2826 -9588
rect -2742 9588 -2708 9604
rect -2742 -9604 -2708 -9588
rect -2628 9588 -2594 9604
rect -2628 -9604 -2594 -9588
rect -2510 9588 -2476 9604
rect -2510 -9604 -2476 -9588
rect -2396 9588 -2362 9604
rect -2396 -9604 -2362 -9588
rect -2278 9588 -2244 9604
rect -2278 -9604 -2244 -9588
rect -2164 9588 -2130 9604
rect -2164 -9604 -2130 -9588
rect -2046 9588 -2012 9604
rect -2046 -9604 -2012 -9588
rect -1932 9588 -1898 9604
rect -1932 -9604 -1898 -9588
rect -1814 9588 -1780 9604
rect -1814 -9604 -1780 -9588
rect -1700 9588 -1666 9604
rect -1700 -9604 -1666 -9588
rect -1582 9588 -1548 9604
rect -1582 -9604 -1548 -9588
rect -1468 9588 -1434 9604
rect -1468 -9604 -1434 -9588
rect -1350 9588 -1316 9604
rect -1350 -9604 -1316 -9588
rect -1236 9588 -1202 9604
rect -1236 -9604 -1202 -9588
rect -1118 9588 -1084 9604
rect -1118 -9604 -1084 -9588
rect -1004 9588 -970 9604
rect -1004 -9604 -970 -9588
rect -886 9588 -852 9604
rect -886 -9604 -852 -9588
rect -772 9588 -738 9604
rect -772 -9604 -738 -9588
rect -654 9588 -620 9604
rect -654 -9604 -620 -9588
rect -540 9588 -506 9604
rect -540 -9604 -506 -9588
rect -422 9588 -388 9604
rect -422 -9604 -388 -9588
rect -308 9588 -274 9604
rect -308 -9604 -274 -9588
rect -190 9588 -156 9604
rect -190 -9604 -156 -9588
rect -76 9588 -42 9604
rect -76 -9604 -42 -9588
rect 42 9588 76 9604
rect 42 -9604 76 -9588
rect 156 9588 190 9604
rect 156 -9604 190 -9588
rect 274 9588 308 9604
rect 274 -9604 308 -9588
rect 388 9588 422 9604
rect 388 -9604 422 -9588
rect 506 9588 540 9604
rect 506 -9604 540 -9588
rect 620 9588 654 9604
rect 620 -9604 654 -9588
rect 738 9588 772 9604
rect 738 -9604 772 -9588
rect 852 9588 886 9604
rect 852 -9604 886 -9588
rect 970 9588 1004 9604
rect 970 -9604 1004 -9588
rect 1084 9588 1118 9604
rect 1084 -9604 1118 -9588
rect 1202 9588 1236 9604
rect 1202 -9604 1236 -9588
rect 1316 9588 1350 9604
rect 1316 -9604 1350 -9588
rect 1434 9588 1468 9604
rect 1434 -9604 1468 -9588
rect 1548 9588 1582 9604
rect 1548 -9604 1582 -9588
rect 1666 9588 1700 9604
rect 1666 -9604 1700 -9588
rect 1780 9588 1814 9604
rect 1780 -9604 1814 -9588
rect 1898 9588 1932 9604
rect 1898 -9604 1932 -9588
rect 2012 9588 2046 9604
rect 2012 -9604 2046 -9588
rect 2130 9588 2164 9604
rect 2130 -9604 2164 -9588
rect 2244 9588 2278 9604
rect 2244 -9604 2278 -9588
rect 2362 9588 2396 9604
rect 2362 -9604 2396 -9588
rect 2476 9588 2510 9604
rect 2476 -9604 2510 -9588
rect 2594 9588 2628 9604
rect 2594 -9604 2628 -9588
rect 2708 9588 2742 9604
rect 2708 -9604 2742 -9588
rect 2826 9588 2860 9604
rect 2826 -9604 2860 -9588
rect -2817 -9672 -2801 -9638
rect -2767 -9672 -2751 -9638
rect -2585 -9672 -2569 -9638
rect -2535 -9672 -2519 -9638
rect -2353 -9672 -2337 -9638
rect -2303 -9672 -2287 -9638
rect -2121 -9672 -2105 -9638
rect -2071 -9672 -2055 -9638
rect -1889 -9672 -1873 -9638
rect -1839 -9672 -1823 -9638
rect -1657 -9672 -1641 -9638
rect -1607 -9672 -1591 -9638
rect -1425 -9672 -1409 -9638
rect -1375 -9672 -1359 -9638
rect -1193 -9672 -1177 -9638
rect -1143 -9672 -1127 -9638
rect -961 -9672 -945 -9638
rect -911 -9672 -895 -9638
rect -729 -9672 -713 -9638
rect -679 -9672 -663 -9638
rect -497 -9672 -481 -9638
rect -447 -9672 -431 -9638
rect -265 -9672 -249 -9638
rect -215 -9672 -199 -9638
rect -33 -9672 -17 -9638
rect 17 -9672 33 -9638
rect 199 -9672 215 -9638
rect 249 -9672 265 -9638
rect 431 -9672 447 -9638
rect 481 -9672 497 -9638
rect 663 -9672 679 -9638
rect 713 -9672 729 -9638
rect 895 -9672 911 -9638
rect 945 -9672 961 -9638
rect 1127 -9672 1143 -9638
rect 1177 -9672 1193 -9638
rect 1359 -9672 1375 -9638
rect 1409 -9672 1425 -9638
rect 1591 -9672 1607 -9638
rect 1641 -9672 1657 -9638
rect 1823 -9672 1839 -9638
rect 1873 -9672 1889 -9638
rect 2055 -9672 2071 -9638
rect 2105 -9672 2121 -9638
rect 2287 -9672 2303 -9638
rect 2337 -9672 2353 -9638
rect 2519 -9672 2535 -9638
rect 2569 -9672 2585 -9638
rect 2751 -9672 2767 -9638
rect 2801 -9672 2817 -9638
<< viali >>
rect -2801 9638 -2767 9672
rect -2569 9638 -2535 9672
rect -2337 9638 -2303 9672
rect -2105 9638 -2071 9672
rect -1873 9638 -1839 9672
rect -1641 9638 -1607 9672
rect -1409 9638 -1375 9672
rect -1177 9638 -1143 9672
rect -945 9638 -911 9672
rect -713 9638 -679 9672
rect -481 9638 -447 9672
rect -249 9638 -215 9672
rect -17 9638 17 9672
rect 215 9638 249 9672
rect 447 9638 481 9672
rect 679 9638 713 9672
rect 911 9638 945 9672
rect 1143 9638 1177 9672
rect 1375 9638 1409 9672
rect 1607 9638 1641 9672
rect 1839 9638 1873 9672
rect 2071 9638 2105 9672
rect 2303 9638 2337 9672
rect 2535 9638 2569 9672
rect 2767 9638 2801 9672
rect -2860 -9588 -2826 9588
rect -2742 -9588 -2708 9588
rect -2628 -9588 -2594 9588
rect -2510 -9588 -2476 9588
rect -2396 -9588 -2362 9588
rect -2278 -9588 -2244 9588
rect -2164 -9588 -2130 9588
rect -2046 -9588 -2012 9588
rect -1932 -9588 -1898 9588
rect -1814 -9588 -1780 9588
rect -1700 -9588 -1666 9588
rect -1582 -9588 -1548 9588
rect -1468 -9588 -1434 9588
rect -1350 -9588 -1316 9588
rect -1236 -9588 -1202 9588
rect -1118 -9588 -1084 9588
rect -1004 -9588 -970 9588
rect -886 -9588 -852 9588
rect -772 -9588 -738 9588
rect -654 -9588 -620 9588
rect -540 -9588 -506 9588
rect -422 -9588 -388 9588
rect -308 -9588 -274 9588
rect -190 -9588 -156 9588
rect -76 -9588 -42 9588
rect 42 -9588 76 9588
rect 156 -9588 190 9588
rect 274 -9588 308 9588
rect 388 -9588 422 9588
rect 506 -9588 540 9588
rect 620 -9588 654 9588
rect 738 -9588 772 9588
rect 852 -9588 886 9588
rect 970 -9588 1004 9588
rect 1084 -9588 1118 9588
rect 1202 -9588 1236 9588
rect 1316 -9588 1350 9588
rect 1434 -9588 1468 9588
rect 1548 -9588 1582 9588
rect 1666 -9588 1700 9588
rect 1780 -9588 1814 9588
rect 1898 -9588 1932 9588
rect 2012 -9588 2046 9588
rect 2130 -9588 2164 9588
rect 2244 -9588 2278 9588
rect 2362 -9588 2396 9588
rect 2476 -9588 2510 9588
rect 2594 -9588 2628 9588
rect 2708 -9588 2742 9588
rect 2826 -9588 2860 9588
rect -2801 -9672 -2767 -9638
rect -2569 -9672 -2535 -9638
rect -2337 -9672 -2303 -9638
rect -2105 -9672 -2071 -9638
rect -1873 -9672 -1839 -9638
rect -1641 -9672 -1607 -9638
rect -1409 -9672 -1375 -9638
rect -1177 -9672 -1143 -9638
rect -945 -9672 -911 -9638
rect -713 -9672 -679 -9638
rect -481 -9672 -447 -9638
rect -249 -9672 -215 -9638
rect -17 -9672 17 -9638
rect 215 -9672 249 -9638
rect 447 -9672 481 -9638
rect 679 -9672 713 -9638
rect 911 -9672 945 -9638
rect 1143 -9672 1177 -9638
rect 1375 -9672 1409 -9638
rect 1607 -9672 1641 -9638
rect 1839 -9672 1873 -9638
rect 2071 -9672 2105 -9638
rect 2303 -9672 2337 -9638
rect 2535 -9672 2569 -9638
rect 2767 -9672 2801 -9638
<< metal1 >>
rect -2813 9672 -2755 9678
rect -2813 9638 -2801 9672
rect -2767 9638 -2755 9672
rect -2813 9632 -2755 9638
rect -2581 9672 -2523 9678
rect -2581 9638 -2569 9672
rect -2535 9638 -2523 9672
rect -2581 9632 -2523 9638
rect -2349 9672 -2291 9678
rect -2349 9638 -2337 9672
rect -2303 9638 -2291 9672
rect -2349 9632 -2291 9638
rect -2117 9672 -2059 9678
rect -2117 9638 -2105 9672
rect -2071 9638 -2059 9672
rect -2117 9632 -2059 9638
rect -1885 9672 -1827 9678
rect -1885 9638 -1873 9672
rect -1839 9638 -1827 9672
rect -1885 9632 -1827 9638
rect -1653 9672 -1595 9678
rect -1653 9638 -1641 9672
rect -1607 9638 -1595 9672
rect -1653 9632 -1595 9638
rect -1421 9672 -1363 9678
rect -1421 9638 -1409 9672
rect -1375 9638 -1363 9672
rect -1421 9632 -1363 9638
rect -1189 9672 -1131 9678
rect -1189 9638 -1177 9672
rect -1143 9638 -1131 9672
rect -1189 9632 -1131 9638
rect -957 9672 -899 9678
rect -957 9638 -945 9672
rect -911 9638 -899 9672
rect -957 9632 -899 9638
rect -725 9672 -667 9678
rect -725 9638 -713 9672
rect -679 9638 -667 9672
rect -725 9632 -667 9638
rect -493 9672 -435 9678
rect -493 9638 -481 9672
rect -447 9638 -435 9672
rect -493 9632 -435 9638
rect -261 9672 -203 9678
rect -261 9638 -249 9672
rect -215 9638 -203 9672
rect -261 9632 -203 9638
rect -29 9672 29 9678
rect -29 9638 -17 9672
rect 17 9638 29 9672
rect -29 9632 29 9638
rect 203 9672 261 9678
rect 203 9638 215 9672
rect 249 9638 261 9672
rect 203 9632 261 9638
rect 435 9672 493 9678
rect 435 9638 447 9672
rect 481 9638 493 9672
rect 435 9632 493 9638
rect 667 9672 725 9678
rect 667 9638 679 9672
rect 713 9638 725 9672
rect 667 9632 725 9638
rect 899 9672 957 9678
rect 899 9638 911 9672
rect 945 9638 957 9672
rect 899 9632 957 9638
rect 1131 9672 1189 9678
rect 1131 9638 1143 9672
rect 1177 9638 1189 9672
rect 1131 9632 1189 9638
rect 1363 9672 1421 9678
rect 1363 9638 1375 9672
rect 1409 9638 1421 9672
rect 1363 9632 1421 9638
rect 1595 9672 1653 9678
rect 1595 9638 1607 9672
rect 1641 9638 1653 9672
rect 1595 9632 1653 9638
rect 1827 9672 1885 9678
rect 1827 9638 1839 9672
rect 1873 9638 1885 9672
rect 1827 9632 1885 9638
rect 2059 9672 2117 9678
rect 2059 9638 2071 9672
rect 2105 9638 2117 9672
rect 2059 9632 2117 9638
rect 2291 9672 2349 9678
rect 2291 9638 2303 9672
rect 2337 9638 2349 9672
rect 2291 9632 2349 9638
rect 2523 9672 2581 9678
rect 2523 9638 2535 9672
rect 2569 9638 2581 9672
rect 2523 9632 2581 9638
rect 2755 9672 2813 9678
rect 2755 9638 2767 9672
rect 2801 9638 2813 9672
rect 2755 9632 2813 9638
rect -2866 9588 -2820 9600
rect -2866 -9588 -2860 9588
rect -2826 -9588 -2820 9588
rect -2866 -9600 -2820 -9588
rect -2748 9588 -2702 9600
rect -2748 -9588 -2742 9588
rect -2708 -9588 -2702 9588
rect -2748 -9600 -2702 -9588
rect -2634 9588 -2588 9600
rect -2634 -9588 -2628 9588
rect -2594 -9588 -2588 9588
rect -2634 -9600 -2588 -9588
rect -2516 9588 -2470 9600
rect -2516 -9588 -2510 9588
rect -2476 -9588 -2470 9588
rect -2516 -9600 -2470 -9588
rect -2402 9588 -2356 9600
rect -2402 -9588 -2396 9588
rect -2362 -9588 -2356 9588
rect -2402 -9600 -2356 -9588
rect -2284 9588 -2238 9600
rect -2284 -9588 -2278 9588
rect -2244 -9588 -2238 9588
rect -2284 -9600 -2238 -9588
rect -2170 9588 -2124 9600
rect -2170 -9588 -2164 9588
rect -2130 -9588 -2124 9588
rect -2170 -9600 -2124 -9588
rect -2052 9588 -2006 9600
rect -2052 -9588 -2046 9588
rect -2012 -9588 -2006 9588
rect -2052 -9600 -2006 -9588
rect -1938 9588 -1892 9600
rect -1938 -9588 -1932 9588
rect -1898 -9588 -1892 9588
rect -1938 -9600 -1892 -9588
rect -1820 9588 -1774 9600
rect -1820 -9588 -1814 9588
rect -1780 -9588 -1774 9588
rect -1820 -9600 -1774 -9588
rect -1706 9588 -1660 9600
rect -1706 -9588 -1700 9588
rect -1666 -9588 -1660 9588
rect -1706 -9600 -1660 -9588
rect -1588 9588 -1542 9600
rect -1588 -9588 -1582 9588
rect -1548 -9588 -1542 9588
rect -1588 -9600 -1542 -9588
rect -1474 9588 -1428 9600
rect -1474 -9588 -1468 9588
rect -1434 -9588 -1428 9588
rect -1474 -9600 -1428 -9588
rect -1356 9588 -1310 9600
rect -1356 -9588 -1350 9588
rect -1316 -9588 -1310 9588
rect -1356 -9600 -1310 -9588
rect -1242 9588 -1196 9600
rect -1242 -9588 -1236 9588
rect -1202 -9588 -1196 9588
rect -1242 -9600 -1196 -9588
rect -1124 9588 -1078 9600
rect -1124 -9588 -1118 9588
rect -1084 -9588 -1078 9588
rect -1124 -9600 -1078 -9588
rect -1010 9588 -964 9600
rect -1010 -9588 -1004 9588
rect -970 -9588 -964 9588
rect -1010 -9600 -964 -9588
rect -892 9588 -846 9600
rect -892 -9588 -886 9588
rect -852 -9588 -846 9588
rect -892 -9600 -846 -9588
rect -778 9588 -732 9600
rect -778 -9588 -772 9588
rect -738 -9588 -732 9588
rect -778 -9600 -732 -9588
rect -660 9588 -614 9600
rect -660 -9588 -654 9588
rect -620 -9588 -614 9588
rect -660 -9600 -614 -9588
rect -546 9588 -500 9600
rect -546 -9588 -540 9588
rect -506 -9588 -500 9588
rect -546 -9600 -500 -9588
rect -428 9588 -382 9600
rect -428 -9588 -422 9588
rect -388 -9588 -382 9588
rect -428 -9600 -382 -9588
rect -314 9588 -268 9600
rect -314 -9588 -308 9588
rect -274 -9588 -268 9588
rect -314 -9600 -268 -9588
rect -196 9588 -150 9600
rect -196 -9588 -190 9588
rect -156 -9588 -150 9588
rect -196 -9600 -150 -9588
rect -82 9588 -36 9600
rect -82 -9588 -76 9588
rect -42 -9588 -36 9588
rect -82 -9600 -36 -9588
rect 36 9588 82 9600
rect 36 -9588 42 9588
rect 76 -9588 82 9588
rect 36 -9600 82 -9588
rect 150 9588 196 9600
rect 150 -9588 156 9588
rect 190 -9588 196 9588
rect 150 -9600 196 -9588
rect 268 9588 314 9600
rect 268 -9588 274 9588
rect 308 -9588 314 9588
rect 268 -9600 314 -9588
rect 382 9588 428 9600
rect 382 -9588 388 9588
rect 422 -9588 428 9588
rect 382 -9600 428 -9588
rect 500 9588 546 9600
rect 500 -9588 506 9588
rect 540 -9588 546 9588
rect 500 -9600 546 -9588
rect 614 9588 660 9600
rect 614 -9588 620 9588
rect 654 -9588 660 9588
rect 614 -9600 660 -9588
rect 732 9588 778 9600
rect 732 -9588 738 9588
rect 772 -9588 778 9588
rect 732 -9600 778 -9588
rect 846 9588 892 9600
rect 846 -9588 852 9588
rect 886 -9588 892 9588
rect 846 -9600 892 -9588
rect 964 9588 1010 9600
rect 964 -9588 970 9588
rect 1004 -9588 1010 9588
rect 964 -9600 1010 -9588
rect 1078 9588 1124 9600
rect 1078 -9588 1084 9588
rect 1118 -9588 1124 9588
rect 1078 -9600 1124 -9588
rect 1196 9588 1242 9600
rect 1196 -9588 1202 9588
rect 1236 -9588 1242 9588
rect 1196 -9600 1242 -9588
rect 1310 9588 1356 9600
rect 1310 -9588 1316 9588
rect 1350 -9588 1356 9588
rect 1310 -9600 1356 -9588
rect 1428 9588 1474 9600
rect 1428 -9588 1434 9588
rect 1468 -9588 1474 9588
rect 1428 -9600 1474 -9588
rect 1542 9588 1588 9600
rect 1542 -9588 1548 9588
rect 1582 -9588 1588 9588
rect 1542 -9600 1588 -9588
rect 1660 9588 1706 9600
rect 1660 -9588 1666 9588
rect 1700 -9588 1706 9588
rect 1660 -9600 1706 -9588
rect 1774 9588 1820 9600
rect 1774 -9588 1780 9588
rect 1814 -9588 1820 9588
rect 1774 -9600 1820 -9588
rect 1892 9588 1938 9600
rect 1892 -9588 1898 9588
rect 1932 -9588 1938 9588
rect 1892 -9600 1938 -9588
rect 2006 9588 2052 9600
rect 2006 -9588 2012 9588
rect 2046 -9588 2052 9588
rect 2006 -9600 2052 -9588
rect 2124 9588 2170 9600
rect 2124 -9588 2130 9588
rect 2164 -9588 2170 9588
rect 2124 -9600 2170 -9588
rect 2238 9588 2284 9600
rect 2238 -9588 2244 9588
rect 2278 -9588 2284 9588
rect 2238 -9600 2284 -9588
rect 2356 9588 2402 9600
rect 2356 -9588 2362 9588
rect 2396 -9588 2402 9588
rect 2356 -9600 2402 -9588
rect 2470 9588 2516 9600
rect 2470 -9588 2476 9588
rect 2510 -9588 2516 9588
rect 2470 -9600 2516 -9588
rect 2588 9588 2634 9600
rect 2588 -9588 2594 9588
rect 2628 -9588 2634 9588
rect 2588 -9600 2634 -9588
rect 2702 9588 2748 9600
rect 2702 -9588 2708 9588
rect 2742 -9588 2748 9588
rect 2702 -9600 2748 -9588
rect 2820 9588 2866 9600
rect 2820 -9588 2826 9588
rect 2860 -9588 2866 9588
rect 2820 -9600 2866 -9588
rect -2813 -9638 -2755 -9632
rect -2813 -9672 -2801 -9638
rect -2767 -9672 -2755 -9638
rect -2813 -9678 -2755 -9672
rect -2581 -9638 -2523 -9632
rect -2581 -9672 -2569 -9638
rect -2535 -9672 -2523 -9638
rect -2581 -9678 -2523 -9672
rect -2349 -9638 -2291 -9632
rect -2349 -9672 -2337 -9638
rect -2303 -9672 -2291 -9638
rect -2349 -9678 -2291 -9672
rect -2117 -9638 -2059 -9632
rect -2117 -9672 -2105 -9638
rect -2071 -9672 -2059 -9638
rect -2117 -9678 -2059 -9672
rect -1885 -9638 -1827 -9632
rect -1885 -9672 -1873 -9638
rect -1839 -9672 -1827 -9638
rect -1885 -9678 -1827 -9672
rect -1653 -9638 -1595 -9632
rect -1653 -9672 -1641 -9638
rect -1607 -9672 -1595 -9638
rect -1653 -9678 -1595 -9672
rect -1421 -9638 -1363 -9632
rect -1421 -9672 -1409 -9638
rect -1375 -9672 -1363 -9638
rect -1421 -9678 -1363 -9672
rect -1189 -9638 -1131 -9632
rect -1189 -9672 -1177 -9638
rect -1143 -9672 -1131 -9638
rect -1189 -9678 -1131 -9672
rect -957 -9638 -899 -9632
rect -957 -9672 -945 -9638
rect -911 -9672 -899 -9638
rect -957 -9678 -899 -9672
rect -725 -9638 -667 -9632
rect -725 -9672 -713 -9638
rect -679 -9672 -667 -9638
rect -725 -9678 -667 -9672
rect -493 -9638 -435 -9632
rect -493 -9672 -481 -9638
rect -447 -9672 -435 -9638
rect -493 -9678 -435 -9672
rect -261 -9638 -203 -9632
rect -261 -9672 -249 -9638
rect -215 -9672 -203 -9638
rect -261 -9678 -203 -9672
rect -29 -9638 29 -9632
rect -29 -9672 -17 -9638
rect 17 -9672 29 -9638
rect -29 -9678 29 -9672
rect 203 -9638 261 -9632
rect 203 -9672 215 -9638
rect 249 -9672 261 -9638
rect 203 -9678 261 -9672
rect 435 -9638 493 -9632
rect 435 -9672 447 -9638
rect 481 -9672 493 -9638
rect 435 -9678 493 -9672
rect 667 -9638 725 -9632
rect 667 -9672 679 -9638
rect 713 -9672 725 -9638
rect 667 -9678 725 -9672
rect 899 -9638 957 -9632
rect 899 -9672 911 -9638
rect 945 -9672 957 -9638
rect 899 -9678 957 -9672
rect 1131 -9638 1189 -9632
rect 1131 -9672 1143 -9638
rect 1177 -9672 1189 -9638
rect 1131 -9678 1189 -9672
rect 1363 -9638 1421 -9632
rect 1363 -9672 1375 -9638
rect 1409 -9672 1421 -9638
rect 1363 -9678 1421 -9672
rect 1595 -9638 1653 -9632
rect 1595 -9672 1607 -9638
rect 1641 -9672 1653 -9638
rect 1595 -9678 1653 -9672
rect 1827 -9638 1885 -9632
rect 1827 -9672 1839 -9638
rect 1873 -9672 1885 -9638
rect 1827 -9678 1885 -9672
rect 2059 -9638 2117 -9632
rect 2059 -9672 2071 -9638
rect 2105 -9672 2117 -9638
rect 2059 -9678 2117 -9672
rect 2291 -9638 2349 -9632
rect 2291 -9672 2303 -9638
rect 2337 -9672 2349 -9638
rect 2291 -9678 2349 -9672
rect 2523 -9638 2581 -9632
rect 2523 -9672 2535 -9638
rect 2569 -9672 2581 -9638
rect 2523 -9678 2581 -9672
rect 2755 -9638 2813 -9632
rect 2755 -9672 2767 -9638
rect 2801 -9672 2813 -9638
rect 2755 -9678 2813 -9672
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 96 l 0.3 m 1 nf 25 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
