magic
tech sky130A
magscale 1 2
timestamp 1666401131
<< error_p >>
rect -29 272 29 278
rect -29 238 -17 272
rect -29 232 29 238
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect -29 -278 29 -272
<< pwell >>
rect -226 -410 226 410
<< nmos >>
rect -30 -200 30 200
<< ndiff >>
rect -88 188 -30 200
rect -88 -188 -76 188
rect -42 -188 -30 188
rect -88 -200 -30 -188
rect 30 188 88 200
rect 30 -188 42 188
rect 76 -188 88 188
rect 30 -200 88 -188
<< ndiffc >>
rect -76 -188 -42 188
rect 42 -188 76 188
<< psubdiff >>
rect -190 340 -94 374
rect 94 340 190 374
rect -190 278 -156 340
rect 156 278 190 340
rect -190 -340 -156 -278
rect 156 -340 190 -278
rect -190 -374 -94 -340
rect 94 -374 190 -340
<< psubdiffcont >>
rect -94 340 94 374
rect -190 -278 -156 278
rect 156 -278 190 278
rect -94 -374 94 -340
<< poly >>
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -33 222 33 238
rect -30 200 30 222
rect -30 -222 30 -200
rect -33 -238 33 -222
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
<< polycont >>
rect -17 238 17 272
rect -17 -272 17 -238
<< locali >>
rect -190 340 -94 374
rect 94 340 190 374
rect -190 278 -156 340
rect 156 278 190 340
rect -33 238 -17 272
rect 17 238 33 272
rect -76 188 -42 204
rect -76 -204 -42 -188
rect 42 188 76 204
rect 42 -204 76 -188
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -190 -340 -156 -278
rect 156 -340 190 -278
rect -190 -374 -94 -340
rect 94 -374 190 -340
<< viali >>
rect -17 238 17 272
rect -76 -188 -42 188
rect 42 -188 76 188
rect -17 -272 17 -238
<< metal1 >>
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect -82 188 -36 200
rect -82 -188 -76 188
rect -42 -188 -36 188
rect -82 -200 -36 -188
rect 36 188 82 200
rect 36 -188 42 188
rect 76 -188 82 188
rect 36 -200 82 -188
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
<< properties >>
string FIXED_BBOX -173 -357 173 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
