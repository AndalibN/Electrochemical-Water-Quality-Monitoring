magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -1489 1332 -550 1360
rect -1489 1268 -634 1332
rect -570 1268 -550 1332
rect -1489 1252 -550 1268
rect -1489 1188 -634 1252
rect -570 1188 -550 1252
rect -1489 1172 -550 1188
rect -1489 1108 -634 1172
rect -570 1108 -550 1172
rect -1489 1092 -550 1108
rect -1489 1028 -634 1092
rect -570 1028 -550 1092
rect -1489 1012 -550 1028
rect -1489 948 -634 1012
rect -570 948 -550 1012
rect -1489 932 -550 948
rect -1489 868 -634 932
rect -570 868 -550 932
rect -1489 852 -550 868
rect -1489 788 -634 852
rect -570 788 -550 852
rect -1489 772 -550 788
rect -1489 708 -634 772
rect -570 708 -550 772
rect -1489 692 -550 708
rect -1489 628 -634 692
rect -570 628 -550 692
rect -1489 612 -550 628
rect -1489 548 -634 612
rect -570 548 -550 612
rect -1489 520 -550 548
rect -430 1332 469 1360
rect -430 1268 385 1332
rect 449 1268 469 1332
rect -430 1252 469 1268
rect -430 1188 385 1252
rect 449 1188 469 1252
rect -430 1172 469 1188
rect -430 1108 385 1172
rect 449 1108 469 1172
rect -430 1092 469 1108
rect -430 1028 385 1092
rect 449 1028 469 1092
rect -430 1012 469 1028
rect -430 948 385 1012
rect 449 948 469 1012
rect -430 932 469 948
rect -430 868 385 932
rect 449 868 469 932
rect -430 852 469 868
rect -430 788 385 852
rect 449 788 469 852
rect -430 772 469 788
rect -430 708 385 772
rect 449 708 469 772
rect -430 692 469 708
rect -430 628 385 692
rect 449 628 469 692
rect -430 612 469 628
rect -430 548 385 612
rect 449 548 469 612
rect -430 520 469 548
rect 549 1332 1488 1360
rect 549 1268 1404 1332
rect 1468 1268 1488 1332
rect 549 1252 1488 1268
rect 549 1188 1404 1252
rect 1468 1188 1488 1252
rect 549 1172 1488 1188
rect 549 1108 1404 1172
rect 1468 1108 1488 1172
rect 549 1092 1488 1108
rect 549 1028 1404 1092
rect 1468 1028 1488 1092
rect 549 1012 1488 1028
rect 549 948 1404 1012
rect 1468 948 1488 1012
rect 549 932 1488 948
rect 549 868 1404 932
rect 1468 868 1488 932
rect 549 852 1488 868
rect 549 788 1404 852
rect 1468 788 1488 852
rect 549 772 1488 788
rect 549 708 1404 772
rect 1468 708 1488 772
rect 549 692 1488 708
rect 549 628 1404 692
rect 1468 628 1488 692
rect 549 612 1488 628
rect 549 548 1404 612
rect 1468 548 1488 612
rect 549 520 1488 548
rect -1489 392 -550 420
rect -1489 328 -634 392
rect -570 328 -550 392
rect -1489 312 -550 328
rect -1489 248 -634 312
rect -570 248 -550 312
rect -1489 232 -550 248
rect -1489 168 -634 232
rect -570 168 -550 232
rect -1489 152 -550 168
rect -1489 88 -634 152
rect -570 88 -550 152
rect -1489 72 -550 88
rect -1489 8 -634 72
rect -570 8 -550 72
rect -1489 -8 -550 8
rect -1489 -72 -634 -8
rect -570 -72 -550 -8
rect -1489 -88 -550 -72
rect -1489 -152 -634 -88
rect -570 -152 -550 -88
rect -1489 -168 -550 -152
rect -1489 -232 -634 -168
rect -570 -232 -550 -168
rect -1489 -248 -550 -232
rect -1489 -312 -634 -248
rect -570 -312 -550 -248
rect -1489 -328 -550 -312
rect -1489 -392 -634 -328
rect -570 -392 -550 -328
rect -1489 -420 -550 -392
rect -430 392 469 420
rect -430 328 385 392
rect 449 328 469 392
rect -430 312 469 328
rect -430 248 385 312
rect 449 248 469 312
rect -430 232 469 248
rect -430 168 385 232
rect 449 168 469 232
rect -430 152 469 168
rect -430 88 385 152
rect 449 88 469 152
rect -430 72 469 88
rect -430 8 385 72
rect 449 8 469 72
rect -430 -8 469 8
rect -430 -72 385 -8
rect 449 -72 469 -8
rect -430 -88 469 -72
rect -430 -152 385 -88
rect 449 -152 469 -88
rect -430 -168 469 -152
rect -430 -232 385 -168
rect 449 -232 469 -168
rect -430 -248 469 -232
rect -430 -312 385 -248
rect 449 -312 469 -248
rect -430 -328 469 -312
rect -430 -392 385 -328
rect 449 -392 469 -328
rect -430 -420 469 -392
rect 549 392 1488 420
rect 549 328 1404 392
rect 1468 328 1488 392
rect 549 312 1488 328
rect 549 248 1404 312
rect 1468 248 1488 312
rect 549 232 1488 248
rect 549 168 1404 232
rect 1468 168 1488 232
rect 549 152 1488 168
rect 549 88 1404 152
rect 1468 88 1488 152
rect 549 72 1488 88
rect 549 8 1404 72
rect 1468 8 1488 72
rect 549 -8 1488 8
rect 549 -72 1404 -8
rect 1468 -72 1488 -8
rect 549 -88 1488 -72
rect 549 -152 1404 -88
rect 1468 -152 1488 -88
rect 549 -168 1488 -152
rect 549 -232 1404 -168
rect 1468 -232 1488 -168
rect 549 -248 1488 -232
rect 549 -312 1404 -248
rect 1468 -312 1488 -248
rect 549 -328 1488 -312
rect 549 -392 1404 -328
rect 1468 -392 1488 -328
rect 549 -420 1488 -392
rect -1489 -548 -550 -520
rect -1489 -612 -634 -548
rect -570 -612 -550 -548
rect -1489 -628 -550 -612
rect -1489 -692 -634 -628
rect -570 -692 -550 -628
rect -1489 -708 -550 -692
rect -1489 -772 -634 -708
rect -570 -772 -550 -708
rect -1489 -788 -550 -772
rect -1489 -852 -634 -788
rect -570 -852 -550 -788
rect -1489 -868 -550 -852
rect -1489 -932 -634 -868
rect -570 -932 -550 -868
rect -1489 -948 -550 -932
rect -1489 -1012 -634 -948
rect -570 -1012 -550 -948
rect -1489 -1028 -550 -1012
rect -1489 -1092 -634 -1028
rect -570 -1092 -550 -1028
rect -1489 -1108 -550 -1092
rect -1489 -1172 -634 -1108
rect -570 -1172 -550 -1108
rect -1489 -1188 -550 -1172
rect -1489 -1252 -634 -1188
rect -570 -1252 -550 -1188
rect -1489 -1268 -550 -1252
rect -1489 -1332 -634 -1268
rect -570 -1332 -550 -1268
rect -1489 -1360 -550 -1332
rect -430 -548 469 -520
rect -430 -612 385 -548
rect 449 -612 469 -548
rect -430 -628 469 -612
rect -430 -692 385 -628
rect 449 -692 469 -628
rect -430 -708 469 -692
rect -430 -772 385 -708
rect 449 -772 469 -708
rect -430 -788 469 -772
rect -430 -852 385 -788
rect 449 -852 469 -788
rect -430 -868 469 -852
rect -430 -932 385 -868
rect 449 -932 469 -868
rect -430 -948 469 -932
rect -430 -1012 385 -948
rect 449 -1012 469 -948
rect -430 -1028 469 -1012
rect -430 -1092 385 -1028
rect 449 -1092 469 -1028
rect -430 -1108 469 -1092
rect -430 -1172 385 -1108
rect 449 -1172 469 -1108
rect -430 -1188 469 -1172
rect -430 -1252 385 -1188
rect 449 -1252 469 -1188
rect -430 -1268 469 -1252
rect -430 -1332 385 -1268
rect 449 -1332 469 -1268
rect -430 -1360 469 -1332
rect 549 -548 1488 -520
rect 549 -612 1404 -548
rect 1468 -612 1488 -548
rect 549 -628 1488 -612
rect 549 -692 1404 -628
rect 1468 -692 1488 -628
rect 549 -708 1488 -692
rect 549 -772 1404 -708
rect 1468 -772 1488 -708
rect 549 -788 1488 -772
rect 549 -852 1404 -788
rect 1468 -852 1488 -788
rect 549 -868 1488 -852
rect 549 -932 1404 -868
rect 1468 -932 1488 -868
rect 549 -948 1488 -932
rect 549 -1012 1404 -948
rect 1468 -1012 1488 -948
rect 549 -1028 1488 -1012
rect 549 -1092 1404 -1028
rect 1468 -1092 1488 -1028
rect 549 -1108 1488 -1092
rect 549 -1172 1404 -1108
rect 1468 -1172 1488 -1108
rect 549 -1188 1488 -1172
rect 549 -1252 1404 -1188
rect 1468 -1252 1488 -1188
rect 549 -1268 1488 -1252
rect 549 -1332 1404 -1268
rect 1468 -1332 1488 -1268
rect 549 -1360 1488 -1332
<< via3 >>
rect -634 1268 -570 1332
rect -634 1188 -570 1252
rect -634 1108 -570 1172
rect -634 1028 -570 1092
rect -634 948 -570 1012
rect -634 868 -570 932
rect -634 788 -570 852
rect -634 708 -570 772
rect -634 628 -570 692
rect -634 548 -570 612
rect 385 1268 449 1332
rect 385 1188 449 1252
rect 385 1108 449 1172
rect 385 1028 449 1092
rect 385 948 449 1012
rect 385 868 449 932
rect 385 788 449 852
rect 385 708 449 772
rect 385 628 449 692
rect 385 548 449 612
rect 1404 1268 1468 1332
rect 1404 1188 1468 1252
rect 1404 1108 1468 1172
rect 1404 1028 1468 1092
rect 1404 948 1468 1012
rect 1404 868 1468 932
rect 1404 788 1468 852
rect 1404 708 1468 772
rect 1404 628 1468 692
rect 1404 548 1468 612
rect -634 328 -570 392
rect -634 248 -570 312
rect -634 168 -570 232
rect -634 88 -570 152
rect -634 8 -570 72
rect -634 -72 -570 -8
rect -634 -152 -570 -88
rect -634 -232 -570 -168
rect -634 -312 -570 -248
rect -634 -392 -570 -328
rect 385 328 449 392
rect 385 248 449 312
rect 385 168 449 232
rect 385 88 449 152
rect 385 8 449 72
rect 385 -72 449 -8
rect 385 -152 449 -88
rect 385 -232 449 -168
rect 385 -312 449 -248
rect 385 -392 449 -328
rect 1404 328 1468 392
rect 1404 248 1468 312
rect 1404 168 1468 232
rect 1404 88 1468 152
rect 1404 8 1468 72
rect 1404 -72 1468 -8
rect 1404 -152 1468 -88
rect 1404 -232 1468 -168
rect 1404 -312 1468 -248
rect 1404 -392 1468 -328
rect -634 -612 -570 -548
rect -634 -692 -570 -628
rect -634 -772 -570 -708
rect -634 -852 -570 -788
rect -634 -932 -570 -868
rect -634 -1012 -570 -948
rect -634 -1092 -570 -1028
rect -634 -1172 -570 -1108
rect -634 -1252 -570 -1188
rect -634 -1332 -570 -1268
rect 385 -612 449 -548
rect 385 -692 449 -628
rect 385 -772 449 -708
rect 385 -852 449 -788
rect 385 -932 449 -868
rect 385 -1012 449 -948
rect 385 -1092 449 -1028
rect 385 -1172 449 -1108
rect 385 -1252 449 -1188
rect 385 -1332 449 -1268
rect 1404 -612 1468 -548
rect 1404 -692 1468 -628
rect 1404 -772 1468 -708
rect 1404 -852 1468 -788
rect 1404 -932 1468 -868
rect 1404 -1012 1468 -948
rect 1404 -1092 1468 -1028
rect 1404 -1172 1468 -1108
rect 1404 -1252 1468 -1188
rect 1404 -1332 1468 -1268
<< mimcap >>
rect -1389 1212 -749 1260
rect -1389 668 -1341 1212
rect -797 668 -749 1212
rect -1389 620 -749 668
rect -370 1212 270 1260
rect -370 668 -322 1212
rect 222 668 270 1212
rect -370 620 270 668
rect 649 1212 1289 1260
rect 649 668 697 1212
rect 1241 668 1289 1212
rect 649 620 1289 668
rect -1389 272 -749 320
rect -1389 -272 -1341 272
rect -797 -272 -749 272
rect -1389 -320 -749 -272
rect -370 272 270 320
rect -370 -272 -322 272
rect 222 -272 270 272
rect -370 -320 270 -272
rect 649 272 1289 320
rect 649 -272 697 272
rect 1241 -272 1289 272
rect 649 -320 1289 -272
rect -1389 -668 -749 -620
rect -1389 -1212 -1341 -668
rect -797 -1212 -749 -668
rect -1389 -1260 -749 -1212
rect -370 -668 270 -620
rect -370 -1212 -322 -668
rect 222 -1212 270 -668
rect -370 -1260 270 -1212
rect 649 -668 1289 -620
rect 649 -1212 697 -668
rect 1241 -1212 1289 -668
rect 649 -1260 1289 -1212
<< mimcapcontact >>
rect -1341 668 -797 1212
rect -322 668 222 1212
rect 697 668 1241 1212
rect -1341 -272 -797 272
rect -322 -272 222 272
rect 697 -272 1241 272
rect -1341 -1212 -797 -668
rect -322 -1212 222 -668
rect 697 -1212 1241 -668
<< metal4 >>
rect -1121 1221 -1017 1410
rect -681 1332 -554 1796
rect -681 1268 -634 1332
rect -570 1268 -554 1332
rect -681 1252 -554 1268
rect -1350 1212 -788 1221
rect -1350 668 -1341 1212
rect -797 668 -788 1212
rect -1350 659 -788 668
rect -681 1188 -634 1252
rect -570 1188 -554 1252
rect -102 1221 2 1410
rect 338 1332 465 1548
rect 338 1268 385 1332
rect 449 1268 465 1332
rect 338 1252 465 1268
rect -681 1172 -554 1188
rect -681 1108 -634 1172
rect -570 1108 -554 1172
rect -681 1092 -554 1108
rect -681 1028 -634 1092
rect -570 1028 -554 1092
rect -681 1012 -554 1028
rect -681 948 -634 1012
rect -570 948 -554 1012
rect -681 932 -554 948
rect -681 868 -634 932
rect -570 868 -554 932
rect -681 852 -554 868
rect -681 788 -634 852
rect -570 788 -554 852
rect -681 772 -554 788
rect -681 708 -634 772
rect -570 708 -554 772
rect -681 692 -554 708
rect -1121 281 -1017 659
rect -681 628 -634 692
rect -570 628 -554 692
rect -331 1212 231 1221
rect -331 668 -322 1212
rect 222 668 231 1212
rect -331 659 231 668
rect 338 1188 385 1252
rect 449 1188 465 1252
rect 917 1221 1021 1410
rect 1357 1332 1484 1549
rect 1357 1268 1404 1332
rect 1468 1268 1484 1332
rect 1357 1252 1484 1268
rect 338 1172 465 1188
rect 338 1108 385 1172
rect 449 1108 465 1172
rect 338 1092 465 1108
rect 338 1028 385 1092
rect 449 1028 465 1092
rect 338 1012 465 1028
rect 338 948 385 1012
rect 449 948 465 1012
rect 338 932 465 948
rect 338 868 385 932
rect 449 868 465 932
rect 338 852 465 868
rect 338 788 385 852
rect 449 788 465 852
rect 338 772 465 788
rect 338 708 385 772
rect 449 708 465 772
rect 338 692 465 708
rect -681 612 -554 628
rect -681 548 -634 612
rect -570 548 -554 612
rect -681 532 -554 548
rect -681 408 -577 532
rect -681 392 -554 408
rect -681 328 -634 392
rect -570 328 -554 392
rect -681 312 -554 328
rect -1350 272 -788 281
rect -1350 -272 -1341 272
rect -797 -272 -788 272
rect -1350 -281 -788 -272
rect -681 248 -634 312
rect -570 248 -554 312
rect -102 281 2 659
rect 338 628 385 692
rect 449 628 465 692
rect 688 1212 1250 1221
rect 688 668 697 1212
rect 1241 668 1250 1212
rect 688 659 1250 668
rect 1357 1188 1404 1252
rect 1468 1188 1484 1252
rect 1357 1172 1484 1188
rect 1357 1108 1404 1172
rect 1468 1108 1484 1172
rect 1357 1092 1484 1108
rect 1357 1028 1404 1092
rect 1468 1028 1484 1092
rect 1357 1012 1484 1028
rect 1357 948 1404 1012
rect 1468 948 1484 1012
rect 1357 932 1484 948
rect 1357 868 1404 932
rect 1468 868 1484 932
rect 1357 852 1484 868
rect 1357 788 1404 852
rect 1468 788 1484 852
rect 1357 772 1484 788
rect 1357 708 1404 772
rect 1468 708 1484 772
rect 1357 692 1484 708
rect 338 612 465 628
rect 338 548 385 612
rect 449 548 465 612
rect 338 532 465 548
rect 338 408 442 532
rect 338 392 465 408
rect 338 328 385 392
rect 449 328 465 392
rect 338 312 465 328
rect -681 232 -554 248
rect -681 168 -634 232
rect -570 168 -554 232
rect -681 152 -554 168
rect -681 88 -634 152
rect -570 88 -554 152
rect -681 72 -554 88
rect -681 8 -634 72
rect -570 8 -554 72
rect -681 -8 -554 8
rect -681 -72 -634 -8
rect -570 -72 -554 -8
rect -681 -88 -554 -72
rect -681 -152 -634 -88
rect -570 -152 -554 -88
rect -681 -168 -554 -152
rect -681 -232 -634 -168
rect -570 -232 -554 -168
rect -681 -248 -554 -232
rect -1121 -659 -1017 -281
rect -681 -312 -634 -248
rect -570 -312 -554 -248
rect -331 272 231 281
rect -331 -272 -322 272
rect 222 -272 231 272
rect -331 -281 231 -272
rect 338 248 385 312
rect 449 248 465 312
rect 917 281 1021 659
rect 1357 628 1404 692
rect 1468 628 1484 692
rect 1357 612 1484 628
rect 1357 548 1404 612
rect 1468 548 1484 612
rect 1357 532 1484 548
rect 1357 408 1461 532
rect 1357 392 1484 408
rect 1357 328 1404 392
rect 1468 328 1484 392
rect 1357 312 1484 328
rect 338 232 465 248
rect 338 168 385 232
rect 449 168 465 232
rect 338 152 465 168
rect 338 88 385 152
rect 449 88 465 152
rect 338 72 465 88
rect 338 8 385 72
rect 449 8 465 72
rect 338 -8 465 8
rect 338 -72 385 -8
rect 449 -72 465 -8
rect 338 -88 465 -72
rect 338 -152 385 -88
rect 449 -152 465 -88
rect 338 -168 465 -152
rect 338 -232 385 -168
rect 449 -232 465 -168
rect 338 -248 465 -232
rect -681 -328 -554 -312
rect -681 -392 -634 -328
rect -570 -392 -554 -328
rect -681 -408 -554 -392
rect -681 -532 -577 -408
rect -681 -548 -554 -532
rect -681 -612 -634 -548
rect -570 -612 -554 -548
rect -681 -628 -554 -612
rect -1350 -668 -788 -659
rect -1350 -1212 -1341 -668
rect -797 -1212 -788 -668
rect -1350 -1224 -788 -1212
rect -681 -692 -634 -628
rect -570 -692 -554 -628
rect -102 -659 2 -281
rect 338 -312 385 -248
rect 449 -312 465 -248
rect 688 272 1250 281
rect 688 -272 697 272
rect 1241 -272 1250 272
rect 688 -281 1250 -272
rect 1357 248 1404 312
rect 1468 248 1484 312
rect 1357 232 1484 248
rect 1357 168 1404 232
rect 1468 168 1484 232
rect 1357 152 1484 168
rect 1357 88 1404 152
rect 1468 88 1484 152
rect 1357 72 1484 88
rect 1357 8 1404 72
rect 1468 8 1484 72
rect 1357 -8 1484 8
rect 1357 -72 1404 -8
rect 1468 -72 1484 -8
rect 1357 -88 1484 -72
rect 1357 -152 1404 -88
rect 1468 -152 1484 -88
rect 1357 -168 1484 -152
rect 1357 -232 1404 -168
rect 1468 -232 1484 -168
rect 1357 -248 1484 -232
rect 338 -328 465 -312
rect 338 -392 385 -328
rect 449 -392 465 -328
rect 338 -408 465 -392
rect 338 -532 442 -408
rect 338 -548 465 -532
rect 338 -612 385 -548
rect 449 -612 465 -548
rect 338 -628 465 -612
rect -681 -708 -554 -692
rect -681 -772 -634 -708
rect -570 -772 -554 -708
rect -681 -788 -554 -772
rect -681 -852 -634 -788
rect -570 -852 -554 -788
rect -681 -868 -554 -852
rect -681 -932 -634 -868
rect -570 -932 -554 -868
rect -681 -948 -554 -932
rect -681 -1012 -634 -948
rect -570 -1012 -554 -948
rect -681 -1028 -554 -1012
rect -681 -1092 -634 -1028
rect -570 -1092 -554 -1028
rect -681 -1108 -554 -1092
rect -681 -1172 -634 -1108
rect -570 -1172 -554 -1108
rect -681 -1188 -554 -1172
rect -681 -1252 -634 -1188
rect -570 -1252 -554 -1188
rect -331 -668 231 -659
rect -331 -1212 -322 -668
rect 222 -1212 231 -668
rect -331 -1220 231 -1212
rect 338 -692 385 -628
rect 449 -692 465 -628
rect 917 -659 1021 -281
rect 1357 -312 1404 -248
rect 1468 -312 1484 -248
rect 1357 -328 1484 -312
rect 1357 -392 1404 -328
rect 1468 -392 1484 -328
rect 1357 -408 1484 -392
rect 1357 -532 1461 -408
rect 1357 -548 1484 -532
rect 1357 -612 1404 -548
rect 1468 -612 1484 -548
rect 1357 -628 1484 -612
rect 338 -708 465 -692
rect 338 -772 385 -708
rect 449 -772 465 -708
rect 338 -788 465 -772
rect 338 -852 385 -788
rect 449 -852 465 -788
rect 338 -868 465 -852
rect 338 -932 385 -868
rect 449 -932 465 -868
rect 338 -948 465 -932
rect 338 -1012 385 -948
rect 449 -1012 465 -948
rect 338 -1028 465 -1012
rect 338 -1092 385 -1028
rect 449 -1092 465 -1028
rect 338 -1108 465 -1092
rect 338 -1172 385 -1108
rect 449 -1172 465 -1108
rect 338 -1188 465 -1172
rect -681 -1268 -554 -1252
rect -681 -1332 -634 -1268
rect -570 -1332 -554 -1268
rect -681 -1348 -554 -1332
rect 338 -1252 385 -1188
rect 449 -1252 465 -1188
rect 688 -668 1250 -659
rect 688 -1212 697 -668
rect 1241 -1212 1250 -668
rect 688 -1231 1250 -1212
rect 1357 -692 1404 -628
rect 1468 -692 1484 -628
rect 1357 -708 1484 -692
rect 1357 -772 1404 -708
rect 1468 -772 1484 -708
rect 1357 -788 1484 -772
rect 1357 -852 1404 -788
rect 1468 -852 1484 -788
rect 1357 -868 1484 -852
rect 1357 -932 1404 -868
rect 1468 -932 1484 -868
rect 1357 -948 1484 -932
rect 1357 -1012 1404 -948
rect 1468 -1012 1484 -948
rect 1357 -1028 1484 -1012
rect 1357 -1092 1404 -1028
rect 1468 -1092 1484 -1028
rect 1357 -1108 1484 -1092
rect 1357 -1172 1404 -1108
rect 1468 -1172 1484 -1108
rect 1357 -1188 1484 -1172
rect 338 -1268 465 -1252
rect 338 -1332 385 -1268
rect 449 -1332 465 -1268
rect 338 -1348 465 -1332
rect 1357 -1252 1404 -1188
rect 1468 -1252 1484 -1188
rect 1357 -1268 1484 -1252
rect 1357 -1332 1404 -1268
rect 1468 -1332 1484 -1268
rect 1357 -1348 1484 -1332
<< properties >>
string FIXED_BBOX 489 520 1329 1360
<< end >>
