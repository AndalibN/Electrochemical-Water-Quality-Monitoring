magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 1600 35 2032
rect -35 -2032 35 -1600
<< xpolyres >>
rect -35 -1600 35 1600
<< viali >>
rect -17 1978 17 2012
rect -17 1906 17 1940
rect -17 1834 17 1868
rect -17 1762 17 1796
rect -17 1690 17 1724
rect -17 1618 17 1652
rect -17 -1653 17 -1619
rect -17 -1725 17 -1691
rect -17 -1797 17 -1763
rect -17 -1869 17 -1835
rect -17 -1941 17 -1907
rect -17 -2013 17 -1979
<< metal1 >>
rect -25 2012 25 2026
rect -25 1978 -17 2012
rect 17 1978 25 2012
rect -25 1940 25 1978
rect -25 1906 -17 1940
rect 17 1906 25 1940
rect -25 1868 25 1906
rect -25 1834 -17 1868
rect 17 1834 25 1868
rect -25 1796 25 1834
rect -25 1762 -17 1796
rect 17 1762 25 1796
rect -25 1724 25 1762
rect -25 1690 -17 1724
rect 17 1690 25 1724
rect -25 1652 25 1690
rect -25 1618 -17 1652
rect 17 1618 25 1652
rect -25 1605 25 1618
rect -25 -1619 25 -1605
rect -25 -1653 -17 -1619
rect 17 -1653 25 -1619
rect -25 -1691 25 -1653
rect -25 -1725 -17 -1691
rect 17 -1725 25 -1691
rect -25 -1763 25 -1725
rect -25 -1797 -17 -1763
rect 17 -1797 25 -1763
rect -25 -1835 25 -1797
rect -25 -1869 -17 -1835
rect 17 -1869 25 -1835
rect -25 -1907 25 -1869
rect -25 -1941 -17 -1907
rect 17 -1941 25 -1907
rect -25 -1979 25 -1941
rect -25 -2013 -17 -1979
rect 17 -2013 25 -1979
rect -25 -2026 25 -2013
<< end >>
