magic
tech sky130A
timestamp 1669522153
<< end >>
