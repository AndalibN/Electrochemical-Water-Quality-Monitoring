magic
tech sky130A
magscale 1 2
timestamp 1669522153
use diffPair  sky130_fd_pr__pfet_01v8_27VBYH_0
timestamp 1669522153
transform 1 0 -2245 0 1 -321
box -1098 -872 948 778
<< end >>
