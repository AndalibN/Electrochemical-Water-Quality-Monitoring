magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -2150 2552 2149 2600
rect -2150 2488 2065 2552
rect 2129 2488 2149 2552
rect -2150 2472 2149 2488
rect -2150 2408 2065 2472
rect 2129 2408 2149 2472
rect -2150 2392 2149 2408
rect -2150 2328 2065 2392
rect 2129 2328 2149 2392
rect -2150 2312 2149 2328
rect -2150 2248 2065 2312
rect 2129 2248 2149 2312
rect -2150 2232 2149 2248
rect -2150 2168 2065 2232
rect 2129 2168 2149 2232
rect -2150 2152 2149 2168
rect -2150 2088 2065 2152
rect 2129 2088 2149 2152
rect -2150 2072 2149 2088
rect -2150 2008 2065 2072
rect 2129 2008 2149 2072
rect -2150 1992 2149 2008
rect -2150 1928 2065 1992
rect 2129 1928 2149 1992
rect -2150 1912 2149 1928
rect -2150 1848 2065 1912
rect 2129 1848 2149 1912
rect -2150 1832 2149 1848
rect -2150 1768 2065 1832
rect 2129 1768 2149 1832
rect -2150 1752 2149 1768
rect -2150 1688 2065 1752
rect 2129 1688 2149 1752
rect -2150 1672 2149 1688
rect -2150 1608 2065 1672
rect 2129 1608 2149 1672
rect -2150 1592 2149 1608
rect -2150 1528 2065 1592
rect 2129 1528 2149 1592
rect -2150 1512 2149 1528
rect -2150 1448 2065 1512
rect 2129 1448 2149 1512
rect -2150 1432 2149 1448
rect -2150 1368 2065 1432
rect 2129 1368 2149 1432
rect -2150 1352 2149 1368
rect -2150 1288 2065 1352
rect 2129 1288 2149 1352
rect -2150 1272 2149 1288
rect -2150 1208 2065 1272
rect 2129 1208 2149 1272
rect -2150 1192 2149 1208
rect -2150 1128 2065 1192
rect 2129 1128 2149 1192
rect -2150 1112 2149 1128
rect -2150 1048 2065 1112
rect 2129 1048 2149 1112
rect -2150 1032 2149 1048
rect -2150 968 2065 1032
rect 2129 968 2149 1032
rect -2150 952 2149 968
rect -2150 888 2065 952
rect 2129 888 2149 952
rect -2150 872 2149 888
rect -2150 808 2065 872
rect 2129 808 2149 872
rect -2150 792 2149 808
rect -2150 728 2065 792
rect 2129 728 2149 792
rect -2150 712 2149 728
rect -2150 648 2065 712
rect 2129 648 2149 712
rect -2150 632 2149 648
rect -2150 568 2065 632
rect 2129 568 2149 632
rect -2150 552 2149 568
rect -2150 488 2065 552
rect 2129 488 2149 552
rect -2150 472 2149 488
rect -2150 408 2065 472
rect 2129 408 2149 472
rect -2150 392 2149 408
rect -2150 328 2065 392
rect 2129 328 2149 392
rect -2150 312 2149 328
rect -2150 248 2065 312
rect 2129 248 2149 312
rect -2150 232 2149 248
rect -2150 168 2065 232
rect 2129 168 2149 232
rect -2150 152 2149 168
rect -2150 88 2065 152
rect 2129 88 2149 152
rect -2150 72 2149 88
rect -2150 8 2065 72
rect 2129 8 2149 72
rect -2150 -8 2149 8
rect -2150 -72 2065 -8
rect 2129 -72 2149 -8
rect -2150 -88 2149 -72
rect -2150 -152 2065 -88
rect 2129 -152 2149 -88
rect -2150 -168 2149 -152
rect -2150 -232 2065 -168
rect 2129 -232 2149 -168
rect -2150 -248 2149 -232
rect -2150 -312 2065 -248
rect 2129 -312 2149 -248
rect -2150 -328 2149 -312
rect -2150 -392 2065 -328
rect 2129 -392 2149 -328
rect -2150 -408 2149 -392
rect -2150 -472 2065 -408
rect 2129 -472 2149 -408
rect -2150 -488 2149 -472
rect -2150 -552 2065 -488
rect 2129 -552 2149 -488
rect -2150 -568 2149 -552
rect -2150 -632 2065 -568
rect 2129 -632 2149 -568
rect -2150 -648 2149 -632
rect -2150 -712 2065 -648
rect 2129 -712 2149 -648
rect -2150 -728 2149 -712
rect -2150 -792 2065 -728
rect 2129 -792 2149 -728
rect -2150 -808 2149 -792
rect -2150 -872 2065 -808
rect 2129 -872 2149 -808
rect -2150 -888 2149 -872
rect -2150 -952 2065 -888
rect 2129 -952 2149 -888
rect -2150 -968 2149 -952
rect -2150 -1032 2065 -968
rect 2129 -1032 2149 -968
rect -2150 -1048 2149 -1032
rect -2150 -1112 2065 -1048
rect 2129 -1112 2149 -1048
rect -2150 -1128 2149 -1112
rect -2150 -1192 2065 -1128
rect 2129 -1192 2149 -1128
rect -2150 -1208 2149 -1192
rect -2150 -1272 2065 -1208
rect 2129 -1272 2149 -1208
rect -2150 -1288 2149 -1272
rect -2150 -1352 2065 -1288
rect 2129 -1352 2149 -1288
rect -2150 -1368 2149 -1352
rect -2150 -1432 2065 -1368
rect 2129 -1432 2149 -1368
rect -2150 -1448 2149 -1432
rect -2150 -1512 2065 -1448
rect 2129 -1512 2149 -1448
rect -2150 -1528 2149 -1512
rect -2150 -1592 2065 -1528
rect 2129 -1592 2149 -1528
rect -2150 -1608 2149 -1592
rect -2150 -1672 2065 -1608
rect 2129 -1672 2149 -1608
rect -2150 -1688 2149 -1672
rect -2150 -1752 2065 -1688
rect 2129 -1752 2149 -1688
rect -2150 -1768 2149 -1752
rect -2150 -1832 2065 -1768
rect 2129 -1832 2149 -1768
rect -2150 -1848 2149 -1832
rect -2150 -1912 2065 -1848
rect 2129 -1912 2149 -1848
rect -2150 -1928 2149 -1912
rect -2150 -1992 2065 -1928
rect 2129 -1992 2149 -1928
rect -2150 -2008 2149 -1992
rect -2150 -2072 2065 -2008
rect 2129 -2072 2149 -2008
rect -2150 -2088 2149 -2072
rect -2150 -2152 2065 -2088
rect 2129 -2152 2149 -2088
rect -2150 -2168 2149 -2152
rect -2150 -2232 2065 -2168
rect 2129 -2232 2149 -2168
rect -2150 -2248 2149 -2232
rect -2150 -2312 2065 -2248
rect 2129 -2312 2149 -2248
rect -2150 -2328 2149 -2312
rect -2150 -2392 2065 -2328
rect 2129 -2392 2149 -2328
rect -2150 -2408 2149 -2392
rect -2150 -2472 2065 -2408
rect 2129 -2472 2149 -2408
rect -2150 -2488 2149 -2472
rect -2150 -2552 2065 -2488
rect 2129 -2552 2149 -2488
rect -2150 -2600 2149 -2552
<< via3 >>
rect 2065 2488 2129 2552
rect 2065 2408 2129 2472
rect 2065 2328 2129 2392
rect 2065 2248 2129 2312
rect 2065 2168 2129 2232
rect 2065 2088 2129 2152
rect 2065 2008 2129 2072
rect 2065 1928 2129 1992
rect 2065 1848 2129 1912
rect 2065 1768 2129 1832
rect 2065 1688 2129 1752
rect 2065 1608 2129 1672
rect 2065 1528 2129 1592
rect 2065 1448 2129 1512
rect 2065 1368 2129 1432
rect 2065 1288 2129 1352
rect 2065 1208 2129 1272
rect 2065 1128 2129 1192
rect 2065 1048 2129 1112
rect 2065 968 2129 1032
rect 2065 888 2129 952
rect 2065 808 2129 872
rect 2065 728 2129 792
rect 2065 648 2129 712
rect 2065 568 2129 632
rect 2065 488 2129 552
rect 2065 408 2129 472
rect 2065 328 2129 392
rect 2065 248 2129 312
rect 2065 168 2129 232
rect 2065 88 2129 152
rect 2065 8 2129 72
rect 2065 -72 2129 -8
rect 2065 -152 2129 -88
rect 2065 -232 2129 -168
rect 2065 -312 2129 -248
rect 2065 -392 2129 -328
rect 2065 -472 2129 -408
rect 2065 -552 2129 -488
rect 2065 -632 2129 -568
rect 2065 -712 2129 -648
rect 2065 -792 2129 -728
rect 2065 -872 2129 -808
rect 2065 -952 2129 -888
rect 2065 -1032 2129 -968
rect 2065 -1112 2129 -1048
rect 2065 -1192 2129 -1128
rect 2065 -1272 2129 -1208
rect 2065 -1352 2129 -1288
rect 2065 -1432 2129 -1368
rect 2065 -1512 2129 -1448
rect 2065 -1592 2129 -1528
rect 2065 -1672 2129 -1608
rect 2065 -1752 2129 -1688
rect 2065 -1832 2129 -1768
rect 2065 -1912 2129 -1848
rect 2065 -1992 2129 -1928
rect 2065 -2072 2129 -2008
rect 2065 -2152 2129 -2088
rect 2065 -2232 2129 -2168
rect 2065 -2312 2129 -2248
rect 2065 -2392 2129 -2328
rect 2065 -2472 2129 -2408
rect 2065 -2552 2129 -2488
<< mimcap >>
rect -2050 2432 1950 2500
rect -2050 -2432 -2002 2432
rect 1902 -2432 1950 2432
rect -2050 -2500 1950 -2432
<< mimcapcontact >>
rect -2002 -2432 1902 2432
<< metal4 >>
rect 2049 2552 2145 2588
rect 2049 2488 2065 2552
rect 2129 2488 2145 2552
rect 2049 2472 2145 2488
rect -2011 2432 1911 2461
rect -2011 -2432 -2002 2432
rect 1902 -2432 1911 2432
rect -2011 -2461 1911 -2432
rect 2049 2408 2065 2472
rect 2129 2408 2145 2472
rect 2049 2392 2145 2408
rect 2049 2328 2065 2392
rect 2129 2328 2145 2392
rect 2049 2312 2145 2328
rect 2049 2248 2065 2312
rect 2129 2248 2145 2312
rect 2049 2232 2145 2248
rect 2049 2168 2065 2232
rect 2129 2168 2145 2232
rect 2049 2152 2145 2168
rect 2049 2088 2065 2152
rect 2129 2088 2145 2152
rect 2049 2072 2145 2088
rect 2049 2008 2065 2072
rect 2129 2008 2145 2072
rect 2049 1992 2145 2008
rect 2049 1928 2065 1992
rect 2129 1928 2145 1992
rect 2049 1912 2145 1928
rect 2049 1848 2065 1912
rect 2129 1848 2145 1912
rect 2049 1832 2145 1848
rect 2049 1768 2065 1832
rect 2129 1768 2145 1832
rect 2049 1752 2145 1768
rect 2049 1688 2065 1752
rect 2129 1688 2145 1752
rect 2049 1672 2145 1688
rect 2049 1608 2065 1672
rect 2129 1608 2145 1672
rect 2049 1592 2145 1608
rect 2049 1528 2065 1592
rect 2129 1528 2145 1592
rect 2049 1512 2145 1528
rect 2049 1448 2065 1512
rect 2129 1448 2145 1512
rect 2049 1432 2145 1448
rect 2049 1368 2065 1432
rect 2129 1368 2145 1432
rect 2049 1352 2145 1368
rect 2049 1288 2065 1352
rect 2129 1288 2145 1352
rect 2049 1272 2145 1288
rect 2049 1208 2065 1272
rect 2129 1208 2145 1272
rect 2049 1192 2145 1208
rect 2049 1128 2065 1192
rect 2129 1128 2145 1192
rect 2049 1112 2145 1128
rect 2049 1048 2065 1112
rect 2129 1048 2145 1112
rect 2049 1032 2145 1048
rect 2049 968 2065 1032
rect 2129 968 2145 1032
rect 2049 952 2145 968
rect 2049 888 2065 952
rect 2129 888 2145 952
rect 2049 872 2145 888
rect 2049 808 2065 872
rect 2129 808 2145 872
rect 2049 792 2145 808
rect 2049 728 2065 792
rect 2129 728 2145 792
rect 2049 712 2145 728
rect 2049 648 2065 712
rect 2129 648 2145 712
rect 2049 632 2145 648
rect 2049 568 2065 632
rect 2129 568 2145 632
rect 2049 552 2145 568
rect 2049 488 2065 552
rect 2129 488 2145 552
rect 2049 472 2145 488
rect 2049 408 2065 472
rect 2129 408 2145 472
rect 2049 392 2145 408
rect 2049 328 2065 392
rect 2129 328 2145 392
rect 2049 312 2145 328
rect 2049 248 2065 312
rect 2129 248 2145 312
rect 2049 232 2145 248
rect 2049 168 2065 232
rect 2129 168 2145 232
rect 2049 152 2145 168
rect 2049 88 2065 152
rect 2129 88 2145 152
rect 2049 72 2145 88
rect 2049 8 2065 72
rect 2129 8 2145 72
rect 2049 -8 2145 8
rect 2049 -72 2065 -8
rect 2129 -72 2145 -8
rect 2049 -88 2145 -72
rect 2049 -152 2065 -88
rect 2129 -152 2145 -88
rect 2049 -168 2145 -152
rect 2049 -232 2065 -168
rect 2129 -232 2145 -168
rect 2049 -248 2145 -232
rect 2049 -312 2065 -248
rect 2129 -312 2145 -248
rect 2049 -328 2145 -312
rect 2049 -392 2065 -328
rect 2129 -392 2145 -328
rect 2049 -408 2145 -392
rect 2049 -472 2065 -408
rect 2129 -472 2145 -408
rect 2049 -488 2145 -472
rect 2049 -552 2065 -488
rect 2129 -552 2145 -488
rect 2049 -568 2145 -552
rect 2049 -632 2065 -568
rect 2129 -632 2145 -568
rect 2049 -648 2145 -632
rect 2049 -712 2065 -648
rect 2129 -712 2145 -648
rect 2049 -728 2145 -712
rect 2049 -792 2065 -728
rect 2129 -792 2145 -728
rect 2049 -808 2145 -792
rect 2049 -872 2065 -808
rect 2129 -872 2145 -808
rect 2049 -888 2145 -872
rect 2049 -952 2065 -888
rect 2129 -952 2145 -888
rect 2049 -968 2145 -952
rect 2049 -1032 2065 -968
rect 2129 -1032 2145 -968
rect 2049 -1048 2145 -1032
rect 2049 -1112 2065 -1048
rect 2129 -1112 2145 -1048
rect 2049 -1128 2145 -1112
rect 2049 -1192 2065 -1128
rect 2129 -1192 2145 -1128
rect 2049 -1208 2145 -1192
rect 2049 -1272 2065 -1208
rect 2129 -1272 2145 -1208
rect 2049 -1288 2145 -1272
rect 2049 -1352 2065 -1288
rect 2129 -1352 2145 -1288
rect 2049 -1368 2145 -1352
rect 2049 -1432 2065 -1368
rect 2129 -1432 2145 -1368
rect 2049 -1448 2145 -1432
rect 2049 -1512 2065 -1448
rect 2129 -1512 2145 -1448
rect 2049 -1528 2145 -1512
rect 2049 -1592 2065 -1528
rect 2129 -1592 2145 -1528
rect 2049 -1608 2145 -1592
rect 2049 -1672 2065 -1608
rect 2129 -1672 2145 -1608
rect 2049 -1688 2145 -1672
rect 2049 -1752 2065 -1688
rect 2129 -1752 2145 -1688
rect 2049 -1768 2145 -1752
rect 2049 -1832 2065 -1768
rect 2129 -1832 2145 -1768
rect 2049 -1848 2145 -1832
rect 2049 -1912 2065 -1848
rect 2129 -1912 2145 -1848
rect 2049 -1928 2145 -1912
rect 2049 -1992 2065 -1928
rect 2129 -1992 2145 -1928
rect 2049 -2008 2145 -1992
rect 2049 -2072 2065 -2008
rect 2129 -2072 2145 -2008
rect 2049 -2088 2145 -2072
rect 2049 -2152 2065 -2088
rect 2129 -2152 2145 -2088
rect 2049 -2168 2145 -2152
rect 2049 -2232 2065 -2168
rect 2129 -2232 2145 -2168
rect 2049 -2248 2145 -2232
rect 2049 -2312 2065 -2248
rect 2129 -2312 2145 -2248
rect 2049 -2328 2145 -2312
rect 2049 -2392 2065 -2328
rect 2129 -2392 2145 -2328
rect 2049 -2408 2145 -2392
rect 2049 -2472 2065 -2408
rect 2129 -2472 2145 -2408
rect 2049 -2488 2145 -2472
rect 2049 -2552 2065 -2488
rect 2129 -2552 2145 -2488
rect 2049 -2588 2145 -2552
<< properties >>
string FIXED_BBOX -2150 -2600 2050 2600
<< end >>
