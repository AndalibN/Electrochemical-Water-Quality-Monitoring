magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -114 -206 114 206
<< nmos >>
rect -30 -180 30 180
<< ndiff >>
rect -88 153 -30 180
rect -88 119 -76 153
rect -42 119 -30 153
rect -88 85 -30 119
rect -88 51 -76 85
rect -42 51 -30 85
rect -88 17 -30 51
rect -88 -17 -76 17
rect -42 -17 -30 17
rect -88 -51 -30 -17
rect -88 -85 -76 -51
rect -42 -85 -30 -51
rect -88 -119 -30 -85
rect -88 -153 -76 -119
rect -42 -153 -30 -119
rect -88 -180 -30 -153
rect 30 153 88 180
rect 30 119 42 153
rect 76 119 88 153
rect 30 85 88 119
rect 30 51 42 85
rect 76 51 88 85
rect 30 17 88 51
rect 30 -17 42 17
rect 76 -17 88 17
rect 30 -51 88 -17
rect 30 -85 42 -51
rect 76 -85 88 -51
rect 30 -119 88 -85
rect 30 -153 42 -119
rect 76 -153 88 -119
rect 30 -180 88 -153
<< ndiffc >>
rect -76 119 -42 153
rect -76 51 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -51
rect -76 -153 -42 -119
rect 42 119 76 153
rect 42 51 76 85
rect 42 -17 76 17
rect 42 -85 76 -51
rect 42 -153 76 -119
<< poly >>
rect -30 180 30 206
rect -30 -206 30 -180
<< locali >>
rect -76 161 -42 184
rect -76 89 -42 119
rect -76 17 -42 51
rect -76 -51 -42 -17
rect -76 -119 -42 -89
rect -76 -184 -42 -161
rect 42 161 76 184
rect 42 89 76 119
rect 42 17 76 51
rect 42 -51 76 -17
rect 42 -119 76 -89
rect 42 -184 76 -161
<< viali >>
rect -76 153 -42 161
rect -76 127 -42 153
rect -76 85 -42 89
rect -76 55 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -55
rect -76 -89 -42 -85
rect -76 -153 -42 -127
rect -76 -161 -42 -153
rect 42 153 76 161
rect 42 127 76 153
rect 42 85 76 89
rect 42 55 76 85
rect 42 -17 76 17
rect 42 -85 76 -55
rect 42 -89 76 -85
rect 42 -153 76 -127
rect 42 -161 76 -153
<< metal1 >>
rect -82 161 -36 180
rect -82 127 -76 161
rect -42 127 -36 161
rect -82 89 -36 127
rect -82 55 -76 89
rect -42 55 -36 89
rect -82 17 -36 55
rect -82 -17 -76 17
rect -42 -17 -36 17
rect -82 -55 -36 -17
rect -82 -89 -76 -55
rect -42 -89 -36 -55
rect -82 -127 -36 -89
rect -82 -161 -76 -127
rect -42 -161 -36 -127
rect -82 -180 -36 -161
rect 36 161 82 180
rect 36 127 42 161
rect 76 127 82 161
rect 36 89 82 127
rect 36 55 42 89
rect 76 55 82 89
rect 36 17 82 55
rect 36 -17 42 17
rect 76 -17 82 17
rect 36 -55 82 -17
rect 36 -89 42 -55
rect 76 -89 82 -55
rect 36 -127 82 -89
rect 36 -161 42 -127
rect 76 -161 82 -127
rect 36 -180 82 -161
<< end >>
