magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -1084 -157 1084 95
<< nmos >>
rect -1000 -131 1000 69
<< ndiff >>
rect -1058 54 -1000 69
rect -1058 20 -1046 54
rect -1012 20 -1000 54
rect -1058 -14 -1000 20
rect -1058 -48 -1046 -14
rect -1012 -48 -1000 -14
rect -1058 -82 -1000 -48
rect -1058 -116 -1046 -82
rect -1012 -116 -1000 -82
rect -1058 -131 -1000 -116
rect 1000 54 1058 69
rect 1000 20 1012 54
rect 1046 20 1058 54
rect 1000 -14 1058 20
rect 1000 -48 1012 -14
rect 1046 -48 1058 -14
rect 1000 -82 1058 -48
rect 1000 -116 1012 -82
rect 1046 -116 1058 -82
rect 1000 -131 1058 -116
<< ndiffc >>
rect -1046 20 -1012 54
rect -1046 -48 -1012 -14
rect -1046 -116 -1012 -82
rect 1012 20 1046 54
rect 1012 -48 1046 -14
rect 1012 -116 1046 -82
<< poly >>
rect -1000 141 1000 157
rect -1000 107 -969 141
rect -935 107 -901 141
rect -867 107 -833 141
rect -799 107 -765 141
rect -731 107 -697 141
rect -663 107 -629 141
rect -595 107 -561 141
rect -527 107 -493 141
rect -459 107 -425 141
rect -391 107 -357 141
rect -323 107 -289 141
rect -255 107 -221 141
rect -187 107 -153 141
rect -119 107 -85 141
rect -51 107 -17 141
rect 17 107 51 141
rect 85 107 119 141
rect 153 107 187 141
rect 221 107 255 141
rect 289 107 323 141
rect 357 107 391 141
rect 425 107 459 141
rect 493 107 527 141
rect 561 107 595 141
rect 629 107 663 141
rect 697 107 731 141
rect 765 107 799 141
rect 833 107 867 141
rect 901 107 935 141
rect 969 107 1000 141
rect -1000 69 1000 107
rect -1000 -157 1000 -131
<< polycont >>
rect -969 107 -935 141
rect -901 107 -867 141
rect -833 107 -799 141
rect -765 107 -731 141
rect -697 107 -663 141
rect -629 107 -595 141
rect -561 107 -527 141
rect -493 107 -459 141
rect -425 107 -391 141
rect -357 107 -323 141
rect -289 107 -255 141
rect -221 107 -187 141
rect -153 107 -119 141
rect -85 107 -51 141
rect -17 107 17 141
rect 51 107 85 141
rect 119 107 153 141
rect 187 107 221 141
rect 255 107 289 141
rect 323 107 357 141
rect 391 107 425 141
rect 459 107 493 141
rect 527 107 561 141
rect 595 107 629 141
rect 663 107 697 141
rect 731 107 765 141
rect 799 107 833 141
rect 867 107 901 141
rect 935 107 969 141
<< locali >>
rect -1000 107 -969 141
rect -919 107 -901 141
rect -847 107 -833 141
rect -775 107 -765 141
rect -703 107 -697 141
rect -631 107 -629 141
rect -595 107 -593 141
rect -527 107 -521 141
rect -459 107 -449 141
rect -391 107 -377 141
rect -323 107 -305 141
rect -255 107 -233 141
rect -187 107 -161 141
rect -119 107 -89 141
rect -51 107 -17 141
rect 17 107 51 141
rect 89 107 119 141
rect 161 107 187 141
rect 233 107 255 141
rect 305 107 323 141
rect 377 107 391 141
rect 449 107 459 141
rect 521 107 527 141
rect 593 107 595 141
rect 629 107 631 141
rect 697 107 703 141
rect 765 107 775 141
rect 833 107 847 141
rect 901 107 919 141
rect 969 107 1000 141
rect -1046 54 -1012 73
rect -1046 -14 -1012 -12
rect -1046 -50 -1012 -48
rect -1046 -135 -1012 -116
rect 1012 54 1046 73
rect 1012 -14 1046 -12
rect 1012 -50 1046 -48
rect 1012 -135 1046 -116
<< viali >>
rect -953 107 -935 141
rect -935 107 -919 141
rect -881 107 -867 141
rect -867 107 -847 141
rect -809 107 -799 141
rect -799 107 -775 141
rect -737 107 -731 141
rect -731 107 -703 141
rect -665 107 -663 141
rect -663 107 -631 141
rect -593 107 -561 141
rect -561 107 -559 141
rect -521 107 -493 141
rect -493 107 -487 141
rect -449 107 -425 141
rect -425 107 -415 141
rect -377 107 -357 141
rect -357 107 -343 141
rect -305 107 -289 141
rect -289 107 -271 141
rect -233 107 -221 141
rect -221 107 -199 141
rect -161 107 -153 141
rect -153 107 -127 141
rect -89 107 -85 141
rect -85 107 -55 141
rect -17 107 17 141
rect 55 107 85 141
rect 85 107 89 141
rect 127 107 153 141
rect 153 107 161 141
rect 199 107 221 141
rect 221 107 233 141
rect 271 107 289 141
rect 289 107 305 141
rect 343 107 357 141
rect 357 107 377 141
rect 415 107 425 141
rect 425 107 449 141
rect 487 107 493 141
rect 493 107 521 141
rect 559 107 561 141
rect 561 107 593 141
rect 631 107 663 141
rect 663 107 665 141
rect 703 107 731 141
rect 731 107 737 141
rect 775 107 799 141
rect 799 107 809 141
rect 847 107 867 141
rect 867 107 881 141
rect 919 107 935 141
rect 935 107 953 141
rect -1046 20 -1012 22
rect -1046 -12 -1012 20
rect -1046 -82 -1012 -50
rect -1046 -84 -1012 -82
rect 1012 20 1046 22
rect 1012 -12 1046 20
rect 1012 -82 1046 -50
rect 1012 -84 1046 -82
<< metal1 >>
rect -996 141 996 147
rect -996 107 -953 141
rect -919 107 -881 141
rect -847 107 -809 141
rect -775 107 -737 141
rect -703 107 -665 141
rect -631 107 -593 141
rect -559 107 -521 141
rect -487 107 -449 141
rect -415 107 -377 141
rect -343 107 -305 141
rect -271 107 -233 141
rect -199 107 -161 141
rect -127 107 -89 141
rect -55 107 -17 141
rect 17 107 55 141
rect 89 107 127 141
rect 161 107 199 141
rect 233 107 271 141
rect 305 107 343 141
rect 377 107 415 141
rect 449 107 487 141
rect 521 107 559 141
rect 593 107 631 141
rect 665 107 703 141
rect 737 107 775 141
rect 809 107 847 141
rect 881 107 919 141
rect 953 107 996 141
rect -996 101 996 107
rect -1052 22 -1006 69
rect -1052 -12 -1046 22
rect -1012 -12 -1006 22
rect -1052 -50 -1006 -12
rect -1052 -84 -1046 -50
rect -1012 -84 -1006 -50
rect -1052 -131 -1006 -84
rect 1006 22 1052 69
rect 1006 -12 1012 22
rect 1046 -12 1052 22
rect 1006 -50 1052 -12
rect 1006 -84 1012 -50
rect 1046 -84 1052 -50
rect 1006 -131 1052 -84
<< end >>
