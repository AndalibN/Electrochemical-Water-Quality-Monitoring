magic
tech sky130A
magscale 1 2
timestamp 1667444884
<< error_s >>
rect 468 6497 503 6531
rect 469 6478 503 6497
rect 488 583 503 6478
rect 522 6444 557 6478
rect 522 583 556 6444
rect 4841 4526 4876 4560
rect 4842 4507 4876 4526
rect 2285 3556 2320 3590
rect 2286 3537 2320 3556
rect 1008 2825 1042 2879
rect 1600 2861 1634 2879
rect 522 549 537 583
rect 1027 530 1042 2825
rect 1061 2791 1096 2825
rect 1061 530 1095 2791
rect 1061 496 1076 530
rect 1564 477 1634 2861
rect 1564 441 1617 477
rect 2305 424 2320 3537
rect 2339 3503 2374 3537
rect 3024 3503 3059 3537
rect 2339 424 2373 3503
rect 3025 3484 3059 3503
rect 2339 390 2354 424
rect 3044 371 3059 3484
rect 3078 3450 3113 3484
rect 3563 3450 3598 3484
rect 4156 3467 4190 3485
rect 3078 371 3112 3450
rect 3564 3431 3598 3450
rect 3078 337 3093 371
rect 3583 318 3598 3431
rect 3617 3397 3652 3431
rect 3617 318 3651 3397
rect 3617 284 3632 318
rect 4120 265 4190 3467
rect 4120 229 4173 265
rect 4861 212 4876 4507
rect 4895 4473 4930 4507
rect 5580 4473 5615 4507
rect 4895 212 4929 4473
rect 5581 4454 5615 4473
rect 4895 178 4910 212
rect 5600 159 5615 4454
rect 5634 4420 5669 4454
rect 6319 4420 6354 4454
rect 5634 159 5668 4420
rect 6320 4401 6354 4420
rect 5634 125 5649 159
rect 6339 106 6354 4401
rect 6373 4367 6408 4401
rect 6373 106 6407 4367
rect 7059 2348 7093 2402
rect 6373 72 6388 106
rect 7078 53 7093 2348
rect 7112 2314 7147 2348
rect 7112 53 7146 2314
rect 7112 19 7127 53
rect 7617 0 7632 2348
rect 7651 0 7685 2402
rect 7651 -34 7666 0
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
use sky130_fd_pr__cap_mim_m3_1_WYFAV5  XC1
timestamp 1666963525
transform 1 0 8557 0 1 211
box -350 -300 349 300
use sky130_fd_pr__cap_mim_m3_1_WYFAV5  XC2
timestamp 1666963525
transform 1 0 9795 0 1 158
box -350 -300 349 300
use sky130_fd_pr__nfet_01v8_U7E5KL  XM1
timestamp 1666963525
transform 1 0 243 0 1 3557
box -296 -3010 296 3010
use sky130_fd_pr__nfet_01v8_U7E5KL  XM2
timestamp 1666963525
transform 1 0 782 0 1 3504
box -296 -3010 296 3010
use sky130_fd_pr__nfet_01v8_6WXQK8  XM3
timestamp 1666877501
transform 1 0 1321 0 1 1651
box -296 -1210 296 1210
use sky130_fd_pr__pfet_01v8_9QH3CS  XM4
timestamp 1666963525
transform 1 0 1960 0 1 2007
box -396 -1619 396 1619
use sky130_fd_pr__pfet_01v8_9QH3CS  XM5
timestamp 1666963525
transform 1 0 2699 0 1 1954
box -396 -1619 396 1619
use sky130_fd_pr__pfet_01v8_GGN3CJ  XM6
timestamp 1666963525
transform 1 0 3338 0 1 1901
box -296 -1619 296 1619
use sky130_fd_pr__pfet_01v8_GGN3CJ  XM7
timestamp 1666963525
transform 1 0 3877 0 1 1848
box -296 -1619 296 1619
use sky130_fd_pr__nfet_01v8_L9BG78  XM8
timestamp 1666963525
transform 1 0 4516 0 1 2386
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM9
timestamp 1666963525
transform 1 0 5255 0 1 2333
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM10
timestamp 1666963525
transform 1 0 5994 0 1 2280
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM11
timestamp 1666963525
transform 1 0 6733 0 1 2227
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_U7E5KL  XM12
timestamp 1666963525
transform 1 0 7911 0 1 2921
box -296 -3010 296 3010
use sky130_fd_pr__pfet_01v8_3HPSVM  XM13
timestamp 1666963525
transform 1 0 9149 0 1 777
box -296 -919 296 919
use sky130_fd_pr__nfet_01v8_6WXQK8  XMB1
timestamp 1666877501
transform 1 0 7372 0 1 1174
box -296 -1210 296 1210
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 Vout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Vinp
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vinm
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VB1
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VB2
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VB3
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 VDD
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 GND
port 7 nsew
<< end >>
