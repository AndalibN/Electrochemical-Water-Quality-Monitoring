magic
tech sky130A
magscale 1 2
timestamp 1666801420
<< error_p >>
rect -32 7623 32 7629
rect -32 7589 -20 7623
rect -32 7583 32 7589
rect -32 3901 32 3907
rect -32 3867 -20 3901
rect -32 3861 32 3867
rect -32 3793 32 3799
rect -32 3759 -20 3793
rect -32 3753 32 3759
rect -32 71 32 77
rect -32 37 -20 71
rect -32 31 32 37
rect -32 -37 32 -31
rect -32 -71 -20 -37
rect -32 -77 32 -71
rect -32 -3759 32 -3753
rect -32 -3793 -20 -3759
rect -32 -3799 32 -3793
rect -32 -3867 32 -3861
rect -32 -3901 -20 -3867
rect -32 -3907 32 -3901
rect -32 -7589 32 -7583
rect -32 -7623 -20 -7589
rect -32 -7629 32 -7623
<< pwell >>
rect -232 -7761 232 7761
<< nmos >>
rect -36 3939 36 7551
rect -36 109 36 3721
rect -36 -3721 36 -109
rect -36 -7551 36 -3939
<< ndiff >>
rect -94 7539 -36 7551
rect -94 3951 -82 7539
rect -48 3951 -36 7539
rect -94 3939 -36 3951
rect 36 7539 94 7551
rect 36 3951 48 7539
rect 82 3951 94 7539
rect 36 3939 94 3951
rect -94 3709 -36 3721
rect -94 121 -82 3709
rect -48 121 -36 3709
rect -94 109 -36 121
rect 36 3709 94 3721
rect 36 121 48 3709
rect 82 121 94 3709
rect 36 109 94 121
rect -94 -121 -36 -109
rect -94 -3709 -82 -121
rect -48 -3709 -36 -121
rect -94 -3721 -36 -3709
rect 36 -121 94 -109
rect 36 -3709 48 -121
rect 82 -3709 94 -121
rect 36 -3721 94 -3709
rect -94 -3951 -36 -3939
rect -94 -7539 -82 -3951
rect -48 -7539 -36 -3951
rect -94 -7551 -36 -7539
rect 36 -3951 94 -3939
rect 36 -7539 48 -3951
rect 82 -7539 94 -3951
rect 36 -7551 94 -7539
<< ndiffc >>
rect -82 3951 -48 7539
rect 48 3951 82 7539
rect -82 121 -48 3709
rect 48 121 82 3709
rect -82 -3709 -48 -121
rect 48 -3709 82 -121
rect -82 -7539 -48 -3951
rect 48 -7539 82 -3951
<< psubdiff >>
rect -196 7691 -100 7725
rect 100 7691 196 7725
rect -196 7629 -162 7691
rect 162 7629 196 7691
rect -196 -7691 -162 -7629
rect 162 -7691 196 -7629
rect -196 -7725 -100 -7691
rect 100 -7725 196 -7691
<< psubdiffcont >>
rect -100 7691 100 7725
rect -196 -7629 -162 7629
rect 162 -7629 196 7629
rect -100 -7725 100 -7691
<< poly >>
rect -36 7623 36 7639
rect -36 7589 -20 7623
rect 20 7589 36 7623
rect -36 7551 36 7589
rect -36 3901 36 3939
rect -36 3867 -20 3901
rect 20 3867 36 3901
rect -36 3851 36 3867
rect -36 3793 36 3809
rect -36 3759 -20 3793
rect 20 3759 36 3793
rect -36 3721 36 3759
rect -36 71 36 109
rect -36 37 -20 71
rect 20 37 36 71
rect -36 21 36 37
rect -36 -37 36 -21
rect -36 -71 -20 -37
rect 20 -71 36 -37
rect -36 -109 36 -71
rect -36 -3759 36 -3721
rect -36 -3793 -20 -3759
rect 20 -3793 36 -3759
rect -36 -3809 36 -3793
rect -36 -3867 36 -3851
rect -36 -3901 -20 -3867
rect 20 -3901 36 -3867
rect -36 -3939 36 -3901
rect -36 -7589 36 -7551
rect -36 -7623 -20 -7589
rect 20 -7623 36 -7589
rect -36 -7639 36 -7623
<< polycont >>
rect -20 7589 20 7623
rect -20 3867 20 3901
rect -20 3759 20 3793
rect -20 37 20 71
rect -20 -71 20 -37
rect -20 -3793 20 -3759
rect -20 -3901 20 -3867
rect -20 -7623 20 -7589
<< locali >>
rect -196 7691 -100 7725
rect 100 7691 196 7725
rect -196 7629 -162 7691
rect 162 7629 196 7691
rect -36 7589 -20 7623
rect 20 7589 36 7623
rect -82 7539 -48 7555
rect -82 3935 -48 3951
rect 48 7539 82 7555
rect 48 3935 82 3951
rect -36 3867 -20 3901
rect 20 3867 36 3901
rect -36 3759 -20 3793
rect 20 3759 36 3793
rect -82 3709 -48 3725
rect -82 105 -48 121
rect 48 3709 82 3725
rect 48 105 82 121
rect -36 37 -20 71
rect 20 37 36 71
rect -36 -71 -20 -37
rect 20 -71 36 -37
rect -82 -121 -48 -105
rect -82 -3725 -48 -3709
rect 48 -121 82 -105
rect 48 -3725 82 -3709
rect -36 -3793 -20 -3759
rect 20 -3793 36 -3759
rect -36 -3901 -20 -3867
rect 20 -3901 36 -3867
rect -82 -3951 -48 -3935
rect -82 -7555 -48 -7539
rect 48 -3951 82 -3935
rect 48 -7555 82 -7539
rect -36 -7623 -20 -7589
rect 20 -7623 36 -7589
rect -196 -7691 -162 -7629
rect 162 -7691 196 -7629
rect -196 -7725 -100 -7691
rect 100 -7725 196 -7691
<< viali >>
rect -20 7589 20 7623
rect -82 3951 -48 7539
rect 48 3951 82 7539
rect -20 3867 20 3901
rect -20 3759 20 3793
rect -82 121 -48 3709
rect 48 121 82 3709
rect -20 37 20 71
rect -20 -71 20 -37
rect -82 -3709 -48 -121
rect 48 -3709 82 -121
rect -20 -3793 20 -3759
rect -20 -3901 20 -3867
rect -82 -7539 -48 -3951
rect 48 -7539 82 -3951
rect -20 -7623 20 -7589
<< metal1 >>
rect -32 7623 32 7629
rect -32 7589 -20 7623
rect 20 7589 32 7623
rect -32 7583 32 7589
rect -88 7539 -42 7551
rect -88 3951 -82 7539
rect -48 3951 -42 7539
rect -88 3939 -42 3951
rect 42 7539 88 7551
rect 42 3951 48 7539
rect 82 3951 88 7539
rect 42 3939 88 3951
rect -32 3901 32 3907
rect -32 3867 -20 3901
rect 20 3867 32 3901
rect -32 3861 32 3867
rect -32 3793 32 3799
rect -32 3759 -20 3793
rect 20 3759 32 3793
rect -32 3753 32 3759
rect -88 3709 -42 3721
rect -88 121 -82 3709
rect -48 121 -42 3709
rect -88 109 -42 121
rect 42 3709 88 3721
rect 42 121 48 3709
rect 82 121 88 3709
rect 42 109 88 121
rect -32 71 32 77
rect -32 37 -20 71
rect 20 37 32 71
rect -32 31 32 37
rect -32 -37 32 -31
rect -32 -71 -20 -37
rect 20 -71 32 -37
rect -32 -77 32 -71
rect -88 -121 -42 -109
rect -88 -3709 -82 -121
rect -48 -3709 -42 -121
rect -88 -3721 -42 -3709
rect 42 -121 88 -109
rect 42 -3709 48 -121
rect 82 -3709 88 -121
rect 42 -3721 88 -3709
rect -32 -3759 32 -3753
rect -32 -3793 -20 -3759
rect 20 -3793 32 -3759
rect -32 -3799 32 -3793
rect -32 -3867 32 -3861
rect -32 -3901 -20 -3867
rect 20 -3901 32 -3867
rect -32 -3907 32 -3901
rect -88 -3951 -42 -3939
rect -88 -7539 -82 -3951
rect -48 -7539 -42 -3951
rect -88 -7551 -42 -7539
rect 42 -3951 88 -3939
rect 42 -7539 48 -3951
rect 82 -7539 88 -3951
rect 42 -7551 88 -7539
rect -32 -7589 32 -7583
rect -32 -7623 -20 -7589
rect 20 -7623 32 -7589
rect -32 -7629 32 -7623
<< properties >>
string FIXED_BBOX -179 -7708 179 7708
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 18.055 l 0.361 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
