magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 70 35 502
rect -35 -502 35 -70
<< xpolyres >>
rect -35 -70 35 70
<< viali >>
rect -17 448 17 482
rect -17 376 17 410
rect -17 304 17 338
rect -17 232 17 266
rect -17 160 17 194
rect -17 88 17 122
rect -17 -123 17 -89
rect -17 -195 17 -161
rect -17 -267 17 -233
rect -17 -339 17 -305
rect -17 -411 17 -377
rect -17 -483 17 -449
<< metal1 >>
rect -25 482 25 496
rect -25 448 -17 482
rect 17 448 25 482
rect -25 410 25 448
rect -25 376 -17 410
rect 17 376 25 410
rect -25 338 25 376
rect -25 304 -17 338
rect 17 304 25 338
rect -25 266 25 304
rect -25 232 -17 266
rect 17 232 25 266
rect -25 194 25 232
rect -25 160 -17 194
rect 17 160 25 194
rect -25 122 25 160
rect -25 88 -17 122
rect 17 88 25 122
rect -25 75 25 88
rect -25 -89 25 -75
rect -25 -123 -17 -89
rect 17 -123 25 -89
rect -25 -161 25 -123
rect -25 -195 -17 -161
rect 17 -195 25 -161
rect -25 -233 25 -195
rect -25 -267 -17 -233
rect 17 -267 25 -233
rect -25 -305 25 -267
rect -25 -339 -17 -305
rect 17 -339 25 -305
rect -25 -377 25 -339
rect -25 -411 -17 -377
rect 17 -411 25 -377
rect -25 -449 25 -411
rect -25 -483 -17 -449
rect 17 -483 25 -449
rect -25 -496 25 -483
<< end >>
