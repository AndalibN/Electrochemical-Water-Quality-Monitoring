magic
tech sky130A
timestamp 1668226541
<< nwell >>
rect -62 -151 62 151
<< pmos >>
rect -15 -120 15 120
<< pdiff >>
rect -44 114 -15 120
rect -44 -114 -38 114
rect -21 -114 -15 114
rect -44 -120 -15 -114
rect 15 114 44 120
rect 15 -114 21 114
rect 38 -114 44 114
rect 15 -120 44 -114
<< pdiffc >>
rect -38 -114 -21 114
rect 21 -114 38 114
<< poly >>
rect -15 120 15 133
rect -15 -133 15 -120
<< locali >>
rect -38 114 -21 122
rect -38 -122 -21 -114
rect 21 114 38 122
rect 21 -122 38 -114
<< viali >>
rect -38 -114 -21 114
rect 21 -114 38 114
<< metal1 >>
rect -41 114 -18 120
rect -41 -114 -38 114
rect -21 -114 -18 114
rect -41 -120 -18 -114
rect 18 114 41 120
rect 18 -114 21 114
rect 38 -114 41 114
rect 18 -120 41 -114
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.4 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
