magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 641 29 647
rect -29 607 -17 641
rect -29 601 29 607
<< pwell >>
rect -114 -657 114 595
<< nmos >>
rect -30 -631 30 569
<< ndiff >>
rect -88 530 -30 569
rect -88 496 -76 530
rect -42 496 -30 530
rect -88 462 -30 496
rect -88 428 -76 462
rect -42 428 -30 462
rect -88 394 -30 428
rect -88 360 -76 394
rect -42 360 -30 394
rect -88 326 -30 360
rect -88 292 -76 326
rect -42 292 -30 326
rect -88 258 -30 292
rect -88 224 -76 258
rect -42 224 -30 258
rect -88 190 -30 224
rect -88 156 -76 190
rect -42 156 -30 190
rect -88 122 -30 156
rect -88 88 -76 122
rect -42 88 -30 122
rect -88 54 -30 88
rect -88 20 -76 54
rect -42 20 -30 54
rect -88 -14 -30 20
rect -88 -48 -76 -14
rect -42 -48 -30 -14
rect -88 -82 -30 -48
rect -88 -116 -76 -82
rect -42 -116 -30 -82
rect -88 -150 -30 -116
rect -88 -184 -76 -150
rect -42 -184 -30 -150
rect -88 -218 -30 -184
rect -88 -252 -76 -218
rect -42 -252 -30 -218
rect -88 -286 -30 -252
rect -88 -320 -76 -286
rect -42 -320 -30 -286
rect -88 -354 -30 -320
rect -88 -388 -76 -354
rect -42 -388 -30 -354
rect -88 -422 -30 -388
rect -88 -456 -76 -422
rect -42 -456 -30 -422
rect -88 -490 -30 -456
rect -88 -524 -76 -490
rect -42 -524 -30 -490
rect -88 -558 -30 -524
rect -88 -592 -76 -558
rect -42 -592 -30 -558
rect -88 -631 -30 -592
rect 30 530 88 569
rect 30 496 42 530
rect 76 496 88 530
rect 30 462 88 496
rect 30 428 42 462
rect 76 428 88 462
rect 30 394 88 428
rect 30 360 42 394
rect 76 360 88 394
rect 30 326 88 360
rect 30 292 42 326
rect 76 292 88 326
rect 30 258 88 292
rect 30 224 42 258
rect 76 224 88 258
rect 30 190 88 224
rect 30 156 42 190
rect 76 156 88 190
rect 30 122 88 156
rect 30 88 42 122
rect 76 88 88 122
rect 30 54 88 88
rect 30 20 42 54
rect 76 20 88 54
rect 30 -14 88 20
rect 30 -48 42 -14
rect 76 -48 88 -14
rect 30 -82 88 -48
rect 30 -116 42 -82
rect 76 -116 88 -82
rect 30 -150 88 -116
rect 30 -184 42 -150
rect 76 -184 88 -150
rect 30 -218 88 -184
rect 30 -252 42 -218
rect 76 -252 88 -218
rect 30 -286 88 -252
rect 30 -320 42 -286
rect 76 -320 88 -286
rect 30 -354 88 -320
rect 30 -388 42 -354
rect 76 -388 88 -354
rect 30 -422 88 -388
rect 30 -456 42 -422
rect 76 -456 88 -422
rect 30 -490 88 -456
rect 30 -524 42 -490
rect 76 -524 88 -490
rect 30 -558 88 -524
rect 30 -592 42 -558
rect 76 -592 88 -558
rect 30 -631 88 -592
<< ndiffc >>
rect -76 496 -42 530
rect -76 428 -42 462
rect -76 360 -42 394
rect -76 292 -42 326
rect -76 224 -42 258
rect -76 156 -42 190
rect -76 88 -42 122
rect -76 20 -42 54
rect -76 -48 -42 -14
rect -76 -116 -42 -82
rect -76 -184 -42 -150
rect -76 -252 -42 -218
rect -76 -320 -42 -286
rect -76 -388 -42 -354
rect -76 -456 -42 -422
rect -76 -524 -42 -490
rect -76 -592 -42 -558
rect 42 496 76 530
rect 42 428 76 462
rect 42 360 76 394
rect 42 292 76 326
rect 42 224 76 258
rect 42 156 76 190
rect 42 88 76 122
rect 42 20 76 54
rect 42 -48 76 -14
rect 42 -116 76 -82
rect 42 -184 76 -150
rect 42 -252 76 -218
rect 42 -320 76 -286
rect 42 -388 76 -354
rect 42 -456 76 -422
rect 42 -524 76 -490
rect 42 -592 76 -558
<< poly >>
rect -33 641 33 657
rect -33 607 -17 641
rect 17 607 33 641
rect -33 591 33 607
rect -30 569 30 591
rect -30 -657 30 -631
<< polycont >>
rect -17 607 17 641
<< locali >>
rect -33 607 -17 641
rect 17 607 33 641
rect -76 530 -42 573
rect -76 462 -42 492
rect -76 394 -42 420
rect -76 326 -42 348
rect -76 258 -42 276
rect -76 190 -42 204
rect -76 122 -42 132
rect -76 54 -42 60
rect -76 -14 -42 -12
rect -76 -50 -42 -48
rect -76 -122 -42 -116
rect -76 -194 -42 -184
rect -76 -266 -42 -252
rect -76 -338 -42 -320
rect -76 -410 -42 -388
rect -76 -482 -42 -456
rect -76 -554 -42 -524
rect -76 -635 -42 -592
rect 42 530 76 573
rect 42 462 76 492
rect 42 394 76 420
rect 42 326 76 348
rect 42 258 76 276
rect 42 190 76 204
rect 42 122 76 132
rect 42 54 76 60
rect 42 -14 76 -12
rect 42 -50 76 -48
rect 42 -122 76 -116
rect 42 -194 76 -184
rect 42 -266 76 -252
rect 42 -338 76 -320
rect 42 -410 76 -388
rect 42 -482 76 -456
rect 42 -554 76 -524
rect 42 -635 76 -592
<< viali >>
rect -17 607 17 641
rect -76 496 -42 526
rect -76 492 -42 496
rect -76 428 -42 454
rect -76 420 -42 428
rect -76 360 -42 382
rect -76 348 -42 360
rect -76 292 -42 310
rect -76 276 -42 292
rect -76 224 -42 238
rect -76 204 -42 224
rect -76 156 -42 166
rect -76 132 -42 156
rect -76 88 -42 94
rect -76 60 -42 88
rect -76 20 -42 22
rect -76 -12 -42 20
rect -76 -82 -42 -50
rect -76 -84 -42 -82
rect -76 -150 -42 -122
rect -76 -156 -42 -150
rect -76 -218 -42 -194
rect -76 -228 -42 -218
rect -76 -286 -42 -266
rect -76 -300 -42 -286
rect -76 -354 -42 -338
rect -76 -372 -42 -354
rect -76 -422 -42 -410
rect -76 -444 -42 -422
rect -76 -490 -42 -482
rect -76 -516 -42 -490
rect -76 -558 -42 -554
rect -76 -588 -42 -558
rect 42 496 76 526
rect 42 492 76 496
rect 42 428 76 454
rect 42 420 76 428
rect 42 360 76 382
rect 42 348 76 360
rect 42 292 76 310
rect 42 276 76 292
rect 42 224 76 238
rect 42 204 76 224
rect 42 156 76 166
rect 42 132 76 156
rect 42 88 76 94
rect 42 60 76 88
rect 42 20 76 22
rect 42 -12 76 20
rect 42 -82 76 -50
rect 42 -84 76 -82
rect 42 -150 76 -122
rect 42 -156 76 -150
rect 42 -218 76 -194
rect 42 -228 76 -218
rect 42 -286 76 -266
rect 42 -300 76 -286
rect 42 -354 76 -338
rect 42 -372 76 -354
rect 42 -422 76 -410
rect 42 -444 76 -422
rect 42 -490 76 -482
rect 42 -516 76 -490
rect 42 -558 76 -554
rect 42 -588 76 -558
<< metal1 >>
rect -29 641 29 647
rect -29 607 -17 641
rect 17 607 29 641
rect -29 601 29 607
rect -82 526 -36 569
rect -82 492 -76 526
rect -42 492 -36 526
rect -82 454 -36 492
rect -82 420 -76 454
rect -42 420 -36 454
rect -82 382 -36 420
rect -82 348 -76 382
rect -42 348 -36 382
rect -82 310 -36 348
rect -82 276 -76 310
rect -42 276 -36 310
rect -82 238 -36 276
rect -82 204 -76 238
rect -42 204 -36 238
rect -82 166 -36 204
rect -82 132 -76 166
rect -42 132 -36 166
rect -82 94 -36 132
rect -82 60 -76 94
rect -42 60 -36 94
rect -82 22 -36 60
rect -82 -12 -76 22
rect -42 -12 -36 22
rect -82 -50 -36 -12
rect -82 -84 -76 -50
rect -42 -84 -36 -50
rect -82 -122 -36 -84
rect -82 -156 -76 -122
rect -42 -156 -36 -122
rect -82 -194 -36 -156
rect -82 -228 -76 -194
rect -42 -228 -36 -194
rect -82 -266 -36 -228
rect -82 -300 -76 -266
rect -42 -300 -36 -266
rect -82 -338 -36 -300
rect -82 -372 -76 -338
rect -42 -372 -36 -338
rect -82 -410 -36 -372
rect -82 -444 -76 -410
rect -42 -444 -36 -410
rect -82 -482 -36 -444
rect -82 -516 -76 -482
rect -42 -516 -36 -482
rect -82 -554 -36 -516
rect -82 -588 -76 -554
rect -42 -588 -36 -554
rect -82 -631 -36 -588
rect 36 526 82 569
rect 36 492 42 526
rect 76 492 82 526
rect 36 454 82 492
rect 36 420 42 454
rect 76 420 82 454
rect 36 382 82 420
rect 36 348 42 382
rect 76 348 82 382
rect 36 310 82 348
rect 36 276 42 310
rect 76 276 82 310
rect 36 238 82 276
rect 36 204 42 238
rect 76 204 82 238
rect 36 166 82 204
rect 36 132 42 166
rect 76 132 82 166
rect 36 94 82 132
rect 36 60 42 94
rect 76 60 82 94
rect 36 22 82 60
rect 36 -12 42 22
rect 76 -12 82 22
rect 36 -50 82 -12
rect 36 -84 42 -50
rect 76 -84 82 -50
rect 36 -122 82 -84
rect 36 -156 42 -122
rect 76 -156 82 -122
rect 36 -194 82 -156
rect 36 -228 42 -194
rect 76 -228 82 -194
rect 36 -266 82 -228
rect 36 -300 42 -266
rect 76 -300 82 -266
rect 36 -338 82 -300
rect 36 -372 42 -338
rect 76 -372 82 -338
rect 36 -410 82 -372
rect 36 -444 42 -410
rect 76 -444 82 -410
rect 36 -482 82 -444
rect 36 -516 42 -482
rect 76 -516 82 -482
rect 36 -554 82 -516
rect 36 -588 42 -554
rect 76 -588 82 -554
rect 36 -631 82 -588
<< end >>
