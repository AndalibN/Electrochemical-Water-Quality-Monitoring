magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -523 -1500 567 1500
<< pmos >>
rect -407 -1400 -7 1400
rect 51 -1400 451 1400
<< pdiff >>
rect -487 1377 -407 1400
rect -487 1343 -475 1377
rect -441 1343 -407 1377
rect -487 1309 -407 1343
rect -487 1275 -475 1309
rect -441 1275 -407 1309
rect -487 1241 -407 1275
rect -487 1207 -475 1241
rect -441 1207 -407 1241
rect -487 1173 -407 1207
rect -487 1139 -475 1173
rect -441 1139 -407 1173
rect -487 1105 -407 1139
rect -487 1071 -475 1105
rect -441 1071 -407 1105
rect -487 1037 -407 1071
rect -487 1003 -475 1037
rect -441 1003 -407 1037
rect -487 969 -407 1003
rect -487 935 -475 969
rect -441 935 -407 969
rect -487 901 -407 935
rect -487 867 -475 901
rect -441 867 -407 901
rect -487 833 -407 867
rect -487 799 -475 833
rect -441 799 -407 833
rect -487 765 -407 799
rect -487 731 -475 765
rect -441 731 -407 765
rect -487 697 -407 731
rect -487 663 -475 697
rect -441 663 -407 697
rect -487 629 -407 663
rect -487 595 -475 629
rect -441 595 -407 629
rect -487 561 -407 595
rect -487 527 -475 561
rect -441 527 -407 561
rect -487 493 -407 527
rect -487 459 -475 493
rect -441 459 -407 493
rect -487 425 -407 459
rect -487 391 -475 425
rect -441 391 -407 425
rect -487 357 -407 391
rect -487 323 -475 357
rect -441 323 -407 357
rect -487 289 -407 323
rect -487 255 -475 289
rect -441 255 -407 289
rect -487 221 -407 255
rect -487 187 -475 221
rect -441 187 -407 221
rect -487 153 -407 187
rect -487 119 -475 153
rect -441 119 -407 153
rect -487 85 -407 119
rect -487 51 -475 85
rect -441 51 -407 85
rect -487 17 -407 51
rect -487 -17 -475 17
rect -441 -17 -407 17
rect -487 -51 -407 -17
rect -487 -85 -475 -51
rect -441 -85 -407 -51
rect -487 -119 -407 -85
rect -487 -153 -475 -119
rect -441 -153 -407 -119
rect -487 -187 -407 -153
rect -487 -221 -475 -187
rect -441 -221 -407 -187
rect -487 -255 -407 -221
rect -487 -289 -475 -255
rect -441 -289 -407 -255
rect -487 -323 -407 -289
rect -487 -357 -475 -323
rect -441 -357 -407 -323
rect -487 -391 -407 -357
rect -487 -425 -475 -391
rect -441 -425 -407 -391
rect -487 -459 -407 -425
rect -487 -493 -475 -459
rect -441 -493 -407 -459
rect -487 -527 -407 -493
rect -487 -561 -475 -527
rect -441 -561 -407 -527
rect -487 -595 -407 -561
rect -487 -629 -475 -595
rect -441 -629 -407 -595
rect -487 -663 -407 -629
rect -487 -697 -475 -663
rect -441 -697 -407 -663
rect -487 -731 -407 -697
rect -487 -765 -475 -731
rect -441 -765 -407 -731
rect -487 -799 -407 -765
rect -487 -833 -475 -799
rect -441 -833 -407 -799
rect -487 -867 -407 -833
rect -487 -901 -475 -867
rect -441 -901 -407 -867
rect -487 -935 -407 -901
rect -487 -969 -475 -935
rect -441 -969 -407 -935
rect -487 -1003 -407 -969
rect -487 -1037 -475 -1003
rect -441 -1037 -407 -1003
rect -487 -1071 -407 -1037
rect -487 -1105 -475 -1071
rect -441 -1105 -407 -1071
rect -487 -1139 -407 -1105
rect -487 -1173 -475 -1139
rect -441 -1173 -407 -1139
rect -487 -1207 -407 -1173
rect -487 -1241 -475 -1207
rect -441 -1241 -407 -1207
rect -487 -1275 -407 -1241
rect -487 -1309 -475 -1275
rect -441 -1309 -407 -1275
rect -487 -1343 -407 -1309
rect -487 -1377 -475 -1343
rect -441 -1377 -407 -1343
rect -487 -1400 -407 -1377
rect -7 1377 51 1400
rect -7 1343 5 1377
rect 39 1343 51 1377
rect -7 1309 51 1343
rect -7 1275 5 1309
rect 39 1275 51 1309
rect -7 1241 51 1275
rect -7 1207 5 1241
rect 39 1207 51 1241
rect -7 1173 51 1207
rect -7 1139 5 1173
rect 39 1139 51 1173
rect -7 1105 51 1139
rect -7 1071 5 1105
rect 39 1071 51 1105
rect -7 1037 51 1071
rect -7 1003 5 1037
rect 39 1003 51 1037
rect -7 969 51 1003
rect -7 935 5 969
rect 39 935 51 969
rect -7 901 51 935
rect -7 867 5 901
rect 39 867 51 901
rect -7 833 51 867
rect -7 799 5 833
rect 39 799 51 833
rect -7 765 51 799
rect -7 731 5 765
rect 39 731 51 765
rect -7 697 51 731
rect -7 663 5 697
rect 39 663 51 697
rect -7 629 51 663
rect -7 595 5 629
rect 39 595 51 629
rect -7 561 51 595
rect -7 527 5 561
rect 39 527 51 561
rect -7 493 51 527
rect -7 459 5 493
rect 39 459 51 493
rect -7 425 51 459
rect -7 391 5 425
rect 39 391 51 425
rect -7 357 51 391
rect -7 323 5 357
rect 39 323 51 357
rect -7 289 51 323
rect -7 255 5 289
rect 39 255 51 289
rect -7 221 51 255
rect -7 187 5 221
rect 39 187 51 221
rect -7 153 51 187
rect -7 119 5 153
rect 39 119 51 153
rect -7 85 51 119
rect -7 51 5 85
rect 39 51 51 85
rect -7 17 51 51
rect -7 -17 5 17
rect 39 -17 51 17
rect -7 -51 51 -17
rect -7 -85 5 -51
rect 39 -85 51 -51
rect -7 -119 51 -85
rect -7 -153 5 -119
rect 39 -153 51 -119
rect -7 -187 51 -153
rect -7 -221 5 -187
rect 39 -221 51 -187
rect -7 -255 51 -221
rect -7 -289 5 -255
rect 39 -289 51 -255
rect -7 -323 51 -289
rect -7 -357 5 -323
rect 39 -357 51 -323
rect -7 -391 51 -357
rect -7 -425 5 -391
rect 39 -425 51 -391
rect -7 -459 51 -425
rect -7 -493 5 -459
rect 39 -493 51 -459
rect -7 -527 51 -493
rect -7 -561 5 -527
rect 39 -561 51 -527
rect -7 -595 51 -561
rect -7 -629 5 -595
rect 39 -629 51 -595
rect -7 -663 51 -629
rect -7 -697 5 -663
rect 39 -697 51 -663
rect -7 -731 51 -697
rect -7 -765 5 -731
rect 39 -765 51 -731
rect -7 -799 51 -765
rect -7 -833 5 -799
rect 39 -833 51 -799
rect -7 -867 51 -833
rect -7 -901 5 -867
rect 39 -901 51 -867
rect -7 -935 51 -901
rect -7 -969 5 -935
rect 39 -969 51 -935
rect -7 -1003 51 -969
rect -7 -1037 5 -1003
rect 39 -1037 51 -1003
rect -7 -1071 51 -1037
rect -7 -1105 5 -1071
rect 39 -1105 51 -1071
rect -7 -1139 51 -1105
rect -7 -1173 5 -1139
rect 39 -1173 51 -1139
rect -7 -1207 51 -1173
rect -7 -1241 5 -1207
rect 39 -1241 51 -1207
rect -7 -1275 51 -1241
rect -7 -1309 5 -1275
rect 39 -1309 51 -1275
rect -7 -1343 51 -1309
rect -7 -1377 5 -1343
rect 39 -1377 51 -1343
rect -7 -1400 51 -1377
rect 451 1377 531 1400
rect 451 1343 474 1377
rect 508 1343 531 1377
rect 451 1309 531 1343
rect 451 1275 474 1309
rect 508 1275 531 1309
rect 451 1241 531 1275
rect 451 1207 474 1241
rect 508 1207 531 1241
rect 451 1173 531 1207
rect 451 1139 474 1173
rect 508 1139 531 1173
rect 451 1105 531 1139
rect 451 1071 474 1105
rect 508 1071 531 1105
rect 451 1037 531 1071
rect 451 1003 474 1037
rect 508 1003 531 1037
rect 451 969 531 1003
rect 451 935 474 969
rect 508 935 531 969
rect 451 901 531 935
rect 451 867 474 901
rect 508 867 531 901
rect 451 833 531 867
rect 451 799 474 833
rect 508 799 531 833
rect 451 765 531 799
rect 451 731 474 765
rect 508 731 531 765
rect 451 697 531 731
rect 451 663 474 697
rect 508 663 531 697
rect 451 629 531 663
rect 451 595 474 629
rect 508 595 531 629
rect 451 561 531 595
rect 451 527 474 561
rect 508 527 531 561
rect 451 493 531 527
rect 451 459 474 493
rect 508 459 531 493
rect 451 425 531 459
rect 451 391 474 425
rect 508 391 531 425
rect 451 357 531 391
rect 451 323 474 357
rect 508 323 531 357
rect 451 289 531 323
rect 451 255 474 289
rect 508 255 531 289
rect 451 221 531 255
rect 451 187 474 221
rect 508 187 531 221
rect 451 153 531 187
rect 451 119 474 153
rect 508 119 531 153
rect 451 85 531 119
rect 451 51 474 85
rect 508 51 531 85
rect 451 17 531 51
rect 451 -17 474 17
rect 508 -17 531 17
rect 451 -51 531 -17
rect 451 -85 474 -51
rect 508 -85 531 -51
rect 451 -119 531 -85
rect 451 -153 474 -119
rect 508 -153 531 -119
rect 451 -187 531 -153
rect 451 -221 474 -187
rect 508 -221 531 -187
rect 451 -255 531 -221
rect 451 -289 474 -255
rect 508 -289 531 -255
rect 451 -323 531 -289
rect 451 -357 474 -323
rect 508 -357 531 -323
rect 451 -391 531 -357
rect 451 -425 474 -391
rect 508 -425 531 -391
rect 451 -459 531 -425
rect 451 -493 474 -459
rect 508 -493 531 -459
rect 451 -527 531 -493
rect 451 -561 474 -527
rect 508 -561 531 -527
rect 451 -595 531 -561
rect 451 -629 474 -595
rect 508 -629 531 -595
rect 451 -663 531 -629
rect 451 -697 474 -663
rect 508 -697 531 -663
rect 451 -731 531 -697
rect 451 -765 474 -731
rect 508 -765 531 -731
rect 451 -799 531 -765
rect 451 -833 474 -799
rect 508 -833 531 -799
rect 451 -867 531 -833
rect 451 -901 474 -867
rect 508 -901 531 -867
rect 451 -935 531 -901
rect 451 -969 474 -935
rect 508 -969 531 -935
rect 451 -1003 531 -969
rect 451 -1037 474 -1003
rect 508 -1037 531 -1003
rect 451 -1071 531 -1037
rect 451 -1105 474 -1071
rect 508 -1105 531 -1071
rect 451 -1139 531 -1105
rect 451 -1173 474 -1139
rect 508 -1173 531 -1139
rect 451 -1207 531 -1173
rect 451 -1241 474 -1207
rect 508 -1241 531 -1207
rect 451 -1275 531 -1241
rect 451 -1309 474 -1275
rect 508 -1309 531 -1275
rect 451 -1343 531 -1309
rect 451 -1377 474 -1343
rect 508 -1377 531 -1343
rect 451 -1400 531 -1377
<< pdiffc >>
rect -475 1343 -441 1377
rect -475 1275 -441 1309
rect -475 1207 -441 1241
rect -475 1139 -441 1173
rect -475 1071 -441 1105
rect -475 1003 -441 1037
rect -475 935 -441 969
rect -475 867 -441 901
rect -475 799 -441 833
rect -475 731 -441 765
rect -475 663 -441 697
rect -475 595 -441 629
rect -475 527 -441 561
rect -475 459 -441 493
rect -475 391 -441 425
rect -475 323 -441 357
rect -475 255 -441 289
rect -475 187 -441 221
rect -475 119 -441 153
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -475 -153 -441 -119
rect -475 -221 -441 -187
rect -475 -289 -441 -255
rect -475 -357 -441 -323
rect -475 -425 -441 -391
rect -475 -493 -441 -459
rect -475 -561 -441 -527
rect -475 -629 -441 -595
rect -475 -697 -441 -663
rect -475 -765 -441 -731
rect -475 -833 -441 -799
rect -475 -901 -441 -867
rect -475 -969 -441 -935
rect -475 -1037 -441 -1003
rect -475 -1105 -441 -1071
rect -475 -1173 -441 -1139
rect -475 -1241 -441 -1207
rect -475 -1309 -441 -1275
rect -475 -1377 -441 -1343
rect 5 1343 39 1377
rect 5 1275 39 1309
rect 5 1207 39 1241
rect 5 1139 39 1173
rect 5 1071 39 1105
rect 5 1003 39 1037
rect 5 935 39 969
rect 5 867 39 901
rect 5 799 39 833
rect 5 731 39 765
rect 5 663 39 697
rect 5 595 39 629
rect 5 527 39 561
rect 5 459 39 493
rect 5 391 39 425
rect 5 323 39 357
rect 5 255 39 289
rect 5 187 39 221
rect 5 119 39 153
rect 5 51 39 85
rect 5 -17 39 17
rect 5 -85 39 -51
rect 5 -153 39 -119
rect 5 -221 39 -187
rect 5 -289 39 -255
rect 5 -357 39 -323
rect 5 -425 39 -391
rect 5 -493 39 -459
rect 5 -561 39 -527
rect 5 -629 39 -595
rect 5 -697 39 -663
rect 5 -765 39 -731
rect 5 -833 39 -799
rect 5 -901 39 -867
rect 5 -969 39 -935
rect 5 -1037 39 -1003
rect 5 -1105 39 -1071
rect 5 -1173 39 -1139
rect 5 -1241 39 -1207
rect 5 -1309 39 -1275
rect 5 -1377 39 -1343
rect 474 1343 508 1377
rect 474 1275 508 1309
rect 474 1207 508 1241
rect 474 1139 508 1173
rect 474 1071 508 1105
rect 474 1003 508 1037
rect 474 935 508 969
rect 474 867 508 901
rect 474 799 508 833
rect 474 731 508 765
rect 474 663 508 697
rect 474 595 508 629
rect 474 527 508 561
rect 474 459 508 493
rect 474 391 508 425
rect 474 323 508 357
rect 474 255 508 289
rect 474 187 508 221
rect 474 119 508 153
rect 474 51 508 85
rect 474 -17 508 17
rect 474 -85 508 -51
rect 474 -153 508 -119
rect 474 -221 508 -187
rect 474 -289 508 -255
rect 474 -357 508 -323
rect 474 -425 508 -391
rect 474 -493 508 -459
rect 474 -561 508 -527
rect 474 -629 508 -595
rect 474 -697 508 -663
rect 474 -765 508 -731
rect 474 -833 508 -799
rect 474 -901 508 -867
rect 474 -969 508 -935
rect 474 -1037 508 -1003
rect 474 -1105 508 -1071
rect 474 -1173 508 -1139
rect 474 -1241 508 -1207
rect 474 -1309 508 -1275
rect 474 -1377 508 -1343
<< poly >>
rect -407 1481 -7 1497
rect -407 1447 -360 1481
rect -326 1447 -292 1481
rect -258 1447 -224 1481
rect -190 1447 -156 1481
rect -122 1447 -88 1481
rect -54 1447 -7 1481
rect -407 1400 -7 1447
rect 51 1400 451 1497
rect -407 -1434 -7 -1400
rect 51 -1434 451 -1400
rect -407 -1497 451 -1434
<< polycont >>
rect -360 1447 -326 1481
rect -292 1447 -258 1481
rect -224 1447 -190 1481
rect -156 1447 -122 1481
rect -88 1447 -54 1481
<< locali >>
rect -407 1447 -368 1481
rect -326 1447 -296 1481
rect -258 1447 -224 1481
rect -190 1447 -156 1481
rect -118 1447 -88 1481
rect -46 1447 -7 1481
rect -475 1385 -441 1404
rect -475 1313 -441 1343
rect -475 1241 -441 1275
rect -475 1173 -441 1207
rect -475 1105 -441 1135
rect -475 1037 -441 1063
rect -475 969 -441 991
rect -475 901 -441 919
rect -475 833 -441 847
rect -475 765 -441 775
rect -475 697 -441 703
rect -475 629 -441 631
rect -475 593 -441 595
rect -475 521 -441 527
rect -475 449 -441 459
rect -475 377 -441 391
rect -475 305 -441 323
rect -475 233 -441 255
rect -475 161 -441 187
rect -475 89 -441 119
rect -475 17 -441 51
rect -475 -51 -441 -17
rect -475 -119 -441 -89
rect -475 -187 -441 -161
rect -475 -255 -441 -233
rect -475 -323 -441 -305
rect -475 -391 -441 -377
rect -475 -459 -441 -449
rect -475 -527 -441 -521
rect -475 -595 -441 -593
rect -475 -631 -441 -629
rect -475 -703 -441 -697
rect -475 -775 -441 -765
rect -475 -847 -441 -833
rect -475 -919 -441 -901
rect -475 -991 -441 -969
rect -475 -1063 -441 -1037
rect -475 -1135 -441 -1105
rect -475 -1207 -441 -1173
rect -475 -1275 -441 -1241
rect -475 -1343 -441 -1313
rect -475 -1404 -441 -1385
rect 5 1385 39 1404
rect 5 1313 39 1343
rect 5 1241 39 1275
rect 5 1173 39 1207
rect 5 1105 39 1135
rect 5 1037 39 1063
rect 5 969 39 991
rect 5 901 39 919
rect 5 833 39 847
rect 5 765 39 775
rect 5 697 39 703
rect 5 629 39 631
rect 5 593 39 595
rect 5 521 39 527
rect 5 449 39 459
rect 5 377 39 391
rect 5 305 39 323
rect 5 233 39 255
rect 5 161 39 187
rect 5 89 39 119
rect 5 17 39 51
rect 5 -51 39 -17
rect 5 -119 39 -89
rect 5 -187 39 -161
rect 5 -255 39 -233
rect 5 -323 39 -305
rect 5 -391 39 -377
rect 5 -459 39 -449
rect 5 -527 39 -521
rect 5 -595 39 -593
rect 5 -631 39 -629
rect 5 -703 39 -697
rect 5 -775 39 -765
rect 5 -847 39 -833
rect 5 -919 39 -901
rect 5 -991 39 -969
rect 5 -1063 39 -1037
rect 5 -1135 39 -1105
rect 5 -1207 39 -1173
rect 5 -1275 39 -1241
rect 5 -1343 39 -1313
rect 5 -1404 39 -1385
rect 474 1385 508 1404
rect 474 1313 508 1343
rect 474 1241 508 1275
rect 474 1173 508 1207
rect 474 1105 508 1135
rect 474 1037 508 1063
rect 474 969 508 991
rect 474 901 508 919
rect 474 833 508 847
rect 474 765 508 775
rect 474 697 508 703
rect 474 629 508 631
rect 474 593 508 595
rect 474 521 508 527
rect 474 449 508 459
rect 474 377 508 391
rect 474 305 508 323
rect 474 233 508 255
rect 474 161 508 187
rect 474 89 508 119
rect 474 17 508 51
rect 474 -51 508 -17
rect 474 -119 508 -89
rect 474 -187 508 -161
rect 474 -255 508 -233
rect 474 -323 508 -305
rect 474 -391 508 -377
rect 474 -459 508 -449
rect 474 -527 508 -521
rect 474 -595 508 -593
rect 474 -631 508 -629
rect 474 -703 508 -697
rect 474 -775 508 -765
rect 474 -847 508 -833
rect 474 -919 508 -901
rect 474 -991 508 -969
rect 474 -1063 508 -1037
rect 474 -1135 508 -1105
rect 474 -1207 508 -1173
rect 474 -1275 508 -1241
rect 474 -1343 508 -1313
rect 474 -1404 508 -1385
<< viali >>
rect -368 1447 -360 1481
rect -360 1447 -334 1481
rect -296 1447 -292 1481
rect -292 1447 -262 1481
rect -224 1447 -190 1481
rect -152 1447 -122 1481
rect -122 1447 -118 1481
rect -80 1447 -54 1481
rect -54 1447 -46 1481
rect -475 1377 -441 1385
rect -475 1351 -441 1377
rect -475 1309 -441 1313
rect -475 1279 -441 1309
rect -475 1207 -441 1241
rect -475 1139 -441 1169
rect -475 1135 -441 1139
rect -475 1071 -441 1097
rect -475 1063 -441 1071
rect -475 1003 -441 1025
rect -475 991 -441 1003
rect -475 935 -441 953
rect -475 919 -441 935
rect -475 867 -441 881
rect -475 847 -441 867
rect -475 799 -441 809
rect -475 775 -441 799
rect -475 731 -441 737
rect -475 703 -441 731
rect -475 663 -441 665
rect -475 631 -441 663
rect -475 561 -441 593
rect -475 559 -441 561
rect -475 493 -441 521
rect -475 487 -441 493
rect -475 425 -441 449
rect -475 415 -441 425
rect -475 357 -441 377
rect -475 343 -441 357
rect -475 289 -441 305
rect -475 271 -441 289
rect -475 221 -441 233
rect -475 199 -441 221
rect -475 153 -441 161
rect -475 127 -441 153
rect -475 85 -441 89
rect -475 55 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -55
rect -475 -89 -441 -85
rect -475 -153 -441 -127
rect -475 -161 -441 -153
rect -475 -221 -441 -199
rect -475 -233 -441 -221
rect -475 -289 -441 -271
rect -475 -305 -441 -289
rect -475 -357 -441 -343
rect -475 -377 -441 -357
rect -475 -425 -441 -415
rect -475 -449 -441 -425
rect -475 -493 -441 -487
rect -475 -521 -441 -493
rect -475 -561 -441 -559
rect -475 -593 -441 -561
rect -475 -663 -441 -631
rect -475 -665 -441 -663
rect -475 -731 -441 -703
rect -475 -737 -441 -731
rect -475 -799 -441 -775
rect -475 -809 -441 -799
rect -475 -867 -441 -847
rect -475 -881 -441 -867
rect -475 -935 -441 -919
rect -475 -953 -441 -935
rect -475 -1003 -441 -991
rect -475 -1025 -441 -1003
rect -475 -1071 -441 -1063
rect -475 -1097 -441 -1071
rect -475 -1139 -441 -1135
rect -475 -1169 -441 -1139
rect -475 -1241 -441 -1207
rect -475 -1309 -441 -1279
rect -475 -1313 -441 -1309
rect -475 -1377 -441 -1351
rect -475 -1385 -441 -1377
rect 5 1377 39 1385
rect 5 1351 39 1377
rect 5 1309 39 1313
rect 5 1279 39 1309
rect 5 1207 39 1241
rect 5 1139 39 1169
rect 5 1135 39 1139
rect 5 1071 39 1097
rect 5 1063 39 1071
rect 5 1003 39 1025
rect 5 991 39 1003
rect 5 935 39 953
rect 5 919 39 935
rect 5 867 39 881
rect 5 847 39 867
rect 5 799 39 809
rect 5 775 39 799
rect 5 731 39 737
rect 5 703 39 731
rect 5 663 39 665
rect 5 631 39 663
rect 5 561 39 593
rect 5 559 39 561
rect 5 493 39 521
rect 5 487 39 493
rect 5 425 39 449
rect 5 415 39 425
rect 5 357 39 377
rect 5 343 39 357
rect 5 289 39 305
rect 5 271 39 289
rect 5 221 39 233
rect 5 199 39 221
rect 5 153 39 161
rect 5 127 39 153
rect 5 85 39 89
rect 5 55 39 85
rect 5 -17 39 17
rect 5 -85 39 -55
rect 5 -89 39 -85
rect 5 -153 39 -127
rect 5 -161 39 -153
rect 5 -221 39 -199
rect 5 -233 39 -221
rect 5 -289 39 -271
rect 5 -305 39 -289
rect 5 -357 39 -343
rect 5 -377 39 -357
rect 5 -425 39 -415
rect 5 -449 39 -425
rect 5 -493 39 -487
rect 5 -521 39 -493
rect 5 -561 39 -559
rect 5 -593 39 -561
rect 5 -663 39 -631
rect 5 -665 39 -663
rect 5 -731 39 -703
rect 5 -737 39 -731
rect 5 -799 39 -775
rect 5 -809 39 -799
rect 5 -867 39 -847
rect 5 -881 39 -867
rect 5 -935 39 -919
rect 5 -953 39 -935
rect 5 -1003 39 -991
rect 5 -1025 39 -1003
rect 5 -1071 39 -1063
rect 5 -1097 39 -1071
rect 5 -1139 39 -1135
rect 5 -1169 39 -1139
rect 5 -1241 39 -1207
rect 5 -1309 39 -1279
rect 5 -1313 39 -1309
rect 5 -1377 39 -1351
rect 5 -1385 39 -1377
rect 474 1377 508 1385
rect 474 1351 508 1377
rect 474 1309 508 1313
rect 474 1279 508 1309
rect 474 1207 508 1241
rect 474 1139 508 1169
rect 474 1135 508 1139
rect 474 1071 508 1097
rect 474 1063 508 1071
rect 474 1003 508 1025
rect 474 991 508 1003
rect 474 935 508 953
rect 474 919 508 935
rect 474 867 508 881
rect 474 847 508 867
rect 474 799 508 809
rect 474 775 508 799
rect 474 731 508 737
rect 474 703 508 731
rect 474 663 508 665
rect 474 631 508 663
rect 474 561 508 593
rect 474 559 508 561
rect 474 493 508 521
rect 474 487 508 493
rect 474 425 508 449
rect 474 415 508 425
rect 474 357 508 377
rect 474 343 508 357
rect 474 289 508 305
rect 474 271 508 289
rect 474 221 508 233
rect 474 199 508 221
rect 474 153 508 161
rect 474 127 508 153
rect 474 85 508 89
rect 474 55 508 85
rect 474 -17 508 17
rect 474 -85 508 -55
rect 474 -89 508 -85
rect 474 -153 508 -127
rect 474 -161 508 -153
rect 474 -221 508 -199
rect 474 -233 508 -221
rect 474 -289 508 -271
rect 474 -305 508 -289
rect 474 -357 508 -343
rect 474 -377 508 -357
rect 474 -425 508 -415
rect 474 -449 508 -425
rect 474 -493 508 -487
rect 474 -521 508 -493
rect 474 -561 508 -559
rect 474 -593 508 -561
rect 474 -663 508 -631
rect 474 -665 508 -663
rect 474 -731 508 -703
rect 474 -737 508 -731
rect 474 -799 508 -775
rect 474 -809 508 -799
rect 474 -867 508 -847
rect 474 -881 508 -867
rect 474 -935 508 -919
rect 474 -953 508 -935
rect 474 -1003 508 -991
rect 474 -1025 508 -1003
rect 474 -1071 508 -1063
rect 474 -1097 508 -1071
rect 474 -1139 508 -1135
rect 474 -1169 508 -1139
rect 474 -1241 508 -1207
rect 474 -1309 508 -1279
rect 474 -1313 508 -1309
rect 474 -1377 508 -1351
rect 474 -1385 508 -1377
<< metal1 >>
rect -403 1481 -11 1487
rect -403 1447 -368 1481
rect -334 1447 -296 1481
rect -262 1447 -224 1481
rect -190 1447 -152 1481
rect -118 1447 -80 1481
rect -46 1447 -11 1481
rect -403 1441 -11 1447
rect -481 1385 -435 1400
rect -481 1351 -475 1385
rect -441 1351 -435 1385
rect -481 1313 -435 1351
rect -481 1279 -475 1313
rect -441 1279 -435 1313
rect -481 1241 -435 1279
rect -481 1207 -475 1241
rect -441 1207 -435 1241
rect -481 1169 -435 1207
rect -481 1135 -475 1169
rect -441 1135 -435 1169
rect -481 1097 -435 1135
rect -481 1063 -475 1097
rect -441 1063 -435 1097
rect -481 1025 -435 1063
rect -481 991 -475 1025
rect -441 991 -435 1025
rect -481 953 -435 991
rect -481 919 -475 953
rect -441 919 -435 953
rect -481 881 -435 919
rect -481 847 -475 881
rect -441 847 -435 881
rect -481 809 -435 847
rect -481 775 -475 809
rect -441 775 -435 809
rect -481 737 -435 775
rect -481 703 -475 737
rect -441 703 -435 737
rect -481 665 -435 703
rect -481 631 -475 665
rect -441 631 -435 665
rect -481 593 -435 631
rect -481 559 -475 593
rect -441 559 -435 593
rect -481 521 -435 559
rect -481 487 -475 521
rect -441 487 -435 521
rect -481 449 -435 487
rect -481 415 -475 449
rect -441 415 -435 449
rect -481 377 -435 415
rect -481 343 -475 377
rect -441 343 -435 377
rect -481 305 -435 343
rect -481 271 -475 305
rect -441 271 -435 305
rect -481 233 -435 271
rect -481 199 -475 233
rect -441 199 -435 233
rect -481 161 -435 199
rect -481 127 -475 161
rect -441 127 -435 161
rect -481 89 -435 127
rect -481 55 -475 89
rect -441 55 -435 89
rect -481 17 -435 55
rect -481 -17 -475 17
rect -441 -17 -435 17
rect -481 -55 -435 -17
rect -481 -89 -475 -55
rect -441 -89 -435 -55
rect -481 -127 -435 -89
rect -481 -161 -475 -127
rect -441 -161 -435 -127
rect -481 -199 -435 -161
rect -481 -233 -475 -199
rect -441 -233 -435 -199
rect -481 -271 -435 -233
rect -481 -305 -475 -271
rect -441 -305 -435 -271
rect -481 -343 -435 -305
rect -481 -377 -475 -343
rect -441 -377 -435 -343
rect -481 -415 -435 -377
rect -481 -449 -475 -415
rect -441 -449 -435 -415
rect -481 -487 -435 -449
rect -481 -521 -475 -487
rect -441 -521 -435 -487
rect -481 -559 -435 -521
rect -481 -593 -475 -559
rect -441 -593 -435 -559
rect -481 -631 -435 -593
rect -481 -665 -475 -631
rect -441 -665 -435 -631
rect -481 -703 -435 -665
rect -481 -737 -475 -703
rect -441 -737 -435 -703
rect -481 -775 -435 -737
rect -481 -809 -475 -775
rect -441 -809 -435 -775
rect -481 -847 -435 -809
rect -481 -881 -475 -847
rect -441 -881 -435 -847
rect -481 -919 -435 -881
rect -481 -953 -475 -919
rect -441 -953 -435 -919
rect -481 -991 -435 -953
rect -481 -1025 -475 -991
rect -441 -1025 -435 -991
rect -481 -1063 -435 -1025
rect -481 -1097 -475 -1063
rect -441 -1097 -435 -1063
rect -481 -1135 -435 -1097
rect -481 -1169 -475 -1135
rect -441 -1169 -435 -1135
rect -481 -1207 -435 -1169
rect -481 -1241 -475 -1207
rect -441 -1241 -435 -1207
rect -481 -1279 -435 -1241
rect -481 -1313 -475 -1279
rect -441 -1313 -435 -1279
rect -481 -1351 -435 -1313
rect -481 -1385 -475 -1351
rect -441 -1385 -435 -1351
rect -481 -1400 -435 -1385
rect -1 1385 45 1400
rect -1 1351 5 1385
rect 39 1351 45 1385
rect -1 1313 45 1351
rect -1 1279 5 1313
rect 39 1279 45 1313
rect -1 1241 45 1279
rect -1 1207 5 1241
rect 39 1207 45 1241
rect -1 1169 45 1207
rect -1 1135 5 1169
rect 39 1135 45 1169
rect -1 1097 45 1135
rect -1 1063 5 1097
rect 39 1063 45 1097
rect -1 1025 45 1063
rect -1 991 5 1025
rect 39 991 45 1025
rect -1 953 45 991
rect -1 919 5 953
rect 39 919 45 953
rect -1 881 45 919
rect -1 847 5 881
rect 39 847 45 881
rect -1 809 45 847
rect -1 775 5 809
rect 39 775 45 809
rect -1 737 45 775
rect -1 703 5 737
rect 39 703 45 737
rect -1 665 45 703
rect -1 631 5 665
rect 39 631 45 665
rect -1 593 45 631
rect -1 559 5 593
rect 39 559 45 593
rect -1 521 45 559
rect -1 487 5 521
rect 39 487 45 521
rect -1 449 45 487
rect -1 415 5 449
rect 39 415 45 449
rect -1 377 45 415
rect -1 343 5 377
rect 39 343 45 377
rect -1 305 45 343
rect -1 271 5 305
rect 39 271 45 305
rect -1 233 45 271
rect -1 199 5 233
rect 39 199 45 233
rect -1 161 45 199
rect -1 127 5 161
rect 39 127 45 161
rect -1 89 45 127
rect -1 55 5 89
rect 39 55 45 89
rect -1 17 45 55
rect -1 -17 5 17
rect 39 -17 45 17
rect -1 -55 45 -17
rect -1 -89 5 -55
rect 39 -89 45 -55
rect -1 -127 45 -89
rect -1 -161 5 -127
rect 39 -161 45 -127
rect -1 -199 45 -161
rect -1 -233 5 -199
rect 39 -233 45 -199
rect -1 -271 45 -233
rect -1 -305 5 -271
rect 39 -305 45 -271
rect -1 -343 45 -305
rect -1 -377 5 -343
rect 39 -377 45 -343
rect -1 -415 45 -377
rect -1 -449 5 -415
rect 39 -449 45 -415
rect -1 -487 45 -449
rect -1 -521 5 -487
rect 39 -521 45 -487
rect -1 -559 45 -521
rect -1 -593 5 -559
rect 39 -593 45 -559
rect -1 -631 45 -593
rect -1 -665 5 -631
rect 39 -665 45 -631
rect -1 -703 45 -665
rect -1 -737 5 -703
rect 39 -737 45 -703
rect -1 -775 45 -737
rect -1 -809 5 -775
rect 39 -809 45 -775
rect -1 -847 45 -809
rect -1 -881 5 -847
rect 39 -881 45 -847
rect -1 -919 45 -881
rect -1 -953 5 -919
rect 39 -953 45 -919
rect -1 -991 45 -953
rect -1 -1025 5 -991
rect 39 -1025 45 -991
rect -1 -1063 45 -1025
rect -1 -1097 5 -1063
rect 39 -1097 45 -1063
rect -1 -1135 45 -1097
rect -1 -1169 5 -1135
rect 39 -1169 45 -1135
rect -1 -1207 45 -1169
rect -1 -1241 5 -1207
rect 39 -1241 45 -1207
rect -1 -1279 45 -1241
rect -1 -1313 5 -1279
rect 39 -1313 45 -1279
rect -1 -1351 45 -1313
rect -1 -1385 5 -1351
rect 39 -1385 45 -1351
rect -1 -1400 45 -1385
rect 468 1385 514 1400
rect 468 1351 474 1385
rect 508 1351 514 1385
rect 468 1313 514 1351
rect 468 1279 474 1313
rect 508 1279 514 1313
rect 468 1241 514 1279
rect 468 1207 474 1241
rect 508 1207 514 1241
rect 468 1169 514 1207
rect 468 1135 474 1169
rect 508 1135 514 1169
rect 468 1097 514 1135
rect 468 1063 474 1097
rect 508 1063 514 1097
rect 468 1025 514 1063
rect 468 991 474 1025
rect 508 991 514 1025
rect 468 953 514 991
rect 468 919 474 953
rect 508 919 514 953
rect 468 881 514 919
rect 468 847 474 881
rect 508 847 514 881
rect 468 809 514 847
rect 468 775 474 809
rect 508 775 514 809
rect 468 737 514 775
rect 468 703 474 737
rect 508 703 514 737
rect 468 665 514 703
rect 468 631 474 665
rect 508 631 514 665
rect 468 593 514 631
rect 468 559 474 593
rect 508 559 514 593
rect 468 521 514 559
rect 468 487 474 521
rect 508 487 514 521
rect 468 449 514 487
rect 468 415 474 449
rect 508 415 514 449
rect 468 377 514 415
rect 468 343 474 377
rect 508 343 514 377
rect 468 305 514 343
rect 468 271 474 305
rect 508 271 514 305
rect 468 233 514 271
rect 468 199 474 233
rect 508 199 514 233
rect 468 161 514 199
rect 468 127 474 161
rect 508 127 514 161
rect 468 89 514 127
rect 468 55 474 89
rect 508 55 514 89
rect 468 17 514 55
rect 468 -17 474 17
rect 508 -17 514 17
rect 468 -55 514 -17
rect 468 -89 474 -55
rect 508 -89 514 -55
rect 468 -127 514 -89
rect 468 -161 474 -127
rect 508 -161 514 -127
rect 468 -199 514 -161
rect 468 -233 474 -199
rect 508 -233 514 -199
rect 468 -271 514 -233
rect 468 -305 474 -271
rect 508 -305 514 -271
rect 468 -343 514 -305
rect 468 -377 474 -343
rect 508 -377 514 -343
rect 468 -415 514 -377
rect 468 -449 474 -415
rect 508 -449 514 -415
rect 468 -487 514 -449
rect 468 -521 474 -487
rect 508 -521 514 -487
rect 468 -559 514 -521
rect 468 -593 474 -559
rect 508 -593 514 -559
rect 468 -631 514 -593
rect 468 -665 474 -631
rect 508 -665 514 -631
rect 468 -703 514 -665
rect 468 -737 474 -703
rect 508 -737 514 -703
rect 468 -775 514 -737
rect 468 -809 474 -775
rect 508 -809 514 -775
rect 468 -847 514 -809
rect 468 -881 474 -847
rect 508 -881 514 -847
rect 468 -919 514 -881
rect 468 -953 474 -919
rect 508 -953 514 -919
rect 468 -991 514 -953
rect 468 -1025 474 -991
rect 508 -1025 514 -991
rect 468 -1063 514 -1025
rect 468 -1097 474 -1063
rect 508 -1097 514 -1063
rect 468 -1135 514 -1097
rect 468 -1169 474 -1135
rect 508 -1169 514 -1135
rect 468 -1207 514 -1169
rect 468 -1241 474 -1207
rect 508 -1241 514 -1207
rect 468 -1279 514 -1241
rect 468 -1313 474 -1279
rect 508 -1313 514 -1279
rect 468 -1351 514 -1313
rect 468 -1385 474 -1351
rect 508 -1385 514 -1351
rect 468 -1400 514 -1385
<< end >>
