magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 300 35 732
rect -35 -732 35 -300
<< xpolyres >>
rect -35 -300 35 300
<< viali >>
rect -17 678 17 712
rect -17 606 17 640
rect -17 534 17 568
rect -17 462 17 496
rect -17 390 17 424
rect -17 318 17 352
rect -17 -353 17 -319
rect -17 -425 17 -391
rect -17 -497 17 -463
rect -17 -569 17 -535
rect -17 -641 17 -607
rect -17 -713 17 -679
<< metal1 >>
rect -25 712 25 726
rect -25 678 -17 712
rect 17 678 25 712
rect -25 640 25 678
rect -25 606 -17 640
rect 17 606 25 640
rect -25 568 25 606
rect -25 534 -17 568
rect 17 534 25 568
rect -25 496 25 534
rect -25 462 -17 496
rect 17 462 25 496
rect -25 424 25 462
rect -25 390 -17 424
rect 17 390 25 424
rect -25 352 25 390
rect -25 318 -17 352
rect 17 318 25 352
rect -25 305 25 318
rect -25 -319 25 -305
rect -25 -353 -17 -319
rect 17 -353 25 -319
rect -25 -391 25 -353
rect -25 -425 -17 -391
rect 17 -425 25 -391
rect -25 -463 25 -425
rect -25 -497 -17 -463
rect 17 -497 25 -463
rect -25 -535 25 -497
rect -25 -569 -17 -535
rect 17 -569 25 -535
rect -25 -607 25 -569
rect -25 -641 -17 -607
rect 17 -641 25 -607
rect -25 -679 25 -641
rect -25 -713 -17 -679
rect 17 -713 25 -679
rect -25 -726 25 -713
<< end >>
