magic
tech sky130A
magscale 1 2
timestamp 1667588522
<< xpolycontact >>
rect -35 9090 35 9522
rect -35 -9522 35 -9090
<< xpolyres >>
rect -35 -9090 35 9090
<< viali >>
rect -19 9107 19 9504
rect -19 -9504 19 -9107
<< metal1 >>
rect -25 9504 25 9516
rect -25 9107 -19 9504
rect 19 9107 25 9504
rect -25 9095 25 9107
rect -25 -9107 25 -9095
rect -25 -9504 -19 -9107
rect 19 -9504 25 -9107
rect -25 -9516 25 -9504
<< res0p35 >>
rect -37 -9092 37 9092
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 90.9 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 520.504k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
