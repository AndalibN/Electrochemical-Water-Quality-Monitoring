magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -850 752 849 800
rect -850 688 765 752
rect 829 688 849 752
rect -850 672 849 688
rect -850 608 765 672
rect 829 608 849 672
rect -850 592 849 608
rect -850 528 765 592
rect 829 528 849 592
rect -850 512 849 528
rect -850 448 765 512
rect 829 448 849 512
rect -850 432 849 448
rect -850 368 765 432
rect 829 368 849 432
rect -850 352 849 368
rect -850 288 765 352
rect 829 288 849 352
rect -850 272 849 288
rect -850 208 765 272
rect 829 208 849 272
rect -850 192 849 208
rect -850 128 765 192
rect 829 128 849 192
rect -850 112 849 128
rect -850 48 765 112
rect 829 48 849 112
rect -850 32 849 48
rect -850 -32 765 32
rect 829 -32 849 32
rect -850 -48 849 -32
rect -850 -112 765 -48
rect 829 -112 849 -48
rect -850 -128 849 -112
rect -850 -192 765 -128
rect 829 -192 849 -128
rect -850 -208 849 -192
rect -850 -272 765 -208
rect 829 -272 849 -208
rect -850 -288 849 -272
rect -850 -352 765 -288
rect 829 -352 849 -288
rect -850 -368 849 -352
rect -850 -432 765 -368
rect 829 -432 849 -368
rect -850 -448 849 -432
rect -850 -512 765 -448
rect 829 -512 849 -448
rect -850 -528 849 -512
rect -850 -592 765 -528
rect 829 -592 849 -528
rect -850 -608 849 -592
rect -850 -672 765 -608
rect 829 -672 849 -608
rect -850 -688 849 -672
rect -850 -752 765 -688
rect 829 -752 849 -688
rect -850 -800 849 -752
<< via3 >>
rect 765 688 829 752
rect 765 608 829 672
rect 765 528 829 592
rect 765 448 829 512
rect 765 368 829 432
rect 765 288 829 352
rect 765 208 829 272
rect 765 128 829 192
rect 765 48 829 112
rect 765 -32 829 32
rect 765 -112 829 -48
rect 765 -192 829 -128
rect 765 -272 829 -208
rect 765 -352 829 -288
rect 765 -432 829 -368
rect 765 -512 829 -448
rect 765 -592 829 -528
rect 765 -672 829 -608
rect 765 -752 829 -688
<< mimcap >>
rect -750 632 650 700
rect -750 -632 -682 632
rect 582 -632 650 632
rect -750 -700 650 -632
<< mimcapcontact >>
rect -682 -632 582 632
<< metal4 >>
rect 749 752 845 788
rect 749 688 765 752
rect 829 688 845 752
rect 749 672 845 688
rect -711 632 611 661
rect -711 -632 -682 632
rect 582 -632 611 632
rect -711 -661 611 -632
rect 749 608 765 672
rect 829 608 845 672
rect 749 592 845 608
rect 749 528 765 592
rect 829 528 845 592
rect 749 512 845 528
rect 749 448 765 512
rect 829 448 845 512
rect 749 432 845 448
rect 749 368 765 432
rect 829 368 845 432
rect 749 352 845 368
rect 749 288 765 352
rect 829 288 845 352
rect 749 272 845 288
rect 749 208 765 272
rect 829 208 845 272
rect 749 192 845 208
rect 749 128 765 192
rect 829 128 845 192
rect 749 112 845 128
rect 749 48 765 112
rect 829 48 845 112
rect 749 32 845 48
rect 749 -32 765 32
rect 829 -32 845 32
rect 749 -48 845 -32
rect 749 -112 765 -48
rect 829 -112 845 -48
rect 749 -128 845 -112
rect 749 -192 765 -128
rect 829 -192 845 -128
rect 749 -208 845 -192
rect 749 -272 765 -208
rect 829 -272 845 -208
rect 749 -288 845 -272
rect 749 -352 765 -288
rect 829 -352 845 -288
rect 749 -368 845 -352
rect 749 -432 765 -368
rect 829 -432 845 -368
rect 749 -448 845 -432
rect 749 -512 765 -448
rect 829 -512 845 -448
rect 749 -528 845 -512
rect 749 -592 765 -528
rect 829 -592 845 -528
rect 749 -608 845 -592
rect 749 -672 765 -608
rect 829 -672 845 -608
rect 749 -688 845 -672
rect 749 -752 765 -688
rect 829 -752 845 -688
rect 749 -788 845 -752
<< properties >>
string FIXED_BBOX -850 -800 750 800
<< end >>
