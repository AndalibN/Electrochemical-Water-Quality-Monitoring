magic
tech sky130A
magscale 1 2
timestamp 1668094110
<< error_p >>
rect -29 672 29 678
rect -29 638 -17 672
rect -29 632 29 638
rect -29 -638 29 -632
rect -29 -672 -17 -638
rect -29 -678 29 -672
<< nmos >>
rect -30 -600 30 600
<< ndiff >>
rect -88 588 -30 600
rect -88 -588 -76 588
rect -42 -588 -30 588
rect -88 -600 -30 -588
rect 30 588 88 600
rect 30 -588 42 588
rect 76 -588 88 588
rect 30 -600 88 -588
<< ndiffc >>
rect -76 -588 -42 588
rect 42 -588 76 588
<< poly >>
rect -33 672 33 688
rect -33 638 -17 672
rect 17 638 33 672
rect -33 622 33 638
rect -30 600 30 622
rect -30 -622 30 -600
rect -33 -638 33 -622
rect -33 -672 -17 -638
rect 17 -672 33 -638
rect -33 -688 33 -672
<< polycont >>
rect -17 638 17 672
rect -17 -672 17 -638
<< locali >>
rect -33 638 -17 672
rect 17 638 33 672
rect -76 588 -42 604
rect -76 -604 -42 -588
rect 42 588 76 604
rect 42 -604 76 -588
rect -33 -672 -17 -638
rect 17 -672 33 -638
<< viali >>
rect -17 638 17 672
rect -76 -588 -42 588
rect 42 -588 76 588
rect -17 -672 17 -638
<< metal1 >>
rect -29 672 29 678
rect -29 638 -17 672
rect 17 638 29 672
rect -29 632 29 638
rect -82 588 -36 600
rect -82 -588 -76 588
rect -42 -588 -36 588
rect -82 -600 -36 -588
rect 36 588 82 600
rect 36 -588 42 588
rect 76 -588 82 588
rect 36 -600 82 -588
rect -29 -638 29 -632
rect -29 -672 -17 -638
rect 17 -672 29 -638
rect -29 -678 29 -672
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
