magic
tech sky130A
magscale 1 2
timestamp 1667408630
<< nwell >>
rect -294 -2064 294 2098
<< pmos >>
rect -200 -1964 200 2036
<< pdiff >>
rect -258 2024 -200 2036
rect -258 -1952 -246 2024
rect -212 -1952 -200 2024
rect -258 -1964 -200 -1952
rect 200 2024 258 2036
rect 200 -1952 212 2024
rect 246 -1952 258 2024
rect 200 -1964 258 -1952
<< pdiffc >>
rect -246 -1952 -212 2024
rect 212 -1952 246 2024
<< poly >>
rect -200 2036 200 2062
rect -200 -2011 200 -1964
rect -200 -2045 -184 -2011
rect 184 -2045 200 -2011
rect -200 -2061 200 -2045
<< polycont >>
rect -184 -2045 184 -2011
<< locali >>
rect -246 2024 -212 2040
rect -246 -1968 -212 -1952
rect 212 2024 246 2040
rect 212 -1968 246 -1952
rect -200 -2045 -184 -2011
rect 184 -2045 200 -2011
<< viali >>
rect -246 -1952 -212 2024
rect 212 -1952 246 2024
rect -184 -2045 184 -2011
<< metal1 >>
rect -252 2024 -206 2036
rect -252 -1952 -246 2024
rect -212 -1952 -206 2024
rect -252 -1964 -206 -1952
rect 206 2024 252 2036
rect 206 -1952 212 2024
rect 246 -1952 252 2024
rect 206 -1964 252 -1952
rect -196 -2011 196 -2005
rect -196 -2045 -184 -2011
rect 184 -2045 196 -2011
rect -196 -2051 196 -2045
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
