magic
tech sky130A
magscale 1 2
timestamp 1668370622
<< nmos >>
rect -561 -6000 -501 6000
rect -443 -6000 -383 6000
rect -325 -6000 -265 6000
rect -207 -6000 -147 6000
rect -89 -6000 -29 6000
rect 29 -6000 89 6000
rect 147 -6000 207 6000
rect 265 -6000 325 6000
rect 383 -6000 443 6000
rect 501 -6000 561 6000
<< ndiff >>
rect -619 5988 -561 6000
rect -619 -5988 -607 5988
rect -573 -5988 -561 5988
rect -619 -6000 -561 -5988
rect -501 5988 -443 6000
rect -501 -5988 -489 5988
rect -455 -5988 -443 5988
rect -501 -6000 -443 -5988
rect -383 5988 -325 6000
rect -383 -5988 -371 5988
rect -337 -5988 -325 5988
rect -383 -6000 -325 -5988
rect -265 5988 -207 6000
rect -265 -5988 -253 5988
rect -219 -5988 -207 5988
rect -265 -6000 -207 -5988
rect -147 5988 -89 6000
rect -147 -5988 -135 5988
rect -101 -5988 -89 5988
rect -147 -6000 -89 -5988
rect -29 5988 29 6000
rect -29 -5988 -17 5988
rect 17 -5988 29 5988
rect -29 -6000 29 -5988
rect 89 5988 147 6000
rect 89 -5988 101 5988
rect 135 -5988 147 5988
rect 89 -6000 147 -5988
rect 207 5988 265 6000
rect 207 -5988 219 5988
rect 253 -5988 265 5988
rect 207 -6000 265 -5988
rect 325 5988 383 6000
rect 325 -5988 337 5988
rect 371 -5988 383 5988
rect 325 -6000 383 -5988
rect 443 5988 501 6000
rect 443 -5988 455 5988
rect 489 -5988 501 5988
rect 443 -6000 501 -5988
rect 561 5988 619 6000
rect 561 -5988 573 5988
rect 607 -5988 619 5988
rect 561 -6000 619 -5988
<< ndiffc >>
rect -607 -5988 -573 5988
rect -489 -5988 -455 5988
rect -371 -5988 -337 5988
rect -253 -5988 -219 5988
rect -135 -5988 -101 5988
rect -17 -5988 17 5988
rect 101 -5988 135 5988
rect 219 -5988 253 5988
rect 337 -5988 371 5988
rect 455 -5988 489 5988
rect 573 -5988 607 5988
<< poly >>
rect -564 6072 -498 6088
rect -564 6038 -548 6072
rect -514 6038 -498 6072
rect -564 6022 -498 6038
rect -446 6072 -380 6088
rect -446 6038 -430 6072
rect -396 6038 -380 6072
rect -446 6022 -380 6038
rect -328 6072 -262 6088
rect -328 6038 -312 6072
rect -278 6038 -262 6072
rect -328 6022 -262 6038
rect -210 6072 -144 6088
rect -210 6038 -194 6072
rect -160 6038 -144 6072
rect -210 6022 -144 6038
rect -92 6072 -26 6088
rect -92 6038 -76 6072
rect -42 6038 -26 6072
rect -92 6022 -26 6038
rect 26 6072 92 6088
rect 26 6038 42 6072
rect 76 6038 92 6072
rect 26 6022 92 6038
rect 144 6072 210 6088
rect 144 6038 160 6072
rect 194 6038 210 6072
rect 144 6022 210 6038
rect 262 6072 328 6088
rect 262 6038 278 6072
rect 312 6038 328 6072
rect 262 6022 328 6038
rect 380 6072 446 6088
rect 380 6038 396 6072
rect 430 6038 446 6072
rect 380 6022 446 6038
rect 498 6072 564 6088
rect 498 6038 514 6072
rect 548 6038 564 6072
rect 498 6022 564 6038
rect -561 6000 -501 6022
rect -443 6000 -383 6022
rect -325 6000 -265 6022
rect -207 6000 -147 6022
rect -89 6000 -29 6022
rect 29 6000 89 6022
rect 147 6000 207 6022
rect 265 6000 325 6022
rect 383 6000 443 6022
rect 501 6000 561 6022
rect -561 -6022 -501 -6000
rect -443 -6022 -383 -6000
rect -325 -6022 -265 -6000
rect -207 -6022 -147 -6000
rect -89 -6022 -29 -6000
rect 29 -6022 89 -6000
rect 147 -6022 207 -6000
rect 265 -6022 325 -6000
rect 383 -6022 443 -6000
rect 501 -6022 561 -6000
rect -564 -6032 -498 -6022
rect -446 -6032 -380 -6022
rect -328 -6032 -262 -6022
rect -210 -6032 -144 -6022
rect -92 -6032 -26 -6022
rect 26 -6032 92 -6022
rect 144 -6032 210 -6022
rect 262 -6032 328 -6022
rect 380 -6032 446 -6022
rect 498 -6032 564 -6022
rect -564 -6078 564 -6032
rect -564 -6088 -498 -6078
rect -446 -6088 -380 -6078
rect -328 -6088 -262 -6078
rect -210 -6088 -144 -6078
rect -92 -6088 -26 -6078
rect 26 -6088 92 -6078
rect 144 -6088 210 -6078
rect 262 -6088 328 -6078
rect 380 -6088 446 -6078
rect 498 -6088 564 -6078
<< polycont >>
rect -548 6038 -514 6072
rect -430 6038 -396 6072
rect -312 6038 -278 6072
rect -194 6038 -160 6072
rect -76 6038 -42 6072
rect 42 6038 76 6072
rect 160 6038 194 6072
rect 278 6038 312 6072
rect 396 6038 430 6072
rect 514 6038 548 6072
<< locali >>
rect -564 6038 -548 6072
rect -514 6038 -498 6072
rect -446 6038 -430 6072
rect -396 6038 -380 6072
rect -328 6038 -312 6072
rect -278 6038 -262 6072
rect -210 6038 -194 6072
rect -160 6038 -144 6072
rect -92 6038 -76 6072
rect -42 6038 -26 6072
rect 26 6038 42 6072
rect 76 6038 92 6072
rect 144 6038 160 6072
rect 194 6038 210 6072
rect 262 6038 278 6072
rect 312 6038 328 6072
rect 380 6038 396 6072
rect 430 6038 446 6072
rect 498 6038 514 6072
rect 548 6038 564 6072
rect -607 5988 -573 6004
rect -607 -6004 -573 -5988
rect -489 5988 -455 6004
rect -489 -6004 -455 -5988
rect -371 5988 -337 6004
rect -371 -6004 -337 -5988
rect -253 5988 -219 6004
rect -253 -6004 -219 -5988
rect -135 5988 -101 6004
rect -135 -6004 -101 -5988
rect -17 5988 17 6004
rect -17 -6004 17 -5988
rect 101 5988 135 6004
rect 101 -6004 135 -5988
rect 219 5988 253 6004
rect 219 -6004 253 -5988
rect 337 5988 371 6004
rect 337 -6004 371 -5988
rect 455 5988 489 6004
rect 455 -6004 489 -5988
rect 573 5988 607 6004
rect 573 -6004 607 -5988
<< viali >>
rect -548 6038 -514 6072
rect -430 6038 -396 6072
rect -312 6038 -278 6072
rect -194 6038 -160 6072
rect -76 6038 -42 6072
rect 42 6038 76 6072
rect 160 6038 194 6072
rect 278 6038 312 6072
rect 396 6038 430 6072
rect 514 6038 548 6072
rect -607 -5988 -573 5988
rect -489 -5988 -455 5988
rect -371 -5988 -337 5988
rect -253 -5988 -219 5988
rect -135 -5988 -101 5988
rect -17 -5988 17 5988
rect 101 -5988 135 5988
rect 219 -5988 253 5988
rect 337 -5988 371 5988
rect 455 -5988 489 5988
rect 573 -5988 607 5988
<< metal1 >>
rect -560 6072 -502 6078
rect -560 6038 -548 6072
rect -514 6038 -502 6072
rect -560 6032 -502 6038
rect -442 6072 -384 6078
rect -442 6038 -430 6072
rect -396 6038 -384 6072
rect -442 6032 -384 6038
rect -324 6072 -266 6078
rect -324 6038 -312 6072
rect -278 6038 -266 6072
rect -324 6032 -266 6038
rect -206 6072 -148 6078
rect -206 6038 -194 6072
rect -160 6038 -148 6072
rect -206 6032 -148 6038
rect -88 6072 -30 6078
rect -88 6038 -76 6072
rect -42 6038 -30 6072
rect -88 6032 -30 6038
rect 30 6072 88 6078
rect 30 6038 42 6072
rect 76 6038 88 6072
rect 30 6032 88 6038
rect 148 6072 206 6078
rect 148 6038 160 6072
rect 194 6038 206 6072
rect 148 6032 206 6038
rect 266 6072 324 6078
rect 266 6038 278 6072
rect 312 6038 324 6072
rect 266 6032 324 6038
rect 384 6072 442 6078
rect 384 6038 396 6072
rect 430 6038 442 6072
rect 384 6032 442 6038
rect 502 6072 560 6078
rect 502 6038 514 6072
rect 548 6038 560 6072
rect 502 6032 560 6038
rect -613 5988 -567 6000
rect -613 -5988 -607 5988
rect -573 -5988 -567 5988
rect -613 -6000 -567 -5988
rect -495 5988 -449 6000
rect -495 -5988 -489 5988
rect -455 -5988 -449 5988
rect -495 -6000 -449 -5988
rect -377 5988 -331 6000
rect -377 -5988 -371 5988
rect -337 -5988 -331 5988
rect -377 -6000 -331 -5988
rect -259 5988 -213 6000
rect -259 -5988 -253 5988
rect -219 -5988 -213 5988
rect -259 -6000 -213 -5988
rect -141 5988 -95 6000
rect -141 -5988 -135 5988
rect -101 -5988 -95 5988
rect -141 -6000 -95 -5988
rect -23 5988 23 6000
rect -23 -5988 -17 5988
rect 17 -5988 23 5988
rect -23 -6000 23 -5988
rect 95 5988 141 6000
rect 95 -5988 101 5988
rect 135 -5988 141 5988
rect 95 -6000 141 -5988
rect 213 5988 259 6000
rect 213 -5988 219 5988
rect 253 -5988 259 5988
rect 213 -6000 259 -5988
rect 331 5988 377 6000
rect 331 -5988 337 5988
rect 371 -5988 377 5988
rect 331 -6000 377 -5988
rect 449 5988 495 6000
rect 449 -5988 455 5988
rect 489 -5988 495 5988
rect 449 -6000 495 -5988
rect 567 5988 613 6000
rect 567 -5988 573 5988
rect 607 -5988 613 5988
rect 567 -6000 613 -5988
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 60 l 0.3 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
