magic
tech sky130A
magscale 1 2
timestamp 1667488624
<< error_p >>
rect 498 2394 556 2400
rect 498 2360 510 2394
rect 498 2354 556 2360
<< error_s >>
rect 352 1067 386 1085
rect 129 929 187 935
rect 129 895 141 929
rect 129 889 187 895
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1067
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__nfet_01v8_L9ESAD  XM3
timestamp 1667488624
transform 1 0 158 0 1 807
box -211 -260 211 260
use sky130_fd_pr__pfet_01v8_UGACMG  XM4
timestamp 1666901446
transform 1 0 527 0 1 1513
box -211 -1019 211 1019
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {}
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 CLK
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vin
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vout
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 CLKinverted
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Vdd!
port 5 nsew
<< end >>
