magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -35 1400 35 1832
rect -35 -1832 35 -1400
<< xpolyres >>
rect -35 -1400 35 1400
<< viali >>
rect -17 1778 17 1812
rect -17 1706 17 1740
rect -17 1634 17 1668
rect -17 1562 17 1596
rect -17 1490 17 1524
rect -17 1418 17 1452
rect -17 -1453 17 -1419
rect -17 -1525 17 -1491
rect -17 -1597 17 -1563
rect -17 -1669 17 -1635
rect -17 -1741 17 -1707
rect -17 -1813 17 -1779
<< metal1 >>
rect -25 1812 25 1826
rect -25 1778 -17 1812
rect 17 1778 25 1812
rect -25 1740 25 1778
rect -25 1706 -17 1740
rect 17 1706 25 1740
rect -25 1668 25 1706
rect -25 1634 -17 1668
rect 17 1634 25 1668
rect -25 1596 25 1634
rect -25 1562 -17 1596
rect 17 1562 25 1596
rect -25 1524 25 1562
rect -25 1490 -17 1524
rect 17 1490 25 1524
rect -25 1452 25 1490
rect -25 1418 -17 1452
rect 17 1418 25 1452
rect -25 1405 25 1418
rect -25 -1419 25 -1405
rect -25 -1453 -17 -1419
rect 17 -1453 25 -1419
rect -25 -1491 25 -1453
rect -25 -1525 -17 -1491
rect 17 -1525 25 -1491
rect -25 -1563 25 -1525
rect -25 -1597 -17 -1563
rect 17 -1597 25 -1563
rect -25 -1635 25 -1597
rect -25 -1669 -17 -1635
rect 17 -1669 25 -1635
rect -25 -1707 25 -1669
rect -25 -1741 -17 -1707
rect 17 -1741 25 -1707
rect -25 -1779 25 -1741
rect -25 -1813 -17 -1779
rect 17 -1813 25 -1779
rect -25 -1826 25 -1813
<< end >>
