magic
tech sky130A
magscale 1 2
timestamp 1666102132
<< nwell >>
rect -246 -12461 246 12461
<< pmos >>
rect -50 11242 50 12242
rect -50 10006 50 11006
rect -50 8770 50 9770
rect -50 7534 50 8534
rect -50 6298 50 7298
rect -50 5062 50 6062
rect -50 3826 50 4826
rect -50 2590 50 3590
rect -50 1354 50 2354
rect -50 118 50 1118
rect -50 -1118 50 -118
rect -50 -2354 50 -1354
rect -50 -3590 50 -2590
rect -50 -4826 50 -3826
rect -50 -6062 50 -5062
rect -50 -7298 50 -6298
rect -50 -8534 50 -7534
rect -50 -9770 50 -8770
rect -50 -11006 50 -10006
rect -50 -12242 50 -11242
<< pdiff >>
rect -108 12230 -50 12242
rect -108 11254 -96 12230
rect -62 11254 -50 12230
rect -108 11242 -50 11254
rect 50 12230 108 12242
rect 50 11254 62 12230
rect 96 11254 108 12230
rect 50 11242 108 11254
rect -108 10994 -50 11006
rect -108 10018 -96 10994
rect -62 10018 -50 10994
rect -108 10006 -50 10018
rect 50 10994 108 11006
rect 50 10018 62 10994
rect 96 10018 108 10994
rect 50 10006 108 10018
rect -108 9758 -50 9770
rect -108 8782 -96 9758
rect -62 8782 -50 9758
rect -108 8770 -50 8782
rect 50 9758 108 9770
rect 50 8782 62 9758
rect 96 8782 108 9758
rect 50 8770 108 8782
rect -108 8522 -50 8534
rect -108 7546 -96 8522
rect -62 7546 -50 8522
rect -108 7534 -50 7546
rect 50 8522 108 8534
rect 50 7546 62 8522
rect 96 7546 108 8522
rect 50 7534 108 7546
rect -108 7286 -50 7298
rect -108 6310 -96 7286
rect -62 6310 -50 7286
rect -108 6298 -50 6310
rect 50 7286 108 7298
rect 50 6310 62 7286
rect 96 6310 108 7286
rect 50 6298 108 6310
rect -108 6050 -50 6062
rect -108 5074 -96 6050
rect -62 5074 -50 6050
rect -108 5062 -50 5074
rect 50 6050 108 6062
rect 50 5074 62 6050
rect 96 5074 108 6050
rect 50 5062 108 5074
rect -108 4814 -50 4826
rect -108 3838 -96 4814
rect -62 3838 -50 4814
rect -108 3826 -50 3838
rect 50 4814 108 4826
rect 50 3838 62 4814
rect 96 3838 108 4814
rect 50 3826 108 3838
rect -108 3578 -50 3590
rect -108 2602 -96 3578
rect -62 2602 -50 3578
rect -108 2590 -50 2602
rect 50 3578 108 3590
rect 50 2602 62 3578
rect 96 2602 108 3578
rect 50 2590 108 2602
rect -108 2342 -50 2354
rect -108 1366 -96 2342
rect -62 1366 -50 2342
rect -108 1354 -50 1366
rect 50 2342 108 2354
rect 50 1366 62 2342
rect 96 1366 108 2342
rect 50 1354 108 1366
rect -108 1106 -50 1118
rect -108 130 -96 1106
rect -62 130 -50 1106
rect -108 118 -50 130
rect 50 1106 108 1118
rect 50 130 62 1106
rect 96 130 108 1106
rect 50 118 108 130
rect -108 -130 -50 -118
rect -108 -1106 -96 -130
rect -62 -1106 -50 -130
rect -108 -1118 -50 -1106
rect 50 -130 108 -118
rect 50 -1106 62 -130
rect 96 -1106 108 -130
rect 50 -1118 108 -1106
rect -108 -1366 -50 -1354
rect -108 -2342 -96 -1366
rect -62 -2342 -50 -1366
rect -108 -2354 -50 -2342
rect 50 -1366 108 -1354
rect 50 -2342 62 -1366
rect 96 -2342 108 -1366
rect 50 -2354 108 -2342
rect -108 -2602 -50 -2590
rect -108 -3578 -96 -2602
rect -62 -3578 -50 -2602
rect -108 -3590 -50 -3578
rect 50 -2602 108 -2590
rect 50 -3578 62 -2602
rect 96 -3578 108 -2602
rect 50 -3590 108 -3578
rect -108 -3838 -50 -3826
rect -108 -4814 -96 -3838
rect -62 -4814 -50 -3838
rect -108 -4826 -50 -4814
rect 50 -3838 108 -3826
rect 50 -4814 62 -3838
rect 96 -4814 108 -3838
rect 50 -4826 108 -4814
rect -108 -5074 -50 -5062
rect -108 -6050 -96 -5074
rect -62 -6050 -50 -5074
rect -108 -6062 -50 -6050
rect 50 -5074 108 -5062
rect 50 -6050 62 -5074
rect 96 -6050 108 -5074
rect 50 -6062 108 -6050
rect -108 -6310 -50 -6298
rect -108 -7286 -96 -6310
rect -62 -7286 -50 -6310
rect -108 -7298 -50 -7286
rect 50 -6310 108 -6298
rect 50 -7286 62 -6310
rect 96 -7286 108 -6310
rect 50 -7298 108 -7286
rect -108 -7546 -50 -7534
rect -108 -8522 -96 -7546
rect -62 -8522 -50 -7546
rect -108 -8534 -50 -8522
rect 50 -7546 108 -7534
rect 50 -8522 62 -7546
rect 96 -8522 108 -7546
rect 50 -8534 108 -8522
rect -108 -8782 -50 -8770
rect -108 -9758 -96 -8782
rect -62 -9758 -50 -8782
rect -108 -9770 -50 -9758
rect 50 -8782 108 -8770
rect 50 -9758 62 -8782
rect 96 -9758 108 -8782
rect 50 -9770 108 -9758
rect -108 -10018 -50 -10006
rect -108 -10994 -96 -10018
rect -62 -10994 -50 -10018
rect -108 -11006 -50 -10994
rect 50 -10018 108 -10006
rect 50 -10994 62 -10018
rect 96 -10994 108 -10018
rect 50 -11006 108 -10994
rect -108 -11254 -50 -11242
rect -108 -12230 -96 -11254
rect -62 -12230 -50 -11254
rect -108 -12242 -50 -12230
rect 50 -11254 108 -11242
rect 50 -12230 62 -11254
rect 96 -12230 108 -11254
rect 50 -12242 108 -12230
<< pdiffc >>
rect -96 11254 -62 12230
rect 62 11254 96 12230
rect -96 10018 -62 10994
rect 62 10018 96 10994
rect -96 8782 -62 9758
rect 62 8782 96 9758
rect -96 7546 -62 8522
rect 62 7546 96 8522
rect -96 6310 -62 7286
rect 62 6310 96 7286
rect -96 5074 -62 6050
rect 62 5074 96 6050
rect -96 3838 -62 4814
rect 62 3838 96 4814
rect -96 2602 -62 3578
rect 62 2602 96 3578
rect -96 1366 -62 2342
rect 62 1366 96 2342
rect -96 130 -62 1106
rect 62 130 96 1106
rect -96 -1106 -62 -130
rect 62 -1106 96 -130
rect -96 -2342 -62 -1366
rect 62 -2342 96 -1366
rect -96 -3578 -62 -2602
rect 62 -3578 96 -2602
rect -96 -4814 -62 -3838
rect 62 -4814 96 -3838
rect -96 -6050 -62 -5074
rect 62 -6050 96 -5074
rect -96 -7286 -62 -6310
rect 62 -7286 96 -6310
rect -96 -8522 -62 -7546
rect 62 -8522 96 -7546
rect -96 -9758 -62 -8782
rect 62 -9758 96 -8782
rect -96 -10994 -62 -10018
rect 62 -10994 96 -10018
rect -96 -12230 -62 -11254
rect 62 -12230 96 -11254
<< nsubdiff >>
rect -210 12391 -114 12425
rect 114 12391 210 12425
rect -210 12329 -176 12391
rect 176 12329 210 12391
rect -210 -12391 -176 -12329
rect 176 -12391 210 -12329
rect -210 -12425 -114 -12391
rect 114 -12425 210 -12391
<< nsubdiffcont >>
rect -114 12391 114 12425
rect -210 -12329 -176 12329
rect 176 -12329 210 12329
rect -114 -12425 114 -12391
<< poly >>
rect -50 12323 50 12339
rect -50 12289 -34 12323
rect 34 12289 50 12323
rect -50 12242 50 12289
rect -50 11195 50 11242
rect -50 11161 -34 11195
rect 34 11161 50 11195
rect -50 11145 50 11161
rect -50 11087 50 11103
rect -50 11053 -34 11087
rect 34 11053 50 11087
rect -50 11006 50 11053
rect -50 9959 50 10006
rect -50 9925 -34 9959
rect 34 9925 50 9959
rect -50 9909 50 9925
rect -50 9851 50 9867
rect -50 9817 -34 9851
rect 34 9817 50 9851
rect -50 9770 50 9817
rect -50 8723 50 8770
rect -50 8689 -34 8723
rect 34 8689 50 8723
rect -50 8673 50 8689
rect -50 8615 50 8631
rect -50 8581 -34 8615
rect 34 8581 50 8615
rect -50 8534 50 8581
rect -50 7487 50 7534
rect -50 7453 -34 7487
rect 34 7453 50 7487
rect -50 7437 50 7453
rect -50 7379 50 7395
rect -50 7345 -34 7379
rect 34 7345 50 7379
rect -50 7298 50 7345
rect -50 6251 50 6298
rect -50 6217 -34 6251
rect 34 6217 50 6251
rect -50 6201 50 6217
rect -50 6143 50 6159
rect -50 6109 -34 6143
rect 34 6109 50 6143
rect -50 6062 50 6109
rect -50 5015 50 5062
rect -50 4981 -34 5015
rect 34 4981 50 5015
rect -50 4965 50 4981
rect -50 4907 50 4923
rect -50 4873 -34 4907
rect 34 4873 50 4907
rect -50 4826 50 4873
rect -50 3779 50 3826
rect -50 3745 -34 3779
rect 34 3745 50 3779
rect -50 3729 50 3745
rect -50 3671 50 3687
rect -50 3637 -34 3671
rect 34 3637 50 3671
rect -50 3590 50 3637
rect -50 2543 50 2590
rect -50 2509 -34 2543
rect 34 2509 50 2543
rect -50 2493 50 2509
rect -50 2435 50 2451
rect -50 2401 -34 2435
rect 34 2401 50 2435
rect -50 2354 50 2401
rect -50 1307 50 1354
rect -50 1273 -34 1307
rect 34 1273 50 1307
rect -50 1257 50 1273
rect -50 1199 50 1215
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -50 1118 50 1165
rect -50 71 50 118
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -118 50 -71
rect -50 -1165 50 -1118
rect -50 -1199 -34 -1165
rect 34 -1199 50 -1165
rect -50 -1215 50 -1199
rect -50 -1273 50 -1257
rect -50 -1307 -34 -1273
rect 34 -1307 50 -1273
rect -50 -1354 50 -1307
rect -50 -2401 50 -2354
rect -50 -2435 -34 -2401
rect 34 -2435 50 -2401
rect -50 -2451 50 -2435
rect -50 -2509 50 -2493
rect -50 -2543 -34 -2509
rect 34 -2543 50 -2509
rect -50 -2590 50 -2543
rect -50 -3637 50 -3590
rect -50 -3671 -34 -3637
rect 34 -3671 50 -3637
rect -50 -3687 50 -3671
rect -50 -3745 50 -3729
rect -50 -3779 -34 -3745
rect 34 -3779 50 -3745
rect -50 -3826 50 -3779
rect -50 -4873 50 -4826
rect -50 -4907 -34 -4873
rect 34 -4907 50 -4873
rect -50 -4923 50 -4907
rect -50 -4981 50 -4965
rect -50 -5015 -34 -4981
rect 34 -5015 50 -4981
rect -50 -5062 50 -5015
rect -50 -6109 50 -6062
rect -50 -6143 -34 -6109
rect 34 -6143 50 -6109
rect -50 -6159 50 -6143
rect -50 -6217 50 -6201
rect -50 -6251 -34 -6217
rect 34 -6251 50 -6217
rect -50 -6298 50 -6251
rect -50 -7345 50 -7298
rect -50 -7379 -34 -7345
rect 34 -7379 50 -7345
rect -50 -7395 50 -7379
rect -50 -7453 50 -7437
rect -50 -7487 -34 -7453
rect 34 -7487 50 -7453
rect -50 -7534 50 -7487
rect -50 -8581 50 -8534
rect -50 -8615 -34 -8581
rect 34 -8615 50 -8581
rect -50 -8631 50 -8615
rect -50 -8689 50 -8673
rect -50 -8723 -34 -8689
rect 34 -8723 50 -8689
rect -50 -8770 50 -8723
rect -50 -9817 50 -9770
rect -50 -9851 -34 -9817
rect 34 -9851 50 -9817
rect -50 -9867 50 -9851
rect -50 -9925 50 -9909
rect -50 -9959 -34 -9925
rect 34 -9959 50 -9925
rect -50 -10006 50 -9959
rect -50 -11053 50 -11006
rect -50 -11087 -34 -11053
rect 34 -11087 50 -11053
rect -50 -11103 50 -11087
rect -50 -11161 50 -11145
rect -50 -11195 -34 -11161
rect 34 -11195 50 -11161
rect -50 -11242 50 -11195
rect -50 -12289 50 -12242
rect -50 -12323 -34 -12289
rect 34 -12323 50 -12289
rect -50 -12339 50 -12323
<< polycont >>
rect -34 12289 34 12323
rect -34 11161 34 11195
rect -34 11053 34 11087
rect -34 9925 34 9959
rect -34 9817 34 9851
rect -34 8689 34 8723
rect -34 8581 34 8615
rect -34 7453 34 7487
rect -34 7345 34 7379
rect -34 6217 34 6251
rect -34 6109 34 6143
rect -34 4981 34 5015
rect -34 4873 34 4907
rect -34 3745 34 3779
rect -34 3637 34 3671
rect -34 2509 34 2543
rect -34 2401 34 2435
rect -34 1273 34 1307
rect -34 1165 34 1199
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1199 34 -1165
rect -34 -1307 34 -1273
rect -34 -2435 34 -2401
rect -34 -2543 34 -2509
rect -34 -3671 34 -3637
rect -34 -3779 34 -3745
rect -34 -4907 34 -4873
rect -34 -5015 34 -4981
rect -34 -6143 34 -6109
rect -34 -6251 34 -6217
rect -34 -7379 34 -7345
rect -34 -7487 34 -7453
rect -34 -8615 34 -8581
rect -34 -8723 34 -8689
rect -34 -9851 34 -9817
rect -34 -9959 34 -9925
rect -34 -11087 34 -11053
rect -34 -11195 34 -11161
rect -34 -12323 34 -12289
<< locali >>
rect -210 12391 -114 12425
rect 114 12391 210 12425
rect -210 12329 -176 12391
rect 176 12329 210 12391
rect -50 12289 -34 12323
rect 34 12289 50 12323
rect -96 12230 -62 12246
rect -96 11238 -62 11254
rect 62 12230 96 12246
rect 62 11238 96 11254
rect -50 11161 -34 11195
rect 34 11161 50 11195
rect -50 11053 -34 11087
rect 34 11053 50 11087
rect -96 10994 -62 11010
rect -96 10002 -62 10018
rect 62 10994 96 11010
rect 62 10002 96 10018
rect -50 9925 -34 9959
rect 34 9925 50 9959
rect -50 9817 -34 9851
rect 34 9817 50 9851
rect -96 9758 -62 9774
rect -96 8766 -62 8782
rect 62 9758 96 9774
rect 62 8766 96 8782
rect -50 8689 -34 8723
rect 34 8689 50 8723
rect -50 8581 -34 8615
rect 34 8581 50 8615
rect -96 8522 -62 8538
rect -96 7530 -62 7546
rect 62 8522 96 8538
rect 62 7530 96 7546
rect -50 7453 -34 7487
rect 34 7453 50 7487
rect -50 7345 -34 7379
rect 34 7345 50 7379
rect -96 7286 -62 7302
rect -96 6294 -62 6310
rect 62 7286 96 7302
rect 62 6294 96 6310
rect -50 6217 -34 6251
rect 34 6217 50 6251
rect -50 6109 -34 6143
rect 34 6109 50 6143
rect -96 6050 -62 6066
rect -96 5058 -62 5074
rect 62 6050 96 6066
rect 62 5058 96 5074
rect -50 4981 -34 5015
rect 34 4981 50 5015
rect -50 4873 -34 4907
rect 34 4873 50 4907
rect -96 4814 -62 4830
rect -96 3822 -62 3838
rect 62 4814 96 4830
rect 62 3822 96 3838
rect -50 3745 -34 3779
rect 34 3745 50 3779
rect -50 3637 -34 3671
rect 34 3637 50 3671
rect -96 3578 -62 3594
rect -96 2586 -62 2602
rect 62 3578 96 3594
rect 62 2586 96 2602
rect -50 2509 -34 2543
rect 34 2509 50 2543
rect -50 2401 -34 2435
rect 34 2401 50 2435
rect -96 2342 -62 2358
rect -96 1350 -62 1366
rect 62 2342 96 2358
rect 62 1350 96 1366
rect -50 1273 -34 1307
rect 34 1273 50 1307
rect -50 1165 -34 1199
rect 34 1165 50 1199
rect -96 1106 -62 1122
rect -96 114 -62 130
rect 62 1106 96 1122
rect 62 114 96 130
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -130 -62 -114
rect -96 -1122 -62 -1106
rect 62 -130 96 -114
rect 62 -1122 96 -1106
rect -50 -1199 -34 -1165
rect 34 -1199 50 -1165
rect -50 -1307 -34 -1273
rect 34 -1307 50 -1273
rect -96 -1366 -62 -1350
rect -96 -2358 -62 -2342
rect 62 -1366 96 -1350
rect 62 -2358 96 -2342
rect -50 -2435 -34 -2401
rect 34 -2435 50 -2401
rect -50 -2543 -34 -2509
rect 34 -2543 50 -2509
rect -96 -2602 -62 -2586
rect -96 -3594 -62 -3578
rect 62 -2602 96 -2586
rect 62 -3594 96 -3578
rect -50 -3671 -34 -3637
rect 34 -3671 50 -3637
rect -50 -3779 -34 -3745
rect 34 -3779 50 -3745
rect -96 -3838 -62 -3822
rect -96 -4830 -62 -4814
rect 62 -3838 96 -3822
rect 62 -4830 96 -4814
rect -50 -4907 -34 -4873
rect 34 -4907 50 -4873
rect -50 -5015 -34 -4981
rect 34 -5015 50 -4981
rect -96 -5074 -62 -5058
rect -96 -6066 -62 -6050
rect 62 -5074 96 -5058
rect 62 -6066 96 -6050
rect -50 -6143 -34 -6109
rect 34 -6143 50 -6109
rect -50 -6251 -34 -6217
rect 34 -6251 50 -6217
rect -96 -6310 -62 -6294
rect -96 -7302 -62 -7286
rect 62 -6310 96 -6294
rect 62 -7302 96 -7286
rect -50 -7379 -34 -7345
rect 34 -7379 50 -7345
rect -50 -7487 -34 -7453
rect 34 -7487 50 -7453
rect -96 -7546 -62 -7530
rect -96 -8538 -62 -8522
rect 62 -7546 96 -7530
rect 62 -8538 96 -8522
rect -50 -8615 -34 -8581
rect 34 -8615 50 -8581
rect -50 -8723 -34 -8689
rect 34 -8723 50 -8689
rect -96 -8782 -62 -8766
rect -96 -9774 -62 -9758
rect 62 -8782 96 -8766
rect 62 -9774 96 -9758
rect -50 -9851 -34 -9817
rect 34 -9851 50 -9817
rect -50 -9959 -34 -9925
rect 34 -9959 50 -9925
rect -96 -10018 -62 -10002
rect -96 -11010 -62 -10994
rect 62 -10018 96 -10002
rect 62 -11010 96 -10994
rect -50 -11087 -34 -11053
rect 34 -11087 50 -11053
rect -50 -11195 -34 -11161
rect 34 -11195 50 -11161
rect -96 -11254 -62 -11238
rect -96 -12246 -62 -12230
rect 62 -11254 96 -11238
rect 62 -12246 96 -12230
rect -50 -12323 -34 -12289
rect 34 -12323 50 -12289
rect -210 -12391 -176 -12329
rect 176 -12391 210 -12329
rect -210 -12425 -114 -12391
rect 114 -12425 210 -12391
<< viali >>
rect -34 12289 34 12323
rect -96 11254 -62 12230
rect 62 11254 96 12230
rect -34 11161 34 11195
rect -34 11053 34 11087
rect -96 10018 -62 10994
rect 62 10018 96 10994
rect -34 9925 34 9959
rect -34 9817 34 9851
rect -96 8782 -62 9758
rect 62 8782 96 9758
rect -34 8689 34 8723
rect -34 8581 34 8615
rect -96 7546 -62 8522
rect 62 7546 96 8522
rect -34 7453 34 7487
rect -34 7345 34 7379
rect -96 6310 -62 7286
rect 62 6310 96 7286
rect -34 6217 34 6251
rect -34 6109 34 6143
rect -96 5074 -62 6050
rect 62 5074 96 6050
rect -34 4981 34 5015
rect -34 4873 34 4907
rect -96 3838 -62 4814
rect 62 3838 96 4814
rect -34 3745 34 3779
rect -34 3637 34 3671
rect -96 2602 -62 3578
rect 62 2602 96 3578
rect -34 2509 34 2543
rect -34 2401 34 2435
rect -96 1366 -62 2342
rect 62 1366 96 2342
rect -34 1273 34 1307
rect -34 1165 34 1199
rect -96 130 -62 1106
rect 62 130 96 1106
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1106 -62 -130
rect 62 -1106 96 -130
rect -34 -1199 34 -1165
rect -34 -1307 34 -1273
rect -96 -2342 -62 -1366
rect 62 -2342 96 -1366
rect -34 -2435 34 -2401
rect -34 -2543 34 -2509
rect -96 -3578 -62 -2602
rect 62 -3578 96 -2602
rect -34 -3671 34 -3637
rect -34 -3779 34 -3745
rect -96 -4814 -62 -3838
rect 62 -4814 96 -3838
rect -34 -4907 34 -4873
rect -34 -5015 34 -4981
rect -96 -6050 -62 -5074
rect 62 -6050 96 -5074
rect -34 -6143 34 -6109
rect -34 -6251 34 -6217
rect -96 -7286 -62 -6310
rect 62 -7286 96 -6310
rect -34 -7379 34 -7345
rect -34 -7487 34 -7453
rect -96 -8522 -62 -7546
rect 62 -8522 96 -7546
rect -34 -8615 34 -8581
rect -34 -8723 34 -8689
rect -96 -9758 -62 -8782
rect 62 -9758 96 -8782
rect -34 -9851 34 -9817
rect -34 -9959 34 -9925
rect -96 -10994 -62 -10018
rect 62 -10994 96 -10018
rect -34 -11087 34 -11053
rect -34 -11195 34 -11161
rect -96 -12230 -62 -11254
rect 62 -12230 96 -11254
rect -34 -12323 34 -12289
<< metal1 >>
rect -46 12323 46 12329
rect -46 12289 -34 12323
rect 34 12289 46 12323
rect -46 12283 46 12289
rect -102 12230 -56 12242
rect -102 11254 -96 12230
rect -62 11254 -56 12230
rect -102 11242 -56 11254
rect 56 12230 102 12242
rect 56 11254 62 12230
rect 96 11254 102 12230
rect 56 11242 102 11254
rect -46 11195 46 11201
rect -46 11161 -34 11195
rect 34 11161 46 11195
rect -46 11155 46 11161
rect -46 11087 46 11093
rect -46 11053 -34 11087
rect 34 11053 46 11087
rect -46 11047 46 11053
rect -102 10994 -56 11006
rect -102 10018 -96 10994
rect -62 10018 -56 10994
rect -102 10006 -56 10018
rect 56 10994 102 11006
rect 56 10018 62 10994
rect 96 10018 102 10994
rect 56 10006 102 10018
rect -46 9959 46 9965
rect -46 9925 -34 9959
rect 34 9925 46 9959
rect -46 9919 46 9925
rect -46 9851 46 9857
rect -46 9817 -34 9851
rect 34 9817 46 9851
rect -46 9811 46 9817
rect -102 9758 -56 9770
rect -102 8782 -96 9758
rect -62 8782 -56 9758
rect -102 8770 -56 8782
rect 56 9758 102 9770
rect 56 8782 62 9758
rect 96 8782 102 9758
rect 56 8770 102 8782
rect -46 8723 46 8729
rect -46 8689 -34 8723
rect 34 8689 46 8723
rect -46 8683 46 8689
rect -46 8615 46 8621
rect -46 8581 -34 8615
rect 34 8581 46 8615
rect -46 8575 46 8581
rect -102 8522 -56 8534
rect -102 7546 -96 8522
rect -62 7546 -56 8522
rect -102 7534 -56 7546
rect 56 8522 102 8534
rect 56 7546 62 8522
rect 96 7546 102 8522
rect 56 7534 102 7546
rect -46 7487 46 7493
rect -46 7453 -34 7487
rect 34 7453 46 7487
rect -46 7447 46 7453
rect -46 7379 46 7385
rect -46 7345 -34 7379
rect 34 7345 46 7379
rect -46 7339 46 7345
rect -102 7286 -56 7298
rect -102 6310 -96 7286
rect -62 6310 -56 7286
rect -102 6298 -56 6310
rect 56 7286 102 7298
rect 56 6310 62 7286
rect 96 6310 102 7286
rect 56 6298 102 6310
rect -46 6251 46 6257
rect -46 6217 -34 6251
rect 34 6217 46 6251
rect -46 6211 46 6217
rect -46 6143 46 6149
rect -46 6109 -34 6143
rect 34 6109 46 6143
rect -46 6103 46 6109
rect -102 6050 -56 6062
rect -102 5074 -96 6050
rect -62 5074 -56 6050
rect -102 5062 -56 5074
rect 56 6050 102 6062
rect 56 5074 62 6050
rect 96 5074 102 6050
rect 56 5062 102 5074
rect -46 5015 46 5021
rect -46 4981 -34 5015
rect 34 4981 46 5015
rect -46 4975 46 4981
rect -46 4907 46 4913
rect -46 4873 -34 4907
rect 34 4873 46 4907
rect -46 4867 46 4873
rect -102 4814 -56 4826
rect -102 3838 -96 4814
rect -62 3838 -56 4814
rect -102 3826 -56 3838
rect 56 4814 102 4826
rect 56 3838 62 4814
rect 96 3838 102 4814
rect 56 3826 102 3838
rect -46 3779 46 3785
rect -46 3745 -34 3779
rect 34 3745 46 3779
rect -46 3739 46 3745
rect -46 3671 46 3677
rect -46 3637 -34 3671
rect 34 3637 46 3671
rect -46 3631 46 3637
rect -102 3578 -56 3590
rect -102 2602 -96 3578
rect -62 2602 -56 3578
rect -102 2590 -56 2602
rect 56 3578 102 3590
rect 56 2602 62 3578
rect 96 2602 102 3578
rect 56 2590 102 2602
rect -46 2543 46 2549
rect -46 2509 -34 2543
rect 34 2509 46 2543
rect -46 2503 46 2509
rect -46 2435 46 2441
rect -46 2401 -34 2435
rect 34 2401 46 2435
rect -46 2395 46 2401
rect -102 2342 -56 2354
rect -102 1366 -96 2342
rect -62 1366 -56 2342
rect -102 1354 -56 1366
rect 56 2342 102 2354
rect 56 1366 62 2342
rect 96 1366 102 2342
rect 56 1354 102 1366
rect -46 1307 46 1313
rect -46 1273 -34 1307
rect 34 1273 46 1307
rect -46 1267 46 1273
rect -46 1199 46 1205
rect -46 1165 -34 1199
rect 34 1165 46 1199
rect -46 1159 46 1165
rect -102 1106 -56 1118
rect -102 130 -96 1106
rect -62 130 -56 1106
rect -102 118 -56 130
rect 56 1106 102 1118
rect 56 130 62 1106
rect 96 130 102 1106
rect 56 118 102 130
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -130 -56 -118
rect -102 -1106 -96 -130
rect -62 -1106 -56 -130
rect -102 -1118 -56 -1106
rect 56 -130 102 -118
rect 56 -1106 62 -130
rect 96 -1106 102 -130
rect 56 -1118 102 -1106
rect -46 -1165 46 -1159
rect -46 -1199 -34 -1165
rect 34 -1199 46 -1165
rect -46 -1205 46 -1199
rect -46 -1273 46 -1267
rect -46 -1307 -34 -1273
rect 34 -1307 46 -1273
rect -46 -1313 46 -1307
rect -102 -1366 -56 -1354
rect -102 -2342 -96 -1366
rect -62 -2342 -56 -1366
rect -102 -2354 -56 -2342
rect 56 -1366 102 -1354
rect 56 -2342 62 -1366
rect 96 -2342 102 -1366
rect 56 -2354 102 -2342
rect -46 -2401 46 -2395
rect -46 -2435 -34 -2401
rect 34 -2435 46 -2401
rect -46 -2441 46 -2435
rect -46 -2509 46 -2503
rect -46 -2543 -34 -2509
rect 34 -2543 46 -2509
rect -46 -2549 46 -2543
rect -102 -2602 -56 -2590
rect -102 -3578 -96 -2602
rect -62 -3578 -56 -2602
rect -102 -3590 -56 -3578
rect 56 -2602 102 -2590
rect 56 -3578 62 -2602
rect 96 -3578 102 -2602
rect 56 -3590 102 -3578
rect -46 -3637 46 -3631
rect -46 -3671 -34 -3637
rect 34 -3671 46 -3637
rect -46 -3677 46 -3671
rect -46 -3745 46 -3739
rect -46 -3779 -34 -3745
rect 34 -3779 46 -3745
rect -46 -3785 46 -3779
rect -102 -3838 -56 -3826
rect -102 -4814 -96 -3838
rect -62 -4814 -56 -3838
rect -102 -4826 -56 -4814
rect 56 -3838 102 -3826
rect 56 -4814 62 -3838
rect 96 -4814 102 -3838
rect 56 -4826 102 -4814
rect -46 -4873 46 -4867
rect -46 -4907 -34 -4873
rect 34 -4907 46 -4873
rect -46 -4913 46 -4907
rect -46 -4981 46 -4975
rect -46 -5015 -34 -4981
rect 34 -5015 46 -4981
rect -46 -5021 46 -5015
rect -102 -5074 -56 -5062
rect -102 -6050 -96 -5074
rect -62 -6050 -56 -5074
rect -102 -6062 -56 -6050
rect 56 -5074 102 -5062
rect 56 -6050 62 -5074
rect 96 -6050 102 -5074
rect 56 -6062 102 -6050
rect -46 -6109 46 -6103
rect -46 -6143 -34 -6109
rect 34 -6143 46 -6109
rect -46 -6149 46 -6143
rect -46 -6217 46 -6211
rect -46 -6251 -34 -6217
rect 34 -6251 46 -6217
rect -46 -6257 46 -6251
rect -102 -6310 -56 -6298
rect -102 -7286 -96 -6310
rect -62 -7286 -56 -6310
rect -102 -7298 -56 -7286
rect 56 -6310 102 -6298
rect 56 -7286 62 -6310
rect 96 -7286 102 -6310
rect 56 -7298 102 -7286
rect -46 -7345 46 -7339
rect -46 -7379 -34 -7345
rect 34 -7379 46 -7345
rect -46 -7385 46 -7379
rect -46 -7453 46 -7447
rect -46 -7487 -34 -7453
rect 34 -7487 46 -7453
rect -46 -7493 46 -7487
rect -102 -7546 -56 -7534
rect -102 -8522 -96 -7546
rect -62 -8522 -56 -7546
rect -102 -8534 -56 -8522
rect 56 -7546 102 -7534
rect 56 -8522 62 -7546
rect 96 -8522 102 -7546
rect 56 -8534 102 -8522
rect -46 -8581 46 -8575
rect -46 -8615 -34 -8581
rect 34 -8615 46 -8581
rect -46 -8621 46 -8615
rect -46 -8689 46 -8683
rect -46 -8723 -34 -8689
rect 34 -8723 46 -8689
rect -46 -8729 46 -8723
rect -102 -8782 -56 -8770
rect -102 -9758 -96 -8782
rect -62 -9758 -56 -8782
rect -102 -9770 -56 -9758
rect 56 -8782 102 -8770
rect 56 -9758 62 -8782
rect 96 -9758 102 -8782
rect 56 -9770 102 -9758
rect -46 -9817 46 -9811
rect -46 -9851 -34 -9817
rect 34 -9851 46 -9817
rect -46 -9857 46 -9851
rect -46 -9925 46 -9919
rect -46 -9959 -34 -9925
rect 34 -9959 46 -9925
rect -46 -9965 46 -9959
rect -102 -10018 -56 -10006
rect -102 -10994 -96 -10018
rect -62 -10994 -56 -10018
rect -102 -11006 -56 -10994
rect 56 -10018 102 -10006
rect 56 -10994 62 -10018
rect 96 -10994 102 -10018
rect 56 -11006 102 -10994
rect -46 -11053 46 -11047
rect -46 -11087 -34 -11053
rect 34 -11087 46 -11053
rect -46 -11093 46 -11087
rect -46 -11161 46 -11155
rect -46 -11195 -34 -11161
rect 34 -11195 46 -11161
rect -46 -11201 46 -11195
rect -102 -11254 -56 -11242
rect -102 -12230 -96 -11254
rect -62 -12230 -56 -11254
rect -102 -12242 -56 -12230
rect 56 -11254 102 -11242
rect 56 -12230 62 -11254
rect 96 -12230 102 -11254
rect 56 -12242 102 -12230
rect -46 -12289 46 -12283
rect -46 -12323 -34 -12289
rect 34 -12323 46 -12289
rect -46 -12329 46 -12323
<< properties >>
string FIXED_BBOX -193 -12408 193 12408
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
