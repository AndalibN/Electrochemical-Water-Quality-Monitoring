magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect 173 68 787 2165
<< metal1 >>
rect 481 2534 547 2594
rect 396 2479 462 2507
rect 396 2427 403 2479
rect 455 2427 462 2479
rect 396 2402 462 2427
rect 494 2480 560 2506
rect 494 2428 499 2480
rect 551 2428 560 2480
rect 494 2402 560 2428
rect 395 1929 461 1967
rect 395 1877 404 1929
rect 456 1877 461 1929
rect 395 1865 461 1877
rect 395 1813 404 1865
rect 456 1813 461 1865
rect 395 1801 461 1813
rect 395 1749 404 1801
rect 456 1749 461 1801
rect 395 1737 461 1749
rect 395 1685 404 1737
rect 456 1685 461 1737
rect 395 1673 461 1685
rect 395 1621 404 1673
rect 456 1621 461 1673
rect 395 1609 461 1621
rect 395 1557 404 1609
rect 456 1557 461 1609
rect 395 1545 461 1557
rect 395 1493 404 1545
rect 456 1493 461 1545
rect 395 1481 461 1493
rect 395 1429 404 1481
rect 456 1429 461 1481
rect 395 1417 461 1429
rect 395 1365 404 1417
rect 456 1365 461 1417
rect 395 1353 461 1365
rect 395 1301 404 1353
rect 456 1301 461 1353
rect 395 1289 461 1301
rect 395 1237 404 1289
rect 456 1237 461 1289
rect 395 1225 461 1237
rect 395 1173 404 1225
rect 456 1173 461 1225
rect 395 1161 461 1173
rect 395 1109 404 1161
rect 456 1109 461 1161
rect 395 1097 461 1109
rect 395 1045 404 1097
rect 456 1045 461 1097
rect 395 1033 461 1045
rect 395 981 404 1033
rect 456 981 461 1033
rect 395 969 461 981
rect 395 917 404 969
rect 456 917 461 969
rect 395 905 461 917
rect 395 853 404 905
rect 456 853 461 905
rect 395 841 461 853
rect 395 789 404 841
rect 456 789 461 841
rect 395 777 461 789
rect 395 725 404 777
rect 456 725 461 777
rect 395 713 461 725
rect 395 661 404 713
rect 456 661 461 713
rect 395 649 461 661
rect 395 597 404 649
rect 456 597 461 649
rect 395 585 461 597
rect 395 533 404 585
rect 456 533 461 585
rect 395 521 461 533
rect 395 469 404 521
rect 456 469 461 521
rect 395 457 461 469
rect 395 405 404 457
rect 456 405 461 457
rect 395 367 461 405
rect 494 1928 560 1967
rect 494 1876 500 1928
rect 552 1876 560 1928
rect 494 1864 560 1876
rect 494 1812 500 1864
rect 552 1812 560 1864
rect 494 1800 560 1812
rect 494 1748 500 1800
rect 552 1748 560 1800
rect 494 1736 560 1748
rect 494 1684 500 1736
rect 552 1684 560 1736
rect 494 1672 560 1684
rect 494 1620 500 1672
rect 552 1620 560 1672
rect 494 1608 560 1620
rect 494 1556 500 1608
rect 552 1556 560 1608
rect 494 1544 560 1556
rect 494 1492 500 1544
rect 552 1492 560 1544
rect 494 1480 560 1492
rect 494 1428 500 1480
rect 552 1428 560 1480
rect 494 1416 560 1428
rect 494 1364 500 1416
rect 552 1364 560 1416
rect 494 1352 560 1364
rect 494 1300 500 1352
rect 552 1300 560 1352
rect 494 1288 560 1300
rect 494 1236 500 1288
rect 552 1236 560 1288
rect 494 1224 560 1236
rect 494 1172 500 1224
rect 552 1172 560 1224
rect 494 1160 560 1172
rect 494 1108 500 1160
rect 552 1108 560 1160
rect 494 1096 560 1108
rect 494 1044 500 1096
rect 552 1044 560 1096
rect 494 1032 560 1044
rect 494 980 500 1032
rect 552 980 560 1032
rect 494 968 560 980
rect 494 916 500 968
rect 552 916 560 968
rect 494 904 560 916
rect 494 852 500 904
rect 552 852 560 904
rect 494 840 560 852
rect 494 788 500 840
rect 552 788 560 840
rect 494 776 560 788
rect 494 724 500 776
rect 552 724 560 776
rect 494 712 560 724
rect 494 660 500 712
rect 552 660 560 712
rect 494 648 560 660
rect 494 596 500 648
rect 552 596 560 648
rect 494 584 560 596
rect 494 532 500 584
rect 552 532 560 584
rect 494 520 560 532
rect 494 468 500 520
rect 552 468 560 520
rect 494 456 560 468
rect 494 404 500 456
rect 552 404 560 456
rect 494 367 560 404
rect 445 270 511 329
<< via1 >>
rect 403 2427 455 2479
rect 499 2428 551 2480
rect 404 1877 456 1929
rect 404 1813 456 1865
rect 404 1749 456 1801
rect 404 1685 456 1737
rect 404 1621 456 1673
rect 404 1557 456 1609
rect 404 1493 456 1545
rect 404 1429 456 1481
rect 404 1365 456 1417
rect 404 1301 456 1353
rect 404 1237 456 1289
rect 404 1173 456 1225
rect 404 1109 456 1161
rect 404 1045 456 1097
rect 404 981 456 1033
rect 404 917 456 969
rect 404 853 456 905
rect 404 789 456 841
rect 404 725 456 777
rect 404 661 456 713
rect 404 597 456 649
rect 404 533 456 585
rect 404 469 456 521
rect 404 405 456 457
rect 500 1876 552 1928
rect 500 1812 552 1864
rect 500 1748 552 1800
rect 500 1684 552 1736
rect 500 1620 552 1672
rect 500 1556 552 1608
rect 500 1492 552 1544
rect 500 1428 552 1480
rect 500 1364 552 1416
rect 500 1300 552 1352
rect 500 1236 552 1288
rect 500 1172 552 1224
rect 500 1108 552 1160
rect 500 1044 552 1096
rect 500 980 552 1032
rect 500 916 552 968
rect 500 852 552 904
rect 500 788 552 840
rect 500 724 552 776
rect 500 660 552 712
rect 500 596 552 648
rect 500 532 552 584
rect 500 468 552 520
rect 500 404 552 456
<< metal2 >>
rect 396 2479 462 2507
rect 396 2427 403 2479
rect 455 2427 462 2479
rect 396 1929 462 2427
rect 396 1877 404 1929
rect 456 1877 462 1929
rect 396 1865 462 1877
rect 396 1813 404 1865
rect 456 1813 462 1865
rect 396 1801 462 1813
rect 396 1749 404 1801
rect 456 1749 462 1801
rect 396 1737 462 1749
rect 396 1685 404 1737
rect 456 1685 462 1737
rect 396 1673 462 1685
rect 396 1621 404 1673
rect 456 1621 462 1673
rect 396 1609 462 1621
rect 396 1557 404 1609
rect 456 1557 462 1609
rect 396 1545 462 1557
rect 396 1493 404 1545
rect 456 1493 462 1545
rect 396 1481 462 1493
rect 396 1429 404 1481
rect 456 1429 462 1481
rect 396 1417 462 1429
rect 396 1365 404 1417
rect 456 1365 462 1417
rect 396 1353 462 1365
rect 396 1301 404 1353
rect 456 1301 462 1353
rect 396 1289 462 1301
rect 396 1237 404 1289
rect 456 1237 462 1289
rect 396 1225 462 1237
rect 396 1173 404 1225
rect 456 1173 462 1225
rect 396 1161 462 1173
rect 396 1109 404 1161
rect 456 1109 462 1161
rect 396 1097 462 1109
rect 396 1045 404 1097
rect 456 1045 462 1097
rect 396 1033 462 1045
rect 396 981 404 1033
rect 456 981 462 1033
rect 396 969 462 981
rect 396 917 404 969
rect 456 917 462 969
rect 396 905 462 917
rect 396 853 404 905
rect 456 853 462 905
rect 396 841 462 853
rect 396 789 404 841
rect 456 789 462 841
rect 396 777 462 789
rect 396 725 404 777
rect 456 725 462 777
rect 396 713 462 725
rect 396 661 404 713
rect 456 661 462 713
rect 396 649 462 661
rect 396 597 404 649
rect 456 597 462 649
rect 396 585 462 597
rect 396 533 404 585
rect 456 533 462 585
rect 396 521 462 533
rect 396 469 404 521
rect 456 469 462 521
rect 396 457 462 469
rect 396 405 404 457
rect 456 405 462 457
rect 396 367 462 405
rect 494 2480 560 2507
rect 494 2428 499 2480
rect 551 2428 560 2480
rect 494 1928 560 2428
rect 494 1876 500 1928
rect 552 1876 560 1928
rect 494 1864 560 1876
rect 494 1812 500 1864
rect 552 1812 560 1864
rect 494 1800 560 1812
rect 494 1748 500 1800
rect 552 1748 560 1800
rect 494 1736 560 1748
rect 494 1684 500 1736
rect 552 1684 560 1736
rect 494 1672 560 1684
rect 494 1620 500 1672
rect 552 1620 560 1672
rect 494 1608 560 1620
rect 494 1556 500 1608
rect 552 1556 560 1608
rect 494 1544 560 1556
rect 494 1492 500 1544
rect 552 1492 560 1544
rect 494 1480 560 1492
rect 494 1428 500 1480
rect 552 1428 560 1480
rect 494 1416 560 1428
rect 494 1364 500 1416
rect 552 1364 560 1416
rect 494 1352 560 1364
rect 494 1300 500 1352
rect 552 1300 560 1352
rect 494 1288 560 1300
rect 494 1236 500 1288
rect 552 1236 560 1288
rect 494 1224 560 1236
rect 494 1172 500 1224
rect 552 1172 560 1224
rect 494 1160 560 1172
rect 494 1108 500 1160
rect 552 1108 560 1160
rect 494 1096 560 1108
rect 494 1044 500 1096
rect 552 1044 560 1096
rect 494 1032 560 1044
rect 494 980 500 1032
rect 552 980 560 1032
rect 494 968 560 980
rect 494 916 500 968
rect 552 916 560 968
rect 494 904 560 916
rect 494 852 500 904
rect 552 852 560 904
rect 494 840 560 852
rect 494 788 500 840
rect 552 788 560 840
rect 494 776 560 788
rect 494 724 500 776
rect 552 724 560 776
rect 494 712 560 724
rect 494 660 500 712
rect 552 660 560 712
rect 494 648 560 660
rect 494 596 500 648
rect 552 596 560 648
rect 494 584 560 596
rect 494 532 500 584
rect 552 532 560 584
rect 494 520 560 532
rect 494 468 500 520
rect 552 468 560 520
rect 494 456 560 468
rect 494 404 500 456
rect 552 404 560 456
rect 494 367 560 404
use sky130_fd_pr__nfet_01v8_JBX99N  XM3
timestamp 1669522153
transform 1 0 478 0 1 2487
box -99 -107 99 107
use sky130_fd_pr__pfet_01v8_MGSTUG  XM4
timestamp 1669522153
transform 1 0 478 0 1 1131
box -109 -864 109 898
<< labels >>
rlabel metal1 s 472 296 472 296 4 CLKinverted
port 1 nsew
rlabel metal1 s 508 2564 508 2564 4 CLK
port 2 nsew
rlabel metal2 s 418 2180 418 2180 4 Vin
port 3 nsew
rlabel metal2 s 530 2180 530 2180 4 Vout
port 4 nsew
<< end >>
