magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -173 -326 173 326
<< nmos >>
rect -89 -300 -29 300
rect 29 -300 89 300
<< ndiff >>
rect -147 255 -89 300
rect -147 221 -135 255
rect -101 221 -89 255
rect -147 187 -89 221
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -221 -89 -187
rect -147 -255 -135 -221
rect -101 -255 -89 -221
rect -147 -300 -89 -255
rect -29 255 29 300
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -300 29 -255
rect 89 255 147 300
rect 89 221 101 255
rect 135 221 147 255
rect 89 187 147 221
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -221 147 -187
rect 89 -255 101 -221
rect 135 -255 147 -221
rect 89 -300 147 -255
<< ndiffc >>
rect -135 221 -101 255
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -135 -255 -101 -221
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect 101 221 135 255
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 101 -255 135 -221
<< poly >>
rect -89 323 89 369
rect -89 300 -29 323
rect 29 300 89 323
rect -89 -326 -29 -300
rect 29 -326 89 -300
<< locali >>
rect -135 269 -101 304
rect -135 197 -101 221
rect -135 125 -101 153
rect -135 53 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -53
rect -135 -153 -101 -125
rect -135 -221 -101 -197
rect -135 -304 -101 -269
rect -17 269 17 304
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -304 17 -269
rect 101 269 135 304
rect 101 197 135 221
rect 101 125 135 153
rect 101 53 135 85
rect 101 -17 135 17
rect 101 -85 135 -53
rect 101 -153 135 -125
rect 101 -221 135 -197
rect 101 -304 135 -269
<< viali >>
rect -135 255 -101 269
rect -135 235 -101 255
rect -135 187 -101 197
rect -135 163 -101 187
rect -135 119 -101 125
rect -135 91 -101 119
rect -135 51 -101 53
rect -135 19 -101 51
rect -135 -51 -101 -19
rect -135 -53 -101 -51
rect -135 -119 -101 -91
rect -135 -125 -101 -119
rect -135 -187 -101 -163
rect -135 -197 -101 -187
rect -135 -255 -101 -235
rect -135 -269 -101 -255
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect 101 255 135 269
rect 101 235 135 255
rect 101 187 135 197
rect 101 163 135 187
rect 101 119 135 125
rect 101 91 135 119
rect 101 51 135 53
rect 101 19 135 51
rect 101 -51 135 -19
rect 101 -53 135 -51
rect 101 -119 135 -91
rect 101 -125 135 -119
rect 101 -187 135 -163
rect 101 -197 135 -187
rect 101 -255 135 -235
rect 101 -269 135 -255
<< metal1 >>
rect -141 269 -95 300
rect -141 235 -135 269
rect -101 235 -95 269
rect -141 197 -95 235
rect -141 163 -135 197
rect -101 163 -95 197
rect -141 125 -95 163
rect -141 91 -135 125
rect -101 91 -95 125
rect -141 53 -95 91
rect -141 19 -135 53
rect -101 19 -95 53
rect -141 -19 -95 19
rect -141 -53 -135 -19
rect -101 -53 -95 -19
rect -141 -91 -95 -53
rect -141 -125 -135 -91
rect -101 -125 -95 -91
rect -141 -163 -95 -125
rect -141 -197 -135 -163
rect -101 -197 -95 -163
rect -141 -235 -95 -197
rect -141 -269 -135 -235
rect -101 -269 -95 -235
rect -141 -300 -95 -269
rect -23 269 23 300
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -300 23 -269
rect 95 269 141 300
rect 95 235 101 269
rect 135 235 141 269
rect 95 197 141 235
rect 95 163 101 197
rect 135 163 141 197
rect 95 125 141 163
rect 95 91 101 125
rect 135 91 141 125
rect 95 53 141 91
rect 95 19 101 53
rect 135 19 141 53
rect 95 -19 141 19
rect 95 -53 101 -19
rect 135 -53 141 -19
rect 95 -91 141 -53
rect 95 -125 101 -91
rect 135 -125 141 -91
rect 95 -163 141 -125
rect 95 -197 101 -163
rect 135 -197 141 -163
rect 95 -235 141 -197
rect 95 -269 101 -235
rect 135 -269 141 -235
rect 95 -300 141 -269
<< end >>
