magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -356 272 355 306
rect -356 208 271 272
rect 335 208 355 272
rect -356 192 355 208
rect -356 128 271 192
rect 335 128 355 192
rect -356 112 355 128
rect -356 48 271 112
rect 335 48 355 112
rect -356 32 355 48
rect -356 -32 271 32
rect 335 -32 355 32
rect -356 -48 355 -32
rect -356 -112 271 -48
rect 335 -112 355 -48
rect -356 -128 355 -112
rect -356 -192 271 -128
rect 335 -192 355 -128
rect -356 -208 355 -192
rect -356 -272 271 -208
rect 335 -272 355 -208
rect -356 -306 355 -272
<< via3 >>
rect 271 208 335 272
rect 271 128 335 192
rect 271 48 335 112
rect 271 -32 335 32
rect 271 -112 335 -48
rect 271 -192 335 -128
rect 271 -272 335 -208
<< mimcap >>
rect -256 152 156 206
rect -256 -152 -202 152
rect 102 -152 156 152
rect -256 -206 156 -152
<< mimcapcontact >>
rect -202 -152 102 152
<< metal4 >>
rect 255 272 351 294
rect 255 208 271 272
rect 335 208 351 272
rect 255 192 351 208
rect -217 152 117 167
rect -217 -152 -202 152
rect 102 -152 117 152
rect -217 -167 117 -152
rect 255 128 271 192
rect 335 128 351 192
rect 255 112 351 128
rect 255 48 271 112
rect 335 48 351 112
rect 255 32 351 48
rect 255 -32 271 32
rect 335 -32 351 32
rect 255 -48 351 -32
rect 255 -112 271 -48
rect 335 -112 351 -48
rect 255 -128 351 -112
rect 255 -192 271 -128
rect 335 -192 351 -128
rect 255 -208 351 -192
rect 255 -272 271 -208
rect 335 -272 351 -208
rect 255 -294 351 -272
<< properties >>
string FIXED_BBOX -356 -306 256 306
<< end >>
