magic
tech sky130A
magscale 1 2
timestamp 1666903823
<< nmos >>
rect -1000 -1031 1000 969
<< ndiff >>
rect -1058 957 -1000 969
rect -1058 -1019 -1046 957
rect -1012 -1019 -1000 957
rect -1058 -1031 -1000 -1019
rect 1000 957 1058 969
rect 1000 -1019 1012 957
rect 1046 -1019 1058 957
rect 1000 -1031 1058 -1019
<< ndiffc >>
rect -1046 -1019 -1012 957
rect 1012 -1019 1046 957
<< poly >>
rect -1000 1041 1000 1057
rect -1000 1007 -984 1041
rect 984 1007 1000 1041
rect -1000 969 1000 1007
rect -1000 -1057 1000 -1031
<< polycont >>
rect -984 1007 984 1041
<< locali >>
rect -1000 1007 -984 1041
rect 984 1007 1000 1041
rect -1046 957 -1012 973
rect -1046 -1035 -1012 -1019
rect 1012 957 1046 973
rect 1012 -1035 1046 -1019
<< viali >>
rect -984 1007 984 1041
rect -1046 -1019 -1012 957
rect 1012 -1019 1046 957
<< metal1 >>
rect -996 1041 996 1047
rect -996 1007 -984 1041
rect 984 1007 996 1041
rect -996 1001 996 1007
rect -1052 957 -1006 969
rect -1052 -1019 -1046 957
rect -1012 -1019 -1006 957
rect -1052 -1031 -1006 -1019
rect 1006 957 1052 969
rect 1006 -1019 1012 957
rect 1046 -1019 1052 957
rect 1006 -1031 1052 -1019
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 10.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
