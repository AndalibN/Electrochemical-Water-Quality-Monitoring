magic
tech sky130A
magscale 1 2
timestamp 1666802528
<< checkpaint >>
rect -1313 2274 1639 2327
rect -1313 -713 2018 2274
rect -1260 -766 2018 -713
rect -1260 -3260 1460 -766
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__nfet_01v8_A83VMN  X0
timestamp 0
transform 1 0 163 0 1 807
box -216 -260 216 260
use sky130_fd_pr__nfet_01v8_A83VMN  X1
timestamp 0
transform 1 0 542 0 1 754
box -216 -260 216 260
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 a_n29_n50#
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 a_n127_n50#
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 a_69_n50#
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 a_n82_72#
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 {}
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VSUBS
port 5 nsew
<< end >>
