magic
tech sky130A
magscale 1 2
timestamp 1666810850
<< nwell >>
rect -194 -1098 194 1064
<< pmos >>
rect -100 -1036 100 964
<< pdiff >>
rect -158 952 -100 964
rect -158 -1024 -146 952
rect -112 -1024 -100 952
rect -158 -1036 -100 -1024
rect 100 952 158 964
rect 100 -1024 112 952
rect 146 -1024 158 952
rect 100 -1036 158 -1024
<< pdiffc >>
rect -146 -1024 -112 952
rect 112 -1024 146 952
<< poly >>
rect -100 1045 100 1061
rect -100 1011 -84 1045
rect 84 1011 100 1045
rect -100 964 100 1011
rect -100 -1062 100 -1036
<< polycont >>
rect -84 1011 84 1045
<< locali >>
rect -100 1011 -84 1045
rect 84 1011 100 1045
rect -146 952 -112 968
rect -146 -1040 -112 -1024
rect 112 952 146 968
rect 112 -1040 146 -1024
<< viali >>
rect -84 1011 84 1045
rect -146 -1024 -112 952
rect 112 -1024 146 952
<< metal1 >>
rect -96 1045 96 1051
rect -96 1011 -84 1045
rect 84 1011 96 1045
rect -96 1005 96 1011
rect -152 952 -106 964
rect -152 -1024 -146 952
rect -112 -1024 -106 952
rect -152 -1036 -106 -1024
rect 106 952 152 964
rect 106 -1024 112 952
rect 146 -1024 152 952
rect 106 -1036 152 -1024
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
