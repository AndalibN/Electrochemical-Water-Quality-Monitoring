magic
tech sky130A
magscale 1 2
timestamp 1666403283
<< error_p >>
rect -265 511 -207 517
rect -147 511 -89 517
rect -29 511 29 517
rect 89 511 147 517
rect 207 511 265 517
rect -265 477 -253 511
rect -147 477 -135 511
rect -29 477 -17 511
rect 89 477 101 511
rect 207 477 219 511
rect -265 471 -207 477
rect -147 471 -89 477
rect -29 471 29 477
rect 89 471 147 477
rect 207 471 265 477
rect -265 -477 -207 -471
rect -147 -477 -89 -471
rect -29 -477 29 -471
rect 89 -477 147 -471
rect 207 -477 265 -471
rect -265 -511 -253 -477
rect -147 -511 -135 -477
rect -29 -511 -17 -477
rect 89 -511 101 -477
rect 207 -511 219 -477
rect -265 -517 -207 -511
rect -147 -517 -89 -511
rect -29 -517 29 -511
rect 89 -517 147 -511
rect 207 -517 265 -511
<< nwell >>
rect -360 -530 360 530
<< pmos >>
rect -266 -430 -206 430
rect -148 -430 -88 430
rect -30 -430 30 430
rect 88 -430 148 430
rect 206 -430 266 430
<< pdiff >>
rect -324 418 -266 430
rect -324 -418 -312 418
rect -278 -418 -266 418
rect -324 -430 -266 -418
rect -206 418 -148 430
rect -206 -418 -194 418
rect -160 -418 -148 418
rect -206 -430 -148 -418
rect -88 418 -30 430
rect -88 -418 -76 418
rect -42 -418 -30 418
rect -88 -430 -30 -418
rect 30 418 88 430
rect 30 -418 42 418
rect 76 -418 88 418
rect 30 -430 88 -418
rect 148 418 206 430
rect 148 -418 160 418
rect 194 -418 206 418
rect 148 -430 206 -418
rect 266 418 324 430
rect 266 -418 278 418
rect 312 -418 324 418
rect 266 -430 324 -418
<< pdiffc >>
rect -312 -418 -278 418
rect -194 -418 -160 418
rect -76 -418 -42 418
rect 42 -418 76 418
rect 160 -418 194 418
rect 278 -418 312 418
<< poly >>
rect -269 511 -203 527
rect -269 477 -253 511
rect -219 477 -203 511
rect -269 461 -203 477
rect -151 511 -85 527
rect -151 477 -135 511
rect -101 477 -85 511
rect -151 461 -85 477
rect -33 511 33 527
rect -33 477 -17 511
rect 17 477 33 511
rect -33 461 33 477
rect 85 511 151 527
rect 85 477 101 511
rect 135 477 151 511
rect 85 461 151 477
rect 203 511 269 527
rect 203 477 219 511
rect 253 477 269 511
rect 203 461 269 477
rect -266 430 -206 461
rect -148 430 -88 461
rect -30 430 30 461
rect 88 430 148 461
rect 206 430 266 461
rect -266 -461 -206 -430
rect -148 -461 -88 -430
rect -30 -461 30 -430
rect 88 -461 148 -430
rect 206 -461 266 -430
rect -269 -477 -203 -461
rect -269 -511 -253 -477
rect -219 -511 -203 -477
rect -269 -527 -203 -511
rect -151 -477 -85 -461
rect -151 -511 -135 -477
rect -101 -511 -85 -477
rect -151 -527 -85 -511
rect -33 -477 33 -461
rect -33 -511 -17 -477
rect 17 -511 33 -477
rect -33 -527 33 -511
rect 85 -477 151 -461
rect 85 -511 101 -477
rect 135 -511 151 -477
rect 85 -527 151 -511
rect 203 -477 269 -461
rect 203 -511 219 -477
rect 253 -511 269 -477
rect 203 -527 269 -511
<< polycont >>
rect -253 477 -219 511
rect -135 477 -101 511
rect -17 477 17 511
rect 101 477 135 511
rect 219 477 253 511
rect -253 -511 -219 -477
rect -135 -511 -101 -477
rect -17 -511 17 -477
rect 101 -511 135 -477
rect 219 -511 253 -477
<< locali >>
rect -269 477 -253 511
rect -219 477 -203 511
rect -151 477 -135 511
rect -101 477 -85 511
rect -33 477 -17 511
rect 17 477 33 511
rect 85 477 101 511
rect 135 477 151 511
rect 203 477 219 511
rect 253 477 269 511
rect -312 418 -278 434
rect -312 -434 -278 -418
rect -194 418 -160 434
rect -194 -434 -160 -418
rect -76 418 -42 434
rect -76 -434 -42 -418
rect 42 418 76 434
rect 42 -434 76 -418
rect 160 418 194 434
rect 160 -434 194 -418
rect 278 418 312 434
rect 278 -434 312 -418
rect -269 -511 -253 -477
rect -219 -511 -203 -477
rect -151 -511 -135 -477
rect -101 -511 -85 -477
rect -33 -511 -17 -477
rect 17 -511 33 -477
rect 85 -511 101 -477
rect 135 -511 151 -477
rect 203 -511 219 -477
rect 253 -511 269 -477
<< viali >>
rect -253 477 -219 511
rect -135 477 -101 511
rect -17 477 17 511
rect 101 477 135 511
rect 219 477 253 511
rect -312 -418 -278 418
rect -194 -418 -160 418
rect -76 -418 -42 418
rect 42 -418 76 418
rect 160 -418 194 418
rect 278 -418 312 418
rect -253 -511 -219 -477
rect -135 -511 -101 -477
rect -17 -511 17 -477
rect 101 -511 135 -477
rect 219 -511 253 -477
<< metal1 >>
rect -265 511 -207 517
rect -265 477 -253 511
rect -219 477 -207 511
rect -265 471 -207 477
rect -147 511 -89 517
rect -147 477 -135 511
rect -101 477 -89 511
rect -147 471 -89 477
rect -29 511 29 517
rect -29 477 -17 511
rect 17 477 29 511
rect -29 471 29 477
rect 89 511 147 517
rect 89 477 101 511
rect 135 477 147 511
rect 89 471 147 477
rect 207 511 265 517
rect 207 477 219 511
rect 253 477 265 511
rect 207 471 265 477
rect -318 418 -272 430
rect -318 -418 -312 418
rect -278 -418 -272 418
rect -318 -430 -272 -418
rect -200 418 -154 430
rect -200 -418 -194 418
rect -160 -418 -154 418
rect -200 -430 -154 -418
rect -82 418 -36 430
rect -82 -418 -76 418
rect -42 -418 -36 418
rect -82 -430 -36 -418
rect 36 418 82 430
rect 36 -418 42 418
rect 76 -418 82 418
rect 36 -430 82 -418
rect 154 418 200 430
rect 154 -418 160 418
rect 194 -418 200 418
rect 154 -430 200 -418
rect 272 418 318 430
rect 272 -418 278 418
rect 312 -418 318 418
rect 272 -430 318 -418
rect -265 -477 -207 -471
rect -265 -511 -253 -477
rect -219 -511 -207 -477
rect -265 -517 -207 -511
rect -147 -477 -89 -471
rect -147 -511 -135 -477
rect -101 -511 -89 -477
rect -147 -517 -89 -511
rect -29 -477 29 -471
rect -29 -511 -17 -477
rect 17 -511 29 -477
rect -29 -517 29 -511
rect 89 -477 147 -471
rect 89 -511 101 -477
rect 135 -511 147 -477
rect 89 -517 147 -511
rect 207 -477 265 -471
rect 207 -511 219 -477
rect 253 -511 265 -477
rect 207 -517 265 -511
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.3 l 0.3 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
