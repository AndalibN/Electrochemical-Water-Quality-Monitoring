magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< xpolycontact >>
rect -671 50 -601 482
rect -671 -482 -601 -50
rect -353 50 -283 482
rect -353 -482 -283 -50
rect -35 50 35 482
rect -35 -482 35 -50
rect 283 50 353 482
rect 283 -482 353 -50
rect 601 50 671 482
rect 601 -482 671 -50
<< xpolyres >>
rect -671 -50 -601 50
rect -353 -50 -283 50
rect -35 -50 35 50
rect 283 -50 353 50
rect 601 -50 671 50
<< viali >>
rect -653 428 -619 462
rect -653 356 -619 390
rect -653 284 -619 318
rect -653 212 -619 246
rect -653 140 -619 174
rect -653 68 -619 102
rect -335 428 -301 462
rect -335 356 -301 390
rect -335 284 -301 318
rect -335 212 -301 246
rect -335 140 -301 174
rect -335 68 -301 102
rect -17 428 17 462
rect -17 356 17 390
rect -17 284 17 318
rect -17 212 17 246
rect -17 140 17 174
rect -17 68 17 102
rect 301 428 335 462
rect 301 356 335 390
rect 301 284 335 318
rect 301 212 335 246
rect 301 140 335 174
rect 301 68 335 102
rect 619 428 653 462
rect 619 356 653 390
rect 619 284 653 318
rect 619 212 653 246
rect 619 140 653 174
rect 619 68 653 102
rect -653 -103 -619 -69
rect -653 -175 -619 -141
rect -653 -247 -619 -213
rect -653 -319 -619 -285
rect -653 -391 -619 -357
rect -653 -463 -619 -429
rect -335 -103 -301 -69
rect -335 -175 -301 -141
rect -335 -247 -301 -213
rect -335 -319 -301 -285
rect -335 -391 -301 -357
rect -335 -463 -301 -429
rect -17 -103 17 -69
rect -17 -175 17 -141
rect -17 -247 17 -213
rect -17 -319 17 -285
rect -17 -391 17 -357
rect -17 -463 17 -429
rect 301 -103 335 -69
rect 301 -175 335 -141
rect 301 -247 335 -213
rect 301 -319 335 -285
rect 301 -391 335 -357
rect 301 -463 335 -429
rect 619 -103 653 -69
rect 619 -175 653 -141
rect 619 -247 653 -213
rect 619 -319 653 -285
rect 619 -391 653 -357
rect 619 -463 653 -429
<< metal1 >>
rect -661 462 -611 476
rect -661 428 -653 462
rect -619 428 -611 462
rect -661 390 -611 428
rect -661 356 -653 390
rect -619 356 -611 390
rect -661 318 -611 356
rect -661 284 -653 318
rect -619 284 -611 318
rect -661 246 -611 284
rect -661 212 -653 246
rect -619 212 -611 246
rect -661 174 -611 212
rect -661 140 -653 174
rect -619 140 -611 174
rect -661 102 -611 140
rect -661 68 -653 102
rect -619 68 -611 102
rect -661 55 -611 68
rect -343 462 -293 476
rect -343 428 -335 462
rect -301 428 -293 462
rect -343 390 -293 428
rect -343 356 -335 390
rect -301 356 -293 390
rect -343 318 -293 356
rect -343 284 -335 318
rect -301 284 -293 318
rect -343 246 -293 284
rect -343 212 -335 246
rect -301 212 -293 246
rect -343 174 -293 212
rect -343 140 -335 174
rect -301 140 -293 174
rect -343 102 -293 140
rect -343 68 -335 102
rect -301 68 -293 102
rect -343 55 -293 68
rect -25 462 25 476
rect -25 428 -17 462
rect 17 428 25 462
rect -25 390 25 428
rect -25 356 -17 390
rect 17 356 25 390
rect -25 318 25 356
rect -25 284 -17 318
rect 17 284 25 318
rect -25 246 25 284
rect -25 212 -17 246
rect 17 212 25 246
rect -25 174 25 212
rect -25 140 -17 174
rect 17 140 25 174
rect -25 102 25 140
rect -25 68 -17 102
rect 17 68 25 102
rect -25 55 25 68
rect 293 462 343 476
rect 293 428 301 462
rect 335 428 343 462
rect 293 390 343 428
rect 293 356 301 390
rect 335 356 343 390
rect 293 318 343 356
rect 293 284 301 318
rect 335 284 343 318
rect 293 246 343 284
rect 293 212 301 246
rect 335 212 343 246
rect 293 174 343 212
rect 293 140 301 174
rect 335 140 343 174
rect 293 102 343 140
rect 293 68 301 102
rect 335 68 343 102
rect 293 55 343 68
rect 611 462 661 476
rect 611 428 619 462
rect 653 428 661 462
rect 611 390 661 428
rect 611 356 619 390
rect 653 356 661 390
rect 611 318 661 356
rect 611 284 619 318
rect 653 284 661 318
rect 611 246 661 284
rect 611 212 619 246
rect 653 212 661 246
rect 611 174 661 212
rect 611 140 619 174
rect 653 140 661 174
rect 611 102 661 140
rect 611 68 619 102
rect 653 68 661 102
rect 611 55 661 68
rect -661 -69 -611 -55
rect -661 -103 -653 -69
rect -619 -103 -611 -69
rect -661 -141 -611 -103
rect -661 -175 -653 -141
rect -619 -175 -611 -141
rect -661 -213 -611 -175
rect -661 -247 -653 -213
rect -619 -247 -611 -213
rect -661 -285 -611 -247
rect -661 -319 -653 -285
rect -619 -319 -611 -285
rect -661 -357 -611 -319
rect -661 -391 -653 -357
rect -619 -391 -611 -357
rect -661 -429 -611 -391
rect -661 -463 -653 -429
rect -619 -463 -611 -429
rect -661 -476 -611 -463
rect -343 -69 -293 -55
rect -343 -103 -335 -69
rect -301 -103 -293 -69
rect -343 -141 -293 -103
rect -343 -175 -335 -141
rect -301 -175 -293 -141
rect -343 -213 -293 -175
rect -343 -247 -335 -213
rect -301 -247 -293 -213
rect -343 -285 -293 -247
rect -343 -319 -335 -285
rect -301 -319 -293 -285
rect -343 -357 -293 -319
rect -343 -391 -335 -357
rect -301 -391 -293 -357
rect -343 -429 -293 -391
rect -343 -463 -335 -429
rect -301 -463 -293 -429
rect -343 -476 -293 -463
rect -25 -69 25 -55
rect -25 -103 -17 -69
rect 17 -103 25 -69
rect -25 -141 25 -103
rect -25 -175 -17 -141
rect 17 -175 25 -141
rect -25 -213 25 -175
rect -25 -247 -17 -213
rect 17 -247 25 -213
rect -25 -285 25 -247
rect -25 -319 -17 -285
rect 17 -319 25 -285
rect -25 -357 25 -319
rect -25 -391 -17 -357
rect 17 -391 25 -357
rect -25 -429 25 -391
rect -25 -463 -17 -429
rect 17 -463 25 -429
rect -25 -476 25 -463
rect 293 -69 343 -55
rect 293 -103 301 -69
rect 335 -103 343 -69
rect 293 -141 343 -103
rect 293 -175 301 -141
rect 335 -175 343 -141
rect 293 -213 343 -175
rect 293 -247 301 -213
rect 335 -247 343 -213
rect 293 -285 343 -247
rect 293 -319 301 -285
rect 335 -319 343 -285
rect 293 -357 343 -319
rect 293 -391 301 -357
rect 335 -391 343 -357
rect 293 -429 343 -391
rect 293 -463 301 -429
rect 335 -463 343 -429
rect 293 -476 343 -463
rect 611 -69 661 -55
rect 611 -103 619 -69
rect 653 -103 661 -69
rect 611 -141 661 -103
rect 611 -175 619 -141
rect 653 -175 661 -141
rect 611 -213 661 -175
rect 611 -247 619 -213
rect 653 -247 661 -213
rect 611 -285 661 -247
rect 611 -319 619 -285
rect 653 -319 661 -285
rect 611 -357 661 -319
rect 611 -391 619 -357
rect 653 -391 661 -357
rect 611 -429 661 -391
rect 611 -463 619 -429
rect 653 -463 661 -429
rect 611 -476 661 -463
<< end >>
