magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 401 29 407
rect -29 367 -17 401
rect -29 361 29 367
<< pwell >>
rect -102 -417 102 355
<< nmos >>
rect -18 -391 18 329
<< ndiff >>
rect -76 292 -18 329
rect -76 258 -64 292
rect -30 258 -18 292
rect -76 224 -18 258
rect -76 190 -64 224
rect -30 190 -18 224
rect -76 156 -18 190
rect -76 122 -64 156
rect -30 122 -18 156
rect -76 88 -18 122
rect -76 54 -64 88
rect -30 54 -18 88
rect -76 20 -18 54
rect -76 -14 -64 20
rect -30 -14 -18 20
rect -76 -48 -18 -14
rect -76 -82 -64 -48
rect -30 -82 -18 -48
rect -76 -116 -18 -82
rect -76 -150 -64 -116
rect -30 -150 -18 -116
rect -76 -184 -18 -150
rect -76 -218 -64 -184
rect -30 -218 -18 -184
rect -76 -252 -18 -218
rect -76 -286 -64 -252
rect -30 -286 -18 -252
rect -76 -320 -18 -286
rect -76 -354 -64 -320
rect -30 -354 -18 -320
rect -76 -391 -18 -354
rect 18 292 76 329
rect 18 258 30 292
rect 64 258 76 292
rect 18 224 76 258
rect 18 190 30 224
rect 64 190 76 224
rect 18 156 76 190
rect 18 122 30 156
rect 64 122 76 156
rect 18 88 76 122
rect 18 54 30 88
rect 64 54 76 88
rect 18 20 76 54
rect 18 -14 30 20
rect 64 -14 76 20
rect 18 -48 76 -14
rect 18 -82 30 -48
rect 64 -82 76 -48
rect 18 -116 76 -82
rect 18 -150 30 -116
rect 64 -150 76 -116
rect 18 -184 76 -150
rect 18 -218 30 -184
rect 64 -218 76 -184
rect 18 -252 76 -218
rect 18 -286 30 -252
rect 64 -286 76 -252
rect 18 -320 76 -286
rect 18 -354 30 -320
rect 64 -354 76 -320
rect 18 -391 76 -354
<< ndiffc >>
rect -64 258 -30 292
rect -64 190 -30 224
rect -64 122 -30 156
rect -64 54 -30 88
rect -64 -14 -30 20
rect -64 -82 -30 -48
rect -64 -150 -30 -116
rect -64 -218 -30 -184
rect -64 -286 -30 -252
rect -64 -354 -30 -320
rect 30 258 64 292
rect 30 190 64 224
rect 30 122 64 156
rect 30 54 64 88
rect 30 -14 64 20
rect 30 -82 64 -48
rect 30 -150 64 -116
rect 30 -218 64 -184
rect 30 -286 64 -252
rect 30 -354 64 -320
<< poly >>
rect -33 401 33 417
rect -33 367 -17 401
rect 17 367 33 401
rect -33 351 33 367
rect -18 329 18 351
rect -18 -417 18 -391
<< polycont >>
rect -17 367 17 401
<< locali >>
rect -33 367 -17 401
rect 17 367 33 401
rect -64 310 -30 333
rect -64 238 -30 258
rect -64 166 -30 190
rect -64 94 -30 122
rect -64 22 -30 54
rect -64 -48 -30 -14
rect -64 -116 -30 -84
rect -64 -184 -30 -156
rect -64 -252 -30 -228
rect -64 -320 -30 -300
rect -64 -395 -30 -372
rect 30 310 64 333
rect 30 238 64 258
rect 30 166 64 190
rect 30 94 64 122
rect 30 22 64 54
rect 30 -48 64 -14
rect 30 -116 64 -84
rect 30 -184 64 -156
rect 30 -252 64 -228
rect 30 -320 64 -300
rect 30 -395 64 -372
<< viali >>
rect -17 367 17 401
rect -64 292 -30 310
rect -64 276 -30 292
rect -64 224 -30 238
rect -64 204 -30 224
rect -64 156 -30 166
rect -64 132 -30 156
rect -64 88 -30 94
rect -64 60 -30 88
rect -64 20 -30 22
rect -64 -12 -30 20
rect -64 -82 -30 -50
rect -64 -84 -30 -82
rect -64 -150 -30 -122
rect -64 -156 -30 -150
rect -64 -218 -30 -194
rect -64 -228 -30 -218
rect -64 -286 -30 -266
rect -64 -300 -30 -286
rect -64 -354 -30 -338
rect -64 -372 -30 -354
rect 30 292 64 310
rect 30 276 64 292
rect 30 224 64 238
rect 30 204 64 224
rect 30 156 64 166
rect 30 132 64 156
rect 30 88 64 94
rect 30 60 64 88
rect 30 20 64 22
rect 30 -12 64 20
rect 30 -82 64 -50
rect 30 -84 64 -82
rect 30 -150 64 -122
rect 30 -156 64 -150
rect 30 -218 64 -194
rect 30 -228 64 -218
rect 30 -286 64 -266
rect 30 -300 64 -286
rect 30 -354 64 -338
rect 30 -372 64 -354
<< metal1 >>
rect -29 401 29 407
rect -29 367 -17 401
rect 17 367 29 401
rect -29 361 29 367
rect -70 310 -24 329
rect -70 276 -64 310
rect -30 276 -24 310
rect -70 238 -24 276
rect -70 204 -64 238
rect -30 204 -24 238
rect -70 166 -24 204
rect -70 132 -64 166
rect -30 132 -24 166
rect -70 94 -24 132
rect -70 60 -64 94
rect -30 60 -24 94
rect -70 22 -24 60
rect -70 -12 -64 22
rect -30 -12 -24 22
rect -70 -50 -24 -12
rect -70 -84 -64 -50
rect -30 -84 -24 -50
rect -70 -122 -24 -84
rect -70 -156 -64 -122
rect -30 -156 -24 -122
rect -70 -194 -24 -156
rect -70 -228 -64 -194
rect -30 -228 -24 -194
rect -70 -266 -24 -228
rect -70 -300 -64 -266
rect -30 -300 -24 -266
rect -70 -338 -24 -300
rect -70 -372 -64 -338
rect -30 -372 -24 -338
rect -70 -391 -24 -372
rect 24 310 70 329
rect 24 276 30 310
rect 64 276 70 310
rect 24 238 70 276
rect 24 204 30 238
rect 64 204 70 238
rect 24 166 70 204
rect 24 132 30 166
rect 64 132 70 166
rect 24 94 70 132
rect 24 60 30 94
rect 64 60 70 94
rect 24 22 70 60
rect 24 -12 30 22
rect 64 -12 70 22
rect 24 -50 70 -12
rect 24 -84 30 -50
rect 64 -84 70 -50
rect 24 -122 70 -84
rect 24 -156 30 -122
rect 64 -156 70 -122
rect 24 -194 70 -156
rect 24 -228 30 -194
rect 64 -228 70 -194
rect 24 -266 70 -228
rect 24 -300 30 -266
rect 64 -300 70 -266
rect 24 -338 70 -300
rect 24 -372 30 -338
rect 64 -372 70 -338
rect 24 -391 70 -372
<< end >>
