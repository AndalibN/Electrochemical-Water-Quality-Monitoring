magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_s >>
rect 523 428 524 684
rect 559 464 560 648
rect 706 464 708 648
rect 742 428 744 684
<< pdiff >>
rect 559 464 611 648
rect 656 464 708 648
<< metal1 >>
rect 596 1240 665 1295
rect 453 1082 520 1212
rect 552 1191 617 1211
rect 552 1139 557 1191
rect 609 1139 617 1191
rect 552 1113 617 1139
rect 649 1192 716 1212
rect 649 1140 656 1192
rect 708 1140 716 1192
rect 649 1082 716 1140
rect 453 1043 716 1082
rect 550 646 615 656
rect 550 594 559 646
rect 611 594 615 646
rect 550 582 615 594
rect 550 530 559 582
rect 611 530 615 582
rect 550 518 615 530
rect 550 466 559 518
rect 611 466 615 518
rect 550 456 615 466
rect 652 646 716 657
rect 652 594 656 646
rect 708 594 716 646
rect 652 582 716 594
rect 652 530 656 582
rect 708 530 716 582
rect 652 518 716 530
rect 652 466 656 518
rect 708 466 716 518
rect 652 457 716 466
rect 599 364 668 419
<< via1 >>
rect 557 1139 609 1191
rect 656 1140 708 1192
rect 559 594 611 646
rect 559 530 611 582
rect 559 466 611 518
rect 656 594 708 646
rect 656 530 708 582
rect 656 466 708 518
<< metal2 >>
rect 551 1191 616 1214
rect 551 1139 557 1191
rect 609 1139 616 1191
rect 551 646 616 1139
rect 551 594 559 646
rect 611 594 616 646
rect 551 582 616 594
rect 551 530 559 582
rect 611 530 616 582
rect 551 518 616 530
rect 551 466 559 518
rect 611 466 616 518
rect 551 457 616 466
rect 652 1192 716 1213
rect 652 1140 656 1192
rect 708 1140 716 1192
rect 652 646 716 1140
rect 652 594 656 646
rect 708 594 716 646
rect 652 582 716 594
rect 652 530 656 582
rect 708 530 716 582
rect 652 518 716 530
rect 652 466 656 518
rect 708 466 716 518
rect 652 457 716 466
rect 568 456 606 457
rect 660 456 698 457
use sky130_fd_pr__pfet_01v8_MGALHN  XM1
timestamp 1669522153
transform 1 0 633 0 -1 520
box -109 -198 109 164
use sky130_fd_pr__nfet_01v8_67HSAK  sky130_fd_pr__nfet_01v8_67HSAK_0
timestamp 1669522153
transform 1 0 585 0 1 1162
box -151 -76 151 138
<< labels >>
rlabel metal1 s 632 398 632 398 4 ENinverted
port 1 nsew
rlabel metal1 s 626 1264 626 1264 4 EN
port 2 nsew
rlabel metal2 s 576 766 576 766 4 Vin
port 3 nsew
rlabel metal2 s 676 766 676 766 4 Vout
port 4 nsew
<< end >>
