magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -1249 1152 1248 1199
rect -1249 1088 1164 1152
rect 1228 1088 1248 1152
rect -1249 1072 1248 1088
rect -1249 1008 1164 1072
rect 1228 1008 1248 1072
rect -1249 992 1248 1008
rect -1249 928 1164 992
rect 1228 928 1248 992
rect -1249 912 1248 928
rect -1249 848 1164 912
rect 1228 848 1248 912
rect -1249 832 1248 848
rect -1249 768 1164 832
rect 1228 768 1248 832
rect -1249 752 1248 768
rect -1249 688 1164 752
rect 1228 688 1248 752
rect -1249 672 1248 688
rect -1249 608 1164 672
rect 1228 608 1248 672
rect -1249 592 1248 608
rect -1249 528 1164 592
rect 1228 528 1248 592
rect -1249 512 1248 528
rect -1249 448 1164 512
rect 1228 448 1248 512
rect -1249 432 1248 448
rect -1249 368 1164 432
rect 1228 368 1248 432
rect -1249 352 1248 368
rect -1249 288 1164 352
rect 1228 288 1248 352
rect -1249 272 1248 288
rect -1249 208 1164 272
rect 1228 208 1248 272
rect -1249 192 1248 208
rect -1249 128 1164 192
rect 1228 128 1248 192
rect -1249 112 1248 128
rect -1249 48 1164 112
rect 1228 48 1248 112
rect -1249 32 1248 48
rect -1249 -32 1164 32
rect 1228 -32 1248 32
rect -1249 -48 1248 -32
rect -1249 -112 1164 -48
rect 1228 -112 1248 -48
rect -1249 -128 1248 -112
rect -1249 -192 1164 -128
rect 1228 -192 1248 -128
rect -1249 -208 1248 -192
rect -1249 -272 1164 -208
rect 1228 -272 1248 -208
rect -1249 -288 1248 -272
rect -1249 -352 1164 -288
rect 1228 -352 1248 -288
rect -1249 -368 1248 -352
rect -1249 -432 1164 -368
rect 1228 -432 1248 -368
rect -1249 -448 1248 -432
rect -1249 -512 1164 -448
rect 1228 -512 1248 -448
rect -1249 -528 1248 -512
rect -1249 -592 1164 -528
rect 1228 -592 1248 -528
rect -1249 -608 1248 -592
rect -1249 -672 1164 -608
rect 1228 -672 1248 -608
rect -1249 -688 1248 -672
rect -1249 -752 1164 -688
rect 1228 -752 1248 -688
rect -1249 -768 1248 -752
rect -1249 -832 1164 -768
rect 1228 -832 1248 -768
rect -1249 -848 1248 -832
rect -1249 -912 1164 -848
rect 1228 -912 1248 -848
rect -1249 -928 1248 -912
rect -1249 -992 1164 -928
rect 1228 -992 1248 -928
rect -1249 -1008 1248 -992
rect -1249 -1072 1164 -1008
rect 1228 -1072 1248 -1008
rect -1249 -1088 1248 -1072
rect -1249 -1152 1164 -1088
rect 1228 -1152 1248 -1088
rect -1249 -1199 1248 -1152
<< via3 >>
rect 1164 1088 1228 1152
rect 1164 1008 1228 1072
rect 1164 928 1228 992
rect 1164 848 1228 912
rect 1164 768 1228 832
rect 1164 688 1228 752
rect 1164 608 1228 672
rect 1164 528 1228 592
rect 1164 448 1228 512
rect 1164 368 1228 432
rect 1164 288 1228 352
rect 1164 208 1228 272
rect 1164 128 1228 192
rect 1164 48 1228 112
rect 1164 -32 1228 32
rect 1164 -112 1228 -48
rect 1164 -192 1228 -128
rect 1164 -272 1228 -208
rect 1164 -352 1228 -288
rect 1164 -432 1228 -368
rect 1164 -512 1228 -448
rect 1164 -592 1228 -528
rect 1164 -672 1228 -608
rect 1164 -752 1228 -688
rect 1164 -832 1228 -768
rect 1164 -912 1228 -848
rect 1164 -992 1228 -928
rect 1164 -1072 1228 -1008
rect 1164 -1152 1228 -1088
<< mimcap >>
rect -1149 1032 1049 1099
rect -1149 -1032 -1082 1032
rect 982 -1032 1049 1032
rect -1149 -1099 1049 -1032
<< mimcapcontact >>
rect -1082 -1032 982 1032
<< metal4 >>
rect 1148 1152 1244 1187
rect 1148 1088 1164 1152
rect 1228 1088 1244 1152
rect 1148 1072 1244 1088
rect -1110 1032 1010 1060
rect -1110 -1032 -1082 1032
rect 982 -1032 1010 1032
rect -1110 -1060 1010 -1032
rect 1148 1008 1164 1072
rect 1228 1008 1244 1072
rect 1148 992 1244 1008
rect 1148 928 1164 992
rect 1228 928 1244 992
rect 1148 912 1244 928
rect 1148 848 1164 912
rect 1228 848 1244 912
rect 1148 832 1244 848
rect 1148 768 1164 832
rect 1228 768 1244 832
rect 1148 752 1244 768
rect 1148 688 1164 752
rect 1228 688 1244 752
rect 1148 672 1244 688
rect 1148 608 1164 672
rect 1228 608 1244 672
rect 1148 592 1244 608
rect 1148 528 1164 592
rect 1228 528 1244 592
rect 1148 512 1244 528
rect 1148 448 1164 512
rect 1228 448 1244 512
rect 1148 432 1244 448
rect 1148 368 1164 432
rect 1228 368 1244 432
rect 1148 352 1244 368
rect 1148 288 1164 352
rect 1228 288 1244 352
rect 1148 272 1244 288
rect 1148 208 1164 272
rect 1228 208 1244 272
rect 1148 192 1244 208
rect 1148 128 1164 192
rect 1228 128 1244 192
rect 1148 112 1244 128
rect 1148 48 1164 112
rect 1228 48 1244 112
rect 1148 32 1244 48
rect 1148 -32 1164 32
rect 1228 -32 1244 32
rect 1148 -48 1244 -32
rect 1148 -112 1164 -48
rect 1228 -112 1244 -48
rect 1148 -128 1244 -112
rect 1148 -192 1164 -128
rect 1228 -192 1244 -128
rect 1148 -208 1244 -192
rect 1148 -272 1164 -208
rect 1228 -272 1244 -208
rect 1148 -288 1244 -272
rect 1148 -352 1164 -288
rect 1228 -352 1244 -288
rect 1148 -368 1244 -352
rect 1148 -432 1164 -368
rect 1228 -432 1244 -368
rect 1148 -448 1244 -432
rect 1148 -512 1164 -448
rect 1228 -512 1244 -448
rect 1148 -528 1244 -512
rect 1148 -592 1164 -528
rect 1228 -592 1244 -528
rect 1148 -608 1244 -592
rect 1148 -672 1164 -608
rect 1228 -672 1244 -608
rect 1148 -688 1244 -672
rect 1148 -752 1164 -688
rect 1228 -752 1244 -688
rect 1148 -768 1244 -752
rect 1148 -832 1164 -768
rect 1228 -832 1244 -768
rect 1148 -848 1244 -832
rect 1148 -912 1164 -848
rect 1228 -912 1244 -848
rect 1148 -928 1244 -912
rect 1148 -992 1164 -928
rect 1228 -992 1244 -928
rect 1148 -1008 1244 -992
rect 1148 -1072 1164 -1008
rect 1228 -1072 1244 -1008
rect 1148 -1088 1244 -1072
rect 1148 -1152 1164 -1088
rect 1228 -1152 1244 -1088
rect 1148 -1187 1244 -1152
<< properties >>
string FIXED_BBOX -1249 -1199 1149 1199
<< end >>
