magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -513 -1426 513 1426
<< nmos >>
rect -429 -1400 -29 1400
rect 29 -1400 429 1400
<< ndiff >>
rect -487 1377 -429 1400
rect -487 1343 -475 1377
rect -441 1343 -429 1377
rect -487 1309 -429 1343
rect -487 1275 -475 1309
rect -441 1275 -429 1309
rect -487 1241 -429 1275
rect -487 1207 -475 1241
rect -441 1207 -429 1241
rect -487 1173 -429 1207
rect -487 1139 -475 1173
rect -441 1139 -429 1173
rect -487 1105 -429 1139
rect -487 1071 -475 1105
rect -441 1071 -429 1105
rect -487 1037 -429 1071
rect -487 1003 -475 1037
rect -441 1003 -429 1037
rect -487 969 -429 1003
rect -487 935 -475 969
rect -441 935 -429 969
rect -487 901 -429 935
rect -487 867 -475 901
rect -441 867 -429 901
rect -487 833 -429 867
rect -487 799 -475 833
rect -441 799 -429 833
rect -487 765 -429 799
rect -487 731 -475 765
rect -441 731 -429 765
rect -487 697 -429 731
rect -487 663 -475 697
rect -441 663 -429 697
rect -487 629 -429 663
rect -487 595 -475 629
rect -441 595 -429 629
rect -487 561 -429 595
rect -487 527 -475 561
rect -441 527 -429 561
rect -487 493 -429 527
rect -487 459 -475 493
rect -441 459 -429 493
rect -487 425 -429 459
rect -487 391 -475 425
rect -441 391 -429 425
rect -487 357 -429 391
rect -487 323 -475 357
rect -441 323 -429 357
rect -487 289 -429 323
rect -487 255 -475 289
rect -441 255 -429 289
rect -487 221 -429 255
rect -487 187 -475 221
rect -441 187 -429 221
rect -487 153 -429 187
rect -487 119 -475 153
rect -441 119 -429 153
rect -487 85 -429 119
rect -487 51 -475 85
rect -441 51 -429 85
rect -487 17 -429 51
rect -487 -17 -475 17
rect -441 -17 -429 17
rect -487 -51 -429 -17
rect -487 -85 -475 -51
rect -441 -85 -429 -51
rect -487 -119 -429 -85
rect -487 -153 -475 -119
rect -441 -153 -429 -119
rect -487 -187 -429 -153
rect -487 -221 -475 -187
rect -441 -221 -429 -187
rect -487 -255 -429 -221
rect -487 -289 -475 -255
rect -441 -289 -429 -255
rect -487 -323 -429 -289
rect -487 -357 -475 -323
rect -441 -357 -429 -323
rect -487 -391 -429 -357
rect -487 -425 -475 -391
rect -441 -425 -429 -391
rect -487 -459 -429 -425
rect -487 -493 -475 -459
rect -441 -493 -429 -459
rect -487 -527 -429 -493
rect -487 -561 -475 -527
rect -441 -561 -429 -527
rect -487 -595 -429 -561
rect -487 -629 -475 -595
rect -441 -629 -429 -595
rect -487 -663 -429 -629
rect -487 -697 -475 -663
rect -441 -697 -429 -663
rect -487 -731 -429 -697
rect -487 -765 -475 -731
rect -441 -765 -429 -731
rect -487 -799 -429 -765
rect -487 -833 -475 -799
rect -441 -833 -429 -799
rect -487 -867 -429 -833
rect -487 -901 -475 -867
rect -441 -901 -429 -867
rect -487 -935 -429 -901
rect -487 -969 -475 -935
rect -441 -969 -429 -935
rect -487 -1003 -429 -969
rect -487 -1037 -475 -1003
rect -441 -1037 -429 -1003
rect -487 -1071 -429 -1037
rect -487 -1105 -475 -1071
rect -441 -1105 -429 -1071
rect -487 -1139 -429 -1105
rect -487 -1173 -475 -1139
rect -441 -1173 -429 -1139
rect -487 -1207 -429 -1173
rect -487 -1241 -475 -1207
rect -441 -1241 -429 -1207
rect -487 -1275 -429 -1241
rect -487 -1309 -475 -1275
rect -441 -1309 -429 -1275
rect -487 -1343 -429 -1309
rect -487 -1377 -475 -1343
rect -441 -1377 -429 -1343
rect -487 -1400 -429 -1377
rect -29 1377 29 1400
rect -29 1343 -17 1377
rect 17 1343 29 1377
rect -29 1309 29 1343
rect -29 1275 -17 1309
rect 17 1275 29 1309
rect -29 1241 29 1275
rect -29 1207 -17 1241
rect 17 1207 29 1241
rect -29 1173 29 1207
rect -29 1139 -17 1173
rect 17 1139 29 1173
rect -29 1105 29 1139
rect -29 1071 -17 1105
rect 17 1071 29 1105
rect -29 1037 29 1071
rect -29 1003 -17 1037
rect 17 1003 29 1037
rect -29 969 29 1003
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1003 29 -969
rect -29 -1037 -17 -1003
rect 17 -1037 29 -1003
rect -29 -1071 29 -1037
rect -29 -1105 -17 -1071
rect 17 -1105 29 -1071
rect -29 -1139 29 -1105
rect -29 -1173 -17 -1139
rect 17 -1173 29 -1139
rect -29 -1207 29 -1173
rect -29 -1241 -17 -1207
rect 17 -1241 29 -1207
rect -29 -1275 29 -1241
rect -29 -1309 -17 -1275
rect 17 -1309 29 -1275
rect -29 -1343 29 -1309
rect -29 -1377 -17 -1343
rect 17 -1377 29 -1343
rect -29 -1400 29 -1377
rect 429 1377 487 1400
rect 429 1343 441 1377
rect 475 1343 487 1377
rect 429 1309 487 1343
rect 429 1275 441 1309
rect 475 1275 487 1309
rect 429 1241 487 1275
rect 429 1207 441 1241
rect 475 1207 487 1241
rect 429 1173 487 1207
rect 429 1139 441 1173
rect 475 1139 487 1173
rect 429 1105 487 1139
rect 429 1071 441 1105
rect 475 1071 487 1105
rect 429 1037 487 1071
rect 429 1003 441 1037
rect 475 1003 487 1037
rect 429 969 487 1003
rect 429 935 441 969
rect 475 935 487 969
rect 429 901 487 935
rect 429 867 441 901
rect 475 867 487 901
rect 429 833 487 867
rect 429 799 441 833
rect 475 799 487 833
rect 429 765 487 799
rect 429 731 441 765
rect 475 731 487 765
rect 429 697 487 731
rect 429 663 441 697
rect 475 663 487 697
rect 429 629 487 663
rect 429 595 441 629
rect 475 595 487 629
rect 429 561 487 595
rect 429 527 441 561
rect 475 527 487 561
rect 429 493 487 527
rect 429 459 441 493
rect 475 459 487 493
rect 429 425 487 459
rect 429 391 441 425
rect 475 391 487 425
rect 429 357 487 391
rect 429 323 441 357
rect 475 323 487 357
rect 429 289 487 323
rect 429 255 441 289
rect 475 255 487 289
rect 429 221 487 255
rect 429 187 441 221
rect 475 187 487 221
rect 429 153 487 187
rect 429 119 441 153
rect 475 119 487 153
rect 429 85 487 119
rect 429 51 441 85
rect 475 51 487 85
rect 429 17 487 51
rect 429 -17 441 17
rect 475 -17 487 17
rect 429 -51 487 -17
rect 429 -85 441 -51
rect 475 -85 487 -51
rect 429 -119 487 -85
rect 429 -153 441 -119
rect 475 -153 487 -119
rect 429 -187 487 -153
rect 429 -221 441 -187
rect 475 -221 487 -187
rect 429 -255 487 -221
rect 429 -289 441 -255
rect 475 -289 487 -255
rect 429 -323 487 -289
rect 429 -357 441 -323
rect 475 -357 487 -323
rect 429 -391 487 -357
rect 429 -425 441 -391
rect 475 -425 487 -391
rect 429 -459 487 -425
rect 429 -493 441 -459
rect 475 -493 487 -459
rect 429 -527 487 -493
rect 429 -561 441 -527
rect 475 -561 487 -527
rect 429 -595 487 -561
rect 429 -629 441 -595
rect 475 -629 487 -595
rect 429 -663 487 -629
rect 429 -697 441 -663
rect 475 -697 487 -663
rect 429 -731 487 -697
rect 429 -765 441 -731
rect 475 -765 487 -731
rect 429 -799 487 -765
rect 429 -833 441 -799
rect 475 -833 487 -799
rect 429 -867 487 -833
rect 429 -901 441 -867
rect 475 -901 487 -867
rect 429 -935 487 -901
rect 429 -969 441 -935
rect 475 -969 487 -935
rect 429 -1003 487 -969
rect 429 -1037 441 -1003
rect 475 -1037 487 -1003
rect 429 -1071 487 -1037
rect 429 -1105 441 -1071
rect 475 -1105 487 -1071
rect 429 -1139 487 -1105
rect 429 -1173 441 -1139
rect 475 -1173 487 -1139
rect 429 -1207 487 -1173
rect 429 -1241 441 -1207
rect 475 -1241 487 -1207
rect 429 -1275 487 -1241
rect 429 -1309 441 -1275
rect 475 -1309 487 -1275
rect 429 -1343 487 -1309
rect 429 -1377 441 -1343
rect 475 -1377 487 -1343
rect 429 -1400 487 -1377
<< ndiffc >>
rect -475 1343 -441 1377
rect -475 1275 -441 1309
rect -475 1207 -441 1241
rect -475 1139 -441 1173
rect -475 1071 -441 1105
rect -475 1003 -441 1037
rect -475 935 -441 969
rect -475 867 -441 901
rect -475 799 -441 833
rect -475 731 -441 765
rect -475 663 -441 697
rect -475 595 -441 629
rect -475 527 -441 561
rect -475 459 -441 493
rect -475 391 -441 425
rect -475 323 -441 357
rect -475 255 -441 289
rect -475 187 -441 221
rect -475 119 -441 153
rect -475 51 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -51
rect -475 -153 -441 -119
rect -475 -221 -441 -187
rect -475 -289 -441 -255
rect -475 -357 -441 -323
rect -475 -425 -441 -391
rect -475 -493 -441 -459
rect -475 -561 -441 -527
rect -475 -629 -441 -595
rect -475 -697 -441 -663
rect -475 -765 -441 -731
rect -475 -833 -441 -799
rect -475 -901 -441 -867
rect -475 -969 -441 -935
rect -475 -1037 -441 -1003
rect -475 -1105 -441 -1071
rect -475 -1173 -441 -1139
rect -475 -1241 -441 -1207
rect -475 -1309 -441 -1275
rect -475 -1377 -441 -1343
rect -17 1343 17 1377
rect -17 1275 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1173
rect -17 1071 17 1105
rect -17 1003 17 1037
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect -17 -1037 17 -1003
rect -17 -1105 17 -1071
rect -17 -1173 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1275
rect -17 -1377 17 -1343
rect 441 1343 475 1377
rect 441 1275 475 1309
rect 441 1207 475 1241
rect 441 1139 475 1173
rect 441 1071 475 1105
rect 441 1003 475 1037
rect 441 935 475 969
rect 441 867 475 901
rect 441 799 475 833
rect 441 731 475 765
rect 441 663 475 697
rect 441 595 475 629
rect 441 527 475 561
rect 441 459 475 493
rect 441 391 475 425
rect 441 323 475 357
rect 441 255 475 289
rect 441 187 475 221
rect 441 119 475 153
rect 441 51 475 85
rect 441 -17 475 17
rect 441 -85 475 -51
rect 441 -153 475 -119
rect 441 -221 475 -187
rect 441 -289 475 -255
rect 441 -357 475 -323
rect 441 -425 475 -391
rect 441 -493 475 -459
rect 441 -561 475 -527
rect 441 -629 475 -595
rect 441 -697 475 -663
rect 441 -765 475 -731
rect 441 -833 475 -799
rect 441 -901 475 -867
rect 441 -969 475 -935
rect 441 -1037 475 -1003
rect 441 -1105 475 -1071
rect 441 -1173 475 -1139
rect 441 -1241 475 -1207
rect 441 -1309 475 -1275
rect 441 -1377 475 -1343
<< poly >>
rect -429 1400 -29 1426
rect 29 1400 429 1426
rect -429 -1426 -29 -1400
rect 29 -1426 429 -1400
<< locali >>
rect -475 1385 -441 1404
rect -475 1313 -441 1343
rect -475 1241 -441 1275
rect -475 1173 -441 1207
rect -475 1105 -441 1135
rect -475 1037 -441 1063
rect -475 969 -441 991
rect -475 901 -441 919
rect -475 833 -441 847
rect -475 765 -441 775
rect -475 697 -441 703
rect -475 629 -441 631
rect -475 593 -441 595
rect -475 521 -441 527
rect -475 449 -441 459
rect -475 377 -441 391
rect -475 305 -441 323
rect -475 233 -441 255
rect -475 161 -441 187
rect -475 89 -441 119
rect -475 17 -441 51
rect -475 -51 -441 -17
rect -475 -119 -441 -89
rect -475 -187 -441 -161
rect -475 -255 -441 -233
rect -475 -323 -441 -305
rect -475 -391 -441 -377
rect -475 -459 -441 -449
rect -475 -527 -441 -521
rect -475 -595 -441 -593
rect -475 -631 -441 -629
rect -475 -703 -441 -697
rect -475 -775 -441 -765
rect -475 -847 -441 -833
rect -475 -919 -441 -901
rect -475 -991 -441 -969
rect -475 -1063 -441 -1037
rect -475 -1135 -441 -1105
rect -475 -1207 -441 -1173
rect -475 -1275 -441 -1241
rect -475 -1343 -441 -1313
rect -475 -1404 -441 -1385
rect -17 1385 17 1404
rect -17 1313 17 1343
rect -17 1241 17 1275
rect -17 1173 17 1207
rect -17 1105 17 1135
rect -17 1037 17 1063
rect -17 969 17 991
rect -17 901 17 919
rect -17 833 17 847
rect -17 765 17 775
rect -17 697 17 703
rect -17 629 17 631
rect -17 593 17 595
rect -17 521 17 527
rect -17 449 17 459
rect -17 377 17 391
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -391 17 -377
rect -17 -459 17 -449
rect -17 -527 17 -521
rect -17 -595 17 -593
rect -17 -631 17 -629
rect -17 -703 17 -697
rect -17 -775 17 -765
rect -17 -847 17 -833
rect -17 -919 17 -901
rect -17 -991 17 -969
rect -17 -1063 17 -1037
rect -17 -1135 17 -1105
rect -17 -1207 17 -1173
rect -17 -1275 17 -1241
rect -17 -1343 17 -1313
rect -17 -1404 17 -1385
rect 441 1385 475 1404
rect 441 1313 475 1343
rect 441 1241 475 1275
rect 441 1173 475 1207
rect 441 1105 475 1135
rect 441 1037 475 1063
rect 441 969 475 991
rect 441 901 475 919
rect 441 833 475 847
rect 441 765 475 775
rect 441 697 475 703
rect 441 629 475 631
rect 441 593 475 595
rect 441 521 475 527
rect 441 449 475 459
rect 441 377 475 391
rect 441 305 475 323
rect 441 233 475 255
rect 441 161 475 187
rect 441 89 475 119
rect 441 17 475 51
rect 441 -51 475 -17
rect 441 -119 475 -89
rect 441 -187 475 -161
rect 441 -255 475 -233
rect 441 -323 475 -305
rect 441 -391 475 -377
rect 441 -459 475 -449
rect 441 -527 475 -521
rect 441 -595 475 -593
rect 441 -631 475 -629
rect 441 -703 475 -697
rect 441 -775 475 -765
rect 441 -847 475 -833
rect 441 -919 475 -901
rect 441 -991 475 -969
rect 441 -1063 475 -1037
rect 441 -1135 475 -1105
rect 441 -1207 475 -1173
rect 441 -1275 475 -1241
rect 441 -1343 475 -1313
rect 441 -1404 475 -1385
<< viali >>
rect -475 1377 -441 1385
rect -475 1351 -441 1377
rect -475 1309 -441 1313
rect -475 1279 -441 1309
rect -475 1207 -441 1241
rect -475 1139 -441 1169
rect -475 1135 -441 1139
rect -475 1071 -441 1097
rect -475 1063 -441 1071
rect -475 1003 -441 1025
rect -475 991 -441 1003
rect -475 935 -441 953
rect -475 919 -441 935
rect -475 867 -441 881
rect -475 847 -441 867
rect -475 799 -441 809
rect -475 775 -441 799
rect -475 731 -441 737
rect -475 703 -441 731
rect -475 663 -441 665
rect -475 631 -441 663
rect -475 561 -441 593
rect -475 559 -441 561
rect -475 493 -441 521
rect -475 487 -441 493
rect -475 425 -441 449
rect -475 415 -441 425
rect -475 357 -441 377
rect -475 343 -441 357
rect -475 289 -441 305
rect -475 271 -441 289
rect -475 221 -441 233
rect -475 199 -441 221
rect -475 153 -441 161
rect -475 127 -441 153
rect -475 85 -441 89
rect -475 55 -441 85
rect -475 -17 -441 17
rect -475 -85 -441 -55
rect -475 -89 -441 -85
rect -475 -153 -441 -127
rect -475 -161 -441 -153
rect -475 -221 -441 -199
rect -475 -233 -441 -221
rect -475 -289 -441 -271
rect -475 -305 -441 -289
rect -475 -357 -441 -343
rect -475 -377 -441 -357
rect -475 -425 -441 -415
rect -475 -449 -441 -425
rect -475 -493 -441 -487
rect -475 -521 -441 -493
rect -475 -561 -441 -559
rect -475 -593 -441 -561
rect -475 -663 -441 -631
rect -475 -665 -441 -663
rect -475 -731 -441 -703
rect -475 -737 -441 -731
rect -475 -799 -441 -775
rect -475 -809 -441 -799
rect -475 -867 -441 -847
rect -475 -881 -441 -867
rect -475 -935 -441 -919
rect -475 -953 -441 -935
rect -475 -1003 -441 -991
rect -475 -1025 -441 -1003
rect -475 -1071 -441 -1063
rect -475 -1097 -441 -1071
rect -475 -1139 -441 -1135
rect -475 -1169 -441 -1139
rect -475 -1241 -441 -1207
rect -475 -1309 -441 -1279
rect -475 -1313 -441 -1309
rect -475 -1377 -441 -1351
rect -475 -1385 -441 -1377
rect -17 1377 17 1385
rect -17 1351 17 1377
rect -17 1309 17 1313
rect -17 1279 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1169
rect -17 1135 17 1139
rect -17 1071 17 1097
rect -17 1063 17 1071
rect -17 1003 17 1025
rect -17 991 17 1003
rect -17 935 17 953
rect -17 919 17 935
rect -17 867 17 881
rect -17 847 17 867
rect -17 799 17 809
rect -17 775 17 799
rect -17 731 17 737
rect -17 703 17 731
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect -17 -731 17 -703
rect -17 -737 17 -731
rect -17 -799 17 -775
rect -17 -809 17 -799
rect -17 -867 17 -847
rect -17 -881 17 -867
rect -17 -935 17 -919
rect -17 -953 17 -935
rect -17 -1003 17 -991
rect -17 -1025 17 -1003
rect -17 -1071 17 -1063
rect -17 -1097 17 -1071
rect -17 -1139 17 -1135
rect -17 -1169 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1279
rect -17 -1313 17 -1309
rect -17 -1377 17 -1351
rect -17 -1385 17 -1377
rect 441 1377 475 1385
rect 441 1351 475 1377
rect 441 1309 475 1313
rect 441 1279 475 1309
rect 441 1207 475 1241
rect 441 1139 475 1169
rect 441 1135 475 1139
rect 441 1071 475 1097
rect 441 1063 475 1071
rect 441 1003 475 1025
rect 441 991 475 1003
rect 441 935 475 953
rect 441 919 475 935
rect 441 867 475 881
rect 441 847 475 867
rect 441 799 475 809
rect 441 775 475 799
rect 441 731 475 737
rect 441 703 475 731
rect 441 663 475 665
rect 441 631 475 663
rect 441 561 475 593
rect 441 559 475 561
rect 441 493 475 521
rect 441 487 475 493
rect 441 425 475 449
rect 441 415 475 425
rect 441 357 475 377
rect 441 343 475 357
rect 441 289 475 305
rect 441 271 475 289
rect 441 221 475 233
rect 441 199 475 221
rect 441 153 475 161
rect 441 127 475 153
rect 441 85 475 89
rect 441 55 475 85
rect 441 -17 475 17
rect 441 -85 475 -55
rect 441 -89 475 -85
rect 441 -153 475 -127
rect 441 -161 475 -153
rect 441 -221 475 -199
rect 441 -233 475 -221
rect 441 -289 475 -271
rect 441 -305 475 -289
rect 441 -357 475 -343
rect 441 -377 475 -357
rect 441 -425 475 -415
rect 441 -449 475 -425
rect 441 -493 475 -487
rect 441 -521 475 -493
rect 441 -561 475 -559
rect 441 -593 475 -561
rect 441 -663 475 -631
rect 441 -665 475 -663
rect 441 -731 475 -703
rect 441 -737 475 -731
rect 441 -799 475 -775
rect 441 -809 475 -799
rect 441 -867 475 -847
rect 441 -881 475 -867
rect 441 -935 475 -919
rect 441 -953 475 -935
rect 441 -1003 475 -991
rect 441 -1025 475 -1003
rect 441 -1071 475 -1063
rect 441 -1097 475 -1071
rect 441 -1139 475 -1135
rect 441 -1169 475 -1139
rect 441 -1241 475 -1207
rect 441 -1309 475 -1279
rect 441 -1313 475 -1309
rect 441 -1377 475 -1351
rect 441 -1385 475 -1377
<< metal1 >>
rect -481 1385 -435 1400
rect -481 1351 -475 1385
rect -441 1351 -435 1385
rect -481 1313 -435 1351
rect -481 1279 -475 1313
rect -441 1279 -435 1313
rect -481 1241 -435 1279
rect -481 1207 -475 1241
rect -441 1207 -435 1241
rect -481 1169 -435 1207
rect -481 1135 -475 1169
rect -441 1135 -435 1169
rect -481 1097 -435 1135
rect -481 1063 -475 1097
rect -441 1063 -435 1097
rect -481 1025 -435 1063
rect -481 991 -475 1025
rect -441 991 -435 1025
rect -481 953 -435 991
rect -481 919 -475 953
rect -441 919 -435 953
rect -481 881 -435 919
rect -481 847 -475 881
rect -441 847 -435 881
rect -481 809 -435 847
rect -481 775 -475 809
rect -441 775 -435 809
rect -481 737 -435 775
rect -481 703 -475 737
rect -441 703 -435 737
rect -481 665 -435 703
rect -481 631 -475 665
rect -441 631 -435 665
rect -481 593 -435 631
rect -481 559 -475 593
rect -441 559 -435 593
rect -481 521 -435 559
rect -481 487 -475 521
rect -441 487 -435 521
rect -481 449 -435 487
rect -481 415 -475 449
rect -441 415 -435 449
rect -481 377 -435 415
rect -481 343 -475 377
rect -441 343 -435 377
rect -481 305 -435 343
rect -481 271 -475 305
rect -441 271 -435 305
rect -481 233 -435 271
rect -481 199 -475 233
rect -441 199 -435 233
rect -481 161 -435 199
rect -481 127 -475 161
rect -441 127 -435 161
rect -481 89 -435 127
rect -481 55 -475 89
rect -441 55 -435 89
rect -481 17 -435 55
rect -481 -17 -475 17
rect -441 -17 -435 17
rect -481 -55 -435 -17
rect -481 -89 -475 -55
rect -441 -89 -435 -55
rect -481 -127 -435 -89
rect -481 -161 -475 -127
rect -441 -161 -435 -127
rect -481 -199 -435 -161
rect -481 -233 -475 -199
rect -441 -233 -435 -199
rect -481 -271 -435 -233
rect -481 -305 -475 -271
rect -441 -305 -435 -271
rect -481 -343 -435 -305
rect -481 -377 -475 -343
rect -441 -377 -435 -343
rect -481 -415 -435 -377
rect -481 -449 -475 -415
rect -441 -449 -435 -415
rect -481 -487 -435 -449
rect -481 -521 -475 -487
rect -441 -521 -435 -487
rect -481 -559 -435 -521
rect -481 -593 -475 -559
rect -441 -593 -435 -559
rect -481 -631 -435 -593
rect -481 -665 -475 -631
rect -441 -665 -435 -631
rect -481 -703 -435 -665
rect -481 -737 -475 -703
rect -441 -737 -435 -703
rect -481 -775 -435 -737
rect -481 -809 -475 -775
rect -441 -809 -435 -775
rect -481 -847 -435 -809
rect -481 -881 -475 -847
rect -441 -881 -435 -847
rect -481 -919 -435 -881
rect -481 -953 -475 -919
rect -441 -953 -435 -919
rect -481 -991 -435 -953
rect -481 -1025 -475 -991
rect -441 -1025 -435 -991
rect -481 -1063 -435 -1025
rect -481 -1097 -475 -1063
rect -441 -1097 -435 -1063
rect -481 -1135 -435 -1097
rect -481 -1169 -475 -1135
rect -441 -1169 -435 -1135
rect -481 -1207 -435 -1169
rect -481 -1241 -475 -1207
rect -441 -1241 -435 -1207
rect -481 -1279 -435 -1241
rect -481 -1313 -475 -1279
rect -441 -1313 -435 -1279
rect -481 -1351 -435 -1313
rect -481 -1385 -475 -1351
rect -441 -1385 -435 -1351
rect -481 -1400 -435 -1385
rect -23 1385 23 1400
rect -23 1351 -17 1385
rect 17 1351 23 1385
rect -23 1313 23 1351
rect -23 1279 -17 1313
rect 17 1279 23 1313
rect -23 1241 23 1279
rect -23 1207 -17 1241
rect 17 1207 23 1241
rect -23 1169 23 1207
rect -23 1135 -17 1169
rect 17 1135 23 1169
rect -23 1097 23 1135
rect -23 1063 -17 1097
rect 17 1063 23 1097
rect -23 1025 23 1063
rect -23 991 -17 1025
rect 17 991 23 1025
rect -23 953 23 991
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -991 23 -953
rect -23 -1025 -17 -991
rect 17 -1025 23 -991
rect -23 -1063 23 -1025
rect -23 -1097 -17 -1063
rect 17 -1097 23 -1063
rect -23 -1135 23 -1097
rect -23 -1169 -17 -1135
rect 17 -1169 23 -1135
rect -23 -1207 23 -1169
rect -23 -1241 -17 -1207
rect 17 -1241 23 -1207
rect -23 -1279 23 -1241
rect -23 -1313 -17 -1279
rect 17 -1313 23 -1279
rect -23 -1351 23 -1313
rect -23 -1385 -17 -1351
rect 17 -1385 23 -1351
rect -23 -1400 23 -1385
rect 435 1385 481 1400
rect 435 1351 441 1385
rect 475 1351 481 1385
rect 435 1313 481 1351
rect 435 1279 441 1313
rect 475 1279 481 1313
rect 435 1241 481 1279
rect 435 1207 441 1241
rect 475 1207 481 1241
rect 435 1169 481 1207
rect 435 1135 441 1169
rect 475 1135 481 1169
rect 435 1097 481 1135
rect 435 1063 441 1097
rect 475 1063 481 1097
rect 435 1025 481 1063
rect 435 991 441 1025
rect 475 991 481 1025
rect 435 953 481 991
rect 435 919 441 953
rect 475 919 481 953
rect 435 881 481 919
rect 435 847 441 881
rect 475 847 481 881
rect 435 809 481 847
rect 435 775 441 809
rect 475 775 481 809
rect 435 737 481 775
rect 435 703 441 737
rect 475 703 481 737
rect 435 665 481 703
rect 435 631 441 665
rect 475 631 481 665
rect 435 593 481 631
rect 435 559 441 593
rect 475 559 481 593
rect 435 521 481 559
rect 435 487 441 521
rect 475 487 481 521
rect 435 449 481 487
rect 435 415 441 449
rect 475 415 481 449
rect 435 377 481 415
rect 435 343 441 377
rect 475 343 481 377
rect 435 305 481 343
rect 435 271 441 305
rect 475 271 481 305
rect 435 233 481 271
rect 435 199 441 233
rect 475 199 481 233
rect 435 161 481 199
rect 435 127 441 161
rect 475 127 481 161
rect 435 89 481 127
rect 435 55 441 89
rect 475 55 481 89
rect 435 17 481 55
rect 435 -17 441 17
rect 475 -17 481 17
rect 435 -55 481 -17
rect 435 -89 441 -55
rect 475 -89 481 -55
rect 435 -127 481 -89
rect 435 -161 441 -127
rect 475 -161 481 -127
rect 435 -199 481 -161
rect 435 -233 441 -199
rect 475 -233 481 -199
rect 435 -271 481 -233
rect 435 -305 441 -271
rect 475 -305 481 -271
rect 435 -343 481 -305
rect 435 -377 441 -343
rect 475 -377 481 -343
rect 435 -415 481 -377
rect 435 -449 441 -415
rect 475 -449 481 -415
rect 435 -487 481 -449
rect 435 -521 441 -487
rect 475 -521 481 -487
rect 435 -559 481 -521
rect 435 -593 441 -559
rect 475 -593 481 -559
rect 435 -631 481 -593
rect 435 -665 441 -631
rect 475 -665 481 -631
rect 435 -703 481 -665
rect 435 -737 441 -703
rect 475 -737 481 -703
rect 435 -775 481 -737
rect 435 -809 441 -775
rect 475 -809 481 -775
rect 435 -847 481 -809
rect 435 -881 441 -847
rect 475 -881 481 -847
rect 435 -919 481 -881
rect 435 -953 441 -919
rect 475 -953 481 -919
rect 435 -991 481 -953
rect 435 -1025 441 -991
rect 475 -1025 481 -991
rect 435 -1063 481 -1025
rect 435 -1097 441 -1063
rect 475 -1097 481 -1063
rect 435 -1135 481 -1097
rect 435 -1169 441 -1135
rect 475 -1169 481 -1135
rect 435 -1207 481 -1169
rect 435 -1241 441 -1207
rect 475 -1241 481 -1207
rect 435 -1279 481 -1241
rect 435 -1313 441 -1279
rect 475 -1313 481 -1279
rect 435 -1351 481 -1313
rect 435 -1385 441 -1351
rect 475 -1385 481 -1351
rect 435 -1400 481 -1385
<< end >>
