magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nwell >>
rect -144 -10100 144 10100
<< pmos >>
rect -50 -10000 50 10000
<< pdiff >>
rect -108 9988 -50 10000
rect -108 -9988 -96 9988
rect -62 -9988 -50 9988
rect -108 -10000 -50 -9988
rect 50 9988 108 10000
rect 50 -9988 62 9988
rect 96 -9988 108 9988
rect 50 -10000 108 -9988
<< pdiffc >>
rect -96 -9988 -62 9988
rect 62 -9988 96 9988
<< poly >>
rect -50 10081 50 10097
rect -50 10047 -34 10081
rect 34 10047 50 10081
rect -50 10000 50 10047
rect -50 -10047 50 -10000
rect -50 -10081 -34 -10047
rect 34 -10081 50 -10047
rect -50 -10097 50 -10081
<< polycont >>
rect -34 10047 34 10081
rect -34 -10081 34 -10047
<< locali >>
rect -50 10047 -34 10081
rect 34 10047 50 10081
rect -96 9988 -62 10004
rect -96 -10004 -62 -9988
rect 62 9988 96 10004
rect 62 -10004 96 -9988
rect -50 -10081 -34 -10047
rect 34 -10081 50 -10047
<< viali >>
rect -34 10047 34 10081
rect -96 -9988 -62 9988
rect 62 -9988 96 9988
rect -34 -10081 34 -10047
<< metal1 >>
rect -46 10081 46 10087
rect -46 10047 -34 10081
rect 34 10047 46 10081
rect -46 10041 46 10047
rect -102 9988 -56 10000
rect -102 -9988 -96 9988
rect -62 -9988 -56 9988
rect -102 -10000 -56 -9988
rect 56 9988 102 10000
rect 56 -9988 62 9988
rect 96 -9988 102 9988
rect 56 -10000 102 -9988
rect -46 -10047 46 -10041
rect -46 -10081 -34 -10047
rect 34 -10081 46 -10047
rect -46 -10087 46 -10081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 100.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
