magic
tech sky130A
magscale 1 2
timestamp 1667322661
<< nmoslvt >>
rect -2961 -9900 -2421 9900
rect -2363 -9900 -1823 9900
rect -1765 -9900 -1225 9900
rect -1167 -9900 -627 9900
rect -569 -9900 -29 9900
rect 29 -9900 569 9900
rect 627 -9900 1167 9900
rect 1225 -9900 1765 9900
rect 1823 -9900 2363 9900
rect 2421 -9900 2961 9900
<< ndiff >>
rect -3019 9888 -2961 9900
rect -3019 -9888 -3007 9888
rect -2973 -9888 -2961 9888
rect -3019 -9900 -2961 -9888
rect -2421 9888 -2363 9900
rect -2421 -9888 -2409 9888
rect -2375 -9888 -2363 9888
rect -2421 -9900 -2363 -9888
rect -1823 9888 -1765 9900
rect -1823 -9888 -1811 9888
rect -1777 -9888 -1765 9888
rect -1823 -9900 -1765 -9888
rect -1225 9888 -1167 9900
rect -1225 -9888 -1213 9888
rect -1179 -9888 -1167 9888
rect -1225 -9900 -1167 -9888
rect -627 9888 -569 9900
rect -627 -9888 -615 9888
rect -581 -9888 -569 9888
rect -627 -9900 -569 -9888
rect -29 9888 29 9900
rect -29 -9888 -17 9888
rect 17 -9888 29 9888
rect -29 -9900 29 -9888
rect 569 9888 627 9900
rect 569 -9888 581 9888
rect 615 -9888 627 9888
rect 569 -9900 627 -9888
rect 1167 9888 1225 9900
rect 1167 -9888 1179 9888
rect 1213 -9888 1225 9888
rect 1167 -9900 1225 -9888
rect 1765 9888 1823 9900
rect 1765 -9888 1777 9888
rect 1811 -9888 1823 9888
rect 1765 -9900 1823 -9888
rect 2363 9888 2421 9900
rect 2363 -9888 2375 9888
rect 2409 -9888 2421 9888
rect 2363 -9900 2421 -9888
rect 2961 9888 3019 9900
rect 2961 -9888 2973 9888
rect 3007 -9888 3019 9888
rect 2961 -9900 3019 -9888
<< ndiffc >>
rect -3007 -9888 -2973 9888
rect -2409 -9888 -2375 9888
rect -1811 -9888 -1777 9888
rect -1213 -9888 -1179 9888
rect -615 -9888 -581 9888
rect -17 -9888 17 9888
rect 581 -9888 615 9888
rect 1179 -9888 1213 9888
rect 1777 -9888 1811 9888
rect 2375 -9888 2409 9888
rect 2973 -9888 3007 9888
<< poly >>
rect -2961 9972 -2421 9988
rect -2961 9938 -2945 9972
rect -2437 9938 -2421 9972
rect -2961 9900 -2421 9938
rect -2363 9972 -1823 9988
rect -2363 9938 -2347 9972
rect -1839 9938 -1823 9972
rect -2363 9900 -1823 9938
rect -1765 9972 -1225 9988
rect -1765 9938 -1749 9972
rect -1241 9938 -1225 9972
rect -1765 9900 -1225 9938
rect -1167 9972 -627 9988
rect -1167 9938 -1151 9972
rect -643 9938 -627 9972
rect -1167 9900 -627 9938
rect -569 9972 -29 9988
rect -569 9938 -553 9972
rect -45 9938 -29 9972
rect -569 9900 -29 9938
rect 29 9972 569 9988
rect 29 9938 45 9972
rect 553 9938 569 9972
rect 29 9900 569 9938
rect 627 9972 1167 9988
rect 627 9938 643 9972
rect 1151 9938 1167 9972
rect 627 9900 1167 9938
rect 1225 9972 1765 9988
rect 1225 9938 1241 9972
rect 1749 9938 1765 9972
rect 1225 9900 1765 9938
rect 1823 9972 2363 9988
rect 1823 9938 1839 9972
rect 2347 9938 2363 9972
rect 1823 9900 2363 9938
rect 2421 9972 2961 9988
rect 2421 9938 2437 9972
rect 2945 9938 2961 9972
rect 2421 9900 2961 9938
rect -2961 -9938 -2421 -9900
rect -2961 -9972 -2945 -9938
rect -2437 -9972 -2421 -9938
rect -2961 -9988 -2421 -9972
rect -2363 -9938 -1823 -9900
rect -2363 -9972 -2347 -9938
rect -1839 -9972 -1823 -9938
rect -2363 -9988 -1823 -9972
rect -1765 -9938 -1225 -9900
rect -1765 -9972 -1749 -9938
rect -1241 -9972 -1225 -9938
rect -1765 -9988 -1225 -9972
rect -1167 -9938 -627 -9900
rect -1167 -9972 -1151 -9938
rect -643 -9972 -627 -9938
rect -1167 -9988 -627 -9972
rect -569 -9938 -29 -9900
rect -569 -9972 -553 -9938
rect -45 -9972 -29 -9938
rect -569 -9988 -29 -9972
rect 29 -9938 569 -9900
rect 29 -9972 45 -9938
rect 553 -9972 569 -9938
rect 29 -9988 569 -9972
rect 627 -9938 1167 -9900
rect 627 -9972 643 -9938
rect 1151 -9972 1167 -9938
rect 627 -9988 1167 -9972
rect 1225 -9938 1765 -9900
rect 1225 -9972 1241 -9938
rect 1749 -9972 1765 -9938
rect 1225 -9988 1765 -9972
rect 1823 -9938 2363 -9900
rect 1823 -9972 1839 -9938
rect 2347 -9972 2363 -9938
rect 1823 -9988 2363 -9972
rect 2421 -9938 2961 -9900
rect 2421 -9972 2437 -9938
rect 2945 -9972 2961 -9938
rect 2421 -9988 2961 -9972
<< polycont >>
rect -2945 9938 -2437 9972
rect -2347 9938 -1839 9972
rect -1749 9938 -1241 9972
rect -1151 9938 -643 9972
rect -553 9938 -45 9972
rect 45 9938 553 9972
rect 643 9938 1151 9972
rect 1241 9938 1749 9972
rect 1839 9938 2347 9972
rect 2437 9938 2945 9972
rect -2945 -9972 -2437 -9938
rect -2347 -9972 -1839 -9938
rect -1749 -9972 -1241 -9938
rect -1151 -9972 -643 -9938
rect -553 -9972 -45 -9938
rect 45 -9972 553 -9938
rect 643 -9972 1151 -9938
rect 1241 -9972 1749 -9938
rect 1839 -9972 2347 -9938
rect 2437 -9972 2945 -9938
<< locali >>
rect -2961 9938 -2945 9972
rect -2437 9938 -2421 9972
rect -2363 9938 -2347 9972
rect -1839 9938 -1823 9972
rect -1765 9938 -1749 9972
rect -1241 9938 -1225 9972
rect -1167 9938 -1151 9972
rect -643 9938 -627 9972
rect -569 9938 -553 9972
rect -45 9938 -29 9972
rect 29 9938 45 9972
rect 553 9938 569 9972
rect 627 9938 643 9972
rect 1151 9938 1167 9972
rect 1225 9938 1241 9972
rect 1749 9938 1765 9972
rect 1823 9938 1839 9972
rect 2347 9938 2363 9972
rect 2421 9938 2437 9972
rect 2945 9938 2961 9972
rect -3007 9888 -2973 9904
rect -3007 -9904 -2973 -9888
rect -2409 9888 -2375 9904
rect -2409 -9904 -2375 -9888
rect -1811 9888 -1777 9904
rect -1811 -9904 -1777 -9888
rect -1213 9888 -1179 9904
rect -1213 -9904 -1179 -9888
rect -615 9888 -581 9904
rect -615 -9904 -581 -9888
rect -17 9888 17 9904
rect -17 -9904 17 -9888
rect 581 9888 615 9904
rect 581 -9904 615 -9888
rect 1179 9888 1213 9904
rect 1179 -9904 1213 -9888
rect 1777 9888 1811 9904
rect 1777 -9904 1811 -9888
rect 2375 9888 2409 9904
rect 2375 -9904 2409 -9888
rect 2973 9888 3007 9904
rect 2973 -9904 3007 -9888
rect -2961 -9972 -2945 -9938
rect -2437 -9972 -2421 -9938
rect -2363 -9972 -2347 -9938
rect -1839 -9972 -1823 -9938
rect -1765 -9972 -1749 -9938
rect -1241 -9972 -1225 -9938
rect -1167 -9972 -1151 -9938
rect -643 -9972 -627 -9938
rect -569 -9972 -553 -9938
rect -45 -9972 -29 -9938
rect 29 -9972 45 -9938
rect 553 -9972 569 -9938
rect 627 -9972 643 -9938
rect 1151 -9972 1167 -9938
rect 1225 -9972 1241 -9938
rect 1749 -9972 1765 -9938
rect 1823 -9972 1839 -9938
rect 2347 -9972 2363 -9938
rect 2421 -9972 2437 -9938
rect 2945 -9972 2961 -9938
<< viali >>
rect -2945 9938 -2437 9972
rect -2347 9938 -1839 9972
rect -1749 9938 -1241 9972
rect -1151 9938 -643 9972
rect -553 9938 -45 9972
rect 45 9938 553 9972
rect 643 9938 1151 9972
rect 1241 9938 1749 9972
rect 1839 9938 2347 9972
rect 2437 9938 2945 9972
rect -3007 -9888 -2973 9888
rect -2409 -9888 -2375 9888
rect -1811 -9888 -1777 9888
rect -1213 -9888 -1179 9888
rect -615 -9888 -581 9888
rect -17 -9888 17 9888
rect 581 -9888 615 9888
rect 1179 -9888 1213 9888
rect 1777 -9888 1811 9888
rect 2375 -9888 2409 9888
rect 2973 -9888 3007 9888
rect -2945 -9972 -2437 -9938
rect -2347 -9972 -1839 -9938
rect -1749 -9972 -1241 -9938
rect -1151 -9972 -643 -9938
rect -553 -9972 -45 -9938
rect 45 -9972 553 -9938
rect 643 -9972 1151 -9938
rect 1241 -9972 1749 -9938
rect 1839 -9972 2347 -9938
rect 2437 -9972 2945 -9938
<< metal1 >>
rect -2957 9972 -2425 9978
rect -2957 9938 -2945 9972
rect -2437 9938 -2425 9972
rect -2957 9932 -2425 9938
rect -2359 9972 -1827 9978
rect -2359 9938 -2347 9972
rect -1839 9938 -1827 9972
rect -2359 9932 -1827 9938
rect -1761 9972 -1229 9978
rect -1761 9938 -1749 9972
rect -1241 9938 -1229 9972
rect -1761 9932 -1229 9938
rect -1163 9972 -631 9978
rect -1163 9938 -1151 9972
rect -643 9938 -631 9972
rect -1163 9932 -631 9938
rect -565 9972 -33 9978
rect -565 9938 -553 9972
rect -45 9938 -33 9972
rect -565 9932 -33 9938
rect 33 9972 565 9978
rect 33 9938 45 9972
rect 553 9938 565 9972
rect 33 9932 565 9938
rect 631 9972 1163 9978
rect 631 9938 643 9972
rect 1151 9938 1163 9972
rect 631 9932 1163 9938
rect 1229 9972 1761 9978
rect 1229 9938 1241 9972
rect 1749 9938 1761 9972
rect 1229 9932 1761 9938
rect 1827 9972 2359 9978
rect 1827 9938 1839 9972
rect 2347 9938 2359 9972
rect 1827 9932 2359 9938
rect 2425 9972 2957 9978
rect 2425 9938 2437 9972
rect 2945 9938 2957 9972
rect 2425 9932 2957 9938
rect -3013 9888 -2967 9900
rect -3013 -9888 -3007 9888
rect -2973 -9888 -2967 9888
rect -3013 -9900 -2967 -9888
rect -2415 9888 -2369 9900
rect -2415 -9888 -2409 9888
rect -2375 -9888 -2369 9888
rect -2415 -9900 -2369 -9888
rect -1817 9888 -1771 9900
rect -1817 -9888 -1811 9888
rect -1777 -9888 -1771 9888
rect -1817 -9900 -1771 -9888
rect -1219 9888 -1173 9900
rect -1219 -9888 -1213 9888
rect -1179 -9888 -1173 9888
rect -1219 -9900 -1173 -9888
rect -621 9888 -575 9900
rect -621 -9888 -615 9888
rect -581 -9888 -575 9888
rect -621 -9900 -575 -9888
rect -23 9888 23 9900
rect -23 -9888 -17 9888
rect 17 -9888 23 9888
rect -23 -9900 23 -9888
rect 575 9888 621 9900
rect 575 -9888 581 9888
rect 615 -9888 621 9888
rect 575 -9900 621 -9888
rect 1173 9888 1219 9900
rect 1173 -9888 1179 9888
rect 1213 -9888 1219 9888
rect 1173 -9900 1219 -9888
rect 1771 9888 1817 9900
rect 1771 -9888 1777 9888
rect 1811 -9888 1817 9888
rect 1771 -9900 1817 -9888
rect 2369 9888 2415 9900
rect 2369 -9888 2375 9888
rect 2409 -9888 2415 9888
rect 2369 -9900 2415 -9888
rect 2967 9888 3013 9900
rect 2967 -9888 2973 9888
rect 3007 -9888 3013 9888
rect 2967 -9900 3013 -9888
rect -2957 -9938 -2425 -9932
rect -2957 -9972 -2945 -9938
rect -2437 -9972 -2425 -9938
rect -2957 -9978 -2425 -9972
rect -2359 -9938 -1827 -9932
rect -2359 -9972 -2347 -9938
rect -1839 -9972 -1827 -9938
rect -2359 -9978 -1827 -9972
rect -1761 -9938 -1229 -9932
rect -1761 -9972 -1749 -9938
rect -1241 -9972 -1229 -9938
rect -1761 -9978 -1229 -9972
rect -1163 -9938 -631 -9932
rect -1163 -9972 -1151 -9938
rect -643 -9972 -631 -9938
rect -1163 -9978 -631 -9972
rect -565 -9938 -33 -9932
rect -565 -9972 -553 -9938
rect -45 -9972 -33 -9938
rect -565 -9978 -33 -9972
rect 33 -9938 565 -9932
rect 33 -9972 45 -9938
rect 553 -9972 565 -9938
rect 33 -9978 565 -9972
rect 631 -9938 1163 -9932
rect 631 -9972 643 -9938
rect 1151 -9972 1163 -9938
rect 631 -9978 1163 -9972
rect 1229 -9938 1761 -9932
rect 1229 -9972 1241 -9938
rect 1749 -9972 1761 -9938
rect 1229 -9978 1761 -9972
rect 1827 -9938 2359 -9932
rect 1827 -9972 1839 -9938
rect 2347 -9972 2359 -9938
rect 1827 -9978 2359 -9972
rect 2425 -9938 2957 -9932
rect 2425 -9972 2437 -9938
rect 2945 -9972 2957 -9938
rect 2425 -9978 2957 -9972
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 99.0 l 2.7 m 1 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
