magic
tech sky130A
magscale 1 2
timestamp 1667048966
<< nwell >>
rect -194 -864 194 898
<< pmos >>
rect -100 -764 100 836
<< pdiff >>
rect -158 824 -100 836
rect -158 -752 -146 824
rect -112 -752 -100 824
rect -158 -764 -100 -752
rect 100 824 158 836
rect 100 -752 112 824
rect 146 -752 158 824
rect 100 -764 158 -752
<< pdiffc >>
rect -146 -752 -112 824
rect 112 -752 146 824
<< poly >>
rect -100 836 100 862
rect -100 -811 100 -764
rect -100 -845 -84 -811
rect 84 -845 100 -811
rect -100 -861 100 -845
<< polycont >>
rect -84 -845 84 -811
<< locali >>
rect -146 824 -112 840
rect -146 -768 -112 -752
rect 112 824 146 840
rect 112 -768 146 -752
rect -100 -845 -84 -811
rect 84 -845 100 -811
<< viali >>
rect -146 -752 -112 824
rect 112 -752 146 824
rect -84 -845 84 -811
<< metal1 >>
rect -152 824 -106 836
rect -152 -752 -146 824
rect -112 -752 -106 824
rect -152 -764 -106 -752
rect 106 824 152 836
rect 106 -752 112 824
rect 146 -752 152 824
rect 106 -764 152 -752
rect -96 -811 96 -805
rect -96 -845 -84 -811
rect 84 -845 96 -811
rect -96 -851 96 -845
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
