magic
tech sky130A
magscale 1 2
timestamp 1667328903
<< psubdiff >>
rect -1134 572 -784 654
rect -1134 -376 -1056 572
rect -866 -376 -784 572
rect -1134 -462 -784 -376
<< psubdiffcont >>
rect -1056 -376 -866 572
<< xpolycontact >>
rect -671 1000 -601 1432
rect -671 -1432 -601 -1000
rect -353 1000 -283 1432
rect -353 -1432 -283 -1000
rect -35 1000 35 1432
rect -35 -1432 35 -1000
rect 283 1000 353 1432
rect 283 -1432 353 -1000
rect 601 1000 671 1432
rect 601 -1432 671 -1000
<< xpolyres >>
rect -671 -1000 -601 1000
rect -353 -1000 -283 1000
rect -35 -1000 35 1000
rect 283 -1000 353 1000
rect 601 -1000 671 1000
<< locali >>
rect -283 1004 -35 1426
rect 353 1004 601 1426
rect -1094 572 -822 614
rect -1094 -376 -1056 572
rect -866 -376 -822 572
rect -1094 -418 -822 -376
rect -601 -1426 -353 -1004
rect 35 -1426 283 -1004
<< viali >>
rect -655 1017 -617 1414
rect -337 1017 -299 1414
rect -19 1017 19 1414
rect 299 1017 337 1414
rect 617 1017 655 1414
rect -655 -1414 -617 -1017
rect -337 -1414 -299 -1017
rect -19 -1414 19 -1017
rect 299 -1414 337 -1017
rect 617 -1414 655 -1017
<< metal1 >>
rect -661 1414 -611 1426
rect -661 1017 -655 1414
rect -617 1017 -611 1414
rect -661 1005 -611 1017
rect -343 1414 -293 1426
rect -343 1017 -337 1414
rect -299 1017 -293 1414
rect -343 1005 -293 1017
rect -25 1414 25 1426
rect -25 1017 -19 1414
rect 19 1017 25 1414
rect -25 1005 25 1017
rect 293 1414 343 1426
rect 293 1017 299 1414
rect 337 1017 343 1414
rect 293 1005 343 1017
rect 611 1414 661 1426
rect 611 1017 617 1414
rect 655 1017 661 1414
rect 611 1005 661 1017
rect -661 -1017 -611 -1005
rect -661 -1414 -655 -1017
rect -617 -1414 -611 -1017
rect -661 -1426 -611 -1414
rect -343 -1017 -293 -1005
rect -343 -1414 -337 -1017
rect -299 -1414 -293 -1017
rect -343 -1426 -293 -1414
rect -25 -1017 25 -1005
rect -25 -1414 -19 -1017
rect 19 -1414 25 -1017
rect -25 -1426 25 -1414
rect 293 -1017 343 -1005
rect 293 -1414 299 -1017
rect 337 -1414 343 -1017
rect 293 -1426 343 -1414
rect 611 -1017 661 -1005
rect 611 -1414 617 -1017
rect 655 -1414 661 -1017
rect 611 -1426 661 -1414
<< res0p35 >>
rect -673 -1002 -599 1002
rect -355 -1002 -281 1002
rect -37 -1002 37 1002
rect 281 -1002 355 1002
rect 599 -1002 673 1002
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 10 m 1 nx 5 wmin 0.350 lmin 0.50 rho 2000 val 58.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
