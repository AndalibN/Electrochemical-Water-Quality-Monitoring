magic
tech sky130A
magscale 1 2
timestamp 1667262629
<< xpolycontact >>
rect -35 95 35 527
rect -35 -527 35 -95
<< ppolyres >>
rect -35 -95 35 95
<< viali >>
rect -19 112 19 509
rect -19 -509 19 -112
<< metal1 >>
rect -25 509 25 521
rect -25 112 -19 509
rect 19 112 25 509
rect -25 100 25 112
rect -25 -112 25 -100
rect -25 -509 -19 -112
rect 19 -509 25 -112
rect -25 -521 25 -509
<< res0p35 >>
rect -37 -97 37 97
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 0.95 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 1.981k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
