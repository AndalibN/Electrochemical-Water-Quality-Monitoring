magic
tech sky130A
magscale 1 2
timestamp 1667414410
<< xpolycontact >>
rect -35 207 35 639
rect -35 -639 35 -207
<< ppolyres >>
rect -35 -207 35 207
<< viali >>
rect -19 224 19 621
rect -19 -621 19 -224
<< metal1 >>
rect -25 621 25 633
rect -25 224 -19 621
rect 19 224 25 621
rect -25 212 25 224
rect -25 -224 25 -212
rect -25 -621 -19 -224
rect 19 -621 25 -224
rect -25 -633 25 -621
<< res0p35 >>
rect -37 -209 37 209
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 2.07 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 3.004k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
