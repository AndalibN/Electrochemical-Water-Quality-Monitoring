magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -194 -798 194 764
<< pmos >>
rect -100 -736 100 664
<< pdiff >>
rect -158 627 -100 664
rect -158 593 -146 627
rect -112 593 -100 627
rect -158 559 -100 593
rect -158 525 -146 559
rect -112 525 -100 559
rect -158 491 -100 525
rect -158 457 -146 491
rect -112 457 -100 491
rect -158 423 -100 457
rect -158 389 -146 423
rect -112 389 -100 423
rect -158 355 -100 389
rect -158 321 -146 355
rect -112 321 -100 355
rect -158 287 -100 321
rect -158 253 -146 287
rect -112 253 -100 287
rect -158 219 -100 253
rect -158 185 -146 219
rect -112 185 -100 219
rect -158 151 -100 185
rect -158 117 -146 151
rect -112 117 -100 151
rect -158 83 -100 117
rect -158 49 -146 83
rect -112 49 -100 83
rect -158 15 -100 49
rect -158 -19 -146 15
rect -112 -19 -100 15
rect -158 -53 -100 -19
rect -158 -87 -146 -53
rect -112 -87 -100 -53
rect -158 -121 -100 -87
rect -158 -155 -146 -121
rect -112 -155 -100 -121
rect -158 -189 -100 -155
rect -158 -223 -146 -189
rect -112 -223 -100 -189
rect -158 -257 -100 -223
rect -158 -291 -146 -257
rect -112 -291 -100 -257
rect -158 -325 -100 -291
rect -158 -359 -146 -325
rect -112 -359 -100 -325
rect -158 -393 -100 -359
rect -158 -427 -146 -393
rect -112 -427 -100 -393
rect -158 -461 -100 -427
rect -158 -495 -146 -461
rect -112 -495 -100 -461
rect -158 -529 -100 -495
rect -158 -563 -146 -529
rect -112 -563 -100 -529
rect -158 -597 -100 -563
rect -158 -631 -146 -597
rect -112 -631 -100 -597
rect -158 -665 -100 -631
rect -158 -699 -146 -665
rect -112 -699 -100 -665
rect -158 -736 -100 -699
rect 100 627 158 664
rect 100 593 112 627
rect 146 593 158 627
rect 100 559 158 593
rect 100 525 112 559
rect 146 525 158 559
rect 100 491 158 525
rect 100 457 112 491
rect 146 457 158 491
rect 100 423 158 457
rect 100 389 112 423
rect 146 389 158 423
rect 100 355 158 389
rect 100 321 112 355
rect 146 321 158 355
rect 100 287 158 321
rect 100 253 112 287
rect 146 253 158 287
rect 100 219 158 253
rect 100 185 112 219
rect 146 185 158 219
rect 100 151 158 185
rect 100 117 112 151
rect 146 117 158 151
rect 100 83 158 117
rect 100 49 112 83
rect 146 49 158 83
rect 100 15 158 49
rect 100 -19 112 15
rect 146 -19 158 15
rect 100 -53 158 -19
rect 100 -87 112 -53
rect 146 -87 158 -53
rect 100 -121 158 -87
rect 100 -155 112 -121
rect 146 -155 158 -121
rect 100 -189 158 -155
rect 100 -223 112 -189
rect 146 -223 158 -189
rect 100 -257 158 -223
rect 100 -291 112 -257
rect 146 -291 158 -257
rect 100 -325 158 -291
rect 100 -359 112 -325
rect 146 -359 158 -325
rect 100 -393 158 -359
rect 100 -427 112 -393
rect 146 -427 158 -393
rect 100 -461 158 -427
rect 100 -495 112 -461
rect 146 -495 158 -461
rect 100 -529 158 -495
rect 100 -563 112 -529
rect 146 -563 158 -529
rect 100 -597 158 -563
rect 100 -631 112 -597
rect 146 -631 158 -597
rect 100 -665 158 -631
rect 100 -699 112 -665
rect 146 -699 158 -665
rect 100 -736 158 -699
<< pdiffc >>
rect -146 593 -112 627
rect -146 525 -112 559
rect -146 457 -112 491
rect -146 389 -112 423
rect -146 321 -112 355
rect -146 253 -112 287
rect -146 185 -112 219
rect -146 117 -112 151
rect -146 49 -112 83
rect -146 -19 -112 15
rect -146 -87 -112 -53
rect -146 -155 -112 -121
rect -146 -223 -112 -189
rect -146 -291 -112 -257
rect -146 -359 -112 -325
rect -146 -427 -112 -393
rect -146 -495 -112 -461
rect -146 -563 -112 -529
rect -146 -631 -112 -597
rect -146 -699 -112 -665
rect 112 593 146 627
rect 112 525 146 559
rect 112 457 146 491
rect 112 389 146 423
rect 112 321 146 355
rect 112 253 146 287
rect 112 185 146 219
rect 112 117 146 151
rect 112 49 146 83
rect 112 -19 146 15
rect 112 -87 146 -53
rect 112 -155 146 -121
rect 112 -223 146 -189
rect 112 -291 146 -257
rect 112 -359 146 -325
rect 112 -427 146 -393
rect 112 -495 146 -461
rect 112 -563 146 -529
rect 112 -631 146 -597
rect 112 -699 146 -665
<< poly >>
rect -100 745 100 761
rect -100 711 -51 745
rect -17 711 17 745
rect 51 711 100 745
rect -100 664 100 711
rect -100 -762 100 -736
<< polycont >>
rect -51 711 -17 745
rect 17 711 51 745
<< locali >>
rect -100 711 -53 745
rect -17 711 17 745
rect 53 711 100 745
rect -146 629 -112 668
rect -146 559 -112 593
rect -146 491 -112 523
rect -146 423 -112 451
rect -146 355 -112 379
rect -146 287 -112 307
rect -146 219 -112 235
rect -146 151 -112 163
rect -146 83 -112 91
rect -146 15 -112 19
rect -146 -91 -112 -87
rect -146 -163 -112 -155
rect -146 -235 -112 -223
rect -146 -307 -112 -291
rect -146 -379 -112 -359
rect -146 -451 -112 -427
rect -146 -523 -112 -495
rect -146 -595 -112 -563
rect -146 -665 -112 -631
rect -146 -740 -112 -701
rect 112 629 146 668
rect 112 559 146 593
rect 112 491 146 523
rect 112 423 146 451
rect 112 355 146 379
rect 112 287 146 307
rect 112 219 146 235
rect 112 151 146 163
rect 112 83 146 91
rect 112 15 146 19
rect 112 -91 146 -87
rect 112 -163 146 -155
rect 112 -235 146 -223
rect 112 -307 146 -291
rect 112 -379 146 -359
rect 112 -451 146 -427
rect 112 -523 146 -495
rect 112 -595 146 -563
rect 112 -665 146 -631
rect 112 -740 146 -701
<< viali >>
rect -53 711 -51 745
rect -51 711 -19 745
rect 19 711 51 745
rect 51 711 53 745
rect -146 627 -112 629
rect -146 595 -112 627
rect -146 525 -112 557
rect -146 523 -112 525
rect -146 457 -112 485
rect -146 451 -112 457
rect -146 389 -112 413
rect -146 379 -112 389
rect -146 321 -112 341
rect -146 307 -112 321
rect -146 253 -112 269
rect -146 235 -112 253
rect -146 185 -112 197
rect -146 163 -112 185
rect -146 117 -112 125
rect -146 91 -112 117
rect -146 49 -112 53
rect -146 19 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -91
rect -146 -125 -112 -121
rect -146 -189 -112 -163
rect -146 -197 -112 -189
rect -146 -257 -112 -235
rect -146 -269 -112 -257
rect -146 -325 -112 -307
rect -146 -341 -112 -325
rect -146 -393 -112 -379
rect -146 -413 -112 -393
rect -146 -461 -112 -451
rect -146 -485 -112 -461
rect -146 -529 -112 -523
rect -146 -557 -112 -529
rect -146 -597 -112 -595
rect -146 -629 -112 -597
rect -146 -699 -112 -667
rect -146 -701 -112 -699
rect 112 627 146 629
rect 112 595 146 627
rect 112 525 146 557
rect 112 523 146 525
rect 112 457 146 485
rect 112 451 146 457
rect 112 389 146 413
rect 112 379 146 389
rect 112 321 146 341
rect 112 307 146 321
rect 112 253 146 269
rect 112 235 146 253
rect 112 185 146 197
rect 112 163 146 185
rect 112 117 146 125
rect 112 91 146 117
rect 112 49 146 53
rect 112 19 146 49
rect 112 -53 146 -19
rect 112 -121 146 -91
rect 112 -125 146 -121
rect 112 -189 146 -163
rect 112 -197 146 -189
rect 112 -257 146 -235
rect 112 -269 146 -257
rect 112 -325 146 -307
rect 112 -341 146 -325
rect 112 -393 146 -379
rect 112 -413 146 -393
rect 112 -461 146 -451
rect 112 -485 146 -461
rect 112 -529 146 -523
rect 112 -557 146 -529
rect 112 -597 146 -595
rect 112 -629 146 -597
rect 112 -699 146 -667
rect 112 -701 146 -699
<< metal1 >>
rect -96 745 96 751
rect -96 711 -53 745
rect -19 711 19 745
rect 53 711 96 745
rect -96 705 96 711
rect -152 629 -106 664
rect -152 595 -146 629
rect -112 595 -106 629
rect -152 557 -106 595
rect -152 523 -146 557
rect -112 523 -106 557
rect -152 485 -106 523
rect -152 451 -146 485
rect -112 451 -106 485
rect -152 413 -106 451
rect -152 379 -146 413
rect -112 379 -106 413
rect -152 341 -106 379
rect -152 307 -146 341
rect -112 307 -106 341
rect -152 269 -106 307
rect -152 235 -146 269
rect -112 235 -106 269
rect -152 197 -106 235
rect -152 163 -146 197
rect -112 163 -106 197
rect -152 125 -106 163
rect -152 91 -146 125
rect -112 91 -106 125
rect -152 53 -106 91
rect -152 19 -146 53
rect -112 19 -106 53
rect -152 -19 -106 19
rect -152 -53 -146 -19
rect -112 -53 -106 -19
rect -152 -91 -106 -53
rect -152 -125 -146 -91
rect -112 -125 -106 -91
rect -152 -163 -106 -125
rect -152 -197 -146 -163
rect -112 -197 -106 -163
rect -152 -235 -106 -197
rect -152 -269 -146 -235
rect -112 -269 -106 -235
rect -152 -307 -106 -269
rect -152 -341 -146 -307
rect -112 -341 -106 -307
rect -152 -379 -106 -341
rect -152 -413 -146 -379
rect -112 -413 -106 -379
rect -152 -451 -106 -413
rect -152 -485 -146 -451
rect -112 -485 -106 -451
rect -152 -523 -106 -485
rect -152 -557 -146 -523
rect -112 -557 -106 -523
rect -152 -595 -106 -557
rect -152 -629 -146 -595
rect -112 -629 -106 -595
rect -152 -667 -106 -629
rect -152 -701 -146 -667
rect -112 -701 -106 -667
rect -152 -736 -106 -701
rect 106 629 152 664
rect 106 595 112 629
rect 146 595 152 629
rect 106 557 152 595
rect 106 523 112 557
rect 146 523 152 557
rect 106 485 152 523
rect 106 451 112 485
rect 146 451 152 485
rect 106 413 152 451
rect 106 379 112 413
rect 146 379 152 413
rect 106 341 152 379
rect 106 307 112 341
rect 146 307 152 341
rect 106 269 152 307
rect 106 235 112 269
rect 146 235 152 269
rect 106 197 152 235
rect 106 163 112 197
rect 146 163 152 197
rect 106 125 152 163
rect 106 91 112 125
rect 146 91 152 125
rect 106 53 152 91
rect 106 19 112 53
rect 146 19 152 53
rect 106 -19 152 19
rect 106 -53 112 -19
rect 146 -53 152 -19
rect 106 -91 152 -53
rect 106 -125 112 -91
rect 146 -125 152 -91
rect 106 -163 152 -125
rect 106 -197 112 -163
rect 146 -197 152 -163
rect 106 -235 152 -197
rect 106 -269 112 -235
rect 146 -269 152 -235
rect 106 -307 152 -269
rect 106 -341 112 -307
rect 146 -341 152 -307
rect 106 -379 152 -341
rect 106 -413 112 -379
rect 146 -413 152 -379
rect 106 -451 152 -413
rect 106 -485 112 -451
rect 146 -485 152 -451
rect 106 -523 152 -485
rect 106 -557 112 -523
rect 146 -557 152 -523
rect 106 -595 152 -557
rect 106 -629 112 -595
rect 146 -629 152 -595
rect 106 -667 152 -629
rect 106 -701 112 -667
rect 146 -701 152 -667
rect 106 -736 152 -701
<< end >>
