magic
tech sky130A
magscale 1 2
timestamp 1666907867
<< error_p >>
rect -372 1053 -314 1059
rect -176 1053 -118 1059
rect 20 1053 78 1059
rect 216 1053 274 1059
rect 412 1053 470 1059
rect -372 1019 -360 1053
rect -176 1019 -164 1053
rect 20 1019 32 1053
rect 216 1019 228 1053
rect 412 1019 424 1053
rect -372 1013 -314 1019
rect -176 1013 -118 1019
rect 20 1013 78 1019
rect 216 1013 274 1019
rect 412 1013 470 1019
rect -555 710 555 890
rect -555 672 457 710
rect -470 617 -412 623
rect -274 617 -216 623
rect -78 617 -20 623
rect 118 617 176 623
rect 314 617 372 623
rect -470 583 -458 617
rect -274 583 -262 617
rect -78 583 -66 617
rect 118 583 130 617
rect 314 583 326 617
rect -470 577 -412 583
rect -274 577 -216 583
rect -78 577 -20 583
rect 118 577 176 583
rect 314 577 372 583
rect -555 274 555 454
rect -457 236 555 274
rect -372 181 -314 187
rect -176 181 -118 187
rect 20 181 78 187
rect 216 181 274 187
rect 412 181 470 187
rect -372 147 -360 181
rect -176 147 -164 181
rect 20 147 32 181
rect 216 147 228 181
rect 412 147 424 181
rect -372 141 -314 147
rect -176 141 -118 147
rect 20 141 78 147
rect 216 141 274 147
rect 412 141 470 147
rect -555 -162 555 18
rect -555 -200 457 -162
rect -470 -255 -412 -249
rect -274 -255 -216 -249
rect -78 -255 -20 -249
rect 118 -255 176 -249
rect 314 -255 372 -249
rect -470 -289 -458 -255
rect -274 -289 -262 -255
rect -78 -289 -66 -255
rect 118 -289 130 -255
rect 314 -289 326 -255
rect -470 -295 -412 -289
rect -274 -295 -216 -289
rect -78 -295 -20 -289
rect 118 -295 176 -289
rect 314 -295 372 -289
rect -555 -598 555 -418
rect -457 -636 555 -598
rect -372 -691 -314 -685
rect -176 -691 -118 -685
rect 20 -691 78 -685
rect 216 -691 274 -685
rect 412 -691 470 -685
rect -372 -725 -360 -691
rect -176 -725 -164 -691
rect 20 -725 32 -691
rect 216 -725 228 -691
rect 412 -725 424 -691
rect -372 -731 -314 -725
rect -176 -731 -118 -725
rect 20 -731 78 -725
rect 216 -731 274 -725
rect 412 -731 470 -725
rect -470 -1019 -412 -1013
rect -274 -1019 -216 -1013
rect -78 -1019 -20 -1013
rect 118 -1019 176 -1013
rect 314 -1019 372 -1013
rect -470 -1053 -458 -1019
rect -274 -1053 -262 -1019
rect -78 -1053 -66 -1019
rect 118 -1053 130 -1019
rect 314 -1053 326 -1019
rect -470 -1059 -412 -1053
rect -274 -1059 -216 -1053
rect -78 -1059 -20 -1053
rect 118 -1059 176 -1053
rect 314 -1059 372 -1053
<< nwell >>
rect -457 1034 555 1072
rect -555 710 555 1034
rect -555 672 457 710
rect -555 598 457 636
rect -555 274 555 598
rect -457 236 555 274
rect -457 162 555 200
rect -555 -162 555 162
rect -555 -200 457 -162
rect -555 -274 457 -236
rect -555 -598 555 -274
rect -457 -636 555 -598
rect -457 -710 555 -672
rect -555 -1034 555 -710
rect -555 -1072 457 -1034
<< pmos >>
rect -461 772 -421 972
rect -363 772 -323 972
rect -265 772 -225 972
rect -167 772 -127 972
rect -69 772 -29 972
rect 29 772 69 972
rect 127 772 167 972
rect 225 772 265 972
rect 323 772 363 972
rect 421 772 461 972
rect -461 336 -421 536
rect -363 336 -323 536
rect -265 336 -225 536
rect -167 336 -127 536
rect -69 336 -29 536
rect 29 336 69 536
rect 127 336 167 536
rect 225 336 265 536
rect 323 336 363 536
rect 421 336 461 536
rect -461 -100 -421 100
rect -363 -100 -323 100
rect -265 -100 -225 100
rect -167 -100 -127 100
rect -69 -100 -29 100
rect 29 -100 69 100
rect 127 -100 167 100
rect 225 -100 265 100
rect 323 -100 363 100
rect 421 -100 461 100
rect -461 -536 -421 -336
rect -363 -536 -323 -336
rect -265 -536 -225 -336
rect -167 -536 -127 -336
rect -69 -536 -29 -336
rect 29 -536 69 -336
rect 127 -536 167 -336
rect 225 -536 265 -336
rect 323 -536 363 -336
rect 421 -536 461 -336
rect -461 -972 -421 -772
rect -363 -972 -323 -772
rect -265 -972 -225 -772
rect -167 -972 -127 -772
rect -69 -972 -29 -772
rect 29 -972 69 -772
rect 127 -972 167 -772
rect 225 -972 265 -772
rect 323 -972 363 -772
rect 421 -972 461 -772
<< pdiff >>
rect -519 960 -461 972
rect -519 784 -507 960
rect -473 784 -461 960
rect -519 772 -461 784
rect -421 960 -363 972
rect -421 784 -409 960
rect -375 784 -363 960
rect -421 772 -363 784
rect -323 960 -265 972
rect -323 784 -311 960
rect -277 784 -265 960
rect -323 772 -265 784
rect -225 960 -167 972
rect -225 784 -213 960
rect -179 784 -167 960
rect -225 772 -167 784
rect -127 960 -69 972
rect -127 784 -115 960
rect -81 784 -69 960
rect -127 772 -69 784
rect -29 960 29 972
rect -29 784 -17 960
rect 17 784 29 960
rect -29 772 29 784
rect 69 960 127 972
rect 69 784 81 960
rect 115 784 127 960
rect 69 772 127 784
rect 167 960 225 972
rect 167 784 179 960
rect 213 784 225 960
rect 167 772 225 784
rect 265 960 323 972
rect 265 784 277 960
rect 311 784 323 960
rect 265 772 323 784
rect 363 960 421 972
rect 363 784 375 960
rect 409 784 421 960
rect 363 772 421 784
rect 461 960 519 972
rect 461 784 473 960
rect 507 784 519 960
rect 461 772 519 784
rect -519 524 -461 536
rect -519 348 -507 524
rect -473 348 -461 524
rect -519 336 -461 348
rect -421 524 -363 536
rect -421 348 -409 524
rect -375 348 -363 524
rect -421 336 -363 348
rect -323 524 -265 536
rect -323 348 -311 524
rect -277 348 -265 524
rect -323 336 -265 348
rect -225 524 -167 536
rect -225 348 -213 524
rect -179 348 -167 524
rect -225 336 -167 348
rect -127 524 -69 536
rect -127 348 -115 524
rect -81 348 -69 524
rect -127 336 -69 348
rect -29 524 29 536
rect -29 348 -17 524
rect 17 348 29 524
rect -29 336 29 348
rect 69 524 127 536
rect 69 348 81 524
rect 115 348 127 524
rect 69 336 127 348
rect 167 524 225 536
rect 167 348 179 524
rect 213 348 225 524
rect 167 336 225 348
rect 265 524 323 536
rect 265 348 277 524
rect 311 348 323 524
rect 265 336 323 348
rect 363 524 421 536
rect 363 348 375 524
rect 409 348 421 524
rect 363 336 421 348
rect 461 524 519 536
rect 461 348 473 524
rect 507 348 519 524
rect 461 336 519 348
rect -519 88 -461 100
rect -519 -88 -507 88
rect -473 -88 -461 88
rect -519 -100 -461 -88
rect -421 88 -363 100
rect -421 -88 -409 88
rect -375 -88 -363 88
rect -421 -100 -363 -88
rect -323 88 -265 100
rect -323 -88 -311 88
rect -277 -88 -265 88
rect -323 -100 -265 -88
rect -225 88 -167 100
rect -225 -88 -213 88
rect -179 -88 -167 88
rect -225 -100 -167 -88
rect -127 88 -69 100
rect -127 -88 -115 88
rect -81 -88 -69 88
rect -127 -100 -69 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 69 88 127 100
rect 69 -88 81 88
rect 115 -88 127 88
rect 69 -100 127 -88
rect 167 88 225 100
rect 167 -88 179 88
rect 213 -88 225 88
rect 167 -100 225 -88
rect 265 88 323 100
rect 265 -88 277 88
rect 311 -88 323 88
rect 265 -100 323 -88
rect 363 88 421 100
rect 363 -88 375 88
rect 409 -88 421 88
rect 363 -100 421 -88
rect 461 88 519 100
rect 461 -88 473 88
rect 507 -88 519 88
rect 461 -100 519 -88
rect -519 -348 -461 -336
rect -519 -524 -507 -348
rect -473 -524 -461 -348
rect -519 -536 -461 -524
rect -421 -348 -363 -336
rect -421 -524 -409 -348
rect -375 -524 -363 -348
rect -421 -536 -363 -524
rect -323 -348 -265 -336
rect -323 -524 -311 -348
rect -277 -524 -265 -348
rect -323 -536 -265 -524
rect -225 -348 -167 -336
rect -225 -524 -213 -348
rect -179 -524 -167 -348
rect -225 -536 -167 -524
rect -127 -348 -69 -336
rect -127 -524 -115 -348
rect -81 -524 -69 -348
rect -127 -536 -69 -524
rect -29 -348 29 -336
rect -29 -524 -17 -348
rect 17 -524 29 -348
rect -29 -536 29 -524
rect 69 -348 127 -336
rect 69 -524 81 -348
rect 115 -524 127 -348
rect 69 -536 127 -524
rect 167 -348 225 -336
rect 167 -524 179 -348
rect 213 -524 225 -348
rect 167 -536 225 -524
rect 265 -348 323 -336
rect 265 -524 277 -348
rect 311 -524 323 -348
rect 265 -536 323 -524
rect 363 -348 421 -336
rect 363 -524 375 -348
rect 409 -524 421 -348
rect 363 -536 421 -524
rect 461 -348 519 -336
rect 461 -524 473 -348
rect 507 -524 519 -348
rect 461 -536 519 -524
rect -519 -784 -461 -772
rect -519 -960 -507 -784
rect -473 -960 -461 -784
rect -519 -972 -461 -960
rect -421 -784 -363 -772
rect -421 -960 -409 -784
rect -375 -960 -363 -784
rect -421 -972 -363 -960
rect -323 -784 -265 -772
rect -323 -960 -311 -784
rect -277 -960 -265 -784
rect -323 -972 -265 -960
rect -225 -784 -167 -772
rect -225 -960 -213 -784
rect -179 -960 -167 -784
rect -225 -972 -167 -960
rect -127 -784 -69 -772
rect -127 -960 -115 -784
rect -81 -960 -69 -784
rect -127 -972 -69 -960
rect -29 -784 29 -772
rect -29 -960 -17 -784
rect 17 -960 29 -784
rect -29 -972 29 -960
rect 69 -784 127 -772
rect 69 -960 81 -784
rect 115 -960 127 -784
rect 69 -972 127 -960
rect 167 -784 225 -772
rect 167 -960 179 -784
rect 213 -960 225 -784
rect 167 -972 225 -960
rect 265 -784 323 -772
rect 265 -960 277 -784
rect 311 -960 323 -784
rect 265 -972 323 -960
rect 363 -784 421 -772
rect 363 -960 375 -784
rect 409 -960 421 -784
rect 363 -972 421 -960
rect 461 -784 519 -772
rect 461 -960 473 -784
rect 507 -960 519 -784
rect 461 -972 519 -960
<< pdiffc >>
rect -507 784 -473 960
rect -409 784 -375 960
rect -311 784 -277 960
rect -213 784 -179 960
rect -115 784 -81 960
rect -17 784 17 960
rect 81 784 115 960
rect 179 784 213 960
rect 277 784 311 960
rect 375 784 409 960
rect 473 784 507 960
rect -507 348 -473 524
rect -409 348 -375 524
rect -311 348 -277 524
rect -213 348 -179 524
rect -115 348 -81 524
rect -17 348 17 524
rect 81 348 115 524
rect 179 348 213 524
rect 277 348 311 524
rect 375 348 409 524
rect 473 348 507 524
rect -507 -88 -473 88
rect -409 -88 -375 88
rect -311 -88 -277 88
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
rect 277 -88 311 88
rect 375 -88 409 88
rect 473 -88 507 88
rect -507 -524 -473 -348
rect -409 -524 -375 -348
rect -311 -524 -277 -348
rect -213 -524 -179 -348
rect -115 -524 -81 -348
rect -17 -524 17 -348
rect 81 -524 115 -348
rect 179 -524 213 -348
rect 277 -524 311 -348
rect 375 -524 409 -348
rect 473 -524 507 -348
rect -507 -960 -473 -784
rect -409 -960 -375 -784
rect -311 -960 -277 -784
rect -213 -960 -179 -784
rect -115 -960 -81 -784
rect -17 -960 17 -784
rect 81 -960 115 -784
rect 179 -960 213 -784
rect 277 -960 311 -784
rect 375 -960 409 -784
rect 473 -960 507 -784
<< poly >>
rect -376 1053 -310 1069
rect -376 1019 -360 1053
rect -326 1019 -310 1053
rect -376 1003 -310 1019
rect -180 1053 -114 1069
rect -180 1019 -164 1053
rect -130 1019 -114 1053
rect -180 1003 -114 1019
rect 16 1053 82 1069
rect 16 1019 32 1053
rect 66 1019 82 1053
rect 16 1003 82 1019
rect 212 1053 278 1069
rect 212 1019 228 1053
rect 262 1019 278 1053
rect 212 1003 278 1019
rect 408 1053 474 1069
rect 408 1019 424 1053
rect 458 1019 474 1053
rect 408 1003 474 1019
rect -461 972 -421 998
rect -363 972 -323 1003
rect -265 972 -225 998
rect -167 972 -127 1003
rect -69 972 -29 998
rect 29 972 69 1003
rect 127 972 167 998
rect 225 972 265 1003
rect 323 972 363 998
rect 421 972 461 1003
rect -461 741 -421 772
rect -363 746 -323 772
rect -265 741 -225 772
rect -167 746 -127 772
rect -69 741 -29 772
rect 29 746 69 772
rect 127 741 167 772
rect 225 746 265 772
rect 323 741 363 772
rect 421 746 461 772
rect -474 725 -408 741
rect -474 691 -458 725
rect -424 691 -408 725
rect -474 675 -408 691
rect -278 725 -212 741
rect -278 691 -262 725
rect -228 691 -212 725
rect -278 675 -212 691
rect -82 725 -16 741
rect -82 691 -66 725
rect -32 691 -16 725
rect -82 675 -16 691
rect 114 725 180 741
rect 114 691 130 725
rect 164 691 180 725
rect 114 675 180 691
rect 310 725 376 741
rect 310 691 326 725
rect 360 691 376 725
rect 310 675 376 691
rect -474 617 -408 633
rect -474 583 -458 617
rect -424 583 -408 617
rect -474 567 -408 583
rect -278 617 -212 633
rect -278 583 -262 617
rect -228 583 -212 617
rect -278 567 -212 583
rect -82 617 -16 633
rect -82 583 -66 617
rect -32 583 -16 617
rect -82 567 -16 583
rect 114 617 180 633
rect 114 583 130 617
rect 164 583 180 617
rect 114 567 180 583
rect 310 617 376 633
rect 310 583 326 617
rect 360 583 376 617
rect 310 567 376 583
rect -461 536 -421 567
rect -363 536 -323 562
rect -265 536 -225 567
rect -167 536 -127 562
rect -69 536 -29 567
rect 29 536 69 562
rect 127 536 167 567
rect 225 536 265 562
rect 323 536 363 567
rect 421 536 461 562
rect -461 310 -421 336
rect -363 305 -323 336
rect -265 310 -225 336
rect -167 305 -127 336
rect -69 310 -29 336
rect 29 305 69 336
rect 127 310 167 336
rect 225 305 265 336
rect 323 310 363 336
rect 421 305 461 336
rect -376 289 -310 305
rect -376 255 -360 289
rect -326 255 -310 289
rect -376 239 -310 255
rect -180 289 -114 305
rect -180 255 -164 289
rect -130 255 -114 289
rect -180 239 -114 255
rect 16 289 82 305
rect 16 255 32 289
rect 66 255 82 289
rect 16 239 82 255
rect 212 289 278 305
rect 212 255 228 289
rect 262 255 278 289
rect 212 239 278 255
rect 408 289 474 305
rect 408 255 424 289
rect 458 255 474 289
rect 408 239 474 255
rect -376 181 -310 197
rect -376 147 -360 181
rect -326 147 -310 181
rect -376 131 -310 147
rect -180 181 -114 197
rect -180 147 -164 181
rect -130 147 -114 181
rect -180 131 -114 147
rect 16 181 82 197
rect 16 147 32 181
rect 66 147 82 181
rect 16 131 82 147
rect 212 181 278 197
rect 212 147 228 181
rect 262 147 278 181
rect 212 131 278 147
rect 408 181 474 197
rect 408 147 424 181
rect 458 147 474 181
rect 408 131 474 147
rect -461 100 -421 126
rect -363 100 -323 131
rect -265 100 -225 126
rect -167 100 -127 131
rect -69 100 -29 126
rect 29 100 69 131
rect 127 100 167 126
rect 225 100 265 131
rect 323 100 363 126
rect 421 100 461 131
rect -461 -131 -421 -100
rect -363 -126 -323 -100
rect -265 -131 -225 -100
rect -167 -126 -127 -100
rect -69 -131 -29 -100
rect 29 -126 69 -100
rect 127 -131 167 -100
rect 225 -126 265 -100
rect 323 -131 363 -100
rect 421 -126 461 -100
rect -474 -147 -408 -131
rect -474 -181 -458 -147
rect -424 -181 -408 -147
rect -474 -197 -408 -181
rect -278 -147 -212 -131
rect -278 -181 -262 -147
rect -228 -181 -212 -147
rect -278 -197 -212 -181
rect -82 -147 -16 -131
rect -82 -181 -66 -147
rect -32 -181 -16 -147
rect -82 -197 -16 -181
rect 114 -147 180 -131
rect 114 -181 130 -147
rect 164 -181 180 -147
rect 114 -197 180 -181
rect 310 -147 376 -131
rect 310 -181 326 -147
rect 360 -181 376 -147
rect 310 -197 376 -181
rect -474 -255 -408 -239
rect -474 -289 -458 -255
rect -424 -289 -408 -255
rect -474 -305 -408 -289
rect -278 -255 -212 -239
rect -278 -289 -262 -255
rect -228 -289 -212 -255
rect -278 -305 -212 -289
rect -82 -255 -16 -239
rect -82 -289 -66 -255
rect -32 -289 -16 -255
rect -82 -305 -16 -289
rect 114 -255 180 -239
rect 114 -289 130 -255
rect 164 -289 180 -255
rect 114 -305 180 -289
rect 310 -255 376 -239
rect 310 -289 326 -255
rect 360 -289 376 -255
rect 310 -305 376 -289
rect -461 -336 -421 -305
rect -363 -336 -323 -310
rect -265 -336 -225 -305
rect -167 -336 -127 -310
rect -69 -336 -29 -305
rect 29 -336 69 -310
rect 127 -336 167 -305
rect 225 -336 265 -310
rect 323 -336 363 -305
rect 421 -336 461 -310
rect -461 -562 -421 -536
rect -363 -567 -323 -536
rect -265 -562 -225 -536
rect -167 -567 -127 -536
rect -69 -562 -29 -536
rect 29 -567 69 -536
rect 127 -562 167 -536
rect 225 -567 265 -536
rect 323 -562 363 -536
rect 421 -567 461 -536
rect -376 -583 -310 -567
rect -376 -617 -360 -583
rect -326 -617 -310 -583
rect -376 -633 -310 -617
rect -180 -583 -114 -567
rect -180 -617 -164 -583
rect -130 -617 -114 -583
rect -180 -633 -114 -617
rect 16 -583 82 -567
rect 16 -617 32 -583
rect 66 -617 82 -583
rect 16 -633 82 -617
rect 212 -583 278 -567
rect 212 -617 228 -583
rect 262 -617 278 -583
rect 212 -633 278 -617
rect 408 -583 474 -567
rect 408 -617 424 -583
rect 458 -617 474 -583
rect 408 -633 474 -617
rect -376 -691 -310 -675
rect -376 -725 -360 -691
rect -326 -725 -310 -691
rect -376 -741 -310 -725
rect -180 -691 -114 -675
rect -180 -725 -164 -691
rect -130 -725 -114 -691
rect -180 -741 -114 -725
rect 16 -691 82 -675
rect 16 -725 32 -691
rect 66 -725 82 -691
rect 16 -741 82 -725
rect 212 -691 278 -675
rect 212 -725 228 -691
rect 262 -725 278 -691
rect 212 -741 278 -725
rect 408 -691 474 -675
rect 408 -725 424 -691
rect 458 -725 474 -691
rect 408 -741 474 -725
rect -461 -772 -421 -746
rect -363 -772 -323 -741
rect -265 -772 -225 -746
rect -167 -772 -127 -741
rect -69 -772 -29 -746
rect 29 -772 69 -741
rect 127 -772 167 -746
rect 225 -772 265 -741
rect 323 -772 363 -746
rect 421 -772 461 -741
rect -461 -1003 -421 -972
rect -363 -998 -323 -972
rect -265 -1003 -225 -972
rect -167 -998 -127 -972
rect -69 -1003 -29 -972
rect 29 -998 69 -972
rect 127 -1003 167 -972
rect 225 -998 265 -972
rect 323 -1003 363 -972
rect 421 -998 461 -972
rect -474 -1019 -408 -1003
rect -474 -1053 -458 -1019
rect -424 -1053 -408 -1019
rect -474 -1069 -408 -1053
rect -278 -1019 -212 -1003
rect -278 -1053 -262 -1019
rect -228 -1053 -212 -1019
rect -278 -1069 -212 -1053
rect -82 -1019 -16 -1003
rect -82 -1053 -66 -1019
rect -32 -1053 -16 -1019
rect -82 -1069 -16 -1053
rect 114 -1019 180 -1003
rect 114 -1053 130 -1019
rect 164 -1053 180 -1019
rect 114 -1069 180 -1053
rect 310 -1019 376 -1003
rect 310 -1053 326 -1019
rect 360 -1053 376 -1019
rect 310 -1069 376 -1053
<< polycont >>
rect -360 1019 -326 1053
rect -164 1019 -130 1053
rect 32 1019 66 1053
rect 228 1019 262 1053
rect 424 1019 458 1053
rect -458 691 -424 725
rect -262 691 -228 725
rect -66 691 -32 725
rect 130 691 164 725
rect 326 691 360 725
rect -458 583 -424 617
rect -262 583 -228 617
rect -66 583 -32 617
rect 130 583 164 617
rect 326 583 360 617
rect -360 255 -326 289
rect -164 255 -130 289
rect 32 255 66 289
rect 228 255 262 289
rect 424 255 458 289
rect -360 147 -326 181
rect -164 147 -130 181
rect 32 147 66 181
rect 228 147 262 181
rect 424 147 458 181
rect -458 -181 -424 -147
rect -262 -181 -228 -147
rect -66 -181 -32 -147
rect 130 -181 164 -147
rect 326 -181 360 -147
rect -458 -289 -424 -255
rect -262 -289 -228 -255
rect -66 -289 -32 -255
rect 130 -289 164 -255
rect 326 -289 360 -255
rect -360 -617 -326 -583
rect -164 -617 -130 -583
rect 32 -617 66 -583
rect 228 -617 262 -583
rect 424 -617 458 -583
rect -360 -725 -326 -691
rect -164 -725 -130 -691
rect 32 -725 66 -691
rect 228 -725 262 -691
rect 424 -725 458 -691
rect -458 -1053 -424 -1019
rect -262 -1053 -228 -1019
rect -66 -1053 -32 -1019
rect 130 -1053 164 -1019
rect 326 -1053 360 -1019
<< locali >>
rect -376 1019 -360 1053
rect -326 1019 -310 1053
rect -180 1019 -164 1053
rect -130 1019 -114 1053
rect 16 1019 32 1053
rect 66 1019 82 1053
rect 212 1019 228 1053
rect 262 1019 278 1053
rect 408 1019 424 1053
rect 458 1019 474 1053
rect -507 960 -473 976
rect -507 768 -473 784
rect -409 960 -375 976
rect -409 768 -375 784
rect -311 960 -277 976
rect -311 768 -277 784
rect -213 960 -179 976
rect -213 768 -179 784
rect -115 960 -81 976
rect -115 768 -81 784
rect -17 960 17 976
rect -17 768 17 784
rect 81 960 115 976
rect 81 768 115 784
rect 179 960 213 976
rect 179 768 213 784
rect 277 960 311 976
rect 277 768 311 784
rect 375 960 409 976
rect 375 768 409 784
rect 473 960 507 976
rect 473 768 507 784
rect -474 691 -458 725
rect -424 691 -408 725
rect -278 691 -262 725
rect -228 691 -212 725
rect -82 691 -66 725
rect -32 691 -16 725
rect 114 691 130 725
rect 164 691 180 725
rect 310 691 326 725
rect 360 691 376 725
rect -474 583 -458 617
rect -424 583 -408 617
rect -278 583 -262 617
rect -228 583 -212 617
rect -82 583 -66 617
rect -32 583 -16 617
rect 114 583 130 617
rect 164 583 180 617
rect 310 583 326 617
rect 360 583 376 617
rect -507 524 -473 540
rect -507 332 -473 348
rect -409 524 -375 540
rect -409 332 -375 348
rect -311 524 -277 540
rect -311 332 -277 348
rect -213 524 -179 540
rect -213 332 -179 348
rect -115 524 -81 540
rect -115 332 -81 348
rect -17 524 17 540
rect -17 332 17 348
rect 81 524 115 540
rect 81 332 115 348
rect 179 524 213 540
rect 179 332 213 348
rect 277 524 311 540
rect 277 332 311 348
rect 375 524 409 540
rect 375 332 409 348
rect 473 524 507 540
rect 473 332 507 348
rect -376 255 -360 289
rect -326 255 -310 289
rect -180 255 -164 289
rect -130 255 -114 289
rect 16 255 32 289
rect 66 255 82 289
rect 212 255 228 289
rect 262 255 278 289
rect 408 255 424 289
rect 458 255 474 289
rect -376 147 -360 181
rect -326 147 -310 181
rect -180 147 -164 181
rect -130 147 -114 181
rect 16 147 32 181
rect 66 147 82 181
rect 212 147 228 181
rect 262 147 278 181
rect 408 147 424 181
rect 458 147 474 181
rect -507 88 -473 104
rect -507 -104 -473 -88
rect -409 88 -375 104
rect -409 -104 -375 -88
rect -311 88 -277 104
rect -311 -104 -277 -88
rect -213 88 -179 104
rect -213 -104 -179 -88
rect -115 88 -81 104
rect -115 -104 -81 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 81 88 115 104
rect 81 -104 115 -88
rect 179 88 213 104
rect 179 -104 213 -88
rect 277 88 311 104
rect 277 -104 311 -88
rect 375 88 409 104
rect 375 -104 409 -88
rect 473 88 507 104
rect 473 -104 507 -88
rect -474 -181 -458 -147
rect -424 -181 -408 -147
rect -278 -181 -262 -147
rect -228 -181 -212 -147
rect -82 -181 -66 -147
rect -32 -181 -16 -147
rect 114 -181 130 -147
rect 164 -181 180 -147
rect 310 -181 326 -147
rect 360 -181 376 -147
rect -474 -289 -458 -255
rect -424 -289 -408 -255
rect -278 -289 -262 -255
rect -228 -289 -212 -255
rect -82 -289 -66 -255
rect -32 -289 -16 -255
rect 114 -289 130 -255
rect 164 -289 180 -255
rect 310 -289 326 -255
rect 360 -289 376 -255
rect -507 -348 -473 -332
rect -507 -540 -473 -524
rect -409 -348 -375 -332
rect -409 -540 -375 -524
rect -311 -348 -277 -332
rect -311 -540 -277 -524
rect -213 -348 -179 -332
rect -213 -540 -179 -524
rect -115 -348 -81 -332
rect -115 -540 -81 -524
rect -17 -348 17 -332
rect -17 -540 17 -524
rect 81 -348 115 -332
rect 81 -540 115 -524
rect 179 -348 213 -332
rect 179 -540 213 -524
rect 277 -348 311 -332
rect 277 -540 311 -524
rect 375 -348 409 -332
rect 375 -540 409 -524
rect 473 -348 507 -332
rect 473 -540 507 -524
rect -376 -617 -360 -583
rect -326 -617 -310 -583
rect -180 -617 -164 -583
rect -130 -617 -114 -583
rect 16 -617 32 -583
rect 66 -617 82 -583
rect 212 -617 228 -583
rect 262 -617 278 -583
rect 408 -617 424 -583
rect 458 -617 474 -583
rect -376 -725 -360 -691
rect -326 -725 -310 -691
rect -180 -725 -164 -691
rect -130 -725 -114 -691
rect 16 -725 32 -691
rect 66 -725 82 -691
rect 212 -725 228 -691
rect 262 -725 278 -691
rect 408 -725 424 -691
rect 458 -725 474 -691
rect -507 -784 -473 -768
rect -507 -976 -473 -960
rect -409 -784 -375 -768
rect -409 -976 -375 -960
rect -311 -784 -277 -768
rect -311 -976 -277 -960
rect -213 -784 -179 -768
rect -213 -976 -179 -960
rect -115 -784 -81 -768
rect -115 -976 -81 -960
rect -17 -784 17 -768
rect -17 -976 17 -960
rect 81 -784 115 -768
rect 81 -976 115 -960
rect 179 -784 213 -768
rect 179 -976 213 -960
rect 277 -784 311 -768
rect 277 -976 311 -960
rect 375 -784 409 -768
rect 375 -976 409 -960
rect 473 -784 507 -768
rect 473 -976 507 -960
rect -474 -1053 -458 -1019
rect -424 -1053 -408 -1019
rect -278 -1053 -262 -1019
rect -228 -1053 -212 -1019
rect -82 -1053 -66 -1019
rect -32 -1053 -16 -1019
rect 114 -1053 130 -1019
rect 164 -1053 180 -1019
rect 310 -1053 326 -1019
rect 360 -1053 376 -1019
<< viali >>
rect -360 1019 -326 1053
rect -164 1019 -130 1053
rect 32 1019 66 1053
rect 228 1019 262 1053
rect 424 1019 458 1053
rect -507 784 -473 960
rect -409 784 -375 960
rect -311 784 -277 960
rect -213 784 -179 960
rect -115 784 -81 960
rect -17 784 17 960
rect 81 784 115 960
rect 179 784 213 960
rect 277 784 311 960
rect 375 784 409 960
rect 473 784 507 960
rect -458 691 -424 725
rect -262 691 -228 725
rect -66 691 -32 725
rect 130 691 164 725
rect 326 691 360 725
rect -458 583 -424 617
rect -262 583 -228 617
rect -66 583 -32 617
rect 130 583 164 617
rect 326 583 360 617
rect -507 348 -473 524
rect -409 348 -375 524
rect -311 348 -277 524
rect -213 348 -179 524
rect -115 348 -81 524
rect -17 348 17 524
rect 81 348 115 524
rect 179 348 213 524
rect 277 348 311 524
rect 375 348 409 524
rect 473 348 507 524
rect -360 255 -326 289
rect -164 255 -130 289
rect 32 255 66 289
rect 228 255 262 289
rect 424 255 458 289
rect -360 147 -326 181
rect -164 147 -130 181
rect 32 147 66 181
rect 228 147 262 181
rect 424 147 458 181
rect -507 -88 -473 88
rect -409 -88 -375 88
rect -311 -88 -277 88
rect -213 -88 -179 88
rect -115 -88 -81 88
rect -17 -88 17 88
rect 81 -88 115 88
rect 179 -88 213 88
rect 277 -88 311 88
rect 375 -88 409 88
rect 473 -88 507 88
rect -458 -181 -424 -147
rect -262 -181 -228 -147
rect -66 -181 -32 -147
rect 130 -181 164 -147
rect 326 -181 360 -147
rect -458 -289 -424 -255
rect -262 -289 -228 -255
rect -66 -289 -32 -255
rect 130 -289 164 -255
rect 326 -289 360 -255
rect -507 -524 -473 -348
rect -409 -524 -375 -348
rect -311 -524 -277 -348
rect -213 -524 -179 -348
rect -115 -524 -81 -348
rect -17 -524 17 -348
rect 81 -524 115 -348
rect 179 -524 213 -348
rect 277 -524 311 -348
rect 375 -524 409 -348
rect 473 -524 507 -348
rect -360 -617 -326 -583
rect -164 -617 -130 -583
rect 32 -617 66 -583
rect 228 -617 262 -583
rect 424 -617 458 -583
rect -360 -725 -326 -691
rect -164 -725 -130 -691
rect 32 -725 66 -691
rect 228 -725 262 -691
rect 424 -725 458 -691
rect -507 -960 -473 -784
rect -409 -960 -375 -784
rect -311 -960 -277 -784
rect -213 -960 -179 -784
rect -115 -960 -81 -784
rect -17 -960 17 -784
rect 81 -960 115 -784
rect 179 -960 213 -784
rect 277 -960 311 -784
rect 375 -960 409 -784
rect 473 -960 507 -784
rect -458 -1053 -424 -1019
rect -262 -1053 -228 -1019
rect -66 -1053 -32 -1019
rect 130 -1053 164 -1019
rect 326 -1053 360 -1019
<< metal1 >>
rect -372 1053 -314 1059
rect -372 1019 -360 1053
rect -326 1019 -314 1053
rect -372 1013 -314 1019
rect -176 1053 -118 1059
rect -176 1019 -164 1053
rect -130 1019 -118 1053
rect -176 1013 -118 1019
rect 20 1053 78 1059
rect 20 1019 32 1053
rect 66 1019 78 1053
rect 20 1013 78 1019
rect 216 1053 274 1059
rect 216 1019 228 1053
rect 262 1019 274 1053
rect 216 1013 274 1019
rect 412 1053 470 1059
rect 412 1019 424 1053
rect 458 1019 470 1053
rect 412 1013 470 1019
rect -513 960 -467 972
rect -513 784 -507 960
rect -473 784 -467 960
rect -513 772 -467 784
rect -415 960 -369 972
rect -415 784 -409 960
rect -375 784 -369 960
rect -415 772 -369 784
rect -317 960 -271 972
rect -317 784 -311 960
rect -277 784 -271 960
rect -317 772 -271 784
rect -219 960 -173 972
rect -219 784 -213 960
rect -179 784 -173 960
rect -219 772 -173 784
rect -121 960 -75 972
rect -121 784 -115 960
rect -81 784 -75 960
rect -121 772 -75 784
rect -23 960 23 972
rect -23 784 -17 960
rect 17 784 23 960
rect -23 772 23 784
rect 75 960 121 972
rect 75 784 81 960
rect 115 784 121 960
rect 75 772 121 784
rect 173 960 219 972
rect 173 784 179 960
rect 213 784 219 960
rect 173 772 219 784
rect 271 960 317 972
rect 271 784 277 960
rect 311 784 317 960
rect 271 772 317 784
rect 369 960 415 972
rect 369 784 375 960
rect 409 784 415 960
rect 369 772 415 784
rect 467 960 513 972
rect 467 784 473 960
rect 507 784 513 960
rect 467 772 513 784
rect -470 725 -412 731
rect -470 691 -458 725
rect -424 691 -412 725
rect -470 685 -412 691
rect -274 725 -216 731
rect -274 691 -262 725
rect -228 691 -216 725
rect -274 685 -216 691
rect -78 725 -20 731
rect -78 691 -66 725
rect -32 691 -20 725
rect -78 685 -20 691
rect 118 725 176 731
rect 118 691 130 725
rect 164 691 176 725
rect 118 685 176 691
rect 314 725 372 731
rect 314 691 326 725
rect 360 691 372 725
rect 314 685 372 691
rect -470 617 -412 623
rect -470 583 -458 617
rect -424 583 -412 617
rect -470 577 -412 583
rect -274 617 -216 623
rect -274 583 -262 617
rect -228 583 -216 617
rect -274 577 -216 583
rect -78 617 -20 623
rect -78 583 -66 617
rect -32 583 -20 617
rect -78 577 -20 583
rect 118 617 176 623
rect 118 583 130 617
rect 164 583 176 617
rect 118 577 176 583
rect 314 617 372 623
rect 314 583 326 617
rect 360 583 372 617
rect 314 577 372 583
rect -513 524 -467 536
rect -513 348 -507 524
rect -473 348 -467 524
rect -513 336 -467 348
rect -415 524 -369 536
rect -415 348 -409 524
rect -375 348 -369 524
rect -415 336 -369 348
rect -317 524 -271 536
rect -317 348 -311 524
rect -277 348 -271 524
rect -317 336 -271 348
rect -219 524 -173 536
rect -219 348 -213 524
rect -179 348 -173 524
rect -219 336 -173 348
rect -121 524 -75 536
rect -121 348 -115 524
rect -81 348 -75 524
rect -121 336 -75 348
rect -23 524 23 536
rect -23 348 -17 524
rect 17 348 23 524
rect -23 336 23 348
rect 75 524 121 536
rect 75 348 81 524
rect 115 348 121 524
rect 75 336 121 348
rect 173 524 219 536
rect 173 348 179 524
rect 213 348 219 524
rect 173 336 219 348
rect 271 524 317 536
rect 271 348 277 524
rect 311 348 317 524
rect 271 336 317 348
rect 369 524 415 536
rect 369 348 375 524
rect 409 348 415 524
rect 369 336 415 348
rect 467 524 513 536
rect 467 348 473 524
rect 507 348 513 524
rect 467 336 513 348
rect -372 289 -314 295
rect -372 255 -360 289
rect -326 255 -314 289
rect -372 249 -314 255
rect -176 289 -118 295
rect -176 255 -164 289
rect -130 255 -118 289
rect -176 249 -118 255
rect 20 289 78 295
rect 20 255 32 289
rect 66 255 78 289
rect 20 249 78 255
rect 216 289 274 295
rect 216 255 228 289
rect 262 255 274 289
rect 216 249 274 255
rect 412 289 470 295
rect 412 255 424 289
rect 458 255 470 289
rect 412 249 470 255
rect -372 181 -314 187
rect -372 147 -360 181
rect -326 147 -314 181
rect -372 141 -314 147
rect -176 181 -118 187
rect -176 147 -164 181
rect -130 147 -118 181
rect -176 141 -118 147
rect 20 181 78 187
rect 20 147 32 181
rect 66 147 78 181
rect 20 141 78 147
rect 216 181 274 187
rect 216 147 228 181
rect 262 147 274 181
rect 216 141 274 147
rect 412 181 470 187
rect 412 147 424 181
rect 458 147 470 181
rect 412 141 470 147
rect -513 88 -467 100
rect -513 -88 -507 88
rect -473 -88 -467 88
rect -513 -100 -467 -88
rect -415 88 -369 100
rect -415 -88 -409 88
rect -375 -88 -369 88
rect -415 -100 -369 -88
rect -317 88 -271 100
rect -317 -88 -311 88
rect -277 -88 -271 88
rect -317 -100 -271 -88
rect -219 88 -173 100
rect -219 -88 -213 88
rect -179 -88 -173 88
rect -219 -100 -173 -88
rect -121 88 -75 100
rect -121 -88 -115 88
rect -81 -88 -75 88
rect -121 -100 -75 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 75 88 121 100
rect 75 -88 81 88
rect 115 -88 121 88
rect 75 -100 121 -88
rect 173 88 219 100
rect 173 -88 179 88
rect 213 -88 219 88
rect 173 -100 219 -88
rect 271 88 317 100
rect 271 -88 277 88
rect 311 -88 317 88
rect 271 -100 317 -88
rect 369 88 415 100
rect 369 -88 375 88
rect 409 -88 415 88
rect 369 -100 415 -88
rect 467 88 513 100
rect 467 -88 473 88
rect 507 -88 513 88
rect 467 -100 513 -88
rect -470 -147 -412 -141
rect -470 -181 -458 -147
rect -424 -181 -412 -147
rect -470 -187 -412 -181
rect -274 -147 -216 -141
rect -274 -181 -262 -147
rect -228 -181 -216 -147
rect -274 -187 -216 -181
rect -78 -147 -20 -141
rect -78 -181 -66 -147
rect -32 -181 -20 -147
rect -78 -187 -20 -181
rect 118 -147 176 -141
rect 118 -181 130 -147
rect 164 -181 176 -147
rect 118 -187 176 -181
rect 314 -147 372 -141
rect 314 -181 326 -147
rect 360 -181 372 -147
rect 314 -187 372 -181
rect -470 -255 -412 -249
rect -470 -289 -458 -255
rect -424 -289 -412 -255
rect -470 -295 -412 -289
rect -274 -255 -216 -249
rect -274 -289 -262 -255
rect -228 -289 -216 -255
rect -274 -295 -216 -289
rect -78 -255 -20 -249
rect -78 -289 -66 -255
rect -32 -289 -20 -255
rect -78 -295 -20 -289
rect 118 -255 176 -249
rect 118 -289 130 -255
rect 164 -289 176 -255
rect 118 -295 176 -289
rect 314 -255 372 -249
rect 314 -289 326 -255
rect 360 -289 372 -255
rect 314 -295 372 -289
rect -513 -348 -467 -336
rect -513 -524 -507 -348
rect -473 -524 -467 -348
rect -513 -536 -467 -524
rect -415 -348 -369 -336
rect -415 -524 -409 -348
rect -375 -524 -369 -348
rect -415 -536 -369 -524
rect -317 -348 -271 -336
rect -317 -524 -311 -348
rect -277 -524 -271 -348
rect -317 -536 -271 -524
rect -219 -348 -173 -336
rect -219 -524 -213 -348
rect -179 -524 -173 -348
rect -219 -536 -173 -524
rect -121 -348 -75 -336
rect -121 -524 -115 -348
rect -81 -524 -75 -348
rect -121 -536 -75 -524
rect -23 -348 23 -336
rect -23 -524 -17 -348
rect 17 -524 23 -348
rect -23 -536 23 -524
rect 75 -348 121 -336
rect 75 -524 81 -348
rect 115 -524 121 -348
rect 75 -536 121 -524
rect 173 -348 219 -336
rect 173 -524 179 -348
rect 213 -524 219 -348
rect 173 -536 219 -524
rect 271 -348 317 -336
rect 271 -524 277 -348
rect 311 -524 317 -348
rect 271 -536 317 -524
rect 369 -348 415 -336
rect 369 -524 375 -348
rect 409 -524 415 -348
rect 369 -536 415 -524
rect 467 -348 513 -336
rect 467 -524 473 -348
rect 507 -524 513 -348
rect 467 -536 513 -524
rect -372 -583 -314 -577
rect -372 -617 -360 -583
rect -326 -617 -314 -583
rect -372 -623 -314 -617
rect -176 -583 -118 -577
rect -176 -617 -164 -583
rect -130 -617 -118 -583
rect -176 -623 -118 -617
rect 20 -583 78 -577
rect 20 -617 32 -583
rect 66 -617 78 -583
rect 20 -623 78 -617
rect 216 -583 274 -577
rect 216 -617 228 -583
rect 262 -617 274 -583
rect 216 -623 274 -617
rect 412 -583 470 -577
rect 412 -617 424 -583
rect 458 -617 470 -583
rect 412 -623 470 -617
rect -372 -691 -314 -685
rect -372 -725 -360 -691
rect -326 -725 -314 -691
rect -372 -731 -314 -725
rect -176 -691 -118 -685
rect -176 -725 -164 -691
rect -130 -725 -118 -691
rect -176 -731 -118 -725
rect 20 -691 78 -685
rect 20 -725 32 -691
rect 66 -725 78 -691
rect 20 -731 78 -725
rect 216 -691 274 -685
rect 216 -725 228 -691
rect 262 -725 274 -691
rect 216 -731 274 -725
rect 412 -691 470 -685
rect 412 -725 424 -691
rect 458 -725 470 -691
rect 412 -731 470 -725
rect -513 -784 -467 -772
rect -513 -960 -507 -784
rect -473 -960 -467 -784
rect -513 -972 -467 -960
rect -415 -784 -369 -772
rect -415 -960 -409 -784
rect -375 -960 -369 -784
rect -415 -972 -369 -960
rect -317 -784 -271 -772
rect -317 -960 -311 -784
rect -277 -960 -271 -784
rect -317 -972 -271 -960
rect -219 -784 -173 -772
rect -219 -960 -213 -784
rect -179 -960 -173 -784
rect -219 -972 -173 -960
rect -121 -784 -75 -772
rect -121 -960 -115 -784
rect -81 -960 -75 -784
rect -121 -972 -75 -960
rect -23 -784 23 -772
rect -23 -960 -17 -784
rect 17 -960 23 -784
rect -23 -972 23 -960
rect 75 -784 121 -772
rect 75 -960 81 -784
rect 115 -960 121 -784
rect 75 -972 121 -960
rect 173 -784 219 -772
rect 173 -960 179 -784
rect 213 -960 219 -784
rect 173 -972 219 -960
rect 271 -784 317 -772
rect 271 -960 277 -784
rect 311 -960 317 -784
rect 271 -972 317 -960
rect 369 -784 415 -772
rect 369 -960 375 -784
rect 409 -960 415 -784
rect 369 -972 415 -960
rect 467 -784 513 -772
rect 467 -960 473 -784
rect 507 -960 513 -784
rect 467 -972 513 -960
rect -470 -1019 -412 -1013
rect -470 -1053 -458 -1019
rect -424 -1053 -412 -1019
rect -470 -1059 -412 -1053
rect -274 -1019 -216 -1013
rect -274 -1053 -262 -1019
rect -228 -1053 -216 -1019
rect -274 -1059 -216 -1053
rect -78 -1019 -20 -1013
rect -78 -1053 -66 -1019
rect -32 -1053 -20 -1019
rect -78 -1059 -20 -1053
rect 118 -1019 176 -1013
rect 118 -1053 130 -1019
rect 164 -1053 176 -1019
rect 118 -1059 176 -1053
rect 314 -1019 372 -1013
rect 314 -1053 326 -1019
rect 360 -1053 372 -1019
rect 314 -1059 372 -1053
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.2 m 5 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
