magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal4 >>
rect 5400 -7132 6400 4717
rect 5400 -7368 5532 -7132
rect 5768 -7368 5932 -7132
rect 6168 -7368 6400 -7132
rect 5400 -7532 6400 -7368
rect 5400 -7768 5632 -7532
rect 5868 -7768 6032 -7532
rect 6268 -7768 6400 -7532
rect 5400 -8000 6400 -7768
<< via4 >>
rect 5532 -7368 5768 -7132
rect 5932 -7368 6168 -7132
rect 5632 -7768 5868 -7532
rect 6032 -7768 6268 -7532
<< metal5 >>
rect -4800 3200 26200 4200
rect -4200 1600 24600 2600
rect -4200 -25200 -3200 1600
rect -2600 0 23000 1000
rect -2600 -23600 -1600 0
rect -1000 -1600 21400 -600
rect -1000 -22000 0 -1600
rect 600 -3200 19800 -2200
rect 600 -20400 1600 -3200
rect 2200 -4800 18200 -3800
rect 2200 -18800 3200 -4800
rect 3800 -6400 16600 -5400
rect 3800 -17200 4800 -6400
rect 5400 -7132 6400 -7000
rect 5400 -7368 5532 -7132
rect 5768 -7368 5932 -7132
rect 6168 -7368 6400 -7132
rect 5400 -7532 6400 -7368
rect 5400 -7768 5632 -7532
rect 5868 -7768 6032 -7532
rect 6268 -7768 6400 -7532
rect 5400 -15600 6400 -7768
rect 15600 -15600 16600 -6400
rect 5400 -16600 16600 -15600
rect 17200 -17200 18200 -4800
rect 3800 -18200 18200 -17200
rect 18800 -18800 19800 -3200
rect 2200 -19800 19800 -18800
rect 20400 -20400 21400 -1600
rect 600 -21400 21400 -20400
rect 22000 -22000 23000 0
rect -1000 -23000 23000 -22000
rect 23600 -23600 24600 1600
rect -2600 -24600 24600 -23600
rect 25200 -25200 26200 3200
rect -4200 -26200 26200 -25200
<< end >>
