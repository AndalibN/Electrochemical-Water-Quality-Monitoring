magic
tech sky130A
timestamp 1668786957
<< metal5 >>
rect -1750 2100 -650 2300
rect 0 2100 1100 2300
rect -1750 -300 -1550 2100
rect -1350 1700 -650 1900
rect 0 1700 700 1900
rect -1350 100 -1150 1700
rect 500 100 700 1700
rect -1350 -100 700 100
rect 900 -300 1100 2100
rect -1750 -500 -650 -300
rect -850 -700 -650 -500
rect 0 -500 1100 -300
rect 0 -700 200 -500
<< end >>
