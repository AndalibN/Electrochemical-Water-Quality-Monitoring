magic
tech sky130A
magscale 1 2
timestamp 1667590084
<< pwell >>
rect -201 -848 201 848
<< psubdiff >>
rect -165 778 -69 812
rect 69 778 165 812
rect -165 716 -131 778
rect 131 716 165 778
rect -165 -778 -131 -716
rect 131 -778 165 -716
rect -165 -812 -69 -778
rect 69 -812 165 -778
<< psubdiffcont >>
rect -69 778 69 812
rect -165 -716 -131 716
rect 131 -716 165 716
rect -69 -812 69 -778
<< xpolycontact >>
rect -35 250 35 682
rect -35 -682 35 -250
<< ppolyres >>
rect -35 -250 35 250
<< locali >>
rect -165 778 -69 812
rect 69 778 165 812
rect -165 716 -131 778
rect 131 716 165 778
rect -165 -778 -131 -716
rect 131 -778 165 -716
rect -165 -812 -69 -778
rect 69 -812 165 -778
<< viali >>
rect -19 267 19 664
rect -19 -664 19 -267
<< metal1 >>
rect -25 664 25 676
rect -25 267 -19 664
rect 19 267 25 664
rect -25 255 25 267
rect -25 -267 25 -255
rect -25 -664 -19 -267
rect 19 -664 25 -267
rect -25 -676 25 -664
<< res0p35 >>
rect -37 -252 37 252
<< properties >>
string FIXED_BBOX -148 -795 148 795
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 2.5 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 3.397k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
