magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< metal3 >>
rect -1711 1532 -632 1590
rect -1711 1468 -716 1532
rect -652 1468 -632 1532
rect -1711 1452 -632 1468
rect -1711 1388 -716 1452
rect -652 1388 -632 1452
rect -1711 1372 -632 1388
rect -1711 1308 -716 1372
rect -652 1308 -632 1372
rect -1711 1292 -632 1308
rect -1711 1228 -716 1292
rect -652 1228 -632 1292
rect -1711 1212 -632 1228
rect -1711 1148 -716 1212
rect -652 1148 -632 1212
rect -1711 1132 -632 1148
rect -1711 1068 -716 1132
rect -652 1068 -632 1132
rect -1711 1052 -632 1068
rect -1711 988 -716 1052
rect -652 988 -632 1052
rect -1711 972 -632 988
rect -1711 908 -716 972
rect -652 908 -632 972
rect -1711 892 -632 908
rect -1711 828 -716 892
rect -652 828 -632 892
rect -1711 812 -632 828
rect -1711 748 -716 812
rect -652 748 -632 812
rect -1711 732 -632 748
rect -1711 668 -716 732
rect -652 668 -632 732
rect -1711 610 -632 668
rect -540 1512 539 1570
rect -540 1448 455 1512
rect 519 1448 539 1512
rect -540 1432 539 1448
rect -540 1368 455 1432
rect 519 1368 539 1432
rect -540 1352 539 1368
rect -540 1288 455 1352
rect 519 1288 539 1352
rect -540 1272 539 1288
rect -540 1208 455 1272
rect 519 1208 539 1272
rect -540 1192 539 1208
rect -540 1128 455 1192
rect 519 1128 539 1192
rect -540 1112 539 1128
rect -540 1048 455 1112
rect 519 1048 539 1112
rect -540 1032 539 1048
rect -540 968 455 1032
rect 519 968 539 1032
rect -540 952 539 968
rect -540 888 455 952
rect 519 888 539 952
rect -540 872 539 888
rect -540 808 455 872
rect 519 808 539 872
rect -540 792 539 808
rect -540 728 455 792
rect 519 728 539 792
rect -540 712 539 728
rect -540 648 455 712
rect 519 648 539 712
rect -540 590 539 648
rect 631 1532 1710 1590
rect 631 1468 1626 1532
rect 1690 1468 1710 1532
rect 631 1452 1710 1468
rect 631 1388 1626 1452
rect 1690 1388 1710 1452
rect 631 1372 1710 1388
rect 631 1308 1626 1372
rect 1690 1308 1710 1372
rect 631 1292 1710 1308
rect 631 1228 1626 1292
rect 1690 1228 1710 1292
rect 631 1212 1710 1228
rect 631 1148 1626 1212
rect 1690 1148 1710 1212
rect 631 1132 1710 1148
rect 631 1068 1626 1132
rect 1690 1068 1710 1132
rect 631 1052 1710 1068
rect 631 988 1626 1052
rect 1690 988 1710 1052
rect 631 972 1710 988
rect 631 908 1626 972
rect 1690 908 1710 972
rect 631 892 1710 908
rect 631 828 1626 892
rect 1690 828 1710 892
rect 631 812 1710 828
rect 631 748 1626 812
rect 1690 748 1710 812
rect 631 732 1710 748
rect 631 668 1626 732
rect 1690 668 1710 732
rect 631 610 1710 668
rect -1711 452 -632 510
rect -1711 388 -716 452
rect -652 388 -632 452
rect -1711 372 -632 388
rect -1711 308 -716 372
rect -652 308 -632 372
rect -1711 292 -632 308
rect -1711 228 -716 292
rect -652 228 -632 292
rect -1711 212 -632 228
rect -1711 148 -716 212
rect -652 148 -632 212
rect -1711 132 -632 148
rect -1711 68 -716 132
rect -652 68 -632 132
rect -1711 52 -632 68
rect -1711 -12 -716 52
rect -652 -12 -632 52
rect -1711 -28 -632 -12
rect -1711 -92 -716 -28
rect -652 -92 -632 -28
rect -1711 -108 -632 -92
rect -1711 -172 -716 -108
rect -652 -172 -632 -108
rect -1711 -188 -632 -172
rect -1711 -252 -716 -188
rect -652 -252 -632 -188
rect -1711 -268 -632 -252
rect -1711 -332 -716 -268
rect -652 -332 -632 -268
rect -1711 -348 -632 -332
rect -1711 -412 -716 -348
rect -652 -412 -632 -348
rect -1711 -470 -632 -412
rect -540 432 539 490
rect -540 368 455 432
rect 519 368 539 432
rect -540 352 539 368
rect -540 288 455 352
rect 519 288 539 352
rect -540 272 539 288
rect -540 208 455 272
rect 519 208 539 272
rect -540 192 539 208
rect -540 128 455 192
rect 519 128 539 192
rect -540 112 539 128
rect -540 48 455 112
rect 519 48 539 112
rect -540 32 539 48
rect -540 -32 455 32
rect 519 -32 539 32
rect -540 -48 539 -32
rect -540 -112 455 -48
rect 519 -112 539 -48
rect -540 -128 539 -112
rect -540 -192 455 -128
rect 519 -192 539 -128
rect -540 -208 539 -192
rect -540 -272 455 -208
rect 519 -272 539 -208
rect -540 -288 539 -272
rect -540 -352 455 -288
rect 519 -352 539 -288
rect -540 -368 539 -352
rect -540 -432 455 -368
rect 519 -432 539 -368
rect -540 -490 539 -432
rect 631 452 1710 510
rect 631 388 1626 452
rect 1690 388 1710 452
rect 631 372 1710 388
rect 631 308 1626 372
rect 1690 308 1710 372
rect 631 292 1710 308
rect 631 228 1626 292
rect 1690 228 1710 292
rect 631 212 1710 228
rect 631 148 1626 212
rect 1690 148 1710 212
rect 631 132 1710 148
rect 631 68 1626 132
rect 1690 68 1710 132
rect 631 52 1710 68
rect 631 -12 1626 52
rect 1690 -12 1710 52
rect 631 -28 1710 -12
rect 631 -92 1626 -28
rect 1690 -92 1710 -28
rect 631 -108 1710 -92
rect 631 -172 1626 -108
rect 1690 -172 1710 -108
rect 631 -188 1710 -172
rect 631 -252 1626 -188
rect 1690 -252 1710 -188
rect 631 -268 1710 -252
rect 631 -332 1626 -268
rect 1690 -332 1710 -268
rect 631 -348 1710 -332
rect 631 -412 1626 -348
rect 1690 -412 1710 -348
rect 631 -470 1710 -412
rect -1711 -628 -632 -570
rect -1711 -692 -716 -628
rect -652 -692 -632 -628
rect -1711 -708 -632 -692
rect -1711 -772 -716 -708
rect -652 -772 -632 -708
rect -1711 -788 -632 -772
rect -1711 -852 -716 -788
rect -652 -852 -632 -788
rect -1711 -868 -632 -852
rect -1711 -932 -716 -868
rect -652 -932 -632 -868
rect -1711 -948 -632 -932
rect -1711 -1012 -716 -948
rect -652 -1012 -632 -948
rect -1711 -1028 -632 -1012
rect -1711 -1092 -716 -1028
rect -652 -1092 -632 -1028
rect -1711 -1108 -632 -1092
rect -1711 -1172 -716 -1108
rect -652 -1172 -632 -1108
rect -1711 -1188 -632 -1172
rect -1711 -1252 -716 -1188
rect -652 -1252 -632 -1188
rect -1711 -1268 -632 -1252
rect -1711 -1332 -716 -1268
rect -652 -1332 -632 -1268
rect -1711 -1348 -632 -1332
rect -1711 -1412 -716 -1348
rect -652 -1412 -632 -1348
rect -1711 -1428 -632 -1412
rect -1711 -1492 -716 -1428
rect -652 -1492 -632 -1428
rect -1711 -1550 -632 -1492
rect -540 -648 539 -590
rect -540 -712 455 -648
rect 519 -712 539 -648
rect -540 -728 539 -712
rect -540 -792 455 -728
rect 519 -792 539 -728
rect -540 -808 539 -792
rect -540 -872 455 -808
rect 519 -872 539 -808
rect -540 -888 539 -872
rect -540 -952 455 -888
rect 519 -952 539 -888
rect -540 -968 539 -952
rect -540 -1032 455 -968
rect 519 -1032 539 -968
rect -540 -1048 539 -1032
rect -540 -1112 455 -1048
rect 519 -1112 539 -1048
rect -540 -1128 539 -1112
rect -540 -1192 455 -1128
rect 519 -1192 539 -1128
rect -540 -1208 539 -1192
rect -540 -1272 455 -1208
rect 519 -1272 539 -1208
rect -540 -1288 539 -1272
rect -540 -1352 455 -1288
rect 519 -1352 539 -1288
rect -540 -1368 539 -1352
rect -540 -1432 455 -1368
rect 519 -1432 539 -1368
rect -540 -1448 539 -1432
rect -540 -1512 455 -1448
rect 519 -1512 539 -1448
rect -540 -1570 539 -1512
rect 631 -628 1710 -570
rect 631 -692 1626 -628
rect 1690 -692 1710 -628
rect 631 -708 1710 -692
rect 631 -772 1626 -708
rect 1690 -772 1710 -708
rect 631 -788 1710 -772
rect 631 -852 1626 -788
rect 1690 -852 1710 -788
rect 631 -868 1710 -852
rect 631 -932 1626 -868
rect 1690 -932 1710 -868
rect 631 -948 1710 -932
rect 631 -1012 1626 -948
rect 1690 -1012 1710 -948
rect 631 -1028 1710 -1012
rect 631 -1092 1626 -1028
rect 1690 -1092 1710 -1028
rect 631 -1108 1710 -1092
rect 631 -1172 1626 -1108
rect 1690 -1172 1710 -1108
rect 631 -1188 1710 -1172
rect 631 -1252 1626 -1188
rect 1690 -1252 1710 -1188
rect 631 -1268 1710 -1252
rect 631 -1332 1626 -1268
rect 1690 -1332 1710 -1268
rect 631 -1348 1710 -1332
rect 631 -1412 1626 -1348
rect 1690 -1412 1710 -1348
rect 631 -1428 1710 -1412
rect 631 -1492 1626 -1428
rect 1690 -1492 1710 -1428
rect 631 -1550 1710 -1492
<< via3 >>
rect -716 1468 -652 1532
rect -716 1388 -652 1452
rect -716 1308 -652 1372
rect -716 1228 -652 1292
rect -716 1148 -652 1212
rect -716 1068 -652 1132
rect -716 988 -652 1052
rect -716 908 -652 972
rect -716 828 -652 892
rect -716 748 -652 812
rect -716 668 -652 732
rect 455 1448 519 1512
rect 455 1368 519 1432
rect 455 1288 519 1352
rect 455 1208 519 1272
rect 455 1128 519 1192
rect 455 1048 519 1112
rect 455 968 519 1032
rect 455 888 519 952
rect 455 808 519 872
rect 455 728 519 792
rect 455 648 519 712
rect 1626 1468 1690 1532
rect 1626 1388 1690 1452
rect 1626 1308 1690 1372
rect 1626 1228 1690 1292
rect 1626 1148 1690 1212
rect 1626 1068 1690 1132
rect 1626 988 1690 1052
rect 1626 908 1690 972
rect 1626 828 1690 892
rect 1626 748 1690 812
rect 1626 668 1690 732
rect -716 388 -652 452
rect -716 308 -652 372
rect -716 228 -652 292
rect -716 148 -652 212
rect -716 68 -652 132
rect -716 -12 -652 52
rect -716 -92 -652 -28
rect -716 -172 -652 -108
rect -716 -252 -652 -188
rect -716 -332 -652 -268
rect -716 -412 -652 -348
rect 455 368 519 432
rect 455 288 519 352
rect 455 208 519 272
rect 455 128 519 192
rect 455 48 519 112
rect 455 -32 519 32
rect 455 -112 519 -48
rect 455 -192 519 -128
rect 455 -272 519 -208
rect 455 -352 519 -288
rect 455 -432 519 -368
rect 1626 388 1690 452
rect 1626 308 1690 372
rect 1626 228 1690 292
rect 1626 148 1690 212
rect 1626 68 1690 132
rect 1626 -12 1690 52
rect 1626 -92 1690 -28
rect 1626 -172 1690 -108
rect 1626 -252 1690 -188
rect 1626 -332 1690 -268
rect 1626 -412 1690 -348
rect -716 -692 -652 -628
rect -716 -772 -652 -708
rect -716 -852 -652 -788
rect -716 -932 -652 -868
rect -716 -1012 -652 -948
rect -716 -1092 -652 -1028
rect -716 -1172 -652 -1108
rect -716 -1252 -652 -1188
rect -716 -1332 -652 -1268
rect -716 -1412 -652 -1348
rect -716 -1492 -652 -1428
rect 455 -712 519 -648
rect 455 -792 519 -728
rect 455 -872 519 -808
rect 455 -952 519 -888
rect 455 -1032 519 -968
rect 455 -1112 519 -1048
rect 455 -1192 519 -1128
rect 455 -1272 519 -1208
rect 455 -1352 519 -1288
rect 455 -1432 519 -1368
rect 455 -1512 519 -1448
rect 1626 -692 1690 -628
rect 1626 -772 1690 -708
rect 1626 -852 1690 -788
rect 1626 -932 1690 -868
rect 1626 -1012 1690 -948
rect 1626 -1092 1690 -1028
rect 1626 -1172 1690 -1108
rect 1626 -1252 1690 -1188
rect 1626 -1332 1690 -1268
rect 1626 -1412 1690 -1348
rect 1626 -1492 1690 -1428
<< mimcap >>
rect -1611 1412 -831 1490
rect -1611 788 -1533 1412
rect -909 788 -831 1412
rect -1611 710 -831 788
rect -440 1392 340 1470
rect -440 768 -362 1392
rect 262 768 340 1392
rect -440 690 340 768
rect 731 1412 1511 1490
rect 731 788 809 1412
rect 1433 788 1511 1412
rect 731 710 1511 788
rect -1611 332 -831 410
rect -1611 -292 -1533 332
rect -909 -292 -831 332
rect -1611 -370 -831 -292
rect -440 312 340 390
rect -440 -312 -362 312
rect 262 -312 340 312
rect -440 -390 340 -312
rect 731 332 1511 410
rect 731 -292 809 332
rect 1433 -292 1511 332
rect 731 -370 1511 -292
rect -1611 -748 -831 -670
rect -1611 -1372 -1533 -748
rect -909 -1372 -831 -748
rect -1611 -1450 -831 -1372
rect -440 -768 340 -690
rect -440 -1392 -362 -768
rect 262 -1392 340 -768
rect -440 -1470 340 -1392
rect 731 -748 1511 -670
rect 731 -1372 809 -748
rect 1433 -1372 1511 -748
rect 731 -1450 1511 -1372
<< mimcapcontact >>
rect -1533 788 -909 1412
rect -362 768 262 1392
rect 809 788 1433 1412
rect -1533 -292 -909 332
rect -362 -312 262 312
rect 809 -292 1433 332
rect -1533 -1372 -909 -748
rect -362 -1392 262 -768
rect 809 -1372 1433 -748
<< metal4 >>
rect -1572 1412 -870 1640
rect -1572 788 -1533 1412
rect -909 788 -870 1412
rect -1572 332 -870 788
rect -1572 -292 -1533 332
rect -909 -292 -870 332
rect -1572 -748 -870 -292
rect -1572 -1372 -1533 -748
rect -909 -1372 -870 -748
rect -1572 -1972 -870 -1372
rect -763 1532 -636 1978
rect -763 1468 -716 1532
rect -652 1468 -636 1532
rect -763 1452 -636 1468
rect -763 1388 -716 1452
rect -652 1388 -636 1452
rect -763 1372 -636 1388
rect -763 1308 -716 1372
rect -652 1308 -636 1372
rect -763 1292 -636 1308
rect -763 1228 -716 1292
rect -652 1228 -636 1292
rect -763 1212 -636 1228
rect -763 1148 -716 1212
rect -652 1148 -636 1212
rect -763 1132 -636 1148
rect -763 1068 -716 1132
rect -652 1068 -636 1132
rect -763 1052 -636 1068
rect -763 988 -716 1052
rect -652 988 -636 1052
rect -763 972 -636 988
rect -763 908 -716 972
rect -652 908 -636 972
rect -763 892 -636 908
rect -763 828 -716 892
rect -652 828 -636 892
rect -763 812 -636 828
rect -763 748 -716 812
rect -652 748 -636 812
rect -763 732 -636 748
rect -763 668 -716 732
rect -652 668 -636 732
rect -763 452 -636 668
rect -763 388 -716 452
rect -652 388 -636 452
rect -763 372 -636 388
rect -763 308 -716 372
rect -652 308 -636 372
rect -763 292 -636 308
rect -763 228 -716 292
rect -652 228 -636 292
rect -763 212 -636 228
rect -763 148 -716 212
rect -652 148 -636 212
rect -763 132 -636 148
rect -763 68 -716 132
rect -652 68 -636 132
rect -763 52 -636 68
rect -763 -12 -716 52
rect -652 -12 -636 52
rect -763 -28 -636 -12
rect -763 -92 -716 -28
rect -652 -92 -636 -28
rect -763 -108 -636 -92
rect -763 -172 -716 -108
rect -652 -172 -636 -108
rect -763 -188 -636 -172
rect -763 -252 -716 -188
rect -652 -252 -636 -188
rect -763 -268 -636 -252
rect -763 -332 -716 -268
rect -652 -332 -636 -268
rect -763 -348 -636 -332
rect -763 -412 -716 -348
rect -652 -412 -636 -348
rect -763 -628 -636 -412
rect -763 -692 -716 -628
rect -652 -692 -636 -628
rect -763 -708 -636 -692
rect -763 -772 -716 -708
rect -652 -772 -636 -708
rect -763 -788 -636 -772
rect -763 -852 -716 -788
rect -652 -852 -636 -788
rect -763 -868 -636 -852
rect -763 -932 -716 -868
rect -652 -932 -636 -868
rect -763 -948 -636 -932
rect -763 -1012 -716 -948
rect -652 -1012 -636 -948
rect -763 -1028 -636 -1012
rect -763 -1092 -716 -1028
rect -652 -1092 -636 -1028
rect -763 -1108 -636 -1092
rect -763 -1172 -716 -1108
rect -652 -1172 -636 -1108
rect -763 -1188 -636 -1172
rect -763 -1252 -716 -1188
rect -652 -1252 -636 -1188
rect -763 -1268 -636 -1252
rect -763 -1332 -716 -1268
rect -652 -1332 -636 -1268
rect -763 -1348 -636 -1332
rect -763 -1412 -716 -1348
rect -652 -1412 -636 -1348
rect -763 -1428 -636 -1412
rect -763 -1492 -716 -1428
rect -652 -1492 -636 -1428
rect -763 -1538 -636 -1492
rect -401 1392 301 1620
rect -401 768 -362 1392
rect 262 768 301 1392
rect -401 312 301 768
rect -401 -312 -362 312
rect 262 -312 301 312
rect -401 -768 301 -312
rect -401 -1392 -362 -768
rect 262 -1392 301 -768
rect -401 -1972 301 -1392
rect 408 1512 535 1995
rect 408 1448 455 1512
rect 519 1448 535 1512
rect 408 1432 535 1448
rect 408 1368 455 1432
rect 519 1368 535 1432
rect 408 1352 535 1368
rect 408 1288 455 1352
rect 519 1288 535 1352
rect 408 1272 535 1288
rect 408 1208 455 1272
rect 519 1208 535 1272
rect 408 1192 535 1208
rect 408 1128 455 1192
rect 519 1128 535 1192
rect 408 1112 535 1128
rect 408 1048 455 1112
rect 519 1048 535 1112
rect 408 1032 535 1048
rect 408 968 455 1032
rect 519 968 535 1032
rect 408 952 535 968
rect 408 888 455 952
rect 519 888 535 952
rect 408 872 535 888
rect 408 808 455 872
rect 519 808 535 872
rect 408 792 535 808
rect 408 728 455 792
rect 519 728 535 792
rect 408 712 535 728
rect 408 648 455 712
rect 519 648 535 712
rect 408 432 535 648
rect 408 368 455 432
rect 519 368 535 432
rect 408 352 535 368
rect 408 288 455 352
rect 519 288 535 352
rect 408 272 535 288
rect 408 208 455 272
rect 519 208 535 272
rect 408 192 535 208
rect 408 128 455 192
rect 519 128 535 192
rect 408 112 535 128
rect 408 48 455 112
rect 519 48 535 112
rect 408 32 535 48
rect 408 -32 455 32
rect 519 -32 535 32
rect 408 -48 535 -32
rect 408 -112 455 -48
rect 519 -112 535 -48
rect 408 -128 535 -112
rect 408 -192 455 -128
rect 519 -192 535 -128
rect 408 -208 535 -192
rect 408 -272 455 -208
rect 519 -272 535 -208
rect 408 -288 535 -272
rect 408 -352 455 -288
rect 519 -352 535 -288
rect 408 -368 535 -352
rect 408 -432 455 -368
rect 519 -432 535 -368
rect 408 -648 535 -432
rect 408 -712 455 -648
rect 519 -712 535 -648
rect 408 -728 535 -712
rect 408 -792 455 -728
rect 519 -792 535 -728
rect 408 -808 535 -792
rect 408 -872 455 -808
rect 519 -872 535 -808
rect 408 -888 535 -872
rect 408 -952 455 -888
rect 519 -952 535 -888
rect 408 -968 535 -952
rect 408 -1032 455 -968
rect 519 -1032 535 -968
rect 408 -1048 535 -1032
rect 408 -1112 455 -1048
rect 519 -1112 535 -1048
rect 408 -1128 535 -1112
rect 408 -1192 455 -1128
rect 519 -1192 535 -1128
rect 408 -1208 535 -1192
rect 408 -1272 455 -1208
rect 519 -1272 535 -1208
rect 408 -1288 535 -1272
rect 408 -1352 455 -1288
rect 519 -1352 535 -1288
rect 408 -1368 535 -1352
rect 408 -1432 455 -1368
rect 519 -1432 535 -1368
rect 408 -1448 535 -1432
rect 408 -1512 455 -1448
rect 519 -1512 535 -1448
rect 408 -1558 535 -1512
rect 770 1412 1472 1640
rect 770 788 809 1412
rect 1433 788 1472 1412
rect 770 332 1472 788
rect 770 -292 809 332
rect 1433 -292 1472 332
rect 770 -748 1472 -292
rect 770 -1372 809 -748
rect 1433 -1372 1472 -748
rect 770 -1972 1472 -1372
rect 1579 1532 1706 1960
rect 1579 1468 1626 1532
rect 1690 1468 1706 1532
rect 1579 1452 1706 1468
rect 1579 1388 1626 1452
rect 1690 1388 1706 1452
rect 1579 1372 1706 1388
rect 1579 1308 1626 1372
rect 1690 1308 1706 1372
rect 1579 1292 1706 1308
rect 1579 1228 1626 1292
rect 1690 1228 1706 1292
rect 1579 1212 1706 1228
rect 1579 1148 1626 1212
rect 1690 1148 1706 1212
rect 1579 1132 1706 1148
rect 1579 1068 1626 1132
rect 1690 1068 1706 1132
rect 1579 1052 1706 1068
rect 1579 988 1626 1052
rect 1690 988 1706 1052
rect 1579 972 1706 988
rect 1579 908 1626 972
rect 1690 908 1706 972
rect 1579 892 1706 908
rect 1579 828 1626 892
rect 1690 828 1706 892
rect 1579 812 1706 828
rect 1579 748 1626 812
rect 1690 748 1706 812
rect 1579 732 1706 748
rect 1579 668 1626 732
rect 1690 668 1706 732
rect 1579 452 1706 668
rect 1579 388 1626 452
rect 1690 388 1706 452
rect 1579 372 1706 388
rect 1579 308 1626 372
rect 1690 308 1706 372
rect 1579 292 1706 308
rect 1579 228 1626 292
rect 1690 228 1706 292
rect 1579 212 1706 228
rect 1579 148 1626 212
rect 1690 148 1706 212
rect 1579 132 1706 148
rect 1579 68 1626 132
rect 1690 68 1706 132
rect 1579 52 1706 68
rect 1579 -12 1626 52
rect 1690 -12 1706 52
rect 1579 -28 1706 -12
rect 1579 -92 1626 -28
rect 1690 -92 1706 -28
rect 1579 -108 1706 -92
rect 1579 -172 1626 -108
rect 1690 -172 1706 -108
rect 1579 -188 1706 -172
rect 1579 -252 1626 -188
rect 1690 -252 1706 -188
rect 1579 -268 1706 -252
rect 1579 -332 1626 -268
rect 1690 -332 1706 -268
rect 1579 -348 1706 -332
rect 1579 -412 1626 -348
rect 1690 -412 1706 -348
rect 1579 -628 1706 -412
rect 1579 -692 1626 -628
rect 1690 -692 1706 -628
rect 1579 -708 1706 -692
rect 1579 -772 1626 -708
rect 1690 -772 1706 -708
rect 1579 -788 1706 -772
rect 1579 -852 1626 -788
rect 1690 -852 1706 -788
rect 1579 -868 1706 -852
rect 1579 -932 1626 -868
rect 1690 -932 1706 -868
rect 1579 -948 1706 -932
rect 1579 -1012 1626 -948
rect 1690 -1012 1706 -948
rect 1579 -1028 1706 -1012
rect 1579 -1092 1626 -1028
rect 1690 -1092 1706 -1028
rect 1579 -1108 1706 -1092
rect 1579 -1172 1626 -1108
rect 1690 -1172 1706 -1108
rect 1579 -1188 1706 -1172
rect 1579 -1252 1626 -1188
rect 1690 -1252 1706 -1188
rect 1579 -1268 1706 -1252
rect 1579 -1332 1626 -1268
rect 1690 -1332 1706 -1268
rect 1579 -1348 1706 -1332
rect 1579 -1412 1626 -1348
rect 1690 -1412 1706 -1348
rect 1579 -1428 1706 -1412
rect 1579 -1492 1626 -1428
rect 1690 -1492 1706 -1428
rect 1579 -1538 1706 -1492
<< properties >>
string FIXED_BBOX 559 590 1539 1570
<< end >>
