magic
tech sky130A
magscale 1 2
timestamp 1666625676
<< xpolycontact >>
rect -7826 5200 -7756 5632
rect -7826 -5632 -7756 -5200
rect -7508 5200 -7438 5632
rect -7508 -5632 -7438 -5200
rect -7190 5200 -7120 5632
rect -7190 -5632 -7120 -5200
rect -6872 5200 -6802 5632
rect -6872 -5632 -6802 -5200
rect -6554 5200 -6484 5632
rect -6554 -5632 -6484 -5200
rect -6236 5200 -6166 5632
rect -6236 -5632 -6166 -5200
rect -5918 5200 -5848 5632
rect -5918 -5632 -5848 -5200
rect -5600 5200 -5530 5632
rect -5600 -5632 -5530 -5200
rect -5282 5200 -5212 5632
rect -5282 -5632 -5212 -5200
rect -4964 5200 -4894 5632
rect -4964 -5632 -4894 -5200
rect -4646 5200 -4576 5632
rect -4646 -5632 -4576 -5200
rect -4328 5200 -4258 5632
rect -4328 -5632 -4258 -5200
rect -4010 5200 -3940 5632
rect -4010 -5632 -3940 -5200
rect -3692 5200 -3622 5632
rect -3692 -5632 -3622 -5200
rect -3374 5200 -3304 5632
rect -3374 -5632 -3304 -5200
rect -3056 5200 -2986 5632
rect -3056 -5632 -2986 -5200
rect -2738 5200 -2668 5632
rect -2738 -5632 -2668 -5200
rect -2420 5200 -2350 5632
rect -2420 -5632 -2350 -5200
rect -2102 5200 -2032 5632
rect -2102 -5632 -2032 -5200
rect -1784 5200 -1714 5632
rect -1784 -5632 -1714 -5200
rect -1466 5200 -1396 5632
rect -1466 -5632 -1396 -5200
rect -1148 5200 -1078 5632
rect -1148 -5632 -1078 -5200
rect -830 5200 -760 5632
rect -830 -5632 -760 -5200
rect -512 5200 -442 5632
rect -512 -5632 -442 -5200
rect -194 5200 -124 5632
rect -194 -5632 -124 -5200
rect 124 5200 194 5632
rect 124 -5632 194 -5200
rect 442 5200 512 5632
rect 442 -5632 512 -5200
rect 760 5200 830 5632
rect 760 -5632 830 -5200
rect 1078 5200 1148 5632
rect 1078 -5632 1148 -5200
rect 1396 5200 1466 5632
rect 1396 -5632 1466 -5200
rect 1714 5200 1784 5632
rect 1714 -5632 1784 -5200
rect 2032 5200 2102 5632
rect 2032 -5632 2102 -5200
rect 2350 5200 2420 5632
rect 2350 -5632 2420 -5200
rect 2668 5200 2738 5632
rect 2668 -5632 2738 -5200
rect 2986 5200 3056 5632
rect 2986 -5632 3056 -5200
rect 3304 5200 3374 5632
rect 3304 -5632 3374 -5200
rect 3622 5200 3692 5632
rect 3622 -5632 3692 -5200
rect 3940 5200 4010 5632
rect 3940 -5632 4010 -5200
rect 4258 5200 4328 5632
rect 4258 -5632 4328 -5200
rect 4576 5200 4646 5632
rect 4576 -5632 4646 -5200
rect 4894 5200 4964 5632
rect 4894 -5632 4964 -5200
rect 5212 5200 5282 5632
rect 5212 -5632 5282 -5200
rect 5530 5200 5600 5632
rect 5530 -5632 5600 -5200
rect 5848 5200 5918 5632
rect 5848 -5632 5918 -5200
rect 6166 5200 6236 5632
rect 6166 -5632 6236 -5200
rect 6484 5200 6554 5632
rect 6484 -5632 6554 -5200
rect 6802 5200 6872 5632
rect 6802 -5632 6872 -5200
rect 7120 5200 7190 5632
rect 7120 -5632 7190 -5200
rect 7438 5200 7508 5632
rect 7438 -5632 7508 -5200
rect 7756 5200 7826 5632
rect 7756 -5632 7826 -5200
<< xpolyres >>
rect -7826 -5200 -7756 5200
rect -7508 -5200 -7438 5200
rect -7190 -5200 -7120 5200
rect -6872 -5200 -6802 5200
rect -6554 -5200 -6484 5200
rect -6236 -5200 -6166 5200
rect -5918 -5200 -5848 5200
rect -5600 -5200 -5530 5200
rect -5282 -5200 -5212 5200
rect -4964 -5200 -4894 5200
rect -4646 -5200 -4576 5200
rect -4328 -5200 -4258 5200
rect -4010 -5200 -3940 5200
rect -3692 -5200 -3622 5200
rect -3374 -5200 -3304 5200
rect -3056 -5200 -2986 5200
rect -2738 -5200 -2668 5200
rect -2420 -5200 -2350 5200
rect -2102 -5200 -2032 5200
rect -1784 -5200 -1714 5200
rect -1466 -5200 -1396 5200
rect -1148 -5200 -1078 5200
rect -830 -5200 -760 5200
rect -512 -5200 -442 5200
rect -194 -5200 -124 5200
rect 124 -5200 194 5200
rect 442 -5200 512 5200
rect 760 -5200 830 5200
rect 1078 -5200 1148 5200
rect 1396 -5200 1466 5200
rect 1714 -5200 1784 5200
rect 2032 -5200 2102 5200
rect 2350 -5200 2420 5200
rect 2668 -5200 2738 5200
rect 2986 -5200 3056 5200
rect 3304 -5200 3374 5200
rect 3622 -5200 3692 5200
rect 3940 -5200 4010 5200
rect 4258 -5200 4328 5200
rect 4576 -5200 4646 5200
rect 4894 -5200 4964 5200
rect 5212 -5200 5282 5200
rect 5530 -5200 5600 5200
rect 5848 -5200 5918 5200
rect 6166 -5200 6236 5200
rect 6484 -5200 6554 5200
rect 6802 -5200 6872 5200
rect 7120 -5200 7190 5200
rect 7438 -5200 7508 5200
rect 7756 -5200 7826 5200
<< viali >>
rect -7810 5217 -7772 5614
rect -7492 5217 -7454 5614
rect -7174 5217 -7136 5614
rect -6856 5217 -6818 5614
rect -6538 5217 -6500 5614
rect -6220 5217 -6182 5614
rect -5902 5217 -5864 5614
rect -5584 5217 -5546 5614
rect -5266 5217 -5228 5614
rect -4948 5217 -4910 5614
rect -4630 5217 -4592 5614
rect -4312 5217 -4274 5614
rect -3994 5217 -3956 5614
rect -3676 5217 -3638 5614
rect -3358 5217 -3320 5614
rect -3040 5217 -3002 5614
rect -2722 5217 -2684 5614
rect -2404 5217 -2366 5614
rect -2086 5217 -2048 5614
rect -1768 5217 -1730 5614
rect -1450 5217 -1412 5614
rect -1132 5217 -1094 5614
rect -814 5217 -776 5614
rect -496 5217 -458 5614
rect -178 5217 -140 5614
rect 140 5217 178 5614
rect 458 5217 496 5614
rect 776 5217 814 5614
rect 1094 5217 1132 5614
rect 1412 5217 1450 5614
rect 1730 5217 1768 5614
rect 2048 5217 2086 5614
rect 2366 5217 2404 5614
rect 2684 5217 2722 5614
rect 3002 5217 3040 5614
rect 3320 5217 3358 5614
rect 3638 5217 3676 5614
rect 3956 5217 3994 5614
rect 4274 5217 4312 5614
rect 4592 5217 4630 5614
rect 4910 5217 4948 5614
rect 5228 5217 5266 5614
rect 5546 5217 5584 5614
rect 5864 5217 5902 5614
rect 6182 5217 6220 5614
rect 6500 5217 6538 5614
rect 6818 5217 6856 5614
rect 7136 5217 7174 5614
rect 7454 5217 7492 5614
rect 7772 5217 7810 5614
rect -7810 -5614 -7772 -5217
rect -7492 -5614 -7454 -5217
rect -7174 -5614 -7136 -5217
rect -6856 -5614 -6818 -5217
rect -6538 -5614 -6500 -5217
rect -6220 -5614 -6182 -5217
rect -5902 -5614 -5864 -5217
rect -5584 -5614 -5546 -5217
rect -5266 -5614 -5228 -5217
rect -4948 -5614 -4910 -5217
rect -4630 -5614 -4592 -5217
rect -4312 -5614 -4274 -5217
rect -3994 -5614 -3956 -5217
rect -3676 -5614 -3638 -5217
rect -3358 -5614 -3320 -5217
rect -3040 -5614 -3002 -5217
rect -2722 -5614 -2684 -5217
rect -2404 -5614 -2366 -5217
rect -2086 -5614 -2048 -5217
rect -1768 -5614 -1730 -5217
rect -1450 -5614 -1412 -5217
rect -1132 -5614 -1094 -5217
rect -814 -5614 -776 -5217
rect -496 -5614 -458 -5217
rect -178 -5614 -140 -5217
rect 140 -5614 178 -5217
rect 458 -5614 496 -5217
rect 776 -5614 814 -5217
rect 1094 -5614 1132 -5217
rect 1412 -5614 1450 -5217
rect 1730 -5614 1768 -5217
rect 2048 -5614 2086 -5217
rect 2366 -5614 2404 -5217
rect 2684 -5614 2722 -5217
rect 3002 -5614 3040 -5217
rect 3320 -5614 3358 -5217
rect 3638 -5614 3676 -5217
rect 3956 -5614 3994 -5217
rect 4274 -5614 4312 -5217
rect 4592 -5614 4630 -5217
rect 4910 -5614 4948 -5217
rect 5228 -5614 5266 -5217
rect 5546 -5614 5584 -5217
rect 5864 -5614 5902 -5217
rect 6182 -5614 6220 -5217
rect 6500 -5614 6538 -5217
rect 6818 -5614 6856 -5217
rect 7136 -5614 7174 -5217
rect 7454 -5614 7492 -5217
rect 7772 -5614 7810 -5217
<< metal1 >>
rect -7816 5614 -7766 5626
rect -7816 5217 -7810 5614
rect -7772 5217 -7766 5614
rect -7816 5205 -7766 5217
rect -7498 5614 -7448 5626
rect -7498 5217 -7492 5614
rect -7454 5217 -7448 5614
rect -7498 5205 -7448 5217
rect -7180 5614 -7130 5626
rect -7180 5217 -7174 5614
rect -7136 5217 -7130 5614
rect -7180 5205 -7130 5217
rect -6862 5614 -6812 5626
rect -6862 5217 -6856 5614
rect -6818 5217 -6812 5614
rect -6862 5205 -6812 5217
rect -6544 5614 -6494 5626
rect -6544 5217 -6538 5614
rect -6500 5217 -6494 5614
rect -6544 5205 -6494 5217
rect -6226 5614 -6176 5626
rect -6226 5217 -6220 5614
rect -6182 5217 -6176 5614
rect -6226 5205 -6176 5217
rect -5908 5614 -5858 5626
rect -5908 5217 -5902 5614
rect -5864 5217 -5858 5614
rect -5908 5205 -5858 5217
rect -5590 5614 -5540 5626
rect -5590 5217 -5584 5614
rect -5546 5217 -5540 5614
rect -5590 5205 -5540 5217
rect -5272 5614 -5222 5626
rect -5272 5217 -5266 5614
rect -5228 5217 -5222 5614
rect -5272 5205 -5222 5217
rect -4954 5614 -4904 5626
rect -4954 5217 -4948 5614
rect -4910 5217 -4904 5614
rect -4954 5205 -4904 5217
rect -4636 5614 -4586 5626
rect -4636 5217 -4630 5614
rect -4592 5217 -4586 5614
rect -4636 5205 -4586 5217
rect -4318 5614 -4268 5626
rect -4318 5217 -4312 5614
rect -4274 5217 -4268 5614
rect -4318 5205 -4268 5217
rect -4000 5614 -3950 5626
rect -4000 5217 -3994 5614
rect -3956 5217 -3950 5614
rect -4000 5205 -3950 5217
rect -3682 5614 -3632 5626
rect -3682 5217 -3676 5614
rect -3638 5217 -3632 5614
rect -3682 5205 -3632 5217
rect -3364 5614 -3314 5626
rect -3364 5217 -3358 5614
rect -3320 5217 -3314 5614
rect -3364 5205 -3314 5217
rect -3046 5614 -2996 5626
rect -3046 5217 -3040 5614
rect -3002 5217 -2996 5614
rect -3046 5205 -2996 5217
rect -2728 5614 -2678 5626
rect -2728 5217 -2722 5614
rect -2684 5217 -2678 5614
rect -2728 5205 -2678 5217
rect -2410 5614 -2360 5626
rect -2410 5217 -2404 5614
rect -2366 5217 -2360 5614
rect -2410 5205 -2360 5217
rect -2092 5614 -2042 5626
rect -2092 5217 -2086 5614
rect -2048 5217 -2042 5614
rect -2092 5205 -2042 5217
rect -1774 5614 -1724 5626
rect -1774 5217 -1768 5614
rect -1730 5217 -1724 5614
rect -1774 5205 -1724 5217
rect -1456 5614 -1406 5626
rect -1456 5217 -1450 5614
rect -1412 5217 -1406 5614
rect -1456 5205 -1406 5217
rect -1138 5614 -1088 5626
rect -1138 5217 -1132 5614
rect -1094 5217 -1088 5614
rect -1138 5205 -1088 5217
rect -820 5614 -770 5626
rect -820 5217 -814 5614
rect -776 5217 -770 5614
rect -820 5205 -770 5217
rect -502 5614 -452 5626
rect -502 5217 -496 5614
rect -458 5217 -452 5614
rect -502 5205 -452 5217
rect -184 5614 -134 5626
rect -184 5217 -178 5614
rect -140 5217 -134 5614
rect -184 5205 -134 5217
rect 134 5614 184 5626
rect 134 5217 140 5614
rect 178 5217 184 5614
rect 134 5205 184 5217
rect 452 5614 502 5626
rect 452 5217 458 5614
rect 496 5217 502 5614
rect 452 5205 502 5217
rect 770 5614 820 5626
rect 770 5217 776 5614
rect 814 5217 820 5614
rect 770 5205 820 5217
rect 1088 5614 1138 5626
rect 1088 5217 1094 5614
rect 1132 5217 1138 5614
rect 1088 5205 1138 5217
rect 1406 5614 1456 5626
rect 1406 5217 1412 5614
rect 1450 5217 1456 5614
rect 1406 5205 1456 5217
rect 1724 5614 1774 5626
rect 1724 5217 1730 5614
rect 1768 5217 1774 5614
rect 1724 5205 1774 5217
rect 2042 5614 2092 5626
rect 2042 5217 2048 5614
rect 2086 5217 2092 5614
rect 2042 5205 2092 5217
rect 2360 5614 2410 5626
rect 2360 5217 2366 5614
rect 2404 5217 2410 5614
rect 2360 5205 2410 5217
rect 2678 5614 2728 5626
rect 2678 5217 2684 5614
rect 2722 5217 2728 5614
rect 2678 5205 2728 5217
rect 2996 5614 3046 5626
rect 2996 5217 3002 5614
rect 3040 5217 3046 5614
rect 2996 5205 3046 5217
rect 3314 5614 3364 5626
rect 3314 5217 3320 5614
rect 3358 5217 3364 5614
rect 3314 5205 3364 5217
rect 3632 5614 3682 5626
rect 3632 5217 3638 5614
rect 3676 5217 3682 5614
rect 3632 5205 3682 5217
rect 3950 5614 4000 5626
rect 3950 5217 3956 5614
rect 3994 5217 4000 5614
rect 3950 5205 4000 5217
rect 4268 5614 4318 5626
rect 4268 5217 4274 5614
rect 4312 5217 4318 5614
rect 4268 5205 4318 5217
rect 4586 5614 4636 5626
rect 4586 5217 4592 5614
rect 4630 5217 4636 5614
rect 4586 5205 4636 5217
rect 4904 5614 4954 5626
rect 4904 5217 4910 5614
rect 4948 5217 4954 5614
rect 4904 5205 4954 5217
rect 5222 5614 5272 5626
rect 5222 5217 5228 5614
rect 5266 5217 5272 5614
rect 5222 5205 5272 5217
rect 5540 5614 5590 5626
rect 5540 5217 5546 5614
rect 5584 5217 5590 5614
rect 5540 5205 5590 5217
rect 5858 5614 5908 5626
rect 5858 5217 5864 5614
rect 5902 5217 5908 5614
rect 5858 5205 5908 5217
rect 6176 5614 6226 5626
rect 6176 5217 6182 5614
rect 6220 5217 6226 5614
rect 6176 5205 6226 5217
rect 6494 5614 6544 5626
rect 6494 5217 6500 5614
rect 6538 5217 6544 5614
rect 6494 5205 6544 5217
rect 6812 5614 6862 5626
rect 6812 5217 6818 5614
rect 6856 5217 6862 5614
rect 6812 5205 6862 5217
rect 7130 5614 7180 5626
rect 7130 5217 7136 5614
rect 7174 5217 7180 5614
rect 7130 5205 7180 5217
rect 7448 5614 7498 5626
rect 7448 5217 7454 5614
rect 7492 5217 7498 5614
rect 7448 5205 7498 5217
rect 7766 5614 7816 5626
rect 7766 5217 7772 5614
rect 7810 5217 7816 5614
rect 7766 5205 7816 5217
rect -7816 -5217 -7766 -5205
rect -7816 -5614 -7810 -5217
rect -7772 -5614 -7766 -5217
rect -7816 -5626 -7766 -5614
rect -7498 -5217 -7448 -5205
rect -7498 -5614 -7492 -5217
rect -7454 -5614 -7448 -5217
rect -7498 -5626 -7448 -5614
rect -7180 -5217 -7130 -5205
rect -7180 -5614 -7174 -5217
rect -7136 -5614 -7130 -5217
rect -7180 -5626 -7130 -5614
rect -6862 -5217 -6812 -5205
rect -6862 -5614 -6856 -5217
rect -6818 -5614 -6812 -5217
rect -6862 -5626 -6812 -5614
rect -6544 -5217 -6494 -5205
rect -6544 -5614 -6538 -5217
rect -6500 -5614 -6494 -5217
rect -6544 -5626 -6494 -5614
rect -6226 -5217 -6176 -5205
rect -6226 -5614 -6220 -5217
rect -6182 -5614 -6176 -5217
rect -6226 -5626 -6176 -5614
rect -5908 -5217 -5858 -5205
rect -5908 -5614 -5902 -5217
rect -5864 -5614 -5858 -5217
rect -5908 -5626 -5858 -5614
rect -5590 -5217 -5540 -5205
rect -5590 -5614 -5584 -5217
rect -5546 -5614 -5540 -5217
rect -5590 -5626 -5540 -5614
rect -5272 -5217 -5222 -5205
rect -5272 -5614 -5266 -5217
rect -5228 -5614 -5222 -5217
rect -5272 -5626 -5222 -5614
rect -4954 -5217 -4904 -5205
rect -4954 -5614 -4948 -5217
rect -4910 -5614 -4904 -5217
rect -4954 -5626 -4904 -5614
rect -4636 -5217 -4586 -5205
rect -4636 -5614 -4630 -5217
rect -4592 -5614 -4586 -5217
rect -4636 -5626 -4586 -5614
rect -4318 -5217 -4268 -5205
rect -4318 -5614 -4312 -5217
rect -4274 -5614 -4268 -5217
rect -4318 -5626 -4268 -5614
rect -4000 -5217 -3950 -5205
rect -4000 -5614 -3994 -5217
rect -3956 -5614 -3950 -5217
rect -4000 -5626 -3950 -5614
rect -3682 -5217 -3632 -5205
rect -3682 -5614 -3676 -5217
rect -3638 -5614 -3632 -5217
rect -3682 -5626 -3632 -5614
rect -3364 -5217 -3314 -5205
rect -3364 -5614 -3358 -5217
rect -3320 -5614 -3314 -5217
rect -3364 -5626 -3314 -5614
rect -3046 -5217 -2996 -5205
rect -3046 -5614 -3040 -5217
rect -3002 -5614 -2996 -5217
rect -3046 -5626 -2996 -5614
rect -2728 -5217 -2678 -5205
rect -2728 -5614 -2722 -5217
rect -2684 -5614 -2678 -5217
rect -2728 -5626 -2678 -5614
rect -2410 -5217 -2360 -5205
rect -2410 -5614 -2404 -5217
rect -2366 -5614 -2360 -5217
rect -2410 -5626 -2360 -5614
rect -2092 -5217 -2042 -5205
rect -2092 -5614 -2086 -5217
rect -2048 -5614 -2042 -5217
rect -2092 -5626 -2042 -5614
rect -1774 -5217 -1724 -5205
rect -1774 -5614 -1768 -5217
rect -1730 -5614 -1724 -5217
rect -1774 -5626 -1724 -5614
rect -1456 -5217 -1406 -5205
rect -1456 -5614 -1450 -5217
rect -1412 -5614 -1406 -5217
rect -1456 -5626 -1406 -5614
rect -1138 -5217 -1088 -5205
rect -1138 -5614 -1132 -5217
rect -1094 -5614 -1088 -5217
rect -1138 -5626 -1088 -5614
rect -820 -5217 -770 -5205
rect -820 -5614 -814 -5217
rect -776 -5614 -770 -5217
rect -820 -5626 -770 -5614
rect -502 -5217 -452 -5205
rect -502 -5614 -496 -5217
rect -458 -5614 -452 -5217
rect -502 -5626 -452 -5614
rect -184 -5217 -134 -5205
rect -184 -5614 -178 -5217
rect -140 -5614 -134 -5217
rect -184 -5626 -134 -5614
rect 134 -5217 184 -5205
rect 134 -5614 140 -5217
rect 178 -5614 184 -5217
rect 134 -5626 184 -5614
rect 452 -5217 502 -5205
rect 452 -5614 458 -5217
rect 496 -5614 502 -5217
rect 452 -5626 502 -5614
rect 770 -5217 820 -5205
rect 770 -5614 776 -5217
rect 814 -5614 820 -5217
rect 770 -5626 820 -5614
rect 1088 -5217 1138 -5205
rect 1088 -5614 1094 -5217
rect 1132 -5614 1138 -5217
rect 1088 -5626 1138 -5614
rect 1406 -5217 1456 -5205
rect 1406 -5614 1412 -5217
rect 1450 -5614 1456 -5217
rect 1406 -5626 1456 -5614
rect 1724 -5217 1774 -5205
rect 1724 -5614 1730 -5217
rect 1768 -5614 1774 -5217
rect 1724 -5626 1774 -5614
rect 2042 -5217 2092 -5205
rect 2042 -5614 2048 -5217
rect 2086 -5614 2092 -5217
rect 2042 -5626 2092 -5614
rect 2360 -5217 2410 -5205
rect 2360 -5614 2366 -5217
rect 2404 -5614 2410 -5217
rect 2360 -5626 2410 -5614
rect 2678 -5217 2728 -5205
rect 2678 -5614 2684 -5217
rect 2722 -5614 2728 -5217
rect 2678 -5626 2728 -5614
rect 2996 -5217 3046 -5205
rect 2996 -5614 3002 -5217
rect 3040 -5614 3046 -5217
rect 2996 -5626 3046 -5614
rect 3314 -5217 3364 -5205
rect 3314 -5614 3320 -5217
rect 3358 -5614 3364 -5217
rect 3314 -5626 3364 -5614
rect 3632 -5217 3682 -5205
rect 3632 -5614 3638 -5217
rect 3676 -5614 3682 -5217
rect 3632 -5626 3682 -5614
rect 3950 -5217 4000 -5205
rect 3950 -5614 3956 -5217
rect 3994 -5614 4000 -5217
rect 3950 -5626 4000 -5614
rect 4268 -5217 4318 -5205
rect 4268 -5614 4274 -5217
rect 4312 -5614 4318 -5217
rect 4268 -5626 4318 -5614
rect 4586 -5217 4636 -5205
rect 4586 -5614 4592 -5217
rect 4630 -5614 4636 -5217
rect 4586 -5626 4636 -5614
rect 4904 -5217 4954 -5205
rect 4904 -5614 4910 -5217
rect 4948 -5614 4954 -5217
rect 4904 -5626 4954 -5614
rect 5222 -5217 5272 -5205
rect 5222 -5614 5228 -5217
rect 5266 -5614 5272 -5217
rect 5222 -5626 5272 -5614
rect 5540 -5217 5590 -5205
rect 5540 -5614 5546 -5217
rect 5584 -5614 5590 -5217
rect 5540 -5626 5590 -5614
rect 5858 -5217 5908 -5205
rect 5858 -5614 5864 -5217
rect 5902 -5614 5908 -5217
rect 5858 -5626 5908 -5614
rect 6176 -5217 6226 -5205
rect 6176 -5614 6182 -5217
rect 6220 -5614 6226 -5217
rect 6176 -5626 6226 -5614
rect 6494 -5217 6544 -5205
rect 6494 -5614 6500 -5217
rect 6538 -5614 6544 -5217
rect 6494 -5626 6544 -5614
rect 6812 -5217 6862 -5205
rect 6812 -5614 6818 -5217
rect 6856 -5614 6862 -5217
rect 6812 -5626 6862 -5614
rect 7130 -5217 7180 -5205
rect 7130 -5614 7136 -5217
rect 7174 -5614 7180 -5217
rect 7130 -5626 7180 -5614
rect 7448 -5217 7498 -5205
rect 7448 -5614 7454 -5217
rect 7492 -5614 7498 -5217
rect 7448 -5626 7498 -5614
rect 7766 -5217 7816 -5205
rect 7766 -5614 7772 -5217
rect 7810 -5614 7816 -5217
rect 7766 -5626 7816 -5614
<< res0p35 >>
rect -7828 -5202 -7754 5202
rect -7510 -5202 -7436 5202
rect -7192 -5202 -7118 5202
rect -6874 -5202 -6800 5202
rect -6556 -5202 -6482 5202
rect -6238 -5202 -6164 5202
rect -5920 -5202 -5846 5202
rect -5602 -5202 -5528 5202
rect -5284 -5202 -5210 5202
rect -4966 -5202 -4892 5202
rect -4648 -5202 -4574 5202
rect -4330 -5202 -4256 5202
rect -4012 -5202 -3938 5202
rect -3694 -5202 -3620 5202
rect -3376 -5202 -3302 5202
rect -3058 -5202 -2984 5202
rect -2740 -5202 -2666 5202
rect -2422 -5202 -2348 5202
rect -2104 -5202 -2030 5202
rect -1786 -5202 -1712 5202
rect -1468 -5202 -1394 5202
rect -1150 -5202 -1076 5202
rect -832 -5202 -758 5202
rect -514 -5202 -440 5202
rect -196 -5202 -122 5202
rect 122 -5202 196 5202
rect 440 -5202 514 5202
rect 758 -5202 832 5202
rect 1076 -5202 1150 5202
rect 1394 -5202 1468 5202
rect 1712 -5202 1786 5202
rect 2030 -5202 2104 5202
rect 2348 -5202 2422 5202
rect 2666 -5202 2740 5202
rect 2984 -5202 3058 5202
rect 3302 -5202 3376 5202
rect 3620 -5202 3694 5202
rect 3938 -5202 4012 5202
rect 4256 -5202 4330 5202
rect 4574 -5202 4648 5202
rect 4892 -5202 4966 5202
rect 5210 -5202 5284 5202
rect 5528 -5202 5602 5202
rect 5846 -5202 5920 5202
rect 6164 -5202 6238 5202
rect 6482 -5202 6556 5202
rect 6800 -5202 6874 5202
rect 7118 -5202 7192 5202
rect 7436 -5202 7510 5202
rect 7754 -5202 7828 5202
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 52 m 1 nx 50 wmin 0.350 lmin 0.50 rho 2000 val 298.218k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
