magic
tech sky130A
magscale 1 2
timestamp 1666839628
<< error_p >>
rect -855 18 855 236
<< nwell >>
rect -855 18 855 1218
rect -855 -1218 855 -18
<< pmos >>
rect -761 118 -661 1118
rect -603 118 -503 1118
rect -445 118 -345 1118
rect -287 118 -187 1118
rect -129 118 -29 1118
rect 29 118 129 1118
rect 187 118 287 1118
rect 345 118 445 1118
rect 503 118 603 1118
rect 661 118 761 1118
rect -761 -1118 -661 -118
rect -603 -1118 -503 -118
rect -445 -1118 -345 -118
rect -287 -1118 -187 -118
rect -129 -1118 -29 -118
rect 29 -1118 129 -118
rect 187 -1118 287 -118
rect 345 -1118 445 -118
rect 503 -1118 603 -118
rect 661 -1118 761 -118
<< pdiff >>
rect -819 1106 -761 1118
rect -819 130 -807 1106
rect -773 130 -761 1106
rect -819 118 -761 130
rect -661 1106 -603 1118
rect -661 130 -649 1106
rect -615 130 -603 1106
rect -661 118 -603 130
rect -503 1106 -445 1118
rect -503 130 -491 1106
rect -457 130 -445 1106
rect -503 118 -445 130
rect -345 1106 -287 1118
rect -345 130 -333 1106
rect -299 130 -287 1106
rect -345 118 -287 130
rect -187 1106 -129 1118
rect -187 130 -175 1106
rect -141 130 -129 1106
rect -187 118 -129 130
rect -29 1106 29 1118
rect -29 130 -17 1106
rect 17 130 29 1106
rect -29 118 29 130
rect 129 1106 187 1118
rect 129 130 141 1106
rect 175 130 187 1106
rect 129 118 187 130
rect 287 1106 345 1118
rect 287 130 299 1106
rect 333 130 345 1106
rect 287 118 345 130
rect 445 1106 503 1118
rect 445 130 457 1106
rect 491 130 503 1106
rect 445 118 503 130
rect 603 1106 661 1118
rect 603 130 615 1106
rect 649 130 661 1106
rect 603 118 661 130
rect 761 1106 819 1118
rect 761 130 773 1106
rect 807 130 819 1106
rect 761 118 819 130
rect -819 -130 -761 -118
rect -819 -1106 -807 -130
rect -773 -1106 -761 -130
rect -819 -1118 -761 -1106
rect -661 -130 -603 -118
rect -661 -1106 -649 -130
rect -615 -1106 -603 -130
rect -661 -1118 -603 -1106
rect -503 -130 -445 -118
rect -503 -1106 -491 -130
rect -457 -1106 -445 -130
rect -503 -1118 -445 -1106
rect -345 -130 -287 -118
rect -345 -1106 -333 -130
rect -299 -1106 -287 -130
rect -345 -1118 -287 -1106
rect -187 -130 -129 -118
rect -187 -1106 -175 -130
rect -141 -1106 -129 -130
rect -187 -1118 -129 -1106
rect -29 -130 29 -118
rect -29 -1106 -17 -130
rect 17 -1106 29 -130
rect -29 -1118 29 -1106
rect 129 -130 187 -118
rect 129 -1106 141 -130
rect 175 -1106 187 -130
rect 129 -1118 187 -1106
rect 287 -130 345 -118
rect 287 -1106 299 -130
rect 333 -1106 345 -130
rect 287 -1118 345 -1106
rect 445 -130 503 -118
rect 445 -1106 457 -130
rect 491 -1106 503 -130
rect 445 -1118 503 -1106
rect 603 -130 661 -118
rect 603 -1106 615 -130
rect 649 -1106 661 -130
rect 603 -1118 661 -1106
rect 761 -130 819 -118
rect 761 -1106 773 -130
rect 807 -1106 819 -130
rect 761 -1118 819 -1106
<< pdiffc >>
rect -807 130 -773 1106
rect -649 130 -615 1106
rect -491 130 -457 1106
rect -333 130 -299 1106
rect -175 130 -141 1106
rect -17 130 17 1106
rect 141 130 175 1106
rect 299 130 333 1106
rect 457 130 491 1106
rect 615 130 649 1106
rect 773 130 807 1106
rect -807 -1106 -773 -130
rect -649 -1106 -615 -130
rect -491 -1106 -457 -130
rect -333 -1106 -299 -130
rect -175 -1106 -141 -130
rect -17 -1106 17 -130
rect 141 -1106 175 -130
rect 299 -1106 333 -130
rect 457 -1106 491 -130
rect 615 -1106 649 -130
rect 773 -1106 807 -130
<< poly >>
rect -761 1199 -661 1215
rect -761 1165 -745 1199
rect -677 1165 -661 1199
rect -761 1118 -661 1165
rect -603 1199 -503 1215
rect -603 1165 -587 1199
rect -519 1165 -503 1199
rect -603 1118 -503 1165
rect -445 1199 -345 1215
rect -445 1165 -429 1199
rect -361 1165 -345 1199
rect -445 1118 -345 1165
rect -287 1199 -187 1215
rect -287 1165 -271 1199
rect -203 1165 -187 1199
rect -287 1118 -187 1165
rect -129 1199 -29 1215
rect -129 1165 -113 1199
rect -45 1165 -29 1199
rect -129 1118 -29 1165
rect 29 1199 129 1215
rect 29 1165 45 1199
rect 113 1165 129 1199
rect 29 1118 129 1165
rect 187 1199 287 1215
rect 187 1165 203 1199
rect 271 1165 287 1199
rect 187 1118 287 1165
rect 345 1199 445 1215
rect 345 1165 361 1199
rect 429 1165 445 1199
rect 345 1118 445 1165
rect 503 1199 603 1215
rect 503 1165 519 1199
rect 587 1165 603 1199
rect 503 1118 603 1165
rect 661 1199 761 1215
rect 661 1165 677 1199
rect 745 1165 761 1199
rect 661 1118 761 1165
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect -761 -1165 -661 -1118
rect -761 -1199 -745 -1165
rect -677 -1199 -661 -1165
rect -761 -1215 -661 -1199
rect -603 -1165 -503 -1118
rect -603 -1199 -587 -1165
rect -519 -1199 -503 -1165
rect -603 -1215 -503 -1199
rect -445 -1165 -345 -1118
rect -445 -1199 -429 -1165
rect -361 -1199 -345 -1165
rect -445 -1215 -345 -1199
rect -287 -1165 -187 -1118
rect -287 -1199 -271 -1165
rect -203 -1199 -187 -1165
rect -287 -1215 -187 -1199
rect -129 -1165 -29 -1118
rect -129 -1199 -113 -1165
rect -45 -1199 -29 -1165
rect -129 -1215 -29 -1199
rect 29 -1165 129 -1118
rect 29 -1199 45 -1165
rect 113 -1199 129 -1165
rect 29 -1215 129 -1199
rect 187 -1165 287 -1118
rect 187 -1199 203 -1165
rect 271 -1199 287 -1165
rect 187 -1215 287 -1199
rect 345 -1165 445 -1118
rect 345 -1199 361 -1165
rect 429 -1199 445 -1165
rect 345 -1215 445 -1199
rect 503 -1165 603 -1118
rect 503 -1199 519 -1165
rect 587 -1199 603 -1165
rect 503 -1215 603 -1199
rect 661 -1165 761 -1118
rect 661 -1199 677 -1165
rect 745 -1199 761 -1165
rect 661 -1215 761 -1199
<< polycont >>
rect -745 1165 -677 1199
rect -587 1165 -519 1199
rect -429 1165 -361 1199
rect -271 1165 -203 1199
rect -113 1165 -45 1199
rect 45 1165 113 1199
rect 203 1165 271 1199
rect 361 1165 429 1199
rect 519 1165 587 1199
rect 677 1165 745 1199
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect -745 -1199 -677 -1165
rect -587 -1199 -519 -1165
rect -429 -1199 -361 -1165
rect -271 -1199 -203 -1165
rect -113 -1199 -45 -1165
rect 45 -1199 113 -1165
rect 203 -1199 271 -1165
rect 361 -1199 429 -1165
rect 519 -1199 587 -1165
rect 677 -1199 745 -1165
<< locali >>
rect -761 1165 -745 1199
rect -677 1165 -661 1199
rect -603 1165 -587 1199
rect -519 1165 -503 1199
rect -445 1165 -429 1199
rect -361 1165 -345 1199
rect -287 1165 -271 1199
rect -203 1165 -187 1199
rect -129 1165 -113 1199
rect -45 1165 -29 1199
rect 29 1165 45 1199
rect 113 1165 129 1199
rect 187 1165 203 1199
rect 271 1165 287 1199
rect 345 1165 361 1199
rect 429 1165 445 1199
rect 503 1165 519 1199
rect 587 1165 603 1199
rect 661 1165 677 1199
rect 745 1165 761 1199
rect -807 1106 -773 1122
rect -807 114 -773 130
rect -649 1106 -615 1122
rect -649 114 -615 130
rect -491 1106 -457 1122
rect -491 114 -457 130
rect -333 1106 -299 1122
rect -333 114 -299 130
rect -175 1106 -141 1122
rect -175 114 -141 130
rect -17 1106 17 1122
rect -17 114 17 130
rect 141 1106 175 1122
rect 141 114 175 130
rect 299 1106 333 1122
rect 299 114 333 130
rect 457 1106 491 1122
rect 457 114 491 130
rect 615 1106 649 1122
rect 615 114 649 130
rect 773 1106 807 1122
rect 773 114 807 130
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect -807 -130 -773 -114
rect -807 -1122 -773 -1106
rect -649 -130 -615 -114
rect -649 -1122 -615 -1106
rect -491 -130 -457 -114
rect -491 -1122 -457 -1106
rect -333 -130 -299 -114
rect -333 -1122 -299 -1106
rect -175 -130 -141 -114
rect -175 -1122 -141 -1106
rect -17 -130 17 -114
rect -17 -1122 17 -1106
rect 141 -130 175 -114
rect 141 -1122 175 -1106
rect 299 -130 333 -114
rect 299 -1122 333 -1106
rect 457 -130 491 -114
rect 457 -1122 491 -1106
rect 615 -130 649 -114
rect 615 -1122 649 -1106
rect 773 -130 807 -114
rect 773 -1122 807 -1106
rect -761 -1199 -745 -1165
rect -677 -1199 -661 -1165
rect -603 -1199 -587 -1165
rect -519 -1199 -503 -1165
rect -445 -1199 -429 -1165
rect -361 -1199 -345 -1165
rect -287 -1199 -271 -1165
rect -203 -1199 -187 -1165
rect -129 -1199 -113 -1165
rect -45 -1199 -29 -1165
rect 29 -1199 45 -1165
rect 113 -1199 129 -1165
rect 187 -1199 203 -1165
rect 271 -1199 287 -1165
rect 345 -1199 361 -1165
rect 429 -1199 445 -1165
rect 503 -1199 519 -1165
rect 587 -1199 603 -1165
rect 661 -1199 677 -1165
rect 745 -1199 761 -1165
<< viali >>
rect -745 1165 -677 1199
rect -587 1165 -519 1199
rect -429 1165 -361 1199
rect -271 1165 -203 1199
rect -113 1165 -45 1199
rect 45 1165 113 1199
rect 203 1165 271 1199
rect 361 1165 429 1199
rect 519 1165 587 1199
rect 677 1165 745 1199
rect -807 130 -773 1106
rect -649 130 -615 1106
rect -491 130 -457 1106
rect -333 130 -299 1106
rect -175 130 -141 1106
rect -17 130 17 1106
rect 141 130 175 1106
rect 299 130 333 1106
rect 457 130 491 1106
rect 615 130 649 1106
rect 773 130 807 1106
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect -807 -1106 -773 -130
rect -649 -1106 -615 -130
rect -491 -1106 -457 -130
rect -333 -1106 -299 -130
rect -175 -1106 -141 -130
rect -17 -1106 17 -130
rect 141 -1106 175 -130
rect 299 -1106 333 -130
rect 457 -1106 491 -130
rect 615 -1106 649 -130
rect 773 -1106 807 -130
rect -745 -1199 -677 -1165
rect -587 -1199 -519 -1165
rect -429 -1199 -361 -1165
rect -271 -1199 -203 -1165
rect -113 -1199 -45 -1165
rect 45 -1199 113 -1165
rect 203 -1199 271 -1165
rect 361 -1199 429 -1165
rect 519 -1199 587 -1165
rect 677 -1199 745 -1165
<< metal1 >>
rect -757 1199 -665 1205
rect -757 1165 -745 1199
rect -677 1165 -665 1199
rect -757 1159 -665 1165
rect -599 1199 -507 1205
rect -599 1165 -587 1199
rect -519 1165 -507 1199
rect -599 1159 -507 1165
rect -441 1199 -349 1205
rect -441 1165 -429 1199
rect -361 1165 -349 1199
rect -441 1159 -349 1165
rect -283 1199 -191 1205
rect -283 1165 -271 1199
rect -203 1165 -191 1199
rect -283 1159 -191 1165
rect -125 1199 -33 1205
rect -125 1165 -113 1199
rect -45 1165 -33 1199
rect -125 1159 -33 1165
rect 33 1199 125 1205
rect 33 1165 45 1199
rect 113 1165 125 1199
rect 33 1159 125 1165
rect 191 1199 283 1205
rect 191 1165 203 1199
rect 271 1165 283 1199
rect 191 1159 283 1165
rect 349 1199 441 1205
rect 349 1165 361 1199
rect 429 1165 441 1199
rect 349 1159 441 1165
rect 507 1199 599 1205
rect 507 1165 519 1199
rect 587 1165 599 1199
rect 507 1159 599 1165
rect 665 1199 757 1205
rect 665 1165 677 1199
rect 745 1165 757 1199
rect 665 1159 757 1165
rect -813 1106 -767 1118
rect -813 130 -807 1106
rect -773 130 -767 1106
rect -813 118 -767 130
rect -655 1106 -609 1118
rect -655 130 -649 1106
rect -615 130 -609 1106
rect -655 118 -609 130
rect -497 1106 -451 1118
rect -497 130 -491 1106
rect -457 130 -451 1106
rect -497 118 -451 130
rect -339 1106 -293 1118
rect -339 130 -333 1106
rect -299 130 -293 1106
rect -339 118 -293 130
rect -181 1106 -135 1118
rect -181 130 -175 1106
rect -141 130 -135 1106
rect -181 118 -135 130
rect -23 1106 23 1118
rect -23 130 -17 1106
rect 17 130 23 1106
rect -23 118 23 130
rect 135 1106 181 1118
rect 135 130 141 1106
rect 175 130 181 1106
rect 135 118 181 130
rect 293 1106 339 1118
rect 293 130 299 1106
rect 333 130 339 1106
rect 293 118 339 130
rect 451 1106 497 1118
rect 451 130 457 1106
rect 491 130 497 1106
rect 451 118 497 130
rect 609 1106 655 1118
rect 609 130 615 1106
rect 649 130 655 1106
rect 609 118 655 130
rect 767 1106 813 1118
rect 767 130 773 1106
rect 807 130 813 1106
rect 767 118 813 130
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect -813 -130 -767 -118
rect -813 -1106 -807 -130
rect -773 -1106 -767 -130
rect -813 -1118 -767 -1106
rect -655 -130 -609 -118
rect -655 -1106 -649 -130
rect -615 -1106 -609 -130
rect -655 -1118 -609 -1106
rect -497 -130 -451 -118
rect -497 -1106 -491 -130
rect -457 -1106 -451 -130
rect -497 -1118 -451 -1106
rect -339 -130 -293 -118
rect -339 -1106 -333 -130
rect -299 -1106 -293 -130
rect -339 -1118 -293 -1106
rect -181 -130 -135 -118
rect -181 -1106 -175 -130
rect -141 -1106 -135 -130
rect -181 -1118 -135 -1106
rect -23 -130 23 -118
rect -23 -1106 -17 -130
rect 17 -1106 23 -130
rect -23 -1118 23 -1106
rect 135 -130 181 -118
rect 135 -1106 141 -130
rect 175 -1106 181 -130
rect 135 -1118 181 -1106
rect 293 -130 339 -118
rect 293 -1106 299 -130
rect 333 -1106 339 -130
rect 293 -1118 339 -1106
rect 451 -130 497 -118
rect 451 -1106 457 -130
rect 491 -1106 497 -130
rect 451 -1118 497 -1106
rect 609 -130 655 -118
rect 609 -1106 615 -130
rect 649 -1106 655 -130
rect 609 -1118 655 -1106
rect 767 -130 813 -118
rect 767 -1106 773 -130
rect 807 -1106 813 -130
rect 767 -1118 813 -1106
rect -757 -1165 -665 -1159
rect -757 -1199 -745 -1165
rect -677 -1199 -665 -1165
rect -757 -1205 -665 -1199
rect -599 -1165 -507 -1159
rect -599 -1199 -587 -1165
rect -519 -1199 -507 -1165
rect -599 -1205 -507 -1199
rect -441 -1165 -349 -1159
rect -441 -1199 -429 -1165
rect -361 -1199 -349 -1165
rect -441 -1205 -349 -1199
rect -283 -1165 -191 -1159
rect -283 -1199 -271 -1165
rect -203 -1199 -191 -1165
rect -283 -1205 -191 -1199
rect -125 -1165 -33 -1159
rect -125 -1199 -113 -1165
rect -45 -1199 -33 -1165
rect -125 -1205 -33 -1199
rect 33 -1165 125 -1159
rect 33 -1199 45 -1165
rect 113 -1199 125 -1165
rect 33 -1205 125 -1199
rect 191 -1165 283 -1159
rect 191 -1199 203 -1165
rect 271 -1199 283 -1165
rect 191 -1205 283 -1199
rect 349 -1165 441 -1159
rect 349 -1199 361 -1165
rect 429 -1199 441 -1165
rect 349 -1205 441 -1199
rect 507 -1165 599 -1159
rect 507 -1199 519 -1165
rect 587 -1199 599 -1165
rect 507 -1205 599 -1199
rect 665 -1165 757 -1159
rect 665 -1199 677 -1165
rect 745 -1199 757 -1165
rect 665 -1205 757 -1199
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
