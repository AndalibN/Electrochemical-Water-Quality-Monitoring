magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nwell >>
rect -697 -1350 697 1350
<< pmos >>
rect -603 -1250 -503 1250
rect -445 -1250 -345 1250
rect -287 -1250 -187 1250
rect -129 -1250 -29 1250
rect 29 -1250 129 1250
rect 187 -1250 287 1250
rect 345 -1250 445 1250
rect 503 -1250 603 1250
<< pdiff >>
rect -661 1238 -603 1250
rect -661 -1238 -649 1238
rect -615 -1238 -603 1238
rect -661 -1250 -603 -1238
rect -503 1238 -445 1250
rect -503 -1238 -491 1238
rect -457 -1238 -445 1238
rect -503 -1250 -445 -1238
rect -345 1238 -287 1250
rect -345 -1238 -333 1238
rect -299 -1238 -287 1238
rect -345 -1250 -287 -1238
rect -187 1238 -129 1250
rect -187 -1238 -175 1238
rect -141 -1238 -129 1238
rect -187 -1250 -129 -1238
rect -29 1238 29 1250
rect -29 -1238 -17 1238
rect 17 -1238 29 1238
rect -29 -1250 29 -1238
rect 129 1238 187 1250
rect 129 -1238 141 1238
rect 175 -1238 187 1238
rect 129 -1250 187 -1238
rect 287 1238 345 1250
rect 287 -1238 299 1238
rect 333 -1238 345 1238
rect 287 -1250 345 -1238
rect 445 1238 503 1250
rect 445 -1238 457 1238
rect 491 -1238 503 1238
rect 445 -1250 503 -1238
rect 603 1238 661 1250
rect 603 -1238 615 1238
rect 649 -1238 661 1238
rect 603 -1250 661 -1238
<< pdiffc >>
rect -649 -1238 -615 1238
rect -491 -1238 -457 1238
rect -333 -1238 -299 1238
rect -175 -1238 -141 1238
rect -17 -1238 17 1238
rect 141 -1238 175 1238
rect 299 -1238 333 1238
rect 457 -1238 491 1238
rect 615 -1238 649 1238
<< poly >>
rect -603 1331 -503 1347
rect -603 1297 -587 1331
rect -519 1297 -503 1331
rect -603 1250 -503 1297
rect -445 1331 -345 1347
rect -445 1297 -429 1331
rect -361 1297 -345 1331
rect -445 1250 -345 1297
rect -287 1331 -187 1347
rect -287 1297 -271 1331
rect -203 1297 -187 1331
rect -287 1250 -187 1297
rect -129 1331 -29 1347
rect -129 1297 -113 1331
rect -45 1297 -29 1331
rect -129 1250 -29 1297
rect 29 1331 129 1347
rect 29 1297 45 1331
rect 113 1297 129 1331
rect 29 1250 129 1297
rect 187 1331 287 1347
rect 187 1297 203 1331
rect 271 1297 287 1331
rect 187 1250 287 1297
rect 345 1331 445 1347
rect 345 1297 361 1331
rect 429 1297 445 1331
rect 345 1250 445 1297
rect 503 1331 603 1347
rect 503 1297 519 1331
rect 587 1297 603 1331
rect 503 1250 603 1297
rect -603 -1297 -503 -1250
rect -603 -1331 -587 -1297
rect -519 -1331 -503 -1297
rect -603 -1347 -503 -1331
rect -445 -1297 -345 -1250
rect -445 -1331 -429 -1297
rect -361 -1331 -345 -1297
rect -445 -1347 -345 -1331
rect -287 -1297 -187 -1250
rect -287 -1331 -271 -1297
rect -203 -1331 -187 -1297
rect -287 -1347 -187 -1331
rect -129 -1297 -29 -1250
rect -129 -1331 -113 -1297
rect -45 -1331 -29 -1297
rect -129 -1347 -29 -1331
rect 29 -1297 129 -1250
rect 29 -1331 45 -1297
rect 113 -1331 129 -1297
rect 29 -1347 129 -1331
rect 187 -1297 287 -1250
rect 187 -1331 203 -1297
rect 271 -1331 287 -1297
rect 187 -1347 287 -1331
rect 345 -1297 445 -1250
rect 345 -1331 361 -1297
rect 429 -1331 445 -1297
rect 345 -1347 445 -1331
rect 503 -1297 603 -1250
rect 503 -1331 519 -1297
rect 587 -1331 603 -1297
rect 503 -1347 603 -1331
<< polycont >>
rect -587 1297 -519 1331
rect -429 1297 -361 1331
rect -271 1297 -203 1331
rect -113 1297 -45 1331
rect 45 1297 113 1331
rect 203 1297 271 1331
rect 361 1297 429 1331
rect 519 1297 587 1331
rect -587 -1331 -519 -1297
rect -429 -1331 -361 -1297
rect -271 -1331 -203 -1297
rect -113 -1331 -45 -1297
rect 45 -1331 113 -1297
rect 203 -1331 271 -1297
rect 361 -1331 429 -1297
rect 519 -1331 587 -1297
<< locali >>
rect -603 1297 -587 1331
rect -519 1297 -503 1331
rect -445 1297 -429 1331
rect -361 1297 -345 1331
rect -287 1297 -271 1331
rect -203 1297 -187 1331
rect -129 1297 -113 1331
rect -45 1297 -29 1331
rect 29 1297 45 1331
rect 113 1297 129 1331
rect 187 1297 203 1331
rect 271 1297 287 1331
rect 345 1297 361 1331
rect 429 1297 445 1331
rect 503 1297 519 1331
rect 587 1297 603 1331
rect -649 1238 -615 1254
rect -649 -1254 -615 -1238
rect -491 1238 -457 1254
rect -491 -1254 -457 -1238
rect -333 1238 -299 1254
rect -333 -1254 -299 -1238
rect -175 1238 -141 1254
rect -175 -1254 -141 -1238
rect -17 1238 17 1254
rect -17 -1254 17 -1238
rect 141 1238 175 1254
rect 141 -1254 175 -1238
rect 299 1238 333 1254
rect 299 -1254 333 -1238
rect 457 1238 491 1254
rect 457 -1254 491 -1238
rect 615 1238 649 1254
rect 615 -1254 649 -1238
rect -603 -1331 -587 -1297
rect -519 -1331 -503 -1297
rect -445 -1331 -429 -1297
rect -361 -1331 -345 -1297
rect -287 -1331 -271 -1297
rect -203 -1331 -187 -1297
rect -129 -1331 -113 -1297
rect -45 -1331 -29 -1297
rect 29 -1331 45 -1297
rect 113 -1331 129 -1297
rect 187 -1331 203 -1297
rect 271 -1331 287 -1297
rect 345 -1331 361 -1297
rect 429 -1331 445 -1297
rect 503 -1331 519 -1297
rect 587 -1331 603 -1297
<< viali >>
rect -587 1297 -519 1331
rect -429 1297 -361 1331
rect -271 1297 -203 1331
rect -113 1297 -45 1331
rect 45 1297 113 1331
rect 203 1297 271 1331
rect 361 1297 429 1331
rect 519 1297 587 1331
rect -649 -1238 -615 1238
rect -491 -1238 -457 1238
rect -333 -1238 -299 1238
rect -175 -1238 -141 1238
rect -17 -1238 17 1238
rect 141 -1238 175 1238
rect 299 -1238 333 1238
rect 457 -1238 491 1238
rect 615 -1238 649 1238
rect -587 -1331 -519 -1297
rect -429 -1331 -361 -1297
rect -271 -1331 -203 -1297
rect -113 -1331 -45 -1297
rect 45 -1331 113 -1297
rect 203 -1331 271 -1297
rect 361 -1331 429 -1297
rect 519 -1331 587 -1297
<< metal1 >>
rect -599 1331 -507 1337
rect -599 1297 -587 1331
rect -519 1297 -507 1331
rect -599 1291 -507 1297
rect -441 1331 -349 1337
rect -441 1297 -429 1331
rect -361 1297 -349 1331
rect -441 1291 -349 1297
rect -283 1331 -191 1337
rect -283 1297 -271 1331
rect -203 1297 -191 1331
rect -283 1291 -191 1297
rect -125 1331 -33 1337
rect -125 1297 -113 1331
rect -45 1297 -33 1331
rect -125 1291 -33 1297
rect 33 1331 125 1337
rect 33 1297 45 1331
rect 113 1297 125 1331
rect 33 1291 125 1297
rect 191 1331 283 1337
rect 191 1297 203 1331
rect 271 1297 283 1331
rect 191 1291 283 1297
rect 349 1331 441 1337
rect 349 1297 361 1331
rect 429 1297 441 1331
rect 349 1291 441 1297
rect 507 1331 599 1337
rect 507 1297 519 1331
rect 587 1297 599 1331
rect 507 1291 599 1297
rect -655 1238 -609 1250
rect -655 -1238 -649 1238
rect -615 -1238 -609 1238
rect -655 -1250 -609 -1238
rect -497 1238 -451 1250
rect -497 -1238 -491 1238
rect -457 -1238 -451 1238
rect -497 -1250 -451 -1238
rect -339 1238 -293 1250
rect -339 -1238 -333 1238
rect -299 -1238 -293 1238
rect -339 -1250 -293 -1238
rect -181 1238 -135 1250
rect -181 -1238 -175 1238
rect -141 -1238 -135 1238
rect -181 -1250 -135 -1238
rect -23 1238 23 1250
rect -23 -1238 -17 1238
rect 17 -1238 23 1238
rect -23 -1250 23 -1238
rect 135 1238 181 1250
rect 135 -1238 141 1238
rect 175 -1238 181 1238
rect 135 -1250 181 -1238
rect 293 1238 339 1250
rect 293 -1238 299 1238
rect 333 -1238 339 1238
rect 293 -1250 339 -1238
rect 451 1238 497 1250
rect 451 -1238 457 1238
rect 491 -1238 497 1238
rect 451 -1250 497 -1238
rect 609 1238 655 1250
rect 609 -1238 615 1238
rect 649 -1238 655 1238
rect 609 -1250 655 -1238
rect -599 -1297 -507 -1291
rect -599 -1331 -587 -1297
rect -519 -1331 -507 -1297
rect -599 -1337 -507 -1331
rect -441 -1297 -349 -1291
rect -441 -1331 -429 -1297
rect -361 -1331 -349 -1297
rect -441 -1337 -349 -1331
rect -283 -1297 -191 -1291
rect -283 -1331 -271 -1297
rect -203 -1331 -191 -1297
rect -283 -1337 -191 -1331
rect -125 -1297 -33 -1291
rect -125 -1331 -113 -1297
rect -45 -1331 -33 -1297
rect -125 -1337 -33 -1331
rect 33 -1297 125 -1291
rect 33 -1331 45 -1297
rect 113 -1331 125 -1297
rect 33 -1337 125 -1331
rect 191 -1297 283 -1291
rect 191 -1331 203 -1297
rect 271 -1331 283 -1297
rect 191 -1337 283 -1331
rect 349 -1297 441 -1291
rect 349 -1331 361 -1297
rect 429 -1331 441 -1297
rect 349 -1337 441 -1331
rect 507 -1297 599 -1291
rect 507 -1331 519 -1297
rect 587 -1331 599 -1297
rect 507 -1337 599 -1331
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 12.5 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
