magic
tech sky130A
magscale 1 2
timestamp 1667488624
<< error_p >>
rect -29 432 29 438
rect -29 398 -17 432
rect -29 392 29 398
rect -29 -398 29 -392
rect -29 -432 -17 -398
rect -29 -438 29 -432
<< pwell >>
rect -214 -570 214 570
<< nmos >>
rect -18 -360 18 360
<< ndiff >>
rect -76 348 -18 360
rect -76 -348 -64 348
rect -30 -348 -18 348
rect -76 -360 -18 -348
rect 18 348 76 360
rect 18 -348 30 348
rect 64 -348 76 348
rect 18 -360 76 -348
<< ndiffc >>
rect -64 -348 -30 348
rect 30 -348 64 348
<< psubdiff >>
rect -178 500 -82 534
rect 82 500 178 534
rect -178 438 -144 500
rect 144 438 178 500
rect -178 -500 -144 -438
rect 144 -500 178 -438
rect -178 -534 -82 -500
rect 82 -534 178 -500
<< psubdiffcont >>
rect -82 500 82 534
rect -178 -438 -144 438
rect 144 -438 178 438
rect -82 -534 82 -500
<< poly >>
rect -33 432 33 448
rect -33 398 -17 432
rect 17 398 33 432
rect -33 382 33 398
rect -18 360 18 382
rect -18 -382 18 -360
rect -33 -398 33 -382
rect -33 -432 -17 -398
rect 17 -432 33 -398
rect -33 -448 33 -432
<< polycont >>
rect -17 398 17 432
rect -17 -432 17 -398
<< locali >>
rect -178 500 -82 534
rect 82 500 178 534
rect -178 438 -144 500
rect 144 438 178 500
rect -33 398 -17 432
rect 17 398 33 432
rect -64 348 -30 364
rect -64 -364 -30 -348
rect 30 348 64 364
rect 30 -364 64 -348
rect -33 -432 -17 -398
rect 17 -432 33 -398
rect -178 -500 -144 -438
rect 144 -500 178 -438
rect -178 -534 -82 -500
rect 82 -534 178 -500
<< viali >>
rect -17 398 17 432
rect -64 -348 -30 348
rect 30 -348 64 348
rect -17 -432 17 -398
<< metal1 >>
rect -29 432 29 438
rect -29 398 -17 432
rect 17 398 29 432
rect -29 392 29 398
rect -70 348 -24 360
rect -70 -348 -64 348
rect -30 -348 -24 348
rect -70 -360 -24 -348
rect 24 348 70 360
rect 24 -348 30 348
rect 64 -348 70 348
rect 24 -360 70 -348
rect -29 -398 29 -392
rect -29 -432 -17 -398
rect 17 -432 29 -398
rect -29 -438 29 -432
<< properties >>
string FIXED_BBOX -161 -517 161 517
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.6 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
