magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect 58 -1844 122 -1838
rect 58 -1878 73 -1844
rect 58 -1884 122 -1878
<< pwell >>
rect -185 -1832 210 1832
<< nmos >>
rect -101 -1806 -29 1806
rect 54 -1806 126 1806
<< ndiff >>
rect -159 1785 -101 1806
rect -159 1751 -147 1785
rect -113 1751 -101 1785
rect -159 1717 -101 1751
rect -159 1683 -147 1717
rect -113 1683 -101 1717
rect -159 1649 -101 1683
rect -159 1615 -147 1649
rect -113 1615 -101 1649
rect -159 1581 -101 1615
rect -159 1547 -147 1581
rect -113 1547 -101 1581
rect -159 1513 -101 1547
rect -159 1479 -147 1513
rect -113 1479 -101 1513
rect -159 1445 -101 1479
rect -159 1411 -147 1445
rect -113 1411 -101 1445
rect -159 1377 -101 1411
rect -159 1343 -147 1377
rect -113 1343 -101 1377
rect -159 1309 -101 1343
rect -159 1275 -147 1309
rect -113 1275 -101 1309
rect -159 1241 -101 1275
rect -159 1207 -147 1241
rect -113 1207 -101 1241
rect -159 1173 -101 1207
rect -159 1139 -147 1173
rect -113 1139 -101 1173
rect -159 1105 -101 1139
rect -159 1071 -147 1105
rect -113 1071 -101 1105
rect -159 1037 -101 1071
rect -159 1003 -147 1037
rect -113 1003 -101 1037
rect -159 969 -101 1003
rect -159 935 -147 969
rect -113 935 -101 969
rect -159 901 -101 935
rect -159 867 -147 901
rect -113 867 -101 901
rect -159 833 -101 867
rect -159 799 -147 833
rect -113 799 -101 833
rect -159 765 -101 799
rect -159 731 -147 765
rect -113 731 -101 765
rect -159 697 -101 731
rect -159 663 -147 697
rect -113 663 -101 697
rect -159 629 -101 663
rect -159 595 -147 629
rect -113 595 -101 629
rect -159 561 -101 595
rect -159 527 -147 561
rect -113 527 -101 561
rect -159 493 -101 527
rect -159 459 -147 493
rect -113 459 -101 493
rect -159 425 -101 459
rect -159 391 -147 425
rect -113 391 -101 425
rect -159 357 -101 391
rect -159 323 -147 357
rect -113 323 -101 357
rect -159 289 -101 323
rect -159 255 -147 289
rect -113 255 -101 289
rect -159 221 -101 255
rect -159 187 -147 221
rect -113 187 -101 221
rect -159 153 -101 187
rect -159 119 -147 153
rect -113 119 -101 153
rect -159 85 -101 119
rect -159 51 -147 85
rect -113 51 -101 85
rect -159 17 -101 51
rect -159 -17 -147 17
rect -113 -17 -101 17
rect -159 -51 -101 -17
rect -159 -85 -147 -51
rect -113 -85 -101 -51
rect -159 -119 -101 -85
rect -159 -153 -147 -119
rect -113 -153 -101 -119
rect -159 -187 -101 -153
rect -159 -221 -147 -187
rect -113 -221 -101 -187
rect -159 -255 -101 -221
rect -159 -289 -147 -255
rect -113 -289 -101 -255
rect -159 -323 -101 -289
rect -159 -357 -147 -323
rect -113 -357 -101 -323
rect -159 -391 -101 -357
rect -159 -425 -147 -391
rect -113 -425 -101 -391
rect -159 -459 -101 -425
rect -159 -493 -147 -459
rect -113 -493 -101 -459
rect -159 -527 -101 -493
rect -159 -561 -147 -527
rect -113 -561 -101 -527
rect -159 -595 -101 -561
rect -159 -629 -147 -595
rect -113 -629 -101 -595
rect -159 -663 -101 -629
rect -159 -697 -147 -663
rect -113 -697 -101 -663
rect -159 -731 -101 -697
rect -159 -765 -147 -731
rect -113 -765 -101 -731
rect -159 -799 -101 -765
rect -159 -833 -147 -799
rect -113 -833 -101 -799
rect -159 -867 -101 -833
rect -159 -901 -147 -867
rect -113 -901 -101 -867
rect -159 -935 -101 -901
rect -159 -969 -147 -935
rect -113 -969 -101 -935
rect -159 -1003 -101 -969
rect -159 -1037 -147 -1003
rect -113 -1037 -101 -1003
rect -159 -1071 -101 -1037
rect -159 -1105 -147 -1071
rect -113 -1105 -101 -1071
rect -159 -1139 -101 -1105
rect -159 -1173 -147 -1139
rect -113 -1173 -101 -1139
rect -159 -1207 -101 -1173
rect -159 -1241 -147 -1207
rect -113 -1241 -101 -1207
rect -159 -1275 -101 -1241
rect -159 -1309 -147 -1275
rect -113 -1309 -101 -1275
rect -159 -1343 -101 -1309
rect -159 -1377 -147 -1343
rect -113 -1377 -101 -1343
rect -159 -1411 -101 -1377
rect -159 -1445 -147 -1411
rect -113 -1445 -101 -1411
rect -159 -1479 -101 -1445
rect -159 -1513 -147 -1479
rect -113 -1513 -101 -1479
rect -159 -1547 -101 -1513
rect -159 -1581 -147 -1547
rect -113 -1581 -101 -1547
rect -159 -1615 -101 -1581
rect -159 -1649 -147 -1615
rect -113 -1649 -101 -1615
rect -159 -1683 -101 -1649
rect -159 -1717 -147 -1683
rect -113 -1717 -101 -1683
rect -159 -1751 -101 -1717
rect -159 -1785 -147 -1751
rect -113 -1785 -101 -1751
rect -159 -1806 -101 -1785
rect -29 1785 54 1806
rect -29 1751 -5 1785
rect 29 1751 54 1785
rect -29 1717 54 1751
rect -29 1683 -5 1717
rect 29 1683 54 1717
rect -29 1649 54 1683
rect -29 1615 -5 1649
rect 29 1615 54 1649
rect -29 1581 54 1615
rect -29 1547 -5 1581
rect 29 1547 54 1581
rect -29 1513 54 1547
rect -29 1479 -5 1513
rect 29 1479 54 1513
rect -29 1445 54 1479
rect -29 1411 -5 1445
rect 29 1411 54 1445
rect -29 1377 54 1411
rect -29 1343 -5 1377
rect 29 1343 54 1377
rect -29 1309 54 1343
rect -29 1275 -5 1309
rect 29 1275 54 1309
rect -29 1241 54 1275
rect -29 1207 -5 1241
rect 29 1207 54 1241
rect -29 1173 54 1207
rect -29 1139 -5 1173
rect 29 1139 54 1173
rect -29 1105 54 1139
rect -29 1071 -5 1105
rect 29 1071 54 1105
rect -29 1037 54 1071
rect -29 1003 -5 1037
rect 29 1003 54 1037
rect -29 969 54 1003
rect -29 935 -5 969
rect 29 935 54 969
rect -29 901 54 935
rect -29 867 -5 901
rect 29 867 54 901
rect -29 833 54 867
rect -29 799 -5 833
rect 29 799 54 833
rect -29 765 54 799
rect -29 731 -5 765
rect 29 731 54 765
rect -29 697 54 731
rect -29 663 -5 697
rect 29 663 54 697
rect -29 629 54 663
rect -29 595 -5 629
rect 29 595 54 629
rect -29 561 54 595
rect -29 527 -5 561
rect 29 527 54 561
rect -29 493 54 527
rect -29 459 -5 493
rect 29 459 54 493
rect -29 425 54 459
rect -29 391 -5 425
rect 29 391 54 425
rect -29 357 54 391
rect -29 323 -5 357
rect 29 323 54 357
rect -29 289 54 323
rect -29 255 -5 289
rect 29 255 54 289
rect -29 221 54 255
rect -29 187 -5 221
rect 29 187 54 221
rect -29 153 54 187
rect -29 119 -5 153
rect 29 119 54 153
rect -29 85 54 119
rect -29 51 -5 85
rect 29 51 54 85
rect -29 17 54 51
rect -29 -17 -5 17
rect 29 -17 54 17
rect -29 -51 54 -17
rect -29 -85 -5 -51
rect 29 -85 54 -51
rect -29 -119 54 -85
rect -29 -153 -5 -119
rect 29 -153 54 -119
rect -29 -187 54 -153
rect -29 -221 -5 -187
rect 29 -221 54 -187
rect -29 -255 54 -221
rect -29 -289 -5 -255
rect 29 -289 54 -255
rect -29 -323 54 -289
rect -29 -357 -5 -323
rect 29 -357 54 -323
rect -29 -391 54 -357
rect -29 -425 -5 -391
rect 29 -425 54 -391
rect -29 -459 54 -425
rect -29 -493 -5 -459
rect 29 -493 54 -459
rect -29 -527 54 -493
rect -29 -561 -5 -527
rect 29 -561 54 -527
rect -29 -595 54 -561
rect -29 -629 -5 -595
rect 29 -629 54 -595
rect -29 -663 54 -629
rect -29 -697 -5 -663
rect 29 -697 54 -663
rect -29 -731 54 -697
rect -29 -765 -5 -731
rect 29 -765 54 -731
rect -29 -799 54 -765
rect -29 -833 -5 -799
rect 29 -833 54 -799
rect -29 -867 54 -833
rect -29 -901 -5 -867
rect 29 -901 54 -867
rect -29 -935 54 -901
rect -29 -969 -5 -935
rect 29 -969 54 -935
rect -29 -1003 54 -969
rect -29 -1037 -5 -1003
rect 29 -1037 54 -1003
rect -29 -1071 54 -1037
rect -29 -1105 -5 -1071
rect 29 -1105 54 -1071
rect -29 -1139 54 -1105
rect -29 -1173 -5 -1139
rect 29 -1173 54 -1139
rect -29 -1207 54 -1173
rect -29 -1241 -5 -1207
rect 29 -1241 54 -1207
rect -29 -1275 54 -1241
rect -29 -1309 -5 -1275
rect 29 -1309 54 -1275
rect -29 -1343 54 -1309
rect -29 -1377 -5 -1343
rect 29 -1377 54 -1343
rect -29 -1411 54 -1377
rect -29 -1445 -5 -1411
rect 29 -1445 54 -1411
rect -29 -1479 54 -1445
rect -29 -1513 -5 -1479
rect 29 -1513 54 -1479
rect -29 -1547 54 -1513
rect -29 -1581 -5 -1547
rect 29 -1581 54 -1547
rect -29 -1615 54 -1581
rect -29 -1649 -5 -1615
rect 29 -1649 54 -1615
rect -29 -1683 54 -1649
rect -29 -1717 -5 -1683
rect 29 -1717 54 -1683
rect -29 -1751 54 -1717
rect -29 -1785 -5 -1751
rect 29 -1785 54 -1751
rect -29 -1806 54 -1785
rect 126 1785 184 1806
rect 126 1751 138 1785
rect 172 1751 184 1785
rect 126 1717 184 1751
rect 126 1683 138 1717
rect 172 1683 184 1717
rect 126 1649 184 1683
rect 126 1615 138 1649
rect 172 1615 184 1649
rect 126 1581 184 1615
rect 126 1547 138 1581
rect 172 1547 184 1581
rect 126 1513 184 1547
rect 126 1479 138 1513
rect 172 1479 184 1513
rect 126 1445 184 1479
rect 126 1411 138 1445
rect 172 1411 184 1445
rect 126 1377 184 1411
rect 126 1343 138 1377
rect 172 1343 184 1377
rect 126 1309 184 1343
rect 126 1275 138 1309
rect 172 1275 184 1309
rect 126 1241 184 1275
rect 126 1207 138 1241
rect 172 1207 184 1241
rect 126 1173 184 1207
rect 126 1139 138 1173
rect 172 1139 184 1173
rect 126 1105 184 1139
rect 126 1071 138 1105
rect 172 1071 184 1105
rect 126 1037 184 1071
rect 126 1003 138 1037
rect 172 1003 184 1037
rect 126 969 184 1003
rect 126 935 138 969
rect 172 935 184 969
rect 126 901 184 935
rect 126 867 138 901
rect 172 867 184 901
rect 126 833 184 867
rect 126 799 138 833
rect 172 799 184 833
rect 126 765 184 799
rect 126 731 138 765
rect 172 731 184 765
rect 126 697 184 731
rect 126 663 138 697
rect 172 663 184 697
rect 126 629 184 663
rect 126 595 138 629
rect 172 595 184 629
rect 126 561 184 595
rect 126 527 138 561
rect 172 527 184 561
rect 126 493 184 527
rect 126 459 138 493
rect 172 459 184 493
rect 126 425 184 459
rect 126 391 138 425
rect 172 391 184 425
rect 126 357 184 391
rect 126 323 138 357
rect 172 323 184 357
rect 126 289 184 323
rect 126 255 138 289
rect 172 255 184 289
rect 126 221 184 255
rect 126 187 138 221
rect 172 187 184 221
rect 126 153 184 187
rect 126 119 138 153
rect 172 119 184 153
rect 126 85 184 119
rect 126 51 138 85
rect 172 51 184 85
rect 126 17 184 51
rect 126 -17 138 17
rect 172 -17 184 17
rect 126 -51 184 -17
rect 126 -85 138 -51
rect 172 -85 184 -51
rect 126 -119 184 -85
rect 126 -153 138 -119
rect 172 -153 184 -119
rect 126 -187 184 -153
rect 126 -221 138 -187
rect 172 -221 184 -187
rect 126 -255 184 -221
rect 126 -289 138 -255
rect 172 -289 184 -255
rect 126 -323 184 -289
rect 126 -357 138 -323
rect 172 -357 184 -323
rect 126 -391 184 -357
rect 126 -425 138 -391
rect 172 -425 184 -391
rect 126 -459 184 -425
rect 126 -493 138 -459
rect 172 -493 184 -459
rect 126 -527 184 -493
rect 126 -561 138 -527
rect 172 -561 184 -527
rect 126 -595 184 -561
rect 126 -629 138 -595
rect 172 -629 184 -595
rect 126 -663 184 -629
rect 126 -697 138 -663
rect 172 -697 184 -663
rect 126 -731 184 -697
rect 126 -765 138 -731
rect 172 -765 184 -731
rect 126 -799 184 -765
rect 126 -833 138 -799
rect 172 -833 184 -799
rect 126 -867 184 -833
rect 126 -901 138 -867
rect 172 -901 184 -867
rect 126 -935 184 -901
rect 126 -969 138 -935
rect 172 -969 184 -935
rect 126 -1003 184 -969
rect 126 -1037 138 -1003
rect 172 -1037 184 -1003
rect 126 -1071 184 -1037
rect 126 -1105 138 -1071
rect 172 -1105 184 -1071
rect 126 -1139 184 -1105
rect 126 -1173 138 -1139
rect 172 -1173 184 -1139
rect 126 -1207 184 -1173
rect 126 -1241 138 -1207
rect 172 -1241 184 -1207
rect 126 -1275 184 -1241
rect 126 -1309 138 -1275
rect 172 -1309 184 -1275
rect 126 -1343 184 -1309
rect 126 -1377 138 -1343
rect 172 -1377 184 -1343
rect 126 -1411 184 -1377
rect 126 -1445 138 -1411
rect 172 -1445 184 -1411
rect 126 -1479 184 -1445
rect 126 -1513 138 -1479
rect 172 -1513 184 -1479
rect 126 -1547 184 -1513
rect 126 -1581 138 -1547
rect 172 -1581 184 -1547
rect 126 -1615 184 -1581
rect 126 -1649 138 -1615
rect 172 -1649 184 -1615
rect 126 -1683 184 -1649
rect 126 -1717 138 -1683
rect 172 -1717 184 -1683
rect 126 -1751 184 -1717
rect 126 -1785 138 -1751
rect 172 -1785 184 -1751
rect 126 -1806 184 -1785
<< ndiffc >>
rect -147 1751 -113 1785
rect -147 1683 -113 1717
rect -147 1615 -113 1649
rect -147 1547 -113 1581
rect -147 1479 -113 1513
rect -147 1411 -113 1445
rect -147 1343 -113 1377
rect -147 1275 -113 1309
rect -147 1207 -113 1241
rect -147 1139 -113 1173
rect -147 1071 -113 1105
rect -147 1003 -113 1037
rect -147 935 -113 969
rect -147 867 -113 901
rect -147 799 -113 833
rect -147 731 -113 765
rect -147 663 -113 697
rect -147 595 -113 629
rect -147 527 -113 561
rect -147 459 -113 493
rect -147 391 -113 425
rect -147 323 -113 357
rect -147 255 -113 289
rect -147 187 -113 221
rect -147 119 -113 153
rect -147 51 -113 85
rect -147 -17 -113 17
rect -147 -85 -113 -51
rect -147 -153 -113 -119
rect -147 -221 -113 -187
rect -147 -289 -113 -255
rect -147 -357 -113 -323
rect -147 -425 -113 -391
rect -147 -493 -113 -459
rect -147 -561 -113 -527
rect -147 -629 -113 -595
rect -147 -697 -113 -663
rect -147 -765 -113 -731
rect -147 -833 -113 -799
rect -147 -901 -113 -867
rect -147 -969 -113 -935
rect -147 -1037 -113 -1003
rect -147 -1105 -113 -1071
rect -147 -1173 -113 -1139
rect -147 -1241 -113 -1207
rect -147 -1309 -113 -1275
rect -147 -1377 -113 -1343
rect -147 -1445 -113 -1411
rect -147 -1513 -113 -1479
rect -147 -1581 -113 -1547
rect -147 -1649 -113 -1615
rect -147 -1717 -113 -1683
rect -147 -1785 -113 -1751
rect -5 1751 29 1785
rect -5 1683 29 1717
rect -5 1615 29 1649
rect -5 1547 29 1581
rect -5 1479 29 1513
rect -5 1411 29 1445
rect -5 1343 29 1377
rect -5 1275 29 1309
rect -5 1207 29 1241
rect -5 1139 29 1173
rect -5 1071 29 1105
rect -5 1003 29 1037
rect -5 935 29 969
rect -5 867 29 901
rect -5 799 29 833
rect -5 731 29 765
rect -5 663 29 697
rect -5 595 29 629
rect -5 527 29 561
rect -5 459 29 493
rect -5 391 29 425
rect -5 323 29 357
rect -5 255 29 289
rect -5 187 29 221
rect -5 119 29 153
rect -5 51 29 85
rect -5 -17 29 17
rect -5 -85 29 -51
rect -5 -153 29 -119
rect -5 -221 29 -187
rect -5 -289 29 -255
rect -5 -357 29 -323
rect -5 -425 29 -391
rect -5 -493 29 -459
rect -5 -561 29 -527
rect -5 -629 29 -595
rect -5 -697 29 -663
rect -5 -765 29 -731
rect -5 -833 29 -799
rect -5 -901 29 -867
rect -5 -969 29 -935
rect -5 -1037 29 -1003
rect -5 -1105 29 -1071
rect -5 -1173 29 -1139
rect -5 -1241 29 -1207
rect -5 -1309 29 -1275
rect -5 -1377 29 -1343
rect -5 -1445 29 -1411
rect -5 -1513 29 -1479
rect -5 -1581 29 -1547
rect -5 -1649 29 -1615
rect -5 -1717 29 -1683
rect -5 -1785 29 -1751
rect 138 1751 172 1785
rect 138 1683 172 1717
rect 138 1615 172 1649
rect 138 1547 172 1581
rect 138 1479 172 1513
rect 138 1411 172 1445
rect 138 1343 172 1377
rect 138 1275 172 1309
rect 138 1207 172 1241
rect 138 1139 172 1173
rect 138 1071 172 1105
rect 138 1003 172 1037
rect 138 935 172 969
rect 138 867 172 901
rect 138 799 172 833
rect 138 731 172 765
rect 138 663 172 697
rect 138 595 172 629
rect 138 527 172 561
rect 138 459 172 493
rect 138 391 172 425
rect 138 323 172 357
rect 138 255 172 289
rect 138 187 172 221
rect 138 119 172 153
rect 138 51 172 85
rect 138 -17 172 17
rect 138 -85 172 -51
rect 138 -153 172 -119
rect 138 -221 172 -187
rect 138 -289 172 -255
rect 138 -357 172 -323
rect 138 -425 172 -391
rect 138 -493 172 -459
rect 138 -561 172 -527
rect 138 -629 172 -595
rect 138 -697 172 -663
rect 138 -765 172 -731
rect 138 -833 172 -799
rect 138 -901 172 -867
rect 138 -969 172 -935
rect 138 -1037 172 -1003
rect 138 -1105 172 -1071
rect 138 -1173 172 -1139
rect 138 -1241 172 -1207
rect 138 -1309 172 -1275
rect 138 -1377 172 -1343
rect 138 -1445 172 -1411
rect 138 -1513 172 -1479
rect 138 -1581 172 -1547
rect 138 -1649 172 -1615
rect 138 -1717 172 -1683
rect 138 -1785 172 -1751
<< poly >>
rect -101 1838 126 1894
rect -101 1806 -29 1838
rect 54 1806 126 1838
rect -101 -1832 -29 -1806
rect 54 -1844 126 -1806
rect 54 -1878 73 -1844
rect 107 -1878 126 -1844
rect 54 -1894 126 -1878
<< polycont >>
rect 73 -1878 107 -1844
<< locali >>
rect -147 1785 -113 1810
rect -147 1717 -113 1747
rect -147 1649 -113 1675
rect -147 1581 -113 1603
rect -147 1513 -113 1531
rect -147 1445 -113 1459
rect -147 1377 -113 1387
rect -147 1309 -113 1315
rect -147 1241 -113 1243
rect -147 1205 -113 1207
rect -147 1133 -113 1139
rect -147 1061 -113 1071
rect -147 989 -113 1003
rect -147 917 -113 935
rect -147 845 -113 867
rect -147 773 -113 799
rect -147 701 -113 731
rect -147 629 -113 663
rect -147 561 -113 595
rect -147 493 -113 523
rect -147 425 -113 451
rect -147 357 -113 379
rect -147 289 -113 307
rect -147 221 -113 235
rect -147 153 -113 163
rect -147 85 -113 91
rect -147 17 -113 19
rect -147 -19 -113 -17
rect -147 -91 -113 -85
rect -147 -163 -113 -153
rect -147 -235 -113 -221
rect -147 -307 -113 -289
rect -147 -379 -113 -357
rect -147 -451 -113 -425
rect -147 -523 -113 -493
rect -147 -595 -113 -561
rect -147 -663 -113 -629
rect -147 -731 -113 -701
rect -147 -799 -113 -773
rect -147 -867 -113 -845
rect -147 -935 -113 -917
rect -147 -1003 -113 -989
rect -147 -1071 -113 -1061
rect -147 -1139 -113 -1133
rect -147 -1207 -113 -1205
rect -147 -1243 -113 -1241
rect -147 -1315 -113 -1309
rect -147 -1387 -113 -1377
rect -147 -1459 -113 -1445
rect -147 -1531 -113 -1513
rect -147 -1603 -113 -1581
rect -147 -1675 -113 -1649
rect -147 -1747 -113 -1717
rect -147 -1810 -113 -1785
rect -17 1785 42 1810
rect -17 1747 -5 1785
rect 29 1747 42 1785
rect -17 1717 42 1747
rect -17 1675 -5 1717
rect 29 1675 42 1717
rect -17 1649 42 1675
rect -17 1603 -5 1649
rect 29 1603 42 1649
rect -17 1581 42 1603
rect -17 1531 -5 1581
rect 29 1531 42 1581
rect -17 1513 42 1531
rect -17 1459 -5 1513
rect 29 1459 42 1513
rect -17 1445 42 1459
rect -17 1387 -5 1445
rect 29 1387 42 1445
rect -17 1377 42 1387
rect -17 1315 -5 1377
rect 29 1315 42 1377
rect -17 1309 42 1315
rect -17 1243 -5 1309
rect 29 1243 42 1309
rect -17 1241 42 1243
rect -17 1207 -5 1241
rect 29 1207 42 1241
rect -17 1205 42 1207
rect -17 1139 -5 1205
rect 29 1139 42 1205
rect -17 1133 42 1139
rect -17 1071 -5 1133
rect 29 1071 42 1133
rect -17 1061 42 1071
rect -17 1003 -5 1061
rect 29 1003 42 1061
rect -17 989 42 1003
rect -17 935 -5 989
rect 29 935 42 989
rect -17 917 42 935
rect -17 867 -5 917
rect 29 867 42 917
rect -17 845 42 867
rect -17 799 -5 845
rect 29 799 42 845
rect -17 773 42 799
rect -17 731 -5 773
rect 29 731 42 773
rect -17 701 42 731
rect -17 663 -5 701
rect 29 663 42 701
rect -17 629 42 663
rect -17 595 -5 629
rect 29 595 42 629
rect -17 561 42 595
rect -17 523 -5 561
rect 29 523 42 561
rect -17 493 42 523
rect -17 451 -5 493
rect 29 451 42 493
rect -17 425 42 451
rect -17 379 -5 425
rect 29 379 42 425
rect -17 357 42 379
rect -17 307 -5 357
rect 29 307 42 357
rect -17 289 42 307
rect -17 235 -5 289
rect 29 235 42 289
rect -17 221 42 235
rect -17 163 -5 221
rect 29 163 42 221
rect -17 153 42 163
rect -17 91 -5 153
rect 29 91 42 153
rect -17 85 42 91
rect -17 19 -5 85
rect 29 19 42 85
rect -17 17 42 19
rect -17 -17 -5 17
rect 29 -17 42 17
rect -17 -19 42 -17
rect -17 -85 -5 -19
rect 29 -85 42 -19
rect -17 -91 42 -85
rect -17 -153 -5 -91
rect 29 -153 42 -91
rect -17 -163 42 -153
rect -17 -221 -5 -163
rect 29 -221 42 -163
rect -17 -235 42 -221
rect -17 -289 -5 -235
rect 29 -289 42 -235
rect -17 -307 42 -289
rect -17 -357 -5 -307
rect 29 -357 42 -307
rect -17 -379 42 -357
rect -17 -425 -5 -379
rect 29 -425 42 -379
rect -17 -451 42 -425
rect -17 -493 -5 -451
rect 29 -493 42 -451
rect -17 -523 42 -493
rect -17 -561 -5 -523
rect 29 -561 42 -523
rect -17 -595 42 -561
rect -17 -629 -5 -595
rect 29 -629 42 -595
rect -17 -663 42 -629
rect -17 -701 -5 -663
rect 29 -701 42 -663
rect -17 -731 42 -701
rect -17 -773 -5 -731
rect 29 -773 42 -731
rect -17 -799 42 -773
rect -17 -845 -5 -799
rect 29 -845 42 -799
rect -17 -867 42 -845
rect -17 -917 -5 -867
rect 29 -917 42 -867
rect -17 -935 42 -917
rect -17 -989 -5 -935
rect 29 -989 42 -935
rect -17 -1003 42 -989
rect -17 -1061 -5 -1003
rect 29 -1061 42 -1003
rect -17 -1071 42 -1061
rect -17 -1133 -5 -1071
rect 29 -1133 42 -1071
rect -17 -1139 42 -1133
rect -17 -1205 -5 -1139
rect 29 -1205 42 -1139
rect -17 -1207 42 -1205
rect -17 -1241 -5 -1207
rect 29 -1241 42 -1207
rect -17 -1243 42 -1241
rect -17 -1309 -5 -1243
rect 29 -1309 42 -1243
rect -17 -1315 42 -1309
rect -17 -1377 -5 -1315
rect 29 -1377 42 -1315
rect -17 -1387 42 -1377
rect -17 -1445 -5 -1387
rect 29 -1445 42 -1387
rect -17 -1459 42 -1445
rect -17 -1513 -5 -1459
rect 29 -1513 42 -1459
rect -17 -1531 42 -1513
rect -17 -1581 -5 -1531
rect 29 -1581 42 -1531
rect -17 -1603 42 -1581
rect -17 -1649 -5 -1603
rect 29 -1649 42 -1603
rect -17 -1675 42 -1649
rect -17 -1717 -5 -1675
rect 29 -1717 42 -1675
rect -17 -1747 42 -1717
rect -17 -1785 -5 -1747
rect 29 -1785 42 -1747
rect -17 -1810 42 -1785
rect 138 1785 172 1810
rect 138 1717 172 1747
rect 138 1649 172 1675
rect 138 1581 172 1603
rect 138 1513 172 1531
rect 138 1445 172 1459
rect 138 1377 172 1387
rect 138 1309 172 1315
rect 138 1241 172 1243
rect 138 1205 172 1207
rect 138 1133 172 1139
rect 138 1061 172 1071
rect 138 989 172 1003
rect 138 917 172 935
rect 138 845 172 867
rect 138 773 172 799
rect 138 701 172 731
rect 138 629 172 663
rect 138 561 172 595
rect 138 493 172 523
rect 138 425 172 451
rect 138 357 172 379
rect 138 289 172 307
rect 138 221 172 235
rect 138 153 172 163
rect 138 85 172 91
rect 138 17 172 19
rect 138 -19 172 -17
rect 138 -91 172 -85
rect 138 -163 172 -153
rect 138 -235 172 -221
rect 138 -307 172 -289
rect 138 -379 172 -357
rect 138 -451 172 -425
rect 138 -523 172 -493
rect 138 -595 172 -561
rect 138 -663 172 -629
rect 138 -731 172 -701
rect 138 -799 172 -773
rect 138 -867 172 -845
rect 138 -935 172 -917
rect 138 -1003 172 -989
rect 138 -1071 172 -1061
rect 138 -1139 172 -1133
rect 138 -1207 172 -1205
rect 138 -1243 172 -1241
rect 138 -1315 172 -1309
rect 138 -1387 172 -1377
rect 138 -1459 172 -1445
rect 138 -1531 172 -1513
rect 138 -1603 172 -1581
rect 138 -1675 172 -1649
rect 138 -1747 172 -1717
rect 138 -1810 172 -1785
rect 54 -1878 73 -1844
rect 107 -1878 126 -1844
<< viali >>
rect -147 1751 -113 1781
rect -147 1747 -113 1751
rect -147 1683 -113 1709
rect -147 1675 -113 1683
rect -147 1615 -113 1637
rect -147 1603 -113 1615
rect -147 1547 -113 1565
rect -147 1531 -113 1547
rect -147 1479 -113 1493
rect -147 1459 -113 1479
rect -147 1411 -113 1421
rect -147 1387 -113 1411
rect -147 1343 -113 1349
rect -147 1315 -113 1343
rect -147 1275 -113 1277
rect -147 1243 -113 1275
rect -147 1173 -113 1205
rect -147 1171 -113 1173
rect -147 1105 -113 1133
rect -147 1099 -113 1105
rect -147 1037 -113 1061
rect -147 1027 -113 1037
rect -147 969 -113 989
rect -147 955 -113 969
rect -147 901 -113 917
rect -147 883 -113 901
rect -147 833 -113 845
rect -147 811 -113 833
rect -147 765 -113 773
rect -147 739 -113 765
rect -147 697 -113 701
rect -147 667 -113 697
rect -147 595 -113 629
rect -147 527 -113 557
rect -147 523 -113 527
rect -147 459 -113 485
rect -147 451 -113 459
rect -147 391 -113 413
rect -147 379 -113 391
rect -147 323 -113 341
rect -147 307 -113 323
rect -147 255 -113 269
rect -147 235 -113 255
rect -147 187 -113 197
rect -147 163 -113 187
rect -147 119 -113 125
rect -147 91 -113 119
rect -147 51 -113 53
rect -147 19 -113 51
rect -147 -51 -113 -19
rect -147 -53 -113 -51
rect -147 -119 -113 -91
rect -147 -125 -113 -119
rect -147 -187 -113 -163
rect -147 -197 -113 -187
rect -147 -255 -113 -235
rect -147 -269 -113 -255
rect -147 -323 -113 -307
rect -147 -341 -113 -323
rect -147 -391 -113 -379
rect -147 -413 -113 -391
rect -147 -459 -113 -451
rect -147 -485 -113 -459
rect -147 -527 -113 -523
rect -147 -557 -113 -527
rect -147 -629 -113 -595
rect -147 -697 -113 -667
rect -147 -701 -113 -697
rect -147 -765 -113 -739
rect -147 -773 -113 -765
rect -147 -833 -113 -811
rect -147 -845 -113 -833
rect -147 -901 -113 -883
rect -147 -917 -113 -901
rect -147 -969 -113 -955
rect -147 -989 -113 -969
rect -147 -1037 -113 -1027
rect -147 -1061 -113 -1037
rect -147 -1105 -113 -1099
rect -147 -1133 -113 -1105
rect -147 -1173 -113 -1171
rect -147 -1205 -113 -1173
rect -147 -1275 -113 -1243
rect -147 -1277 -113 -1275
rect -147 -1343 -113 -1315
rect -147 -1349 -113 -1343
rect -147 -1411 -113 -1387
rect -147 -1421 -113 -1411
rect -147 -1479 -113 -1459
rect -147 -1493 -113 -1479
rect -147 -1547 -113 -1531
rect -147 -1565 -113 -1547
rect -147 -1615 -113 -1603
rect -147 -1637 -113 -1615
rect -147 -1683 -113 -1675
rect -147 -1709 -113 -1683
rect -147 -1751 -113 -1747
rect -147 -1781 -113 -1751
rect -5 1751 29 1781
rect -5 1747 29 1751
rect -5 1683 29 1709
rect -5 1675 29 1683
rect -5 1615 29 1637
rect -5 1603 29 1615
rect -5 1547 29 1565
rect -5 1531 29 1547
rect -5 1479 29 1493
rect -5 1459 29 1479
rect -5 1411 29 1421
rect -5 1387 29 1411
rect -5 1343 29 1349
rect -5 1315 29 1343
rect -5 1275 29 1277
rect -5 1243 29 1275
rect -5 1173 29 1205
rect -5 1171 29 1173
rect -5 1105 29 1133
rect -5 1099 29 1105
rect -5 1037 29 1061
rect -5 1027 29 1037
rect -5 969 29 989
rect -5 955 29 969
rect -5 901 29 917
rect -5 883 29 901
rect -5 833 29 845
rect -5 811 29 833
rect -5 765 29 773
rect -5 739 29 765
rect -5 697 29 701
rect -5 667 29 697
rect -5 595 29 629
rect -5 527 29 557
rect -5 523 29 527
rect -5 459 29 485
rect -5 451 29 459
rect -5 391 29 413
rect -5 379 29 391
rect -5 323 29 341
rect -5 307 29 323
rect -5 255 29 269
rect -5 235 29 255
rect -5 187 29 197
rect -5 163 29 187
rect -5 119 29 125
rect -5 91 29 119
rect -5 51 29 53
rect -5 19 29 51
rect -5 -51 29 -19
rect -5 -53 29 -51
rect -5 -119 29 -91
rect -5 -125 29 -119
rect -5 -187 29 -163
rect -5 -197 29 -187
rect -5 -255 29 -235
rect -5 -269 29 -255
rect -5 -323 29 -307
rect -5 -341 29 -323
rect -5 -391 29 -379
rect -5 -413 29 -391
rect -5 -459 29 -451
rect -5 -485 29 -459
rect -5 -527 29 -523
rect -5 -557 29 -527
rect -5 -629 29 -595
rect -5 -697 29 -667
rect -5 -701 29 -697
rect -5 -765 29 -739
rect -5 -773 29 -765
rect -5 -833 29 -811
rect -5 -845 29 -833
rect -5 -901 29 -883
rect -5 -917 29 -901
rect -5 -969 29 -955
rect -5 -989 29 -969
rect -5 -1037 29 -1027
rect -5 -1061 29 -1037
rect -5 -1105 29 -1099
rect -5 -1133 29 -1105
rect -5 -1173 29 -1171
rect -5 -1205 29 -1173
rect -5 -1275 29 -1243
rect -5 -1277 29 -1275
rect -5 -1343 29 -1315
rect -5 -1349 29 -1343
rect -5 -1411 29 -1387
rect -5 -1421 29 -1411
rect -5 -1479 29 -1459
rect -5 -1493 29 -1479
rect -5 -1547 29 -1531
rect -5 -1565 29 -1547
rect -5 -1615 29 -1603
rect -5 -1637 29 -1615
rect -5 -1683 29 -1675
rect -5 -1709 29 -1683
rect -5 -1751 29 -1747
rect -5 -1781 29 -1751
rect 138 1751 172 1781
rect 138 1747 172 1751
rect 138 1683 172 1709
rect 138 1675 172 1683
rect 138 1615 172 1637
rect 138 1603 172 1615
rect 138 1547 172 1565
rect 138 1531 172 1547
rect 138 1479 172 1493
rect 138 1459 172 1479
rect 138 1411 172 1421
rect 138 1387 172 1411
rect 138 1343 172 1349
rect 138 1315 172 1343
rect 138 1275 172 1277
rect 138 1243 172 1275
rect 138 1173 172 1205
rect 138 1171 172 1173
rect 138 1105 172 1133
rect 138 1099 172 1105
rect 138 1037 172 1061
rect 138 1027 172 1037
rect 138 969 172 989
rect 138 955 172 969
rect 138 901 172 917
rect 138 883 172 901
rect 138 833 172 845
rect 138 811 172 833
rect 138 765 172 773
rect 138 739 172 765
rect 138 697 172 701
rect 138 667 172 697
rect 138 595 172 629
rect 138 527 172 557
rect 138 523 172 527
rect 138 459 172 485
rect 138 451 172 459
rect 138 391 172 413
rect 138 379 172 391
rect 138 323 172 341
rect 138 307 172 323
rect 138 255 172 269
rect 138 235 172 255
rect 138 187 172 197
rect 138 163 172 187
rect 138 119 172 125
rect 138 91 172 119
rect 138 51 172 53
rect 138 19 172 51
rect 138 -51 172 -19
rect 138 -53 172 -51
rect 138 -119 172 -91
rect 138 -125 172 -119
rect 138 -187 172 -163
rect 138 -197 172 -187
rect 138 -255 172 -235
rect 138 -269 172 -255
rect 138 -323 172 -307
rect 138 -341 172 -323
rect 138 -391 172 -379
rect 138 -413 172 -391
rect 138 -459 172 -451
rect 138 -485 172 -459
rect 138 -527 172 -523
rect 138 -557 172 -527
rect 138 -629 172 -595
rect 138 -697 172 -667
rect 138 -701 172 -697
rect 138 -765 172 -739
rect 138 -773 172 -765
rect 138 -833 172 -811
rect 138 -845 172 -833
rect 138 -901 172 -883
rect 138 -917 172 -901
rect 138 -969 172 -955
rect 138 -989 172 -969
rect 138 -1037 172 -1027
rect 138 -1061 172 -1037
rect 138 -1105 172 -1099
rect 138 -1133 172 -1105
rect 138 -1173 172 -1171
rect 138 -1205 172 -1173
rect 138 -1275 172 -1243
rect 138 -1277 172 -1275
rect 138 -1343 172 -1315
rect 138 -1349 172 -1343
rect 138 -1411 172 -1387
rect 138 -1421 172 -1411
rect 138 -1479 172 -1459
rect 138 -1493 172 -1479
rect 138 -1547 172 -1531
rect 138 -1565 172 -1547
rect 138 -1615 172 -1603
rect 138 -1637 172 -1615
rect 138 -1683 172 -1675
rect 138 -1709 172 -1683
rect 138 -1751 172 -1747
rect 138 -1781 172 -1751
rect 73 -1878 107 -1844
<< metal1 >>
rect -153 1781 -107 1806
rect -153 1747 -147 1781
rect -113 1747 -107 1781
rect -153 1709 -107 1747
rect -153 1675 -147 1709
rect -113 1675 -107 1709
rect -153 1637 -107 1675
rect -153 1603 -147 1637
rect -113 1603 -107 1637
rect -153 1565 -107 1603
rect -153 1531 -147 1565
rect -113 1531 -107 1565
rect -153 1493 -107 1531
rect -153 1459 -147 1493
rect -113 1459 -107 1493
rect -153 1421 -107 1459
rect -153 1387 -147 1421
rect -113 1387 -107 1421
rect -153 1349 -107 1387
rect -153 1315 -147 1349
rect -113 1315 -107 1349
rect -153 1277 -107 1315
rect -153 1243 -147 1277
rect -113 1243 -107 1277
rect -153 1205 -107 1243
rect -153 1171 -147 1205
rect -113 1171 -107 1205
rect -153 1133 -107 1171
rect -153 1099 -147 1133
rect -113 1099 -107 1133
rect -153 1061 -107 1099
rect -153 1027 -147 1061
rect -113 1027 -107 1061
rect -153 989 -107 1027
rect -153 955 -147 989
rect -113 955 -107 989
rect -153 917 -107 955
rect -153 883 -147 917
rect -113 883 -107 917
rect -153 845 -107 883
rect -153 811 -147 845
rect -113 811 -107 845
rect -153 773 -107 811
rect -153 739 -147 773
rect -113 739 -107 773
rect -153 701 -107 739
rect -153 667 -147 701
rect -113 667 -107 701
rect -153 629 -107 667
rect -153 595 -147 629
rect -113 595 -107 629
rect -153 557 -107 595
rect -153 523 -147 557
rect -113 523 -107 557
rect -153 485 -107 523
rect -153 451 -147 485
rect -113 451 -107 485
rect -153 413 -107 451
rect -153 379 -147 413
rect -113 379 -107 413
rect -153 341 -107 379
rect -153 307 -147 341
rect -113 307 -107 341
rect -153 269 -107 307
rect -153 235 -147 269
rect -113 235 -107 269
rect -153 197 -107 235
rect -153 163 -147 197
rect -113 163 -107 197
rect -153 125 -107 163
rect -153 91 -147 125
rect -113 91 -107 125
rect -153 53 -107 91
rect -153 19 -147 53
rect -113 19 -107 53
rect -153 -19 -107 19
rect -153 -53 -147 -19
rect -113 -53 -107 -19
rect -153 -91 -107 -53
rect -153 -125 -147 -91
rect -113 -125 -107 -91
rect -153 -163 -107 -125
rect -153 -197 -147 -163
rect -113 -197 -107 -163
rect -153 -235 -107 -197
rect -153 -269 -147 -235
rect -113 -269 -107 -235
rect -153 -307 -107 -269
rect -153 -341 -147 -307
rect -113 -341 -107 -307
rect -153 -379 -107 -341
rect -153 -413 -147 -379
rect -113 -413 -107 -379
rect -153 -451 -107 -413
rect -153 -485 -147 -451
rect -113 -485 -107 -451
rect -153 -523 -107 -485
rect -153 -557 -147 -523
rect -113 -557 -107 -523
rect -153 -595 -107 -557
rect -153 -629 -147 -595
rect -113 -629 -107 -595
rect -153 -667 -107 -629
rect -153 -701 -147 -667
rect -113 -701 -107 -667
rect -153 -739 -107 -701
rect -153 -773 -147 -739
rect -113 -773 -107 -739
rect -153 -811 -107 -773
rect -153 -845 -147 -811
rect -113 -845 -107 -811
rect -153 -883 -107 -845
rect -153 -917 -147 -883
rect -113 -917 -107 -883
rect -153 -955 -107 -917
rect -153 -989 -147 -955
rect -113 -989 -107 -955
rect -153 -1027 -107 -989
rect -153 -1061 -147 -1027
rect -113 -1061 -107 -1027
rect -153 -1099 -107 -1061
rect -153 -1133 -147 -1099
rect -113 -1133 -107 -1099
rect -153 -1171 -107 -1133
rect -153 -1205 -147 -1171
rect -113 -1205 -107 -1171
rect -153 -1243 -107 -1205
rect -153 -1277 -147 -1243
rect -113 -1277 -107 -1243
rect -153 -1315 -107 -1277
rect -153 -1349 -147 -1315
rect -113 -1349 -107 -1315
rect -153 -1387 -107 -1349
rect -153 -1421 -147 -1387
rect -113 -1421 -107 -1387
rect -153 -1459 -107 -1421
rect -153 -1493 -147 -1459
rect -113 -1493 -107 -1459
rect -153 -1531 -107 -1493
rect -153 -1565 -147 -1531
rect -113 -1565 -107 -1531
rect -153 -1603 -107 -1565
rect -153 -1637 -147 -1603
rect -113 -1637 -107 -1603
rect -153 -1675 -107 -1637
rect -153 -1709 -147 -1675
rect -113 -1709 -107 -1675
rect -153 -1747 -107 -1709
rect -153 -1781 -147 -1747
rect -113 -1781 -107 -1747
rect -153 -1806 -107 -1781
rect -23 1781 48 1806
rect -23 1747 -5 1781
rect 29 1747 48 1781
rect -23 1709 48 1747
rect -23 1675 -5 1709
rect 29 1675 48 1709
rect -23 1637 48 1675
rect -23 1603 -5 1637
rect 29 1603 48 1637
rect -23 1565 48 1603
rect -23 1531 -5 1565
rect 29 1531 48 1565
rect -23 1493 48 1531
rect -23 1459 -5 1493
rect 29 1459 48 1493
rect -23 1421 48 1459
rect -23 1387 -5 1421
rect 29 1387 48 1421
rect -23 1349 48 1387
rect -23 1315 -5 1349
rect 29 1315 48 1349
rect -23 1277 48 1315
rect -23 1243 -5 1277
rect 29 1243 48 1277
rect -23 1205 48 1243
rect -23 1171 -5 1205
rect 29 1171 48 1205
rect -23 1133 48 1171
rect -23 1099 -5 1133
rect 29 1099 48 1133
rect -23 1061 48 1099
rect -23 1027 -5 1061
rect 29 1027 48 1061
rect -23 989 48 1027
rect -23 955 -5 989
rect 29 955 48 989
rect -23 917 48 955
rect -23 883 -5 917
rect 29 883 48 917
rect -23 845 48 883
rect -23 811 -5 845
rect 29 811 48 845
rect -23 773 48 811
rect -23 739 -5 773
rect 29 739 48 773
rect -23 701 48 739
rect -23 667 -5 701
rect 29 667 48 701
rect -23 629 48 667
rect -23 595 -5 629
rect 29 595 48 629
rect -23 557 48 595
rect -23 523 -5 557
rect 29 523 48 557
rect -23 485 48 523
rect -23 451 -5 485
rect 29 451 48 485
rect -23 413 48 451
rect -23 379 -5 413
rect 29 379 48 413
rect -23 341 48 379
rect -23 307 -5 341
rect 29 307 48 341
rect -23 269 48 307
rect -23 235 -5 269
rect 29 235 48 269
rect -23 197 48 235
rect -23 163 -5 197
rect 29 163 48 197
rect -23 125 48 163
rect -23 91 -5 125
rect 29 91 48 125
rect -23 53 48 91
rect -23 19 -5 53
rect 29 19 48 53
rect -23 -19 48 19
rect -23 -53 -5 -19
rect 29 -53 48 -19
rect -23 -91 48 -53
rect -23 -125 -5 -91
rect 29 -125 48 -91
rect -23 -163 48 -125
rect -23 -197 -5 -163
rect 29 -197 48 -163
rect -23 -235 48 -197
rect -23 -269 -5 -235
rect 29 -269 48 -235
rect -23 -307 48 -269
rect -23 -341 -5 -307
rect 29 -341 48 -307
rect -23 -379 48 -341
rect -23 -413 -5 -379
rect 29 -413 48 -379
rect -23 -451 48 -413
rect -23 -485 -5 -451
rect 29 -485 48 -451
rect -23 -523 48 -485
rect -23 -557 -5 -523
rect 29 -557 48 -523
rect -23 -595 48 -557
rect -23 -629 -5 -595
rect 29 -629 48 -595
rect -23 -667 48 -629
rect -23 -701 -5 -667
rect 29 -701 48 -667
rect -23 -739 48 -701
rect -23 -773 -5 -739
rect 29 -773 48 -739
rect -23 -811 48 -773
rect -23 -845 -5 -811
rect 29 -845 48 -811
rect -23 -883 48 -845
rect -23 -917 -5 -883
rect 29 -917 48 -883
rect -23 -955 48 -917
rect -23 -989 -5 -955
rect 29 -989 48 -955
rect -23 -1027 48 -989
rect -23 -1061 -5 -1027
rect 29 -1061 48 -1027
rect -23 -1099 48 -1061
rect -23 -1133 -5 -1099
rect 29 -1133 48 -1099
rect -23 -1171 48 -1133
rect -23 -1205 -5 -1171
rect 29 -1205 48 -1171
rect -23 -1243 48 -1205
rect -23 -1277 -5 -1243
rect 29 -1277 48 -1243
rect -23 -1315 48 -1277
rect -23 -1349 -5 -1315
rect 29 -1349 48 -1315
rect -23 -1387 48 -1349
rect -23 -1421 -5 -1387
rect 29 -1421 48 -1387
rect -23 -1459 48 -1421
rect -23 -1493 -5 -1459
rect 29 -1493 48 -1459
rect -23 -1531 48 -1493
rect -23 -1565 -5 -1531
rect 29 -1565 48 -1531
rect -23 -1603 48 -1565
rect -23 -1637 -5 -1603
rect 29 -1637 48 -1603
rect -23 -1675 48 -1637
rect -23 -1709 -5 -1675
rect 29 -1709 48 -1675
rect -23 -1747 48 -1709
rect -23 -1781 -5 -1747
rect 29 -1781 48 -1747
rect -23 -1806 48 -1781
rect 132 1781 178 1806
rect 132 1747 138 1781
rect 172 1747 178 1781
rect 132 1709 178 1747
rect 132 1675 138 1709
rect 172 1675 178 1709
rect 132 1637 178 1675
rect 132 1603 138 1637
rect 172 1603 178 1637
rect 132 1565 178 1603
rect 132 1531 138 1565
rect 172 1531 178 1565
rect 132 1493 178 1531
rect 132 1459 138 1493
rect 172 1459 178 1493
rect 132 1421 178 1459
rect 132 1387 138 1421
rect 172 1387 178 1421
rect 132 1349 178 1387
rect 132 1315 138 1349
rect 172 1315 178 1349
rect 132 1277 178 1315
rect 132 1243 138 1277
rect 172 1243 178 1277
rect 132 1205 178 1243
rect 132 1171 138 1205
rect 172 1171 178 1205
rect 132 1133 178 1171
rect 132 1099 138 1133
rect 172 1099 178 1133
rect 132 1061 178 1099
rect 132 1027 138 1061
rect 172 1027 178 1061
rect 132 989 178 1027
rect 132 955 138 989
rect 172 955 178 989
rect 132 917 178 955
rect 132 883 138 917
rect 172 883 178 917
rect 132 845 178 883
rect 132 811 138 845
rect 172 811 178 845
rect 132 773 178 811
rect 132 739 138 773
rect 172 739 178 773
rect 132 701 178 739
rect 132 667 138 701
rect 172 667 178 701
rect 132 629 178 667
rect 132 595 138 629
rect 172 595 178 629
rect 132 557 178 595
rect 132 523 138 557
rect 172 523 178 557
rect 132 485 178 523
rect 132 451 138 485
rect 172 451 178 485
rect 132 413 178 451
rect 132 379 138 413
rect 172 379 178 413
rect 132 341 178 379
rect 132 307 138 341
rect 172 307 178 341
rect 132 269 178 307
rect 132 235 138 269
rect 172 235 178 269
rect 132 197 178 235
rect 132 163 138 197
rect 172 163 178 197
rect 132 125 178 163
rect 132 91 138 125
rect 172 91 178 125
rect 132 53 178 91
rect 132 19 138 53
rect 172 19 178 53
rect 132 -19 178 19
rect 132 -53 138 -19
rect 172 -53 178 -19
rect 132 -91 178 -53
rect 132 -125 138 -91
rect 172 -125 178 -91
rect 132 -163 178 -125
rect 132 -197 138 -163
rect 172 -197 178 -163
rect 132 -235 178 -197
rect 132 -269 138 -235
rect 172 -269 178 -235
rect 132 -307 178 -269
rect 132 -341 138 -307
rect 172 -341 178 -307
rect 132 -379 178 -341
rect 132 -413 138 -379
rect 172 -413 178 -379
rect 132 -451 178 -413
rect 132 -485 138 -451
rect 172 -485 178 -451
rect 132 -523 178 -485
rect 132 -557 138 -523
rect 172 -557 178 -523
rect 132 -595 178 -557
rect 132 -629 138 -595
rect 172 -629 178 -595
rect 132 -667 178 -629
rect 132 -701 138 -667
rect 172 -701 178 -667
rect 132 -739 178 -701
rect 132 -773 138 -739
rect 172 -773 178 -739
rect 132 -811 178 -773
rect 132 -845 138 -811
rect 172 -845 178 -811
rect 132 -883 178 -845
rect 132 -917 138 -883
rect 172 -917 178 -883
rect 132 -955 178 -917
rect 132 -989 138 -955
rect 172 -989 178 -955
rect 132 -1027 178 -989
rect 132 -1061 138 -1027
rect 172 -1061 178 -1027
rect 132 -1099 178 -1061
rect 132 -1133 138 -1099
rect 172 -1133 178 -1099
rect 132 -1171 178 -1133
rect 132 -1205 138 -1171
rect 172 -1205 178 -1171
rect 132 -1243 178 -1205
rect 132 -1277 138 -1243
rect 172 -1277 178 -1243
rect 132 -1315 178 -1277
rect 132 -1349 138 -1315
rect 172 -1349 178 -1315
rect 132 -1387 178 -1349
rect 132 -1421 138 -1387
rect 172 -1421 178 -1387
rect 132 -1459 178 -1421
rect 132 -1493 138 -1459
rect 172 -1493 178 -1459
rect 132 -1531 178 -1493
rect 132 -1565 138 -1531
rect 172 -1565 178 -1531
rect 132 -1603 178 -1565
rect 132 -1637 138 -1603
rect 172 -1637 178 -1603
rect 132 -1675 178 -1637
rect 132 -1709 138 -1675
rect 172 -1709 178 -1675
rect 132 -1747 178 -1709
rect 132 -1781 138 -1747
rect 172 -1781 178 -1747
rect 132 -1806 178 -1781
rect 58 -1844 122 -1838
rect 58 -1878 73 -1844
rect 107 -1878 122 -1844
rect 58 -1884 122 -1878
<< end >>
