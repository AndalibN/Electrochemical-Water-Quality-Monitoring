magic
tech sky130A
magscale 1 2
timestamp 1666402782
<< metal3 >>
rect -2650 2072 2649 2100
rect -2650 -2072 2565 2072
rect 2629 -2072 2649 2072
rect -2650 -2100 2649 -2072
<< via3 >>
rect 2565 -2072 2629 2072
<< mimcap >>
rect -2550 1960 2450 2000
rect -2550 -1960 -2510 1960
rect 2410 -1960 2450 1960
rect -2550 -2000 2450 -1960
<< mimcapcontact >>
rect -2510 -1960 2410 1960
<< metal4 >>
rect 2549 2072 2645 2088
rect -2511 1960 2411 1961
rect -2511 -1960 -2510 1960
rect 2410 -1960 2411 1960
rect -2511 -1961 2411 -1960
rect 2549 -2072 2565 2072
rect 2629 -2072 2645 2072
rect 2549 -2088 2645 -2072
<< properties >>
string FIXED_BBOX -2650 -2100 2550 2100
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25.0 l 20.0 val 1.017k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
