magic
tech sky130A
timestamp 1668049386
<< nmos >>
rect -15 -150 15 150
<< ndiff >>
rect -44 144 -15 150
rect -44 -144 -38 144
rect -21 -144 -15 144
rect -44 -150 -15 -144
rect 15 144 44 150
rect 15 -144 21 144
rect 38 -144 44 144
rect 15 -150 44 -144
<< ndiffc >>
rect -38 -144 -21 144
rect 21 -144 38 144
<< poly >>
rect -15 150 15 163
rect -15 -163 15 -150
<< locali >>
rect -38 144 -21 152
rect -38 -152 -21 -144
rect 21 144 38 152
rect 21 -152 38 -144
<< viali >>
rect -38 -144 -21 144
rect 21 -144 38 144
<< metal1 >>
rect -41 144 -18 150
rect -41 -144 -38 144
rect -21 -144 -18 144
rect -41 -150 -18 -144
rect 18 144 41 150
rect 18 -144 21 144
rect 38 -144 41 144
rect 18 -150 41 -144
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
