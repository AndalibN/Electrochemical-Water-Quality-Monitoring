magic
tech sky130A
magscale 1 2
timestamp 1666105618
<< error_p >>
rect -29 10863 29 10869
rect -29 10829 -17 10863
rect -29 10823 29 10829
rect -114 10482 114 10700
rect -29 10427 29 10433
rect -29 10393 -17 10427
rect -29 10387 29 10393
rect -114 10046 114 10264
rect -29 9991 29 9997
rect -29 9957 -17 9991
rect -29 9951 29 9957
rect -114 9610 114 9828
rect -29 9555 29 9561
rect -29 9521 -17 9555
rect -29 9515 29 9521
rect -114 9174 114 9392
rect -29 9119 29 9125
rect -29 9085 -17 9119
rect -29 9079 29 9085
rect -114 8738 114 8956
rect -29 8683 29 8689
rect -29 8649 -17 8683
rect -29 8643 29 8649
rect -114 8302 114 8520
rect -29 8247 29 8253
rect -29 8213 -17 8247
rect -29 8207 29 8213
rect -114 7866 114 8084
rect -29 7811 29 7817
rect -29 7777 -17 7811
rect -29 7771 29 7777
rect -114 7430 114 7648
rect -29 7375 29 7381
rect -29 7341 -17 7375
rect -29 7335 29 7341
rect -114 6994 114 7212
rect -29 6939 29 6945
rect -29 6905 -17 6939
rect -29 6899 29 6905
rect -114 6558 114 6776
rect -29 6503 29 6509
rect -29 6469 -17 6503
rect -29 6463 29 6469
rect -114 6122 114 6340
rect -29 6067 29 6073
rect -29 6033 -17 6067
rect -29 6027 29 6033
rect -114 5686 114 5904
rect -29 5631 29 5637
rect -29 5597 -17 5631
rect -29 5591 29 5597
rect -114 5250 114 5468
rect -29 5195 29 5201
rect -29 5161 -17 5195
rect -29 5155 29 5161
rect -114 4814 114 5032
rect -29 4759 29 4765
rect -29 4725 -17 4759
rect -29 4719 29 4725
rect -114 4378 114 4596
rect -29 4323 29 4329
rect -29 4289 -17 4323
rect -29 4283 29 4289
rect -114 3942 114 4160
rect -29 3887 29 3893
rect -29 3853 -17 3887
rect -29 3847 29 3853
rect -114 3506 114 3724
rect -29 3451 29 3457
rect -29 3417 -17 3451
rect -29 3411 29 3417
rect -114 3070 114 3288
rect -29 3015 29 3021
rect -29 2981 -17 3015
rect -29 2975 29 2981
rect -114 2634 114 2852
rect -29 2579 29 2585
rect -29 2545 -17 2579
rect -29 2539 29 2545
rect -114 2198 114 2416
rect -29 2143 29 2149
rect -29 2109 -17 2143
rect -29 2103 29 2109
rect -114 1762 114 1980
rect -29 1707 29 1713
rect -29 1673 -17 1707
rect -29 1667 29 1673
rect -114 1326 114 1544
rect -29 1271 29 1277
rect -29 1237 -17 1271
rect -29 1231 29 1237
rect -114 890 114 1108
rect -29 835 29 841
rect -29 801 -17 835
rect -29 795 29 801
rect -114 454 114 672
rect -29 399 29 405
rect -29 365 -17 399
rect -29 359 29 365
rect -114 18 114 236
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -114 -418 114 -200
rect -29 -473 29 -467
rect -29 -507 -17 -473
rect -29 -513 29 -507
rect -114 -854 114 -636
rect -29 -909 29 -903
rect -29 -943 -17 -909
rect -29 -949 29 -943
rect -114 -1290 114 -1072
rect -29 -1345 29 -1339
rect -29 -1379 -17 -1345
rect -29 -1385 29 -1379
rect -114 -1726 114 -1508
rect -29 -1781 29 -1775
rect -29 -1815 -17 -1781
rect -29 -1821 29 -1815
rect -114 -2162 114 -1944
rect -29 -2217 29 -2211
rect -29 -2251 -17 -2217
rect -29 -2257 29 -2251
rect -114 -2598 114 -2380
rect -29 -2653 29 -2647
rect -29 -2687 -17 -2653
rect -29 -2693 29 -2687
rect -114 -3034 114 -2816
rect -29 -3089 29 -3083
rect -29 -3123 -17 -3089
rect -29 -3129 29 -3123
rect -114 -3470 114 -3252
rect -29 -3525 29 -3519
rect -29 -3559 -17 -3525
rect -29 -3565 29 -3559
rect -114 -3906 114 -3688
rect -29 -3961 29 -3955
rect -29 -3995 -17 -3961
rect -29 -4001 29 -3995
rect -114 -4342 114 -4124
rect -29 -4397 29 -4391
rect -29 -4431 -17 -4397
rect -29 -4437 29 -4431
rect -114 -4778 114 -4560
rect -29 -4833 29 -4827
rect -29 -4867 -17 -4833
rect -29 -4873 29 -4867
rect -114 -5214 114 -4996
rect -29 -5269 29 -5263
rect -29 -5303 -17 -5269
rect -29 -5309 29 -5303
rect -114 -5650 114 -5432
rect -29 -5705 29 -5699
rect -29 -5739 -17 -5705
rect -29 -5745 29 -5739
rect -114 -6086 114 -5868
rect -29 -6141 29 -6135
rect -29 -6175 -17 -6141
rect -29 -6181 29 -6175
rect -114 -6522 114 -6304
rect -29 -6577 29 -6571
rect -29 -6611 -17 -6577
rect -29 -6617 29 -6611
rect -114 -6958 114 -6740
rect -29 -7013 29 -7007
rect -29 -7047 -17 -7013
rect -29 -7053 29 -7047
rect -114 -7394 114 -7176
rect -29 -7449 29 -7443
rect -29 -7483 -17 -7449
rect -29 -7489 29 -7483
rect -114 -7830 114 -7612
rect -29 -7885 29 -7879
rect -29 -7919 -17 -7885
rect -29 -7925 29 -7919
rect -114 -8266 114 -8048
rect -29 -8321 29 -8315
rect -29 -8355 -17 -8321
rect -29 -8361 29 -8355
rect -114 -8702 114 -8484
rect -29 -8757 29 -8751
rect -29 -8791 -17 -8757
rect -29 -8797 29 -8791
rect -114 -9138 114 -8920
rect -29 -9193 29 -9187
rect -29 -9227 -17 -9193
rect -29 -9233 29 -9227
rect -114 -9574 114 -9356
rect -29 -9629 29 -9623
rect -29 -9663 -17 -9629
rect -29 -9669 29 -9663
rect -114 -10010 114 -9792
rect -29 -10065 29 -10059
rect -29 -10099 -17 -10065
rect -29 -10105 29 -10099
rect -114 -10446 114 -10228
rect -29 -10501 29 -10495
rect -29 -10535 -17 -10501
rect -29 -10541 29 -10535
rect -29 -10829 29 -10823
rect -29 -10863 -17 -10829
rect -29 -10869 29 -10863
<< nwell >>
rect -114 10482 114 10882
rect -114 10046 114 10446
rect -114 9610 114 10010
rect -114 9174 114 9574
rect -114 8738 114 9138
rect -114 8302 114 8702
rect -114 7866 114 8266
rect -114 7430 114 7830
rect -114 6994 114 7394
rect -114 6558 114 6958
rect -114 6122 114 6522
rect -114 5686 114 6086
rect -114 5250 114 5650
rect -114 4814 114 5214
rect -114 4378 114 4778
rect -114 3942 114 4342
rect -114 3506 114 3906
rect -114 3070 114 3470
rect -114 2634 114 3034
rect -114 2198 114 2598
rect -114 1762 114 2162
rect -114 1326 114 1726
rect -114 890 114 1290
rect -114 454 114 854
rect -114 18 114 418
rect -114 -418 114 -18
rect -114 -854 114 -454
rect -114 -1290 114 -890
rect -114 -1726 114 -1326
rect -114 -2162 114 -1762
rect -114 -2598 114 -2198
rect -114 -3034 114 -2634
rect -114 -3470 114 -3070
rect -114 -3906 114 -3506
rect -114 -4342 114 -3942
rect -114 -4778 114 -4378
rect -114 -5214 114 -4814
rect -114 -5650 114 -5250
rect -114 -6086 114 -5686
rect -114 -6522 114 -6122
rect -114 -6958 114 -6558
rect -114 -7394 114 -6994
rect -114 -7830 114 -7430
rect -114 -8266 114 -7866
rect -114 -8702 114 -8302
rect -114 -9138 114 -8738
rect -114 -9574 114 -9174
rect -114 -10010 114 -9610
rect -114 -10446 114 -10046
rect -114 -10882 114 -10482
<< pmos >>
rect -20 10582 20 10782
rect -20 10146 20 10346
rect -20 9710 20 9910
rect -20 9274 20 9474
rect -20 8838 20 9038
rect -20 8402 20 8602
rect -20 7966 20 8166
rect -20 7530 20 7730
rect -20 7094 20 7294
rect -20 6658 20 6858
rect -20 6222 20 6422
rect -20 5786 20 5986
rect -20 5350 20 5550
rect -20 4914 20 5114
rect -20 4478 20 4678
rect -20 4042 20 4242
rect -20 3606 20 3806
rect -20 3170 20 3370
rect -20 2734 20 2934
rect -20 2298 20 2498
rect -20 1862 20 2062
rect -20 1426 20 1626
rect -20 990 20 1190
rect -20 554 20 754
rect -20 118 20 318
rect -20 -318 20 -118
rect -20 -754 20 -554
rect -20 -1190 20 -990
rect -20 -1626 20 -1426
rect -20 -2062 20 -1862
rect -20 -2498 20 -2298
rect -20 -2934 20 -2734
rect -20 -3370 20 -3170
rect -20 -3806 20 -3606
rect -20 -4242 20 -4042
rect -20 -4678 20 -4478
rect -20 -5114 20 -4914
rect -20 -5550 20 -5350
rect -20 -5986 20 -5786
rect -20 -6422 20 -6222
rect -20 -6858 20 -6658
rect -20 -7294 20 -7094
rect -20 -7730 20 -7530
rect -20 -8166 20 -7966
rect -20 -8602 20 -8402
rect -20 -9038 20 -8838
rect -20 -9474 20 -9274
rect -20 -9910 20 -9710
rect -20 -10346 20 -10146
rect -20 -10782 20 -10582
<< pdiff >>
rect -78 10770 -20 10782
rect -78 10594 -66 10770
rect -32 10594 -20 10770
rect -78 10582 -20 10594
rect 20 10770 78 10782
rect 20 10594 32 10770
rect 66 10594 78 10770
rect 20 10582 78 10594
rect -78 10334 -20 10346
rect -78 10158 -66 10334
rect -32 10158 -20 10334
rect -78 10146 -20 10158
rect 20 10334 78 10346
rect 20 10158 32 10334
rect 66 10158 78 10334
rect 20 10146 78 10158
rect -78 9898 -20 9910
rect -78 9722 -66 9898
rect -32 9722 -20 9898
rect -78 9710 -20 9722
rect 20 9898 78 9910
rect 20 9722 32 9898
rect 66 9722 78 9898
rect 20 9710 78 9722
rect -78 9462 -20 9474
rect -78 9286 -66 9462
rect -32 9286 -20 9462
rect -78 9274 -20 9286
rect 20 9462 78 9474
rect 20 9286 32 9462
rect 66 9286 78 9462
rect 20 9274 78 9286
rect -78 9026 -20 9038
rect -78 8850 -66 9026
rect -32 8850 -20 9026
rect -78 8838 -20 8850
rect 20 9026 78 9038
rect 20 8850 32 9026
rect 66 8850 78 9026
rect 20 8838 78 8850
rect -78 8590 -20 8602
rect -78 8414 -66 8590
rect -32 8414 -20 8590
rect -78 8402 -20 8414
rect 20 8590 78 8602
rect 20 8414 32 8590
rect 66 8414 78 8590
rect 20 8402 78 8414
rect -78 8154 -20 8166
rect -78 7978 -66 8154
rect -32 7978 -20 8154
rect -78 7966 -20 7978
rect 20 8154 78 8166
rect 20 7978 32 8154
rect 66 7978 78 8154
rect 20 7966 78 7978
rect -78 7718 -20 7730
rect -78 7542 -66 7718
rect -32 7542 -20 7718
rect -78 7530 -20 7542
rect 20 7718 78 7730
rect 20 7542 32 7718
rect 66 7542 78 7718
rect 20 7530 78 7542
rect -78 7282 -20 7294
rect -78 7106 -66 7282
rect -32 7106 -20 7282
rect -78 7094 -20 7106
rect 20 7282 78 7294
rect 20 7106 32 7282
rect 66 7106 78 7282
rect 20 7094 78 7106
rect -78 6846 -20 6858
rect -78 6670 -66 6846
rect -32 6670 -20 6846
rect -78 6658 -20 6670
rect 20 6846 78 6858
rect 20 6670 32 6846
rect 66 6670 78 6846
rect 20 6658 78 6670
rect -78 6410 -20 6422
rect -78 6234 -66 6410
rect -32 6234 -20 6410
rect -78 6222 -20 6234
rect 20 6410 78 6422
rect 20 6234 32 6410
rect 66 6234 78 6410
rect 20 6222 78 6234
rect -78 5974 -20 5986
rect -78 5798 -66 5974
rect -32 5798 -20 5974
rect -78 5786 -20 5798
rect 20 5974 78 5986
rect 20 5798 32 5974
rect 66 5798 78 5974
rect 20 5786 78 5798
rect -78 5538 -20 5550
rect -78 5362 -66 5538
rect -32 5362 -20 5538
rect -78 5350 -20 5362
rect 20 5538 78 5550
rect 20 5362 32 5538
rect 66 5362 78 5538
rect 20 5350 78 5362
rect -78 5102 -20 5114
rect -78 4926 -66 5102
rect -32 4926 -20 5102
rect -78 4914 -20 4926
rect 20 5102 78 5114
rect 20 4926 32 5102
rect 66 4926 78 5102
rect 20 4914 78 4926
rect -78 4666 -20 4678
rect -78 4490 -66 4666
rect -32 4490 -20 4666
rect -78 4478 -20 4490
rect 20 4666 78 4678
rect 20 4490 32 4666
rect 66 4490 78 4666
rect 20 4478 78 4490
rect -78 4230 -20 4242
rect -78 4054 -66 4230
rect -32 4054 -20 4230
rect -78 4042 -20 4054
rect 20 4230 78 4242
rect 20 4054 32 4230
rect 66 4054 78 4230
rect 20 4042 78 4054
rect -78 3794 -20 3806
rect -78 3618 -66 3794
rect -32 3618 -20 3794
rect -78 3606 -20 3618
rect 20 3794 78 3806
rect 20 3618 32 3794
rect 66 3618 78 3794
rect 20 3606 78 3618
rect -78 3358 -20 3370
rect -78 3182 -66 3358
rect -32 3182 -20 3358
rect -78 3170 -20 3182
rect 20 3358 78 3370
rect 20 3182 32 3358
rect 66 3182 78 3358
rect 20 3170 78 3182
rect -78 2922 -20 2934
rect -78 2746 -66 2922
rect -32 2746 -20 2922
rect -78 2734 -20 2746
rect 20 2922 78 2934
rect 20 2746 32 2922
rect 66 2746 78 2922
rect 20 2734 78 2746
rect -78 2486 -20 2498
rect -78 2310 -66 2486
rect -32 2310 -20 2486
rect -78 2298 -20 2310
rect 20 2486 78 2498
rect 20 2310 32 2486
rect 66 2310 78 2486
rect 20 2298 78 2310
rect -78 2050 -20 2062
rect -78 1874 -66 2050
rect -32 1874 -20 2050
rect -78 1862 -20 1874
rect 20 2050 78 2062
rect 20 1874 32 2050
rect 66 1874 78 2050
rect 20 1862 78 1874
rect -78 1614 -20 1626
rect -78 1438 -66 1614
rect -32 1438 -20 1614
rect -78 1426 -20 1438
rect 20 1614 78 1626
rect 20 1438 32 1614
rect 66 1438 78 1614
rect 20 1426 78 1438
rect -78 1178 -20 1190
rect -78 1002 -66 1178
rect -32 1002 -20 1178
rect -78 990 -20 1002
rect 20 1178 78 1190
rect 20 1002 32 1178
rect 66 1002 78 1178
rect 20 990 78 1002
rect -78 742 -20 754
rect -78 566 -66 742
rect -32 566 -20 742
rect -78 554 -20 566
rect 20 742 78 754
rect 20 566 32 742
rect 66 566 78 742
rect 20 554 78 566
rect -78 306 -20 318
rect -78 130 -66 306
rect -32 130 -20 306
rect -78 118 -20 130
rect 20 306 78 318
rect 20 130 32 306
rect 66 130 78 306
rect 20 118 78 130
rect -78 -130 -20 -118
rect -78 -306 -66 -130
rect -32 -306 -20 -130
rect -78 -318 -20 -306
rect 20 -130 78 -118
rect 20 -306 32 -130
rect 66 -306 78 -130
rect 20 -318 78 -306
rect -78 -566 -20 -554
rect -78 -742 -66 -566
rect -32 -742 -20 -566
rect -78 -754 -20 -742
rect 20 -566 78 -554
rect 20 -742 32 -566
rect 66 -742 78 -566
rect 20 -754 78 -742
rect -78 -1002 -20 -990
rect -78 -1178 -66 -1002
rect -32 -1178 -20 -1002
rect -78 -1190 -20 -1178
rect 20 -1002 78 -990
rect 20 -1178 32 -1002
rect 66 -1178 78 -1002
rect 20 -1190 78 -1178
rect -78 -1438 -20 -1426
rect -78 -1614 -66 -1438
rect -32 -1614 -20 -1438
rect -78 -1626 -20 -1614
rect 20 -1438 78 -1426
rect 20 -1614 32 -1438
rect 66 -1614 78 -1438
rect 20 -1626 78 -1614
rect -78 -1874 -20 -1862
rect -78 -2050 -66 -1874
rect -32 -2050 -20 -1874
rect -78 -2062 -20 -2050
rect 20 -1874 78 -1862
rect 20 -2050 32 -1874
rect 66 -2050 78 -1874
rect 20 -2062 78 -2050
rect -78 -2310 -20 -2298
rect -78 -2486 -66 -2310
rect -32 -2486 -20 -2310
rect -78 -2498 -20 -2486
rect 20 -2310 78 -2298
rect 20 -2486 32 -2310
rect 66 -2486 78 -2310
rect 20 -2498 78 -2486
rect -78 -2746 -20 -2734
rect -78 -2922 -66 -2746
rect -32 -2922 -20 -2746
rect -78 -2934 -20 -2922
rect 20 -2746 78 -2734
rect 20 -2922 32 -2746
rect 66 -2922 78 -2746
rect 20 -2934 78 -2922
rect -78 -3182 -20 -3170
rect -78 -3358 -66 -3182
rect -32 -3358 -20 -3182
rect -78 -3370 -20 -3358
rect 20 -3182 78 -3170
rect 20 -3358 32 -3182
rect 66 -3358 78 -3182
rect 20 -3370 78 -3358
rect -78 -3618 -20 -3606
rect -78 -3794 -66 -3618
rect -32 -3794 -20 -3618
rect -78 -3806 -20 -3794
rect 20 -3618 78 -3606
rect 20 -3794 32 -3618
rect 66 -3794 78 -3618
rect 20 -3806 78 -3794
rect -78 -4054 -20 -4042
rect -78 -4230 -66 -4054
rect -32 -4230 -20 -4054
rect -78 -4242 -20 -4230
rect 20 -4054 78 -4042
rect 20 -4230 32 -4054
rect 66 -4230 78 -4054
rect 20 -4242 78 -4230
rect -78 -4490 -20 -4478
rect -78 -4666 -66 -4490
rect -32 -4666 -20 -4490
rect -78 -4678 -20 -4666
rect 20 -4490 78 -4478
rect 20 -4666 32 -4490
rect 66 -4666 78 -4490
rect 20 -4678 78 -4666
rect -78 -4926 -20 -4914
rect -78 -5102 -66 -4926
rect -32 -5102 -20 -4926
rect -78 -5114 -20 -5102
rect 20 -4926 78 -4914
rect 20 -5102 32 -4926
rect 66 -5102 78 -4926
rect 20 -5114 78 -5102
rect -78 -5362 -20 -5350
rect -78 -5538 -66 -5362
rect -32 -5538 -20 -5362
rect -78 -5550 -20 -5538
rect 20 -5362 78 -5350
rect 20 -5538 32 -5362
rect 66 -5538 78 -5362
rect 20 -5550 78 -5538
rect -78 -5798 -20 -5786
rect -78 -5974 -66 -5798
rect -32 -5974 -20 -5798
rect -78 -5986 -20 -5974
rect 20 -5798 78 -5786
rect 20 -5974 32 -5798
rect 66 -5974 78 -5798
rect 20 -5986 78 -5974
rect -78 -6234 -20 -6222
rect -78 -6410 -66 -6234
rect -32 -6410 -20 -6234
rect -78 -6422 -20 -6410
rect 20 -6234 78 -6222
rect 20 -6410 32 -6234
rect 66 -6410 78 -6234
rect 20 -6422 78 -6410
rect -78 -6670 -20 -6658
rect -78 -6846 -66 -6670
rect -32 -6846 -20 -6670
rect -78 -6858 -20 -6846
rect 20 -6670 78 -6658
rect 20 -6846 32 -6670
rect 66 -6846 78 -6670
rect 20 -6858 78 -6846
rect -78 -7106 -20 -7094
rect -78 -7282 -66 -7106
rect -32 -7282 -20 -7106
rect -78 -7294 -20 -7282
rect 20 -7106 78 -7094
rect 20 -7282 32 -7106
rect 66 -7282 78 -7106
rect 20 -7294 78 -7282
rect -78 -7542 -20 -7530
rect -78 -7718 -66 -7542
rect -32 -7718 -20 -7542
rect -78 -7730 -20 -7718
rect 20 -7542 78 -7530
rect 20 -7718 32 -7542
rect 66 -7718 78 -7542
rect 20 -7730 78 -7718
rect -78 -7978 -20 -7966
rect -78 -8154 -66 -7978
rect -32 -8154 -20 -7978
rect -78 -8166 -20 -8154
rect 20 -7978 78 -7966
rect 20 -8154 32 -7978
rect 66 -8154 78 -7978
rect 20 -8166 78 -8154
rect -78 -8414 -20 -8402
rect -78 -8590 -66 -8414
rect -32 -8590 -20 -8414
rect -78 -8602 -20 -8590
rect 20 -8414 78 -8402
rect 20 -8590 32 -8414
rect 66 -8590 78 -8414
rect 20 -8602 78 -8590
rect -78 -8850 -20 -8838
rect -78 -9026 -66 -8850
rect -32 -9026 -20 -8850
rect -78 -9038 -20 -9026
rect 20 -8850 78 -8838
rect 20 -9026 32 -8850
rect 66 -9026 78 -8850
rect 20 -9038 78 -9026
rect -78 -9286 -20 -9274
rect -78 -9462 -66 -9286
rect -32 -9462 -20 -9286
rect -78 -9474 -20 -9462
rect 20 -9286 78 -9274
rect 20 -9462 32 -9286
rect 66 -9462 78 -9286
rect 20 -9474 78 -9462
rect -78 -9722 -20 -9710
rect -78 -9898 -66 -9722
rect -32 -9898 -20 -9722
rect -78 -9910 -20 -9898
rect 20 -9722 78 -9710
rect 20 -9898 32 -9722
rect 66 -9898 78 -9722
rect 20 -9910 78 -9898
rect -78 -10158 -20 -10146
rect -78 -10334 -66 -10158
rect -32 -10334 -20 -10158
rect -78 -10346 -20 -10334
rect 20 -10158 78 -10146
rect 20 -10334 32 -10158
rect 66 -10334 78 -10158
rect 20 -10346 78 -10334
rect -78 -10594 -20 -10582
rect -78 -10770 -66 -10594
rect -32 -10770 -20 -10594
rect -78 -10782 -20 -10770
rect 20 -10594 78 -10582
rect 20 -10770 32 -10594
rect 66 -10770 78 -10594
rect 20 -10782 78 -10770
<< pdiffc >>
rect -66 10594 -32 10770
rect 32 10594 66 10770
rect -66 10158 -32 10334
rect 32 10158 66 10334
rect -66 9722 -32 9898
rect 32 9722 66 9898
rect -66 9286 -32 9462
rect 32 9286 66 9462
rect -66 8850 -32 9026
rect 32 8850 66 9026
rect -66 8414 -32 8590
rect 32 8414 66 8590
rect -66 7978 -32 8154
rect 32 7978 66 8154
rect -66 7542 -32 7718
rect 32 7542 66 7718
rect -66 7106 -32 7282
rect 32 7106 66 7282
rect -66 6670 -32 6846
rect 32 6670 66 6846
rect -66 6234 -32 6410
rect 32 6234 66 6410
rect -66 5798 -32 5974
rect 32 5798 66 5974
rect -66 5362 -32 5538
rect 32 5362 66 5538
rect -66 4926 -32 5102
rect 32 4926 66 5102
rect -66 4490 -32 4666
rect 32 4490 66 4666
rect -66 4054 -32 4230
rect 32 4054 66 4230
rect -66 3618 -32 3794
rect 32 3618 66 3794
rect -66 3182 -32 3358
rect 32 3182 66 3358
rect -66 2746 -32 2922
rect 32 2746 66 2922
rect -66 2310 -32 2486
rect 32 2310 66 2486
rect -66 1874 -32 2050
rect 32 1874 66 2050
rect -66 1438 -32 1614
rect 32 1438 66 1614
rect -66 1002 -32 1178
rect 32 1002 66 1178
rect -66 566 -32 742
rect 32 566 66 742
rect -66 130 -32 306
rect 32 130 66 306
rect -66 -306 -32 -130
rect 32 -306 66 -130
rect -66 -742 -32 -566
rect 32 -742 66 -566
rect -66 -1178 -32 -1002
rect 32 -1178 66 -1002
rect -66 -1614 -32 -1438
rect 32 -1614 66 -1438
rect -66 -2050 -32 -1874
rect 32 -2050 66 -1874
rect -66 -2486 -32 -2310
rect 32 -2486 66 -2310
rect -66 -2922 -32 -2746
rect 32 -2922 66 -2746
rect -66 -3358 -32 -3182
rect 32 -3358 66 -3182
rect -66 -3794 -32 -3618
rect 32 -3794 66 -3618
rect -66 -4230 -32 -4054
rect 32 -4230 66 -4054
rect -66 -4666 -32 -4490
rect 32 -4666 66 -4490
rect -66 -5102 -32 -4926
rect 32 -5102 66 -4926
rect -66 -5538 -32 -5362
rect 32 -5538 66 -5362
rect -66 -5974 -32 -5798
rect 32 -5974 66 -5798
rect -66 -6410 -32 -6234
rect 32 -6410 66 -6234
rect -66 -6846 -32 -6670
rect 32 -6846 66 -6670
rect -66 -7282 -32 -7106
rect 32 -7282 66 -7106
rect -66 -7718 -32 -7542
rect 32 -7718 66 -7542
rect -66 -8154 -32 -7978
rect 32 -8154 66 -7978
rect -66 -8590 -32 -8414
rect 32 -8590 66 -8414
rect -66 -9026 -32 -8850
rect 32 -9026 66 -8850
rect -66 -9462 -32 -9286
rect 32 -9462 66 -9286
rect -66 -9898 -32 -9722
rect 32 -9898 66 -9722
rect -66 -10334 -32 -10158
rect 32 -10334 66 -10158
rect -66 -10770 -32 -10594
rect 32 -10770 66 -10594
<< poly >>
rect -33 10863 33 10879
rect -33 10829 -17 10863
rect 17 10829 33 10863
rect -33 10813 33 10829
rect -20 10782 20 10813
rect -20 10551 20 10582
rect -33 10535 33 10551
rect -33 10501 -17 10535
rect 17 10501 33 10535
rect -33 10485 33 10501
rect -33 10427 33 10443
rect -33 10393 -17 10427
rect 17 10393 33 10427
rect -33 10377 33 10393
rect -20 10346 20 10377
rect -20 10115 20 10146
rect -33 10099 33 10115
rect -33 10065 -17 10099
rect 17 10065 33 10099
rect -33 10049 33 10065
rect -33 9991 33 10007
rect -33 9957 -17 9991
rect 17 9957 33 9991
rect -33 9941 33 9957
rect -20 9910 20 9941
rect -20 9679 20 9710
rect -33 9663 33 9679
rect -33 9629 -17 9663
rect 17 9629 33 9663
rect -33 9613 33 9629
rect -33 9555 33 9571
rect -33 9521 -17 9555
rect 17 9521 33 9555
rect -33 9505 33 9521
rect -20 9474 20 9505
rect -20 9243 20 9274
rect -33 9227 33 9243
rect -33 9193 -17 9227
rect 17 9193 33 9227
rect -33 9177 33 9193
rect -33 9119 33 9135
rect -33 9085 -17 9119
rect 17 9085 33 9119
rect -33 9069 33 9085
rect -20 9038 20 9069
rect -20 8807 20 8838
rect -33 8791 33 8807
rect -33 8757 -17 8791
rect 17 8757 33 8791
rect -33 8741 33 8757
rect -33 8683 33 8699
rect -33 8649 -17 8683
rect 17 8649 33 8683
rect -33 8633 33 8649
rect -20 8602 20 8633
rect -20 8371 20 8402
rect -33 8355 33 8371
rect -33 8321 -17 8355
rect 17 8321 33 8355
rect -33 8305 33 8321
rect -33 8247 33 8263
rect -33 8213 -17 8247
rect 17 8213 33 8247
rect -33 8197 33 8213
rect -20 8166 20 8197
rect -20 7935 20 7966
rect -33 7919 33 7935
rect -33 7885 -17 7919
rect 17 7885 33 7919
rect -33 7869 33 7885
rect -33 7811 33 7827
rect -33 7777 -17 7811
rect 17 7777 33 7811
rect -33 7761 33 7777
rect -20 7730 20 7761
rect -20 7499 20 7530
rect -33 7483 33 7499
rect -33 7449 -17 7483
rect 17 7449 33 7483
rect -33 7433 33 7449
rect -33 7375 33 7391
rect -33 7341 -17 7375
rect 17 7341 33 7375
rect -33 7325 33 7341
rect -20 7294 20 7325
rect -20 7063 20 7094
rect -33 7047 33 7063
rect -33 7013 -17 7047
rect 17 7013 33 7047
rect -33 6997 33 7013
rect -33 6939 33 6955
rect -33 6905 -17 6939
rect 17 6905 33 6939
rect -33 6889 33 6905
rect -20 6858 20 6889
rect -20 6627 20 6658
rect -33 6611 33 6627
rect -33 6577 -17 6611
rect 17 6577 33 6611
rect -33 6561 33 6577
rect -33 6503 33 6519
rect -33 6469 -17 6503
rect 17 6469 33 6503
rect -33 6453 33 6469
rect -20 6422 20 6453
rect -20 6191 20 6222
rect -33 6175 33 6191
rect -33 6141 -17 6175
rect 17 6141 33 6175
rect -33 6125 33 6141
rect -33 6067 33 6083
rect -33 6033 -17 6067
rect 17 6033 33 6067
rect -33 6017 33 6033
rect -20 5986 20 6017
rect -20 5755 20 5786
rect -33 5739 33 5755
rect -33 5705 -17 5739
rect 17 5705 33 5739
rect -33 5689 33 5705
rect -33 5631 33 5647
rect -33 5597 -17 5631
rect 17 5597 33 5631
rect -33 5581 33 5597
rect -20 5550 20 5581
rect -20 5319 20 5350
rect -33 5303 33 5319
rect -33 5269 -17 5303
rect 17 5269 33 5303
rect -33 5253 33 5269
rect -33 5195 33 5211
rect -33 5161 -17 5195
rect 17 5161 33 5195
rect -33 5145 33 5161
rect -20 5114 20 5145
rect -20 4883 20 4914
rect -33 4867 33 4883
rect -33 4833 -17 4867
rect 17 4833 33 4867
rect -33 4817 33 4833
rect -33 4759 33 4775
rect -33 4725 -17 4759
rect 17 4725 33 4759
rect -33 4709 33 4725
rect -20 4678 20 4709
rect -20 4447 20 4478
rect -33 4431 33 4447
rect -33 4397 -17 4431
rect 17 4397 33 4431
rect -33 4381 33 4397
rect -33 4323 33 4339
rect -33 4289 -17 4323
rect 17 4289 33 4323
rect -33 4273 33 4289
rect -20 4242 20 4273
rect -20 4011 20 4042
rect -33 3995 33 4011
rect -33 3961 -17 3995
rect 17 3961 33 3995
rect -33 3945 33 3961
rect -33 3887 33 3903
rect -33 3853 -17 3887
rect 17 3853 33 3887
rect -33 3837 33 3853
rect -20 3806 20 3837
rect -20 3575 20 3606
rect -33 3559 33 3575
rect -33 3525 -17 3559
rect 17 3525 33 3559
rect -33 3509 33 3525
rect -33 3451 33 3467
rect -33 3417 -17 3451
rect 17 3417 33 3451
rect -33 3401 33 3417
rect -20 3370 20 3401
rect -20 3139 20 3170
rect -33 3123 33 3139
rect -33 3089 -17 3123
rect 17 3089 33 3123
rect -33 3073 33 3089
rect -33 3015 33 3031
rect -33 2981 -17 3015
rect 17 2981 33 3015
rect -33 2965 33 2981
rect -20 2934 20 2965
rect -20 2703 20 2734
rect -33 2687 33 2703
rect -33 2653 -17 2687
rect 17 2653 33 2687
rect -33 2637 33 2653
rect -33 2579 33 2595
rect -33 2545 -17 2579
rect 17 2545 33 2579
rect -33 2529 33 2545
rect -20 2498 20 2529
rect -20 2267 20 2298
rect -33 2251 33 2267
rect -33 2217 -17 2251
rect 17 2217 33 2251
rect -33 2201 33 2217
rect -33 2143 33 2159
rect -33 2109 -17 2143
rect 17 2109 33 2143
rect -33 2093 33 2109
rect -20 2062 20 2093
rect -20 1831 20 1862
rect -33 1815 33 1831
rect -33 1781 -17 1815
rect 17 1781 33 1815
rect -33 1765 33 1781
rect -33 1707 33 1723
rect -33 1673 -17 1707
rect 17 1673 33 1707
rect -33 1657 33 1673
rect -20 1626 20 1657
rect -20 1395 20 1426
rect -33 1379 33 1395
rect -33 1345 -17 1379
rect 17 1345 33 1379
rect -33 1329 33 1345
rect -33 1271 33 1287
rect -33 1237 -17 1271
rect 17 1237 33 1271
rect -33 1221 33 1237
rect -20 1190 20 1221
rect -20 959 20 990
rect -33 943 33 959
rect -33 909 -17 943
rect 17 909 33 943
rect -33 893 33 909
rect -33 835 33 851
rect -33 801 -17 835
rect 17 801 33 835
rect -33 785 33 801
rect -20 754 20 785
rect -20 523 20 554
rect -33 507 33 523
rect -33 473 -17 507
rect 17 473 33 507
rect -33 457 33 473
rect -33 399 33 415
rect -33 365 -17 399
rect 17 365 33 399
rect -33 349 33 365
rect -20 318 20 349
rect -20 87 20 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -20 -118 20 -87
rect -20 -349 20 -318
rect -33 -365 33 -349
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -415 33 -399
rect -33 -473 33 -457
rect -33 -507 -17 -473
rect 17 -507 33 -473
rect -33 -523 33 -507
rect -20 -554 20 -523
rect -20 -785 20 -754
rect -33 -801 33 -785
rect -33 -835 -17 -801
rect 17 -835 33 -801
rect -33 -851 33 -835
rect -33 -909 33 -893
rect -33 -943 -17 -909
rect 17 -943 33 -909
rect -33 -959 33 -943
rect -20 -990 20 -959
rect -20 -1221 20 -1190
rect -33 -1237 33 -1221
rect -33 -1271 -17 -1237
rect 17 -1271 33 -1237
rect -33 -1287 33 -1271
rect -33 -1345 33 -1329
rect -33 -1379 -17 -1345
rect 17 -1379 33 -1345
rect -33 -1395 33 -1379
rect -20 -1426 20 -1395
rect -20 -1657 20 -1626
rect -33 -1673 33 -1657
rect -33 -1707 -17 -1673
rect 17 -1707 33 -1673
rect -33 -1723 33 -1707
rect -33 -1781 33 -1765
rect -33 -1815 -17 -1781
rect 17 -1815 33 -1781
rect -33 -1831 33 -1815
rect -20 -1862 20 -1831
rect -20 -2093 20 -2062
rect -33 -2109 33 -2093
rect -33 -2143 -17 -2109
rect 17 -2143 33 -2109
rect -33 -2159 33 -2143
rect -33 -2217 33 -2201
rect -33 -2251 -17 -2217
rect 17 -2251 33 -2217
rect -33 -2267 33 -2251
rect -20 -2298 20 -2267
rect -20 -2529 20 -2498
rect -33 -2545 33 -2529
rect -33 -2579 -17 -2545
rect 17 -2579 33 -2545
rect -33 -2595 33 -2579
rect -33 -2653 33 -2637
rect -33 -2687 -17 -2653
rect 17 -2687 33 -2653
rect -33 -2703 33 -2687
rect -20 -2734 20 -2703
rect -20 -2965 20 -2934
rect -33 -2981 33 -2965
rect -33 -3015 -17 -2981
rect 17 -3015 33 -2981
rect -33 -3031 33 -3015
rect -33 -3089 33 -3073
rect -33 -3123 -17 -3089
rect 17 -3123 33 -3089
rect -33 -3139 33 -3123
rect -20 -3170 20 -3139
rect -20 -3401 20 -3370
rect -33 -3417 33 -3401
rect -33 -3451 -17 -3417
rect 17 -3451 33 -3417
rect -33 -3467 33 -3451
rect -33 -3525 33 -3509
rect -33 -3559 -17 -3525
rect 17 -3559 33 -3525
rect -33 -3575 33 -3559
rect -20 -3606 20 -3575
rect -20 -3837 20 -3806
rect -33 -3853 33 -3837
rect -33 -3887 -17 -3853
rect 17 -3887 33 -3853
rect -33 -3903 33 -3887
rect -33 -3961 33 -3945
rect -33 -3995 -17 -3961
rect 17 -3995 33 -3961
rect -33 -4011 33 -3995
rect -20 -4042 20 -4011
rect -20 -4273 20 -4242
rect -33 -4289 33 -4273
rect -33 -4323 -17 -4289
rect 17 -4323 33 -4289
rect -33 -4339 33 -4323
rect -33 -4397 33 -4381
rect -33 -4431 -17 -4397
rect 17 -4431 33 -4397
rect -33 -4447 33 -4431
rect -20 -4478 20 -4447
rect -20 -4709 20 -4678
rect -33 -4725 33 -4709
rect -33 -4759 -17 -4725
rect 17 -4759 33 -4725
rect -33 -4775 33 -4759
rect -33 -4833 33 -4817
rect -33 -4867 -17 -4833
rect 17 -4867 33 -4833
rect -33 -4883 33 -4867
rect -20 -4914 20 -4883
rect -20 -5145 20 -5114
rect -33 -5161 33 -5145
rect -33 -5195 -17 -5161
rect 17 -5195 33 -5161
rect -33 -5211 33 -5195
rect -33 -5269 33 -5253
rect -33 -5303 -17 -5269
rect 17 -5303 33 -5269
rect -33 -5319 33 -5303
rect -20 -5350 20 -5319
rect -20 -5581 20 -5550
rect -33 -5597 33 -5581
rect -33 -5631 -17 -5597
rect 17 -5631 33 -5597
rect -33 -5647 33 -5631
rect -33 -5705 33 -5689
rect -33 -5739 -17 -5705
rect 17 -5739 33 -5705
rect -33 -5755 33 -5739
rect -20 -5786 20 -5755
rect -20 -6017 20 -5986
rect -33 -6033 33 -6017
rect -33 -6067 -17 -6033
rect 17 -6067 33 -6033
rect -33 -6083 33 -6067
rect -33 -6141 33 -6125
rect -33 -6175 -17 -6141
rect 17 -6175 33 -6141
rect -33 -6191 33 -6175
rect -20 -6222 20 -6191
rect -20 -6453 20 -6422
rect -33 -6469 33 -6453
rect -33 -6503 -17 -6469
rect 17 -6503 33 -6469
rect -33 -6519 33 -6503
rect -33 -6577 33 -6561
rect -33 -6611 -17 -6577
rect 17 -6611 33 -6577
rect -33 -6627 33 -6611
rect -20 -6658 20 -6627
rect -20 -6889 20 -6858
rect -33 -6905 33 -6889
rect -33 -6939 -17 -6905
rect 17 -6939 33 -6905
rect -33 -6955 33 -6939
rect -33 -7013 33 -6997
rect -33 -7047 -17 -7013
rect 17 -7047 33 -7013
rect -33 -7063 33 -7047
rect -20 -7094 20 -7063
rect -20 -7325 20 -7294
rect -33 -7341 33 -7325
rect -33 -7375 -17 -7341
rect 17 -7375 33 -7341
rect -33 -7391 33 -7375
rect -33 -7449 33 -7433
rect -33 -7483 -17 -7449
rect 17 -7483 33 -7449
rect -33 -7499 33 -7483
rect -20 -7530 20 -7499
rect -20 -7761 20 -7730
rect -33 -7777 33 -7761
rect -33 -7811 -17 -7777
rect 17 -7811 33 -7777
rect -33 -7827 33 -7811
rect -33 -7885 33 -7869
rect -33 -7919 -17 -7885
rect 17 -7919 33 -7885
rect -33 -7935 33 -7919
rect -20 -7966 20 -7935
rect -20 -8197 20 -8166
rect -33 -8213 33 -8197
rect -33 -8247 -17 -8213
rect 17 -8247 33 -8213
rect -33 -8263 33 -8247
rect -33 -8321 33 -8305
rect -33 -8355 -17 -8321
rect 17 -8355 33 -8321
rect -33 -8371 33 -8355
rect -20 -8402 20 -8371
rect -20 -8633 20 -8602
rect -33 -8649 33 -8633
rect -33 -8683 -17 -8649
rect 17 -8683 33 -8649
rect -33 -8699 33 -8683
rect -33 -8757 33 -8741
rect -33 -8791 -17 -8757
rect 17 -8791 33 -8757
rect -33 -8807 33 -8791
rect -20 -8838 20 -8807
rect -20 -9069 20 -9038
rect -33 -9085 33 -9069
rect -33 -9119 -17 -9085
rect 17 -9119 33 -9085
rect -33 -9135 33 -9119
rect -33 -9193 33 -9177
rect -33 -9227 -17 -9193
rect 17 -9227 33 -9193
rect -33 -9243 33 -9227
rect -20 -9274 20 -9243
rect -20 -9505 20 -9474
rect -33 -9521 33 -9505
rect -33 -9555 -17 -9521
rect 17 -9555 33 -9521
rect -33 -9571 33 -9555
rect -33 -9629 33 -9613
rect -33 -9663 -17 -9629
rect 17 -9663 33 -9629
rect -33 -9679 33 -9663
rect -20 -9710 20 -9679
rect -20 -9941 20 -9910
rect -33 -9957 33 -9941
rect -33 -9991 -17 -9957
rect 17 -9991 33 -9957
rect -33 -10007 33 -9991
rect -33 -10065 33 -10049
rect -33 -10099 -17 -10065
rect 17 -10099 33 -10065
rect -33 -10115 33 -10099
rect -20 -10146 20 -10115
rect -20 -10377 20 -10346
rect -33 -10393 33 -10377
rect -33 -10427 -17 -10393
rect 17 -10427 33 -10393
rect -33 -10443 33 -10427
rect -33 -10501 33 -10485
rect -33 -10535 -17 -10501
rect 17 -10535 33 -10501
rect -33 -10551 33 -10535
rect -20 -10582 20 -10551
rect -20 -10813 20 -10782
rect -33 -10829 33 -10813
rect -33 -10863 -17 -10829
rect 17 -10863 33 -10829
rect -33 -10879 33 -10863
<< polycont >>
rect -17 10829 17 10863
rect -17 10501 17 10535
rect -17 10393 17 10427
rect -17 10065 17 10099
rect -17 9957 17 9991
rect -17 9629 17 9663
rect -17 9521 17 9555
rect -17 9193 17 9227
rect -17 9085 17 9119
rect -17 8757 17 8791
rect -17 8649 17 8683
rect -17 8321 17 8355
rect -17 8213 17 8247
rect -17 7885 17 7919
rect -17 7777 17 7811
rect -17 7449 17 7483
rect -17 7341 17 7375
rect -17 7013 17 7047
rect -17 6905 17 6939
rect -17 6577 17 6611
rect -17 6469 17 6503
rect -17 6141 17 6175
rect -17 6033 17 6067
rect -17 5705 17 5739
rect -17 5597 17 5631
rect -17 5269 17 5303
rect -17 5161 17 5195
rect -17 4833 17 4867
rect -17 4725 17 4759
rect -17 4397 17 4431
rect -17 4289 17 4323
rect -17 3961 17 3995
rect -17 3853 17 3887
rect -17 3525 17 3559
rect -17 3417 17 3451
rect -17 3089 17 3123
rect -17 2981 17 3015
rect -17 2653 17 2687
rect -17 2545 17 2579
rect -17 2217 17 2251
rect -17 2109 17 2143
rect -17 1781 17 1815
rect -17 1673 17 1707
rect -17 1345 17 1379
rect -17 1237 17 1271
rect -17 909 17 943
rect -17 801 17 835
rect -17 473 17 507
rect -17 365 17 399
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -399 17 -365
rect -17 -507 17 -473
rect -17 -835 17 -801
rect -17 -943 17 -909
rect -17 -1271 17 -1237
rect -17 -1379 17 -1345
rect -17 -1707 17 -1673
rect -17 -1815 17 -1781
rect -17 -2143 17 -2109
rect -17 -2251 17 -2217
rect -17 -2579 17 -2545
rect -17 -2687 17 -2653
rect -17 -3015 17 -2981
rect -17 -3123 17 -3089
rect -17 -3451 17 -3417
rect -17 -3559 17 -3525
rect -17 -3887 17 -3853
rect -17 -3995 17 -3961
rect -17 -4323 17 -4289
rect -17 -4431 17 -4397
rect -17 -4759 17 -4725
rect -17 -4867 17 -4833
rect -17 -5195 17 -5161
rect -17 -5303 17 -5269
rect -17 -5631 17 -5597
rect -17 -5739 17 -5705
rect -17 -6067 17 -6033
rect -17 -6175 17 -6141
rect -17 -6503 17 -6469
rect -17 -6611 17 -6577
rect -17 -6939 17 -6905
rect -17 -7047 17 -7013
rect -17 -7375 17 -7341
rect -17 -7483 17 -7449
rect -17 -7811 17 -7777
rect -17 -7919 17 -7885
rect -17 -8247 17 -8213
rect -17 -8355 17 -8321
rect -17 -8683 17 -8649
rect -17 -8791 17 -8757
rect -17 -9119 17 -9085
rect -17 -9227 17 -9193
rect -17 -9555 17 -9521
rect -17 -9663 17 -9629
rect -17 -9991 17 -9957
rect -17 -10099 17 -10065
rect -17 -10427 17 -10393
rect -17 -10535 17 -10501
rect -17 -10863 17 -10829
<< locali >>
rect -33 10829 -17 10863
rect 17 10829 33 10863
rect -66 10770 -32 10786
rect -66 10578 -32 10594
rect 32 10770 66 10786
rect 32 10578 66 10594
rect -33 10501 -17 10535
rect 17 10501 33 10535
rect -33 10393 -17 10427
rect 17 10393 33 10427
rect -66 10334 -32 10350
rect -66 10142 -32 10158
rect 32 10334 66 10350
rect 32 10142 66 10158
rect -33 10065 -17 10099
rect 17 10065 33 10099
rect -33 9957 -17 9991
rect 17 9957 33 9991
rect -66 9898 -32 9914
rect -66 9706 -32 9722
rect 32 9898 66 9914
rect 32 9706 66 9722
rect -33 9629 -17 9663
rect 17 9629 33 9663
rect -33 9521 -17 9555
rect 17 9521 33 9555
rect -66 9462 -32 9478
rect -66 9270 -32 9286
rect 32 9462 66 9478
rect 32 9270 66 9286
rect -33 9193 -17 9227
rect 17 9193 33 9227
rect -33 9085 -17 9119
rect 17 9085 33 9119
rect -66 9026 -32 9042
rect -66 8834 -32 8850
rect 32 9026 66 9042
rect 32 8834 66 8850
rect -33 8757 -17 8791
rect 17 8757 33 8791
rect -33 8649 -17 8683
rect 17 8649 33 8683
rect -66 8590 -32 8606
rect -66 8398 -32 8414
rect 32 8590 66 8606
rect 32 8398 66 8414
rect -33 8321 -17 8355
rect 17 8321 33 8355
rect -33 8213 -17 8247
rect 17 8213 33 8247
rect -66 8154 -32 8170
rect -66 7962 -32 7978
rect 32 8154 66 8170
rect 32 7962 66 7978
rect -33 7885 -17 7919
rect 17 7885 33 7919
rect -33 7777 -17 7811
rect 17 7777 33 7811
rect -66 7718 -32 7734
rect -66 7526 -32 7542
rect 32 7718 66 7734
rect 32 7526 66 7542
rect -33 7449 -17 7483
rect 17 7449 33 7483
rect -33 7341 -17 7375
rect 17 7341 33 7375
rect -66 7282 -32 7298
rect -66 7090 -32 7106
rect 32 7282 66 7298
rect 32 7090 66 7106
rect -33 7013 -17 7047
rect 17 7013 33 7047
rect -33 6905 -17 6939
rect 17 6905 33 6939
rect -66 6846 -32 6862
rect -66 6654 -32 6670
rect 32 6846 66 6862
rect 32 6654 66 6670
rect -33 6577 -17 6611
rect 17 6577 33 6611
rect -33 6469 -17 6503
rect 17 6469 33 6503
rect -66 6410 -32 6426
rect -66 6218 -32 6234
rect 32 6410 66 6426
rect 32 6218 66 6234
rect -33 6141 -17 6175
rect 17 6141 33 6175
rect -33 6033 -17 6067
rect 17 6033 33 6067
rect -66 5974 -32 5990
rect -66 5782 -32 5798
rect 32 5974 66 5990
rect 32 5782 66 5798
rect -33 5705 -17 5739
rect 17 5705 33 5739
rect -33 5597 -17 5631
rect 17 5597 33 5631
rect -66 5538 -32 5554
rect -66 5346 -32 5362
rect 32 5538 66 5554
rect 32 5346 66 5362
rect -33 5269 -17 5303
rect 17 5269 33 5303
rect -33 5161 -17 5195
rect 17 5161 33 5195
rect -66 5102 -32 5118
rect -66 4910 -32 4926
rect 32 5102 66 5118
rect 32 4910 66 4926
rect -33 4833 -17 4867
rect 17 4833 33 4867
rect -33 4725 -17 4759
rect 17 4725 33 4759
rect -66 4666 -32 4682
rect -66 4474 -32 4490
rect 32 4666 66 4682
rect 32 4474 66 4490
rect -33 4397 -17 4431
rect 17 4397 33 4431
rect -33 4289 -17 4323
rect 17 4289 33 4323
rect -66 4230 -32 4246
rect -66 4038 -32 4054
rect 32 4230 66 4246
rect 32 4038 66 4054
rect -33 3961 -17 3995
rect 17 3961 33 3995
rect -33 3853 -17 3887
rect 17 3853 33 3887
rect -66 3794 -32 3810
rect -66 3602 -32 3618
rect 32 3794 66 3810
rect 32 3602 66 3618
rect -33 3525 -17 3559
rect 17 3525 33 3559
rect -33 3417 -17 3451
rect 17 3417 33 3451
rect -66 3358 -32 3374
rect -66 3166 -32 3182
rect 32 3358 66 3374
rect 32 3166 66 3182
rect -33 3089 -17 3123
rect 17 3089 33 3123
rect -33 2981 -17 3015
rect 17 2981 33 3015
rect -66 2922 -32 2938
rect -66 2730 -32 2746
rect 32 2922 66 2938
rect 32 2730 66 2746
rect -33 2653 -17 2687
rect 17 2653 33 2687
rect -33 2545 -17 2579
rect 17 2545 33 2579
rect -66 2486 -32 2502
rect -66 2294 -32 2310
rect 32 2486 66 2502
rect 32 2294 66 2310
rect -33 2217 -17 2251
rect 17 2217 33 2251
rect -33 2109 -17 2143
rect 17 2109 33 2143
rect -66 2050 -32 2066
rect -66 1858 -32 1874
rect 32 2050 66 2066
rect 32 1858 66 1874
rect -33 1781 -17 1815
rect 17 1781 33 1815
rect -33 1673 -17 1707
rect 17 1673 33 1707
rect -66 1614 -32 1630
rect -66 1422 -32 1438
rect 32 1614 66 1630
rect 32 1422 66 1438
rect -33 1345 -17 1379
rect 17 1345 33 1379
rect -33 1237 -17 1271
rect 17 1237 33 1271
rect -66 1178 -32 1194
rect -66 986 -32 1002
rect 32 1178 66 1194
rect 32 986 66 1002
rect -33 909 -17 943
rect 17 909 33 943
rect -33 801 -17 835
rect 17 801 33 835
rect -66 742 -32 758
rect -66 550 -32 566
rect 32 742 66 758
rect 32 550 66 566
rect -33 473 -17 507
rect 17 473 33 507
rect -33 365 -17 399
rect 17 365 33 399
rect -66 306 -32 322
rect -66 114 -32 130
rect 32 306 66 322
rect 32 114 66 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -66 -130 -32 -114
rect -66 -322 -32 -306
rect 32 -130 66 -114
rect 32 -322 66 -306
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -507 -17 -473
rect 17 -507 33 -473
rect -66 -566 -32 -550
rect -66 -758 -32 -742
rect 32 -566 66 -550
rect 32 -758 66 -742
rect -33 -835 -17 -801
rect 17 -835 33 -801
rect -33 -943 -17 -909
rect 17 -943 33 -909
rect -66 -1002 -32 -986
rect -66 -1194 -32 -1178
rect 32 -1002 66 -986
rect 32 -1194 66 -1178
rect -33 -1271 -17 -1237
rect 17 -1271 33 -1237
rect -33 -1379 -17 -1345
rect 17 -1379 33 -1345
rect -66 -1438 -32 -1422
rect -66 -1630 -32 -1614
rect 32 -1438 66 -1422
rect 32 -1630 66 -1614
rect -33 -1707 -17 -1673
rect 17 -1707 33 -1673
rect -33 -1815 -17 -1781
rect 17 -1815 33 -1781
rect -66 -1874 -32 -1858
rect -66 -2066 -32 -2050
rect 32 -1874 66 -1858
rect 32 -2066 66 -2050
rect -33 -2143 -17 -2109
rect 17 -2143 33 -2109
rect -33 -2251 -17 -2217
rect 17 -2251 33 -2217
rect -66 -2310 -32 -2294
rect -66 -2502 -32 -2486
rect 32 -2310 66 -2294
rect 32 -2502 66 -2486
rect -33 -2579 -17 -2545
rect 17 -2579 33 -2545
rect -33 -2687 -17 -2653
rect 17 -2687 33 -2653
rect -66 -2746 -32 -2730
rect -66 -2938 -32 -2922
rect 32 -2746 66 -2730
rect 32 -2938 66 -2922
rect -33 -3015 -17 -2981
rect 17 -3015 33 -2981
rect -33 -3123 -17 -3089
rect 17 -3123 33 -3089
rect -66 -3182 -32 -3166
rect -66 -3374 -32 -3358
rect 32 -3182 66 -3166
rect 32 -3374 66 -3358
rect -33 -3451 -17 -3417
rect 17 -3451 33 -3417
rect -33 -3559 -17 -3525
rect 17 -3559 33 -3525
rect -66 -3618 -32 -3602
rect -66 -3810 -32 -3794
rect 32 -3618 66 -3602
rect 32 -3810 66 -3794
rect -33 -3887 -17 -3853
rect 17 -3887 33 -3853
rect -33 -3995 -17 -3961
rect 17 -3995 33 -3961
rect -66 -4054 -32 -4038
rect -66 -4246 -32 -4230
rect 32 -4054 66 -4038
rect 32 -4246 66 -4230
rect -33 -4323 -17 -4289
rect 17 -4323 33 -4289
rect -33 -4431 -17 -4397
rect 17 -4431 33 -4397
rect -66 -4490 -32 -4474
rect -66 -4682 -32 -4666
rect 32 -4490 66 -4474
rect 32 -4682 66 -4666
rect -33 -4759 -17 -4725
rect 17 -4759 33 -4725
rect -33 -4867 -17 -4833
rect 17 -4867 33 -4833
rect -66 -4926 -32 -4910
rect -66 -5118 -32 -5102
rect 32 -4926 66 -4910
rect 32 -5118 66 -5102
rect -33 -5195 -17 -5161
rect 17 -5195 33 -5161
rect -33 -5303 -17 -5269
rect 17 -5303 33 -5269
rect -66 -5362 -32 -5346
rect -66 -5554 -32 -5538
rect 32 -5362 66 -5346
rect 32 -5554 66 -5538
rect -33 -5631 -17 -5597
rect 17 -5631 33 -5597
rect -33 -5739 -17 -5705
rect 17 -5739 33 -5705
rect -66 -5798 -32 -5782
rect -66 -5990 -32 -5974
rect 32 -5798 66 -5782
rect 32 -5990 66 -5974
rect -33 -6067 -17 -6033
rect 17 -6067 33 -6033
rect -33 -6175 -17 -6141
rect 17 -6175 33 -6141
rect -66 -6234 -32 -6218
rect -66 -6426 -32 -6410
rect 32 -6234 66 -6218
rect 32 -6426 66 -6410
rect -33 -6503 -17 -6469
rect 17 -6503 33 -6469
rect -33 -6611 -17 -6577
rect 17 -6611 33 -6577
rect -66 -6670 -32 -6654
rect -66 -6862 -32 -6846
rect 32 -6670 66 -6654
rect 32 -6862 66 -6846
rect -33 -6939 -17 -6905
rect 17 -6939 33 -6905
rect -33 -7047 -17 -7013
rect 17 -7047 33 -7013
rect -66 -7106 -32 -7090
rect -66 -7298 -32 -7282
rect 32 -7106 66 -7090
rect 32 -7298 66 -7282
rect -33 -7375 -17 -7341
rect 17 -7375 33 -7341
rect -33 -7483 -17 -7449
rect 17 -7483 33 -7449
rect -66 -7542 -32 -7526
rect -66 -7734 -32 -7718
rect 32 -7542 66 -7526
rect 32 -7734 66 -7718
rect -33 -7811 -17 -7777
rect 17 -7811 33 -7777
rect -33 -7919 -17 -7885
rect 17 -7919 33 -7885
rect -66 -7978 -32 -7962
rect -66 -8170 -32 -8154
rect 32 -7978 66 -7962
rect 32 -8170 66 -8154
rect -33 -8247 -17 -8213
rect 17 -8247 33 -8213
rect -33 -8355 -17 -8321
rect 17 -8355 33 -8321
rect -66 -8414 -32 -8398
rect -66 -8606 -32 -8590
rect 32 -8414 66 -8398
rect 32 -8606 66 -8590
rect -33 -8683 -17 -8649
rect 17 -8683 33 -8649
rect -33 -8791 -17 -8757
rect 17 -8791 33 -8757
rect -66 -8850 -32 -8834
rect -66 -9042 -32 -9026
rect 32 -8850 66 -8834
rect 32 -9042 66 -9026
rect -33 -9119 -17 -9085
rect 17 -9119 33 -9085
rect -33 -9227 -17 -9193
rect 17 -9227 33 -9193
rect -66 -9286 -32 -9270
rect -66 -9478 -32 -9462
rect 32 -9286 66 -9270
rect 32 -9478 66 -9462
rect -33 -9555 -17 -9521
rect 17 -9555 33 -9521
rect -33 -9663 -17 -9629
rect 17 -9663 33 -9629
rect -66 -9722 -32 -9706
rect -66 -9914 -32 -9898
rect 32 -9722 66 -9706
rect 32 -9914 66 -9898
rect -33 -9991 -17 -9957
rect 17 -9991 33 -9957
rect -33 -10099 -17 -10065
rect 17 -10099 33 -10065
rect -66 -10158 -32 -10142
rect -66 -10350 -32 -10334
rect 32 -10158 66 -10142
rect 32 -10350 66 -10334
rect -33 -10427 -17 -10393
rect 17 -10427 33 -10393
rect -33 -10535 -17 -10501
rect 17 -10535 33 -10501
rect -66 -10594 -32 -10578
rect -66 -10786 -32 -10770
rect 32 -10594 66 -10578
rect 32 -10786 66 -10770
rect -33 -10863 -17 -10829
rect 17 -10863 33 -10829
<< viali >>
rect -17 10829 17 10863
rect -66 10594 -32 10770
rect 32 10594 66 10770
rect -17 10501 17 10535
rect -17 10393 17 10427
rect -66 10158 -32 10334
rect 32 10158 66 10334
rect -17 10065 17 10099
rect -17 9957 17 9991
rect -66 9722 -32 9898
rect 32 9722 66 9898
rect -17 9629 17 9663
rect -17 9521 17 9555
rect -66 9286 -32 9462
rect 32 9286 66 9462
rect -17 9193 17 9227
rect -17 9085 17 9119
rect -66 8850 -32 9026
rect 32 8850 66 9026
rect -17 8757 17 8791
rect -17 8649 17 8683
rect -66 8414 -32 8590
rect 32 8414 66 8590
rect -17 8321 17 8355
rect -17 8213 17 8247
rect -66 7978 -32 8154
rect 32 7978 66 8154
rect -17 7885 17 7919
rect -17 7777 17 7811
rect -66 7542 -32 7718
rect 32 7542 66 7718
rect -17 7449 17 7483
rect -17 7341 17 7375
rect -66 7106 -32 7282
rect 32 7106 66 7282
rect -17 7013 17 7047
rect -17 6905 17 6939
rect -66 6670 -32 6846
rect 32 6670 66 6846
rect -17 6577 17 6611
rect -17 6469 17 6503
rect -66 6234 -32 6410
rect 32 6234 66 6410
rect -17 6141 17 6175
rect -17 6033 17 6067
rect -66 5798 -32 5974
rect 32 5798 66 5974
rect -17 5705 17 5739
rect -17 5597 17 5631
rect -66 5362 -32 5538
rect 32 5362 66 5538
rect -17 5269 17 5303
rect -17 5161 17 5195
rect -66 4926 -32 5102
rect 32 4926 66 5102
rect -17 4833 17 4867
rect -17 4725 17 4759
rect -66 4490 -32 4666
rect 32 4490 66 4666
rect -17 4397 17 4431
rect -17 4289 17 4323
rect -66 4054 -32 4230
rect 32 4054 66 4230
rect -17 3961 17 3995
rect -17 3853 17 3887
rect -66 3618 -32 3794
rect 32 3618 66 3794
rect -17 3525 17 3559
rect -17 3417 17 3451
rect -66 3182 -32 3358
rect 32 3182 66 3358
rect -17 3089 17 3123
rect -17 2981 17 3015
rect -66 2746 -32 2922
rect 32 2746 66 2922
rect -17 2653 17 2687
rect -17 2545 17 2579
rect -66 2310 -32 2486
rect 32 2310 66 2486
rect -17 2217 17 2251
rect -17 2109 17 2143
rect -66 1874 -32 2050
rect 32 1874 66 2050
rect -17 1781 17 1815
rect -17 1673 17 1707
rect -66 1438 -32 1614
rect 32 1438 66 1614
rect -17 1345 17 1379
rect -17 1237 17 1271
rect -66 1002 -32 1178
rect 32 1002 66 1178
rect -17 909 17 943
rect -17 801 17 835
rect -66 566 -32 742
rect 32 566 66 742
rect -17 473 17 507
rect -17 365 17 399
rect -66 130 -32 306
rect 32 130 66 306
rect -17 37 17 71
rect -17 -71 17 -37
rect -66 -306 -32 -130
rect 32 -306 66 -130
rect -17 -399 17 -365
rect -17 -507 17 -473
rect -66 -742 -32 -566
rect 32 -742 66 -566
rect -17 -835 17 -801
rect -17 -943 17 -909
rect -66 -1178 -32 -1002
rect 32 -1178 66 -1002
rect -17 -1271 17 -1237
rect -17 -1379 17 -1345
rect -66 -1614 -32 -1438
rect 32 -1614 66 -1438
rect -17 -1707 17 -1673
rect -17 -1815 17 -1781
rect -66 -2050 -32 -1874
rect 32 -2050 66 -1874
rect -17 -2143 17 -2109
rect -17 -2251 17 -2217
rect -66 -2486 -32 -2310
rect 32 -2486 66 -2310
rect -17 -2579 17 -2545
rect -17 -2687 17 -2653
rect -66 -2922 -32 -2746
rect 32 -2922 66 -2746
rect -17 -3015 17 -2981
rect -17 -3123 17 -3089
rect -66 -3358 -32 -3182
rect 32 -3358 66 -3182
rect -17 -3451 17 -3417
rect -17 -3559 17 -3525
rect -66 -3794 -32 -3618
rect 32 -3794 66 -3618
rect -17 -3887 17 -3853
rect -17 -3995 17 -3961
rect -66 -4230 -32 -4054
rect 32 -4230 66 -4054
rect -17 -4323 17 -4289
rect -17 -4431 17 -4397
rect -66 -4666 -32 -4490
rect 32 -4666 66 -4490
rect -17 -4759 17 -4725
rect -17 -4867 17 -4833
rect -66 -5102 -32 -4926
rect 32 -5102 66 -4926
rect -17 -5195 17 -5161
rect -17 -5303 17 -5269
rect -66 -5538 -32 -5362
rect 32 -5538 66 -5362
rect -17 -5631 17 -5597
rect -17 -5739 17 -5705
rect -66 -5974 -32 -5798
rect 32 -5974 66 -5798
rect -17 -6067 17 -6033
rect -17 -6175 17 -6141
rect -66 -6410 -32 -6234
rect 32 -6410 66 -6234
rect -17 -6503 17 -6469
rect -17 -6611 17 -6577
rect -66 -6846 -32 -6670
rect 32 -6846 66 -6670
rect -17 -6939 17 -6905
rect -17 -7047 17 -7013
rect -66 -7282 -32 -7106
rect 32 -7282 66 -7106
rect -17 -7375 17 -7341
rect -17 -7483 17 -7449
rect -66 -7718 -32 -7542
rect 32 -7718 66 -7542
rect -17 -7811 17 -7777
rect -17 -7919 17 -7885
rect -66 -8154 -32 -7978
rect 32 -8154 66 -7978
rect -17 -8247 17 -8213
rect -17 -8355 17 -8321
rect -66 -8590 -32 -8414
rect 32 -8590 66 -8414
rect -17 -8683 17 -8649
rect -17 -8791 17 -8757
rect -66 -9026 -32 -8850
rect 32 -9026 66 -8850
rect -17 -9119 17 -9085
rect -17 -9227 17 -9193
rect -66 -9462 -32 -9286
rect 32 -9462 66 -9286
rect -17 -9555 17 -9521
rect -17 -9663 17 -9629
rect -66 -9898 -32 -9722
rect 32 -9898 66 -9722
rect -17 -9991 17 -9957
rect -17 -10099 17 -10065
rect -66 -10334 -32 -10158
rect 32 -10334 66 -10158
rect -17 -10427 17 -10393
rect -17 -10535 17 -10501
rect -66 -10770 -32 -10594
rect 32 -10770 66 -10594
rect -17 -10863 17 -10829
<< metal1 >>
rect -29 10863 29 10869
rect -29 10829 -17 10863
rect 17 10829 29 10863
rect -29 10823 29 10829
rect -72 10770 -26 10782
rect -72 10594 -66 10770
rect -32 10594 -26 10770
rect -72 10582 -26 10594
rect 26 10770 72 10782
rect 26 10594 32 10770
rect 66 10594 72 10770
rect 26 10582 72 10594
rect -29 10535 29 10541
rect -29 10501 -17 10535
rect 17 10501 29 10535
rect -29 10495 29 10501
rect -29 10427 29 10433
rect -29 10393 -17 10427
rect 17 10393 29 10427
rect -29 10387 29 10393
rect -72 10334 -26 10346
rect -72 10158 -66 10334
rect -32 10158 -26 10334
rect -72 10146 -26 10158
rect 26 10334 72 10346
rect 26 10158 32 10334
rect 66 10158 72 10334
rect 26 10146 72 10158
rect -29 10099 29 10105
rect -29 10065 -17 10099
rect 17 10065 29 10099
rect -29 10059 29 10065
rect -29 9991 29 9997
rect -29 9957 -17 9991
rect 17 9957 29 9991
rect -29 9951 29 9957
rect -72 9898 -26 9910
rect -72 9722 -66 9898
rect -32 9722 -26 9898
rect -72 9710 -26 9722
rect 26 9898 72 9910
rect 26 9722 32 9898
rect 66 9722 72 9898
rect 26 9710 72 9722
rect -29 9663 29 9669
rect -29 9629 -17 9663
rect 17 9629 29 9663
rect -29 9623 29 9629
rect -29 9555 29 9561
rect -29 9521 -17 9555
rect 17 9521 29 9555
rect -29 9515 29 9521
rect -72 9462 -26 9474
rect -72 9286 -66 9462
rect -32 9286 -26 9462
rect -72 9274 -26 9286
rect 26 9462 72 9474
rect 26 9286 32 9462
rect 66 9286 72 9462
rect 26 9274 72 9286
rect -29 9227 29 9233
rect -29 9193 -17 9227
rect 17 9193 29 9227
rect -29 9187 29 9193
rect -29 9119 29 9125
rect -29 9085 -17 9119
rect 17 9085 29 9119
rect -29 9079 29 9085
rect -72 9026 -26 9038
rect -72 8850 -66 9026
rect -32 8850 -26 9026
rect -72 8838 -26 8850
rect 26 9026 72 9038
rect 26 8850 32 9026
rect 66 8850 72 9026
rect 26 8838 72 8850
rect -29 8791 29 8797
rect -29 8757 -17 8791
rect 17 8757 29 8791
rect -29 8751 29 8757
rect -29 8683 29 8689
rect -29 8649 -17 8683
rect 17 8649 29 8683
rect -29 8643 29 8649
rect -72 8590 -26 8602
rect -72 8414 -66 8590
rect -32 8414 -26 8590
rect -72 8402 -26 8414
rect 26 8590 72 8602
rect 26 8414 32 8590
rect 66 8414 72 8590
rect 26 8402 72 8414
rect -29 8355 29 8361
rect -29 8321 -17 8355
rect 17 8321 29 8355
rect -29 8315 29 8321
rect -29 8247 29 8253
rect -29 8213 -17 8247
rect 17 8213 29 8247
rect -29 8207 29 8213
rect -72 8154 -26 8166
rect -72 7978 -66 8154
rect -32 7978 -26 8154
rect -72 7966 -26 7978
rect 26 8154 72 8166
rect 26 7978 32 8154
rect 66 7978 72 8154
rect 26 7966 72 7978
rect -29 7919 29 7925
rect -29 7885 -17 7919
rect 17 7885 29 7919
rect -29 7879 29 7885
rect -29 7811 29 7817
rect -29 7777 -17 7811
rect 17 7777 29 7811
rect -29 7771 29 7777
rect -72 7718 -26 7730
rect -72 7542 -66 7718
rect -32 7542 -26 7718
rect -72 7530 -26 7542
rect 26 7718 72 7730
rect 26 7542 32 7718
rect 66 7542 72 7718
rect 26 7530 72 7542
rect -29 7483 29 7489
rect -29 7449 -17 7483
rect 17 7449 29 7483
rect -29 7443 29 7449
rect -29 7375 29 7381
rect -29 7341 -17 7375
rect 17 7341 29 7375
rect -29 7335 29 7341
rect -72 7282 -26 7294
rect -72 7106 -66 7282
rect -32 7106 -26 7282
rect -72 7094 -26 7106
rect 26 7282 72 7294
rect 26 7106 32 7282
rect 66 7106 72 7282
rect 26 7094 72 7106
rect -29 7047 29 7053
rect -29 7013 -17 7047
rect 17 7013 29 7047
rect -29 7007 29 7013
rect -29 6939 29 6945
rect -29 6905 -17 6939
rect 17 6905 29 6939
rect -29 6899 29 6905
rect -72 6846 -26 6858
rect -72 6670 -66 6846
rect -32 6670 -26 6846
rect -72 6658 -26 6670
rect 26 6846 72 6858
rect 26 6670 32 6846
rect 66 6670 72 6846
rect 26 6658 72 6670
rect -29 6611 29 6617
rect -29 6577 -17 6611
rect 17 6577 29 6611
rect -29 6571 29 6577
rect -29 6503 29 6509
rect -29 6469 -17 6503
rect 17 6469 29 6503
rect -29 6463 29 6469
rect -72 6410 -26 6422
rect -72 6234 -66 6410
rect -32 6234 -26 6410
rect -72 6222 -26 6234
rect 26 6410 72 6422
rect 26 6234 32 6410
rect 66 6234 72 6410
rect 26 6222 72 6234
rect -29 6175 29 6181
rect -29 6141 -17 6175
rect 17 6141 29 6175
rect -29 6135 29 6141
rect -29 6067 29 6073
rect -29 6033 -17 6067
rect 17 6033 29 6067
rect -29 6027 29 6033
rect -72 5974 -26 5986
rect -72 5798 -66 5974
rect -32 5798 -26 5974
rect -72 5786 -26 5798
rect 26 5974 72 5986
rect 26 5798 32 5974
rect 66 5798 72 5974
rect 26 5786 72 5798
rect -29 5739 29 5745
rect -29 5705 -17 5739
rect 17 5705 29 5739
rect -29 5699 29 5705
rect -29 5631 29 5637
rect -29 5597 -17 5631
rect 17 5597 29 5631
rect -29 5591 29 5597
rect -72 5538 -26 5550
rect -72 5362 -66 5538
rect -32 5362 -26 5538
rect -72 5350 -26 5362
rect 26 5538 72 5550
rect 26 5362 32 5538
rect 66 5362 72 5538
rect 26 5350 72 5362
rect -29 5303 29 5309
rect -29 5269 -17 5303
rect 17 5269 29 5303
rect -29 5263 29 5269
rect -29 5195 29 5201
rect -29 5161 -17 5195
rect 17 5161 29 5195
rect -29 5155 29 5161
rect -72 5102 -26 5114
rect -72 4926 -66 5102
rect -32 4926 -26 5102
rect -72 4914 -26 4926
rect 26 5102 72 5114
rect 26 4926 32 5102
rect 66 4926 72 5102
rect 26 4914 72 4926
rect -29 4867 29 4873
rect -29 4833 -17 4867
rect 17 4833 29 4867
rect -29 4827 29 4833
rect -29 4759 29 4765
rect -29 4725 -17 4759
rect 17 4725 29 4759
rect -29 4719 29 4725
rect -72 4666 -26 4678
rect -72 4490 -66 4666
rect -32 4490 -26 4666
rect -72 4478 -26 4490
rect 26 4666 72 4678
rect 26 4490 32 4666
rect 66 4490 72 4666
rect 26 4478 72 4490
rect -29 4431 29 4437
rect -29 4397 -17 4431
rect 17 4397 29 4431
rect -29 4391 29 4397
rect -29 4323 29 4329
rect -29 4289 -17 4323
rect 17 4289 29 4323
rect -29 4283 29 4289
rect -72 4230 -26 4242
rect -72 4054 -66 4230
rect -32 4054 -26 4230
rect -72 4042 -26 4054
rect 26 4230 72 4242
rect 26 4054 32 4230
rect 66 4054 72 4230
rect 26 4042 72 4054
rect -29 3995 29 4001
rect -29 3961 -17 3995
rect 17 3961 29 3995
rect -29 3955 29 3961
rect -29 3887 29 3893
rect -29 3853 -17 3887
rect 17 3853 29 3887
rect -29 3847 29 3853
rect -72 3794 -26 3806
rect -72 3618 -66 3794
rect -32 3618 -26 3794
rect -72 3606 -26 3618
rect 26 3794 72 3806
rect 26 3618 32 3794
rect 66 3618 72 3794
rect 26 3606 72 3618
rect -29 3559 29 3565
rect -29 3525 -17 3559
rect 17 3525 29 3559
rect -29 3519 29 3525
rect -29 3451 29 3457
rect -29 3417 -17 3451
rect 17 3417 29 3451
rect -29 3411 29 3417
rect -72 3358 -26 3370
rect -72 3182 -66 3358
rect -32 3182 -26 3358
rect -72 3170 -26 3182
rect 26 3358 72 3370
rect 26 3182 32 3358
rect 66 3182 72 3358
rect 26 3170 72 3182
rect -29 3123 29 3129
rect -29 3089 -17 3123
rect 17 3089 29 3123
rect -29 3083 29 3089
rect -29 3015 29 3021
rect -29 2981 -17 3015
rect 17 2981 29 3015
rect -29 2975 29 2981
rect -72 2922 -26 2934
rect -72 2746 -66 2922
rect -32 2746 -26 2922
rect -72 2734 -26 2746
rect 26 2922 72 2934
rect 26 2746 32 2922
rect 66 2746 72 2922
rect 26 2734 72 2746
rect -29 2687 29 2693
rect -29 2653 -17 2687
rect 17 2653 29 2687
rect -29 2647 29 2653
rect -29 2579 29 2585
rect -29 2545 -17 2579
rect 17 2545 29 2579
rect -29 2539 29 2545
rect -72 2486 -26 2498
rect -72 2310 -66 2486
rect -32 2310 -26 2486
rect -72 2298 -26 2310
rect 26 2486 72 2498
rect 26 2310 32 2486
rect 66 2310 72 2486
rect 26 2298 72 2310
rect -29 2251 29 2257
rect -29 2217 -17 2251
rect 17 2217 29 2251
rect -29 2211 29 2217
rect -29 2143 29 2149
rect -29 2109 -17 2143
rect 17 2109 29 2143
rect -29 2103 29 2109
rect -72 2050 -26 2062
rect -72 1874 -66 2050
rect -32 1874 -26 2050
rect -72 1862 -26 1874
rect 26 2050 72 2062
rect 26 1874 32 2050
rect 66 1874 72 2050
rect 26 1862 72 1874
rect -29 1815 29 1821
rect -29 1781 -17 1815
rect 17 1781 29 1815
rect -29 1775 29 1781
rect -29 1707 29 1713
rect -29 1673 -17 1707
rect 17 1673 29 1707
rect -29 1667 29 1673
rect -72 1614 -26 1626
rect -72 1438 -66 1614
rect -32 1438 -26 1614
rect -72 1426 -26 1438
rect 26 1614 72 1626
rect 26 1438 32 1614
rect 66 1438 72 1614
rect 26 1426 72 1438
rect -29 1379 29 1385
rect -29 1345 -17 1379
rect 17 1345 29 1379
rect -29 1339 29 1345
rect -29 1271 29 1277
rect -29 1237 -17 1271
rect 17 1237 29 1271
rect -29 1231 29 1237
rect -72 1178 -26 1190
rect -72 1002 -66 1178
rect -32 1002 -26 1178
rect -72 990 -26 1002
rect 26 1178 72 1190
rect 26 1002 32 1178
rect 66 1002 72 1178
rect 26 990 72 1002
rect -29 943 29 949
rect -29 909 -17 943
rect 17 909 29 943
rect -29 903 29 909
rect -29 835 29 841
rect -29 801 -17 835
rect 17 801 29 835
rect -29 795 29 801
rect -72 742 -26 754
rect -72 566 -66 742
rect -32 566 -26 742
rect -72 554 -26 566
rect 26 742 72 754
rect 26 566 32 742
rect 66 566 72 742
rect 26 554 72 566
rect -29 507 29 513
rect -29 473 -17 507
rect 17 473 29 507
rect -29 467 29 473
rect -29 399 29 405
rect -29 365 -17 399
rect 17 365 29 399
rect -29 359 29 365
rect -72 306 -26 318
rect -72 130 -66 306
rect -32 130 -26 306
rect -72 118 -26 130
rect 26 306 72 318
rect 26 130 32 306
rect 66 130 72 306
rect 26 118 72 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -72 -130 -26 -118
rect -72 -306 -66 -130
rect -32 -306 -26 -130
rect -72 -318 -26 -306
rect 26 -130 72 -118
rect 26 -306 32 -130
rect 66 -306 72 -130
rect 26 -318 72 -306
rect -29 -365 29 -359
rect -29 -399 -17 -365
rect 17 -399 29 -365
rect -29 -405 29 -399
rect -29 -473 29 -467
rect -29 -507 -17 -473
rect 17 -507 29 -473
rect -29 -513 29 -507
rect -72 -566 -26 -554
rect -72 -742 -66 -566
rect -32 -742 -26 -566
rect -72 -754 -26 -742
rect 26 -566 72 -554
rect 26 -742 32 -566
rect 66 -742 72 -566
rect 26 -754 72 -742
rect -29 -801 29 -795
rect -29 -835 -17 -801
rect 17 -835 29 -801
rect -29 -841 29 -835
rect -29 -909 29 -903
rect -29 -943 -17 -909
rect 17 -943 29 -909
rect -29 -949 29 -943
rect -72 -1002 -26 -990
rect -72 -1178 -66 -1002
rect -32 -1178 -26 -1002
rect -72 -1190 -26 -1178
rect 26 -1002 72 -990
rect 26 -1178 32 -1002
rect 66 -1178 72 -1002
rect 26 -1190 72 -1178
rect -29 -1237 29 -1231
rect -29 -1271 -17 -1237
rect 17 -1271 29 -1237
rect -29 -1277 29 -1271
rect -29 -1345 29 -1339
rect -29 -1379 -17 -1345
rect 17 -1379 29 -1345
rect -29 -1385 29 -1379
rect -72 -1438 -26 -1426
rect -72 -1614 -66 -1438
rect -32 -1614 -26 -1438
rect -72 -1626 -26 -1614
rect 26 -1438 72 -1426
rect 26 -1614 32 -1438
rect 66 -1614 72 -1438
rect 26 -1626 72 -1614
rect -29 -1673 29 -1667
rect -29 -1707 -17 -1673
rect 17 -1707 29 -1673
rect -29 -1713 29 -1707
rect -29 -1781 29 -1775
rect -29 -1815 -17 -1781
rect 17 -1815 29 -1781
rect -29 -1821 29 -1815
rect -72 -1874 -26 -1862
rect -72 -2050 -66 -1874
rect -32 -2050 -26 -1874
rect -72 -2062 -26 -2050
rect 26 -1874 72 -1862
rect 26 -2050 32 -1874
rect 66 -2050 72 -1874
rect 26 -2062 72 -2050
rect -29 -2109 29 -2103
rect -29 -2143 -17 -2109
rect 17 -2143 29 -2109
rect -29 -2149 29 -2143
rect -29 -2217 29 -2211
rect -29 -2251 -17 -2217
rect 17 -2251 29 -2217
rect -29 -2257 29 -2251
rect -72 -2310 -26 -2298
rect -72 -2486 -66 -2310
rect -32 -2486 -26 -2310
rect -72 -2498 -26 -2486
rect 26 -2310 72 -2298
rect 26 -2486 32 -2310
rect 66 -2486 72 -2310
rect 26 -2498 72 -2486
rect -29 -2545 29 -2539
rect -29 -2579 -17 -2545
rect 17 -2579 29 -2545
rect -29 -2585 29 -2579
rect -29 -2653 29 -2647
rect -29 -2687 -17 -2653
rect 17 -2687 29 -2653
rect -29 -2693 29 -2687
rect -72 -2746 -26 -2734
rect -72 -2922 -66 -2746
rect -32 -2922 -26 -2746
rect -72 -2934 -26 -2922
rect 26 -2746 72 -2734
rect 26 -2922 32 -2746
rect 66 -2922 72 -2746
rect 26 -2934 72 -2922
rect -29 -2981 29 -2975
rect -29 -3015 -17 -2981
rect 17 -3015 29 -2981
rect -29 -3021 29 -3015
rect -29 -3089 29 -3083
rect -29 -3123 -17 -3089
rect 17 -3123 29 -3089
rect -29 -3129 29 -3123
rect -72 -3182 -26 -3170
rect -72 -3358 -66 -3182
rect -32 -3358 -26 -3182
rect -72 -3370 -26 -3358
rect 26 -3182 72 -3170
rect 26 -3358 32 -3182
rect 66 -3358 72 -3182
rect 26 -3370 72 -3358
rect -29 -3417 29 -3411
rect -29 -3451 -17 -3417
rect 17 -3451 29 -3417
rect -29 -3457 29 -3451
rect -29 -3525 29 -3519
rect -29 -3559 -17 -3525
rect 17 -3559 29 -3525
rect -29 -3565 29 -3559
rect -72 -3618 -26 -3606
rect -72 -3794 -66 -3618
rect -32 -3794 -26 -3618
rect -72 -3806 -26 -3794
rect 26 -3618 72 -3606
rect 26 -3794 32 -3618
rect 66 -3794 72 -3618
rect 26 -3806 72 -3794
rect -29 -3853 29 -3847
rect -29 -3887 -17 -3853
rect 17 -3887 29 -3853
rect -29 -3893 29 -3887
rect -29 -3961 29 -3955
rect -29 -3995 -17 -3961
rect 17 -3995 29 -3961
rect -29 -4001 29 -3995
rect -72 -4054 -26 -4042
rect -72 -4230 -66 -4054
rect -32 -4230 -26 -4054
rect -72 -4242 -26 -4230
rect 26 -4054 72 -4042
rect 26 -4230 32 -4054
rect 66 -4230 72 -4054
rect 26 -4242 72 -4230
rect -29 -4289 29 -4283
rect -29 -4323 -17 -4289
rect 17 -4323 29 -4289
rect -29 -4329 29 -4323
rect -29 -4397 29 -4391
rect -29 -4431 -17 -4397
rect 17 -4431 29 -4397
rect -29 -4437 29 -4431
rect -72 -4490 -26 -4478
rect -72 -4666 -66 -4490
rect -32 -4666 -26 -4490
rect -72 -4678 -26 -4666
rect 26 -4490 72 -4478
rect 26 -4666 32 -4490
rect 66 -4666 72 -4490
rect 26 -4678 72 -4666
rect -29 -4725 29 -4719
rect -29 -4759 -17 -4725
rect 17 -4759 29 -4725
rect -29 -4765 29 -4759
rect -29 -4833 29 -4827
rect -29 -4867 -17 -4833
rect 17 -4867 29 -4833
rect -29 -4873 29 -4867
rect -72 -4926 -26 -4914
rect -72 -5102 -66 -4926
rect -32 -5102 -26 -4926
rect -72 -5114 -26 -5102
rect 26 -4926 72 -4914
rect 26 -5102 32 -4926
rect 66 -5102 72 -4926
rect 26 -5114 72 -5102
rect -29 -5161 29 -5155
rect -29 -5195 -17 -5161
rect 17 -5195 29 -5161
rect -29 -5201 29 -5195
rect -29 -5269 29 -5263
rect -29 -5303 -17 -5269
rect 17 -5303 29 -5269
rect -29 -5309 29 -5303
rect -72 -5362 -26 -5350
rect -72 -5538 -66 -5362
rect -32 -5538 -26 -5362
rect -72 -5550 -26 -5538
rect 26 -5362 72 -5350
rect 26 -5538 32 -5362
rect 66 -5538 72 -5362
rect 26 -5550 72 -5538
rect -29 -5597 29 -5591
rect -29 -5631 -17 -5597
rect 17 -5631 29 -5597
rect -29 -5637 29 -5631
rect -29 -5705 29 -5699
rect -29 -5739 -17 -5705
rect 17 -5739 29 -5705
rect -29 -5745 29 -5739
rect -72 -5798 -26 -5786
rect -72 -5974 -66 -5798
rect -32 -5974 -26 -5798
rect -72 -5986 -26 -5974
rect 26 -5798 72 -5786
rect 26 -5974 32 -5798
rect 66 -5974 72 -5798
rect 26 -5986 72 -5974
rect -29 -6033 29 -6027
rect -29 -6067 -17 -6033
rect 17 -6067 29 -6033
rect -29 -6073 29 -6067
rect -29 -6141 29 -6135
rect -29 -6175 -17 -6141
rect 17 -6175 29 -6141
rect -29 -6181 29 -6175
rect -72 -6234 -26 -6222
rect -72 -6410 -66 -6234
rect -32 -6410 -26 -6234
rect -72 -6422 -26 -6410
rect 26 -6234 72 -6222
rect 26 -6410 32 -6234
rect 66 -6410 72 -6234
rect 26 -6422 72 -6410
rect -29 -6469 29 -6463
rect -29 -6503 -17 -6469
rect 17 -6503 29 -6469
rect -29 -6509 29 -6503
rect -29 -6577 29 -6571
rect -29 -6611 -17 -6577
rect 17 -6611 29 -6577
rect -29 -6617 29 -6611
rect -72 -6670 -26 -6658
rect -72 -6846 -66 -6670
rect -32 -6846 -26 -6670
rect -72 -6858 -26 -6846
rect 26 -6670 72 -6658
rect 26 -6846 32 -6670
rect 66 -6846 72 -6670
rect 26 -6858 72 -6846
rect -29 -6905 29 -6899
rect -29 -6939 -17 -6905
rect 17 -6939 29 -6905
rect -29 -6945 29 -6939
rect -29 -7013 29 -7007
rect -29 -7047 -17 -7013
rect 17 -7047 29 -7013
rect -29 -7053 29 -7047
rect -72 -7106 -26 -7094
rect -72 -7282 -66 -7106
rect -32 -7282 -26 -7106
rect -72 -7294 -26 -7282
rect 26 -7106 72 -7094
rect 26 -7282 32 -7106
rect 66 -7282 72 -7106
rect 26 -7294 72 -7282
rect -29 -7341 29 -7335
rect -29 -7375 -17 -7341
rect 17 -7375 29 -7341
rect -29 -7381 29 -7375
rect -29 -7449 29 -7443
rect -29 -7483 -17 -7449
rect 17 -7483 29 -7449
rect -29 -7489 29 -7483
rect -72 -7542 -26 -7530
rect -72 -7718 -66 -7542
rect -32 -7718 -26 -7542
rect -72 -7730 -26 -7718
rect 26 -7542 72 -7530
rect 26 -7718 32 -7542
rect 66 -7718 72 -7542
rect 26 -7730 72 -7718
rect -29 -7777 29 -7771
rect -29 -7811 -17 -7777
rect 17 -7811 29 -7777
rect -29 -7817 29 -7811
rect -29 -7885 29 -7879
rect -29 -7919 -17 -7885
rect 17 -7919 29 -7885
rect -29 -7925 29 -7919
rect -72 -7978 -26 -7966
rect -72 -8154 -66 -7978
rect -32 -8154 -26 -7978
rect -72 -8166 -26 -8154
rect 26 -7978 72 -7966
rect 26 -8154 32 -7978
rect 66 -8154 72 -7978
rect 26 -8166 72 -8154
rect -29 -8213 29 -8207
rect -29 -8247 -17 -8213
rect 17 -8247 29 -8213
rect -29 -8253 29 -8247
rect -29 -8321 29 -8315
rect -29 -8355 -17 -8321
rect 17 -8355 29 -8321
rect -29 -8361 29 -8355
rect -72 -8414 -26 -8402
rect -72 -8590 -66 -8414
rect -32 -8590 -26 -8414
rect -72 -8602 -26 -8590
rect 26 -8414 72 -8402
rect 26 -8590 32 -8414
rect 66 -8590 72 -8414
rect 26 -8602 72 -8590
rect -29 -8649 29 -8643
rect -29 -8683 -17 -8649
rect 17 -8683 29 -8649
rect -29 -8689 29 -8683
rect -29 -8757 29 -8751
rect -29 -8791 -17 -8757
rect 17 -8791 29 -8757
rect -29 -8797 29 -8791
rect -72 -8850 -26 -8838
rect -72 -9026 -66 -8850
rect -32 -9026 -26 -8850
rect -72 -9038 -26 -9026
rect 26 -8850 72 -8838
rect 26 -9026 32 -8850
rect 66 -9026 72 -8850
rect 26 -9038 72 -9026
rect -29 -9085 29 -9079
rect -29 -9119 -17 -9085
rect 17 -9119 29 -9085
rect -29 -9125 29 -9119
rect -29 -9193 29 -9187
rect -29 -9227 -17 -9193
rect 17 -9227 29 -9193
rect -29 -9233 29 -9227
rect -72 -9286 -26 -9274
rect -72 -9462 -66 -9286
rect -32 -9462 -26 -9286
rect -72 -9474 -26 -9462
rect 26 -9286 72 -9274
rect 26 -9462 32 -9286
rect 66 -9462 72 -9286
rect 26 -9474 72 -9462
rect -29 -9521 29 -9515
rect -29 -9555 -17 -9521
rect 17 -9555 29 -9521
rect -29 -9561 29 -9555
rect -29 -9629 29 -9623
rect -29 -9663 -17 -9629
rect 17 -9663 29 -9629
rect -29 -9669 29 -9663
rect -72 -9722 -26 -9710
rect -72 -9898 -66 -9722
rect -32 -9898 -26 -9722
rect -72 -9910 -26 -9898
rect 26 -9722 72 -9710
rect 26 -9898 32 -9722
rect 66 -9898 72 -9722
rect 26 -9910 72 -9898
rect -29 -9957 29 -9951
rect -29 -9991 -17 -9957
rect 17 -9991 29 -9957
rect -29 -9997 29 -9991
rect -29 -10065 29 -10059
rect -29 -10099 -17 -10065
rect 17 -10099 29 -10065
rect -29 -10105 29 -10099
rect -72 -10158 -26 -10146
rect -72 -10334 -66 -10158
rect -32 -10334 -26 -10158
rect -72 -10346 -26 -10334
rect 26 -10158 72 -10146
rect 26 -10334 32 -10158
rect 66 -10334 72 -10158
rect 26 -10346 72 -10334
rect -29 -10393 29 -10387
rect -29 -10427 -17 -10393
rect 17 -10427 29 -10393
rect -29 -10433 29 -10427
rect -29 -10501 29 -10495
rect -29 -10535 -17 -10501
rect 17 -10535 29 -10501
rect -29 -10541 29 -10535
rect -72 -10594 -26 -10582
rect -72 -10770 -66 -10594
rect -32 -10770 -26 -10594
rect -72 -10782 -26 -10770
rect 26 -10594 72 -10582
rect 26 -10770 32 -10594
rect 66 -10770 72 -10594
rect 26 -10782 72 -10770
rect -29 -10829 29 -10823
rect -29 -10863 -17 -10829
rect 17 -10863 29 -10829
rect -29 -10869 29 -10863
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.2 m 50 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
