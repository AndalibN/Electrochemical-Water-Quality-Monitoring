magic
tech sky130A
magscale 1 2
timestamp 1667325005
<< nmoslvt >>
rect -2411 -4950 -1871 4950
rect -1765 -4950 -1225 4950
rect -1167 -4950 -627 4950
rect -569 -4950 -29 4950
rect 29 -4950 569 4950
rect 627 -4950 1167 4950
rect 1225 -4950 1765 4950
rect 1823 -4950 2363 4950
<< ndiff >>
rect -2469 4938 -2411 4950
rect -2469 -4938 -2457 4938
rect -2423 -4938 -2411 4938
rect -2469 -4950 -2411 -4938
rect -1871 4938 -1765 4950
rect -1871 -4938 -1859 4938
rect -1781 -4938 -1765 4938
rect -1871 -4950 -1765 -4938
rect -1225 4938 -1167 4950
rect -1225 -4938 -1213 4938
rect -1179 -4938 -1167 4938
rect -1225 -4950 -1167 -4938
rect -627 4938 -569 4950
rect -627 -4938 -615 4938
rect -581 -4938 -569 4938
rect -627 -4950 -569 -4938
rect -29 4938 29 4950
rect -29 -4938 -17 4938
rect 17 -4938 29 4938
rect -29 -4950 29 -4938
rect 569 4938 627 4950
rect 569 -4938 581 4938
rect 615 -4938 627 4938
rect 569 -4950 627 -4938
rect 1167 4938 1225 4950
rect 1167 -4938 1179 4938
rect 1213 -4938 1225 4938
rect 1167 -4950 1225 -4938
rect 1765 4938 1823 4950
rect 1765 -4938 1777 4938
rect 1811 -4938 1823 4938
rect 1765 -4950 1823 -4938
rect 2363 4938 2421 4950
rect 2363 -4938 2375 4938
rect 2409 -4938 2421 4938
rect 2363 -4950 2421 -4938
<< ndiffc >>
rect -2457 -4938 -2423 4938
rect -1859 -4938 -1781 4938
rect -1213 -4938 -1179 4938
rect -615 -4938 -581 4938
rect -17 -4938 17 4938
rect 581 -4938 615 4938
rect 1179 -4938 1213 4938
rect 1777 -4938 1811 4938
rect 2375 -4938 2409 4938
<< poly >>
rect -1765 4982 -627 5038
rect -2411 4950 -1871 4982
rect -1765 4950 -1225 4982
rect -1167 4950 -627 4982
rect -569 4982 569 5038
rect -569 4950 -29 4982
rect 29 4950 569 4982
rect 627 4982 1765 5038
rect 627 4950 1167 4982
rect 1225 4950 1765 4982
rect 1823 4950 2363 5038
rect -2411 -4982 -1871 -4950
rect -1765 -4982 -1225 -4950
rect -2411 -5038 -1225 -4982
rect -1167 -4982 -627 -4950
rect -569 -4982 -29 -4950
rect -1167 -5038 -29 -4982
rect 29 -4982 569 -4950
rect 627 -4982 1167 -4950
rect 29 -5038 1167 -4982
rect 1225 -4982 1765 -4950
rect 1823 -4982 2363 -4950
rect 1225 -5038 2363 -4982
<< locali >>
rect -2457 4938 -2423 4954
rect -2457 -4954 -2423 -4938
rect -1859 4938 -1781 4954
rect -1859 -4954 -1781 -4938
rect -1213 4938 -1179 4954
rect -1213 -4954 -1179 -4938
rect -615 4938 -581 4954
rect -615 -4954 -581 -4938
rect -17 4938 17 4954
rect -17 -4954 17 -4938
rect 581 4938 615 4954
rect 581 -4954 615 -4938
rect 1179 4938 1213 4954
rect 1179 -4954 1213 -4938
rect 1777 4938 1811 4954
rect 1777 -4954 1811 -4938
rect 2375 4938 2409 4954
rect 2375 -4954 2409 -4938
<< viali >>
rect -2457 -4938 -2423 4938
rect -1859 -4938 -1781 4938
rect -1213 -4938 -1179 4938
rect -615 -4938 -581 4938
rect -17 -4938 17 4938
rect 581 -4938 615 4938
rect 1179 -4938 1213 4938
rect 1777 -4938 1811 4938
rect 2375 -4938 2409 4938
<< metal1 >>
rect -2463 4938 -2417 4950
rect -2463 -4938 -2457 4938
rect -2423 -4938 -2417 4938
rect -2463 -4950 -2417 -4938
rect -1865 4938 -1772 4950
rect -1865 -4938 -1859 4938
rect -1781 -4938 -1772 4938
rect -1865 -4950 -1772 -4938
rect -1219 4938 -1173 4950
rect -1219 -4938 -1213 4938
rect -1179 -4938 -1173 4938
rect -1219 -4950 -1173 -4938
rect -621 4938 -575 4950
rect -621 -4938 -615 4938
rect -581 -4938 -575 4938
rect -621 -4950 -575 -4938
rect -23 4938 23 4950
rect -23 -4938 -17 4938
rect 17 -4938 23 4938
rect -23 -4950 23 -4938
rect 575 4938 621 4950
rect 575 -4938 581 4938
rect 615 -4938 621 4938
rect 575 -4950 621 -4938
rect 1173 4938 1219 4950
rect 1173 -4938 1179 4938
rect 1213 -4938 1219 4938
rect 1173 -4950 1219 -4938
rect 1771 4938 1817 4950
rect 1771 -4938 1777 4938
rect 1811 -4938 1817 4938
rect 1771 -4950 1817 -4938
rect 2369 4938 2415 4950
rect 2369 -4938 2375 4938
rect 2409 -4938 2415 4938
rect 2369 -4950 2415 -4938
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 49.5 l 2.7 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
