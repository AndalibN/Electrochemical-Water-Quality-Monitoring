magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -513 -1457 513 1395
<< nmos >>
rect -429 -1431 -29 1369
rect 29 -1431 429 1369
<< ndiff >>
rect -487 1346 -429 1369
rect -487 1312 -475 1346
rect -441 1312 -429 1346
rect -487 1278 -429 1312
rect -487 1244 -475 1278
rect -441 1244 -429 1278
rect -487 1210 -429 1244
rect -487 1176 -475 1210
rect -441 1176 -429 1210
rect -487 1142 -429 1176
rect -487 1108 -475 1142
rect -441 1108 -429 1142
rect -487 1074 -429 1108
rect -487 1040 -475 1074
rect -441 1040 -429 1074
rect -487 1006 -429 1040
rect -487 972 -475 1006
rect -441 972 -429 1006
rect -487 938 -429 972
rect -487 904 -475 938
rect -441 904 -429 938
rect -487 870 -429 904
rect -487 836 -475 870
rect -441 836 -429 870
rect -487 802 -429 836
rect -487 768 -475 802
rect -441 768 -429 802
rect -487 734 -429 768
rect -487 700 -475 734
rect -441 700 -429 734
rect -487 666 -429 700
rect -487 632 -475 666
rect -441 632 -429 666
rect -487 598 -429 632
rect -487 564 -475 598
rect -441 564 -429 598
rect -487 530 -429 564
rect -487 496 -475 530
rect -441 496 -429 530
rect -487 462 -429 496
rect -487 428 -475 462
rect -441 428 -429 462
rect -487 394 -429 428
rect -487 360 -475 394
rect -441 360 -429 394
rect -487 326 -429 360
rect -487 292 -475 326
rect -441 292 -429 326
rect -487 258 -429 292
rect -487 224 -475 258
rect -441 224 -429 258
rect -487 190 -429 224
rect -487 156 -475 190
rect -441 156 -429 190
rect -487 122 -429 156
rect -487 88 -475 122
rect -441 88 -429 122
rect -487 54 -429 88
rect -487 20 -475 54
rect -441 20 -429 54
rect -487 -14 -429 20
rect -487 -48 -475 -14
rect -441 -48 -429 -14
rect -487 -82 -429 -48
rect -487 -116 -475 -82
rect -441 -116 -429 -82
rect -487 -150 -429 -116
rect -487 -184 -475 -150
rect -441 -184 -429 -150
rect -487 -218 -429 -184
rect -487 -252 -475 -218
rect -441 -252 -429 -218
rect -487 -286 -429 -252
rect -487 -320 -475 -286
rect -441 -320 -429 -286
rect -487 -354 -429 -320
rect -487 -388 -475 -354
rect -441 -388 -429 -354
rect -487 -422 -429 -388
rect -487 -456 -475 -422
rect -441 -456 -429 -422
rect -487 -490 -429 -456
rect -487 -524 -475 -490
rect -441 -524 -429 -490
rect -487 -558 -429 -524
rect -487 -592 -475 -558
rect -441 -592 -429 -558
rect -487 -626 -429 -592
rect -487 -660 -475 -626
rect -441 -660 -429 -626
rect -487 -694 -429 -660
rect -487 -728 -475 -694
rect -441 -728 -429 -694
rect -487 -762 -429 -728
rect -487 -796 -475 -762
rect -441 -796 -429 -762
rect -487 -830 -429 -796
rect -487 -864 -475 -830
rect -441 -864 -429 -830
rect -487 -898 -429 -864
rect -487 -932 -475 -898
rect -441 -932 -429 -898
rect -487 -966 -429 -932
rect -487 -1000 -475 -966
rect -441 -1000 -429 -966
rect -487 -1034 -429 -1000
rect -487 -1068 -475 -1034
rect -441 -1068 -429 -1034
rect -487 -1102 -429 -1068
rect -487 -1136 -475 -1102
rect -441 -1136 -429 -1102
rect -487 -1170 -429 -1136
rect -487 -1204 -475 -1170
rect -441 -1204 -429 -1170
rect -487 -1238 -429 -1204
rect -487 -1272 -475 -1238
rect -441 -1272 -429 -1238
rect -487 -1306 -429 -1272
rect -487 -1340 -475 -1306
rect -441 -1340 -429 -1306
rect -487 -1374 -429 -1340
rect -487 -1408 -475 -1374
rect -441 -1408 -429 -1374
rect -487 -1431 -429 -1408
rect -29 1346 29 1369
rect -29 1312 -17 1346
rect 17 1312 29 1346
rect -29 1278 29 1312
rect -29 1244 -17 1278
rect 17 1244 29 1278
rect -29 1210 29 1244
rect -29 1176 -17 1210
rect 17 1176 29 1210
rect -29 1142 29 1176
rect -29 1108 -17 1142
rect 17 1108 29 1142
rect -29 1074 29 1108
rect -29 1040 -17 1074
rect 17 1040 29 1074
rect -29 1006 29 1040
rect -29 972 -17 1006
rect 17 972 29 1006
rect -29 938 29 972
rect -29 904 -17 938
rect 17 904 29 938
rect -29 870 29 904
rect -29 836 -17 870
rect 17 836 29 870
rect -29 802 29 836
rect -29 768 -17 802
rect 17 768 29 802
rect -29 734 29 768
rect -29 700 -17 734
rect 17 700 29 734
rect -29 666 29 700
rect -29 632 -17 666
rect 17 632 29 666
rect -29 598 29 632
rect -29 564 -17 598
rect 17 564 29 598
rect -29 530 29 564
rect -29 496 -17 530
rect 17 496 29 530
rect -29 462 29 496
rect -29 428 -17 462
rect 17 428 29 462
rect -29 394 29 428
rect -29 360 -17 394
rect 17 360 29 394
rect -29 326 29 360
rect -29 292 -17 326
rect 17 292 29 326
rect -29 258 29 292
rect -29 224 -17 258
rect 17 224 29 258
rect -29 190 29 224
rect -29 156 -17 190
rect 17 156 29 190
rect -29 122 29 156
rect -29 88 -17 122
rect 17 88 29 122
rect -29 54 29 88
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -150 29 -116
rect -29 -184 -17 -150
rect 17 -184 29 -150
rect -29 -218 29 -184
rect -29 -252 -17 -218
rect 17 -252 29 -218
rect -29 -286 29 -252
rect -29 -320 -17 -286
rect 17 -320 29 -286
rect -29 -354 29 -320
rect -29 -388 -17 -354
rect 17 -388 29 -354
rect -29 -422 29 -388
rect -29 -456 -17 -422
rect 17 -456 29 -422
rect -29 -490 29 -456
rect -29 -524 -17 -490
rect 17 -524 29 -490
rect -29 -558 29 -524
rect -29 -592 -17 -558
rect 17 -592 29 -558
rect -29 -626 29 -592
rect -29 -660 -17 -626
rect 17 -660 29 -626
rect -29 -694 29 -660
rect -29 -728 -17 -694
rect 17 -728 29 -694
rect -29 -762 29 -728
rect -29 -796 -17 -762
rect 17 -796 29 -762
rect -29 -830 29 -796
rect -29 -864 -17 -830
rect 17 -864 29 -830
rect -29 -898 29 -864
rect -29 -932 -17 -898
rect 17 -932 29 -898
rect -29 -966 29 -932
rect -29 -1000 -17 -966
rect 17 -1000 29 -966
rect -29 -1034 29 -1000
rect -29 -1068 -17 -1034
rect 17 -1068 29 -1034
rect -29 -1102 29 -1068
rect -29 -1136 -17 -1102
rect 17 -1136 29 -1102
rect -29 -1170 29 -1136
rect -29 -1204 -17 -1170
rect 17 -1204 29 -1170
rect -29 -1238 29 -1204
rect -29 -1272 -17 -1238
rect 17 -1272 29 -1238
rect -29 -1306 29 -1272
rect -29 -1340 -17 -1306
rect 17 -1340 29 -1306
rect -29 -1374 29 -1340
rect -29 -1408 -17 -1374
rect 17 -1408 29 -1374
rect -29 -1431 29 -1408
rect 429 1346 487 1369
rect 429 1312 441 1346
rect 475 1312 487 1346
rect 429 1278 487 1312
rect 429 1244 441 1278
rect 475 1244 487 1278
rect 429 1210 487 1244
rect 429 1176 441 1210
rect 475 1176 487 1210
rect 429 1142 487 1176
rect 429 1108 441 1142
rect 475 1108 487 1142
rect 429 1074 487 1108
rect 429 1040 441 1074
rect 475 1040 487 1074
rect 429 1006 487 1040
rect 429 972 441 1006
rect 475 972 487 1006
rect 429 938 487 972
rect 429 904 441 938
rect 475 904 487 938
rect 429 870 487 904
rect 429 836 441 870
rect 475 836 487 870
rect 429 802 487 836
rect 429 768 441 802
rect 475 768 487 802
rect 429 734 487 768
rect 429 700 441 734
rect 475 700 487 734
rect 429 666 487 700
rect 429 632 441 666
rect 475 632 487 666
rect 429 598 487 632
rect 429 564 441 598
rect 475 564 487 598
rect 429 530 487 564
rect 429 496 441 530
rect 475 496 487 530
rect 429 462 487 496
rect 429 428 441 462
rect 475 428 487 462
rect 429 394 487 428
rect 429 360 441 394
rect 475 360 487 394
rect 429 326 487 360
rect 429 292 441 326
rect 475 292 487 326
rect 429 258 487 292
rect 429 224 441 258
rect 475 224 487 258
rect 429 190 487 224
rect 429 156 441 190
rect 475 156 487 190
rect 429 122 487 156
rect 429 88 441 122
rect 475 88 487 122
rect 429 54 487 88
rect 429 20 441 54
rect 475 20 487 54
rect 429 -14 487 20
rect 429 -48 441 -14
rect 475 -48 487 -14
rect 429 -82 487 -48
rect 429 -116 441 -82
rect 475 -116 487 -82
rect 429 -150 487 -116
rect 429 -184 441 -150
rect 475 -184 487 -150
rect 429 -218 487 -184
rect 429 -252 441 -218
rect 475 -252 487 -218
rect 429 -286 487 -252
rect 429 -320 441 -286
rect 475 -320 487 -286
rect 429 -354 487 -320
rect 429 -388 441 -354
rect 475 -388 487 -354
rect 429 -422 487 -388
rect 429 -456 441 -422
rect 475 -456 487 -422
rect 429 -490 487 -456
rect 429 -524 441 -490
rect 475 -524 487 -490
rect 429 -558 487 -524
rect 429 -592 441 -558
rect 475 -592 487 -558
rect 429 -626 487 -592
rect 429 -660 441 -626
rect 475 -660 487 -626
rect 429 -694 487 -660
rect 429 -728 441 -694
rect 475 -728 487 -694
rect 429 -762 487 -728
rect 429 -796 441 -762
rect 475 -796 487 -762
rect 429 -830 487 -796
rect 429 -864 441 -830
rect 475 -864 487 -830
rect 429 -898 487 -864
rect 429 -932 441 -898
rect 475 -932 487 -898
rect 429 -966 487 -932
rect 429 -1000 441 -966
rect 475 -1000 487 -966
rect 429 -1034 487 -1000
rect 429 -1068 441 -1034
rect 475 -1068 487 -1034
rect 429 -1102 487 -1068
rect 429 -1136 441 -1102
rect 475 -1136 487 -1102
rect 429 -1170 487 -1136
rect 429 -1204 441 -1170
rect 475 -1204 487 -1170
rect 429 -1238 487 -1204
rect 429 -1272 441 -1238
rect 475 -1272 487 -1238
rect 429 -1306 487 -1272
rect 429 -1340 441 -1306
rect 475 -1340 487 -1306
rect 429 -1374 487 -1340
rect 429 -1408 441 -1374
rect 475 -1408 487 -1374
rect 429 -1431 487 -1408
<< ndiffc >>
rect -475 1312 -441 1346
rect -475 1244 -441 1278
rect -475 1176 -441 1210
rect -475 1108 -441 1142
rect -475 1040 -441 1074
rect -475 972 -441 1006
rect -475 904 -441 938
rect -475 836 -441 870
rect -475 768 -441 802
rect -475 700 -441 734
rect -475 632 -441 666
rect -475 564 -441 598
rect -475 496 -441 530
rect -475 428 -441 462
rect -475 360 -441 394
rect -475 292 -441 326
rect -475 224 -441 258
rect -475 156 -441 190
rect -475 88 -441 122
rect -475 20 -441 54
rect -475 -48 -441 -14
rect -475 -116 -441 -82
rect -475 -184 -441 -150
rect -475 -252 -441 -218
rect -475 -320 -441 -286
rect -475 -388 -441 -354
rect -475 -456 -441 -422
rect -475 -524 -441 -490
rect -475 -592 -441 -558
rect -475 -660 -441 -626
rect -475 -728 -441 -694
rect -475 -796 -441 -762
rect -475 -864 -441 -830
rect -475 -932 -441 -898
rect -475 -1000 -441 -966
rect -475 -1068 -441 -1034
rect -475 -1136 -441 -1102
rect -475 -1204 -441 -1170
rect -475 -1272 -441 -1238
rect -475 -1340 -441 -1306
rect -475 -1408 -441 -1374
rect -17 1312 17 1346
rect -17 1244 17 1278
rect -17 1176 17 1210
rect -17 1108 17 1142
rect -17 1040 17 1074
rect -17 972 17 1006
rect -17 904 17 938
rect -17 836 17 870
rect -17 768 17 802
rect -17 700 17 734
rect -17 632 17 666
rect -17 564 17 598
rect -17 496 17 530
rect -17 428 17 462
rect -17 360 17 394
rect -17 292 17 326
rect -17 224 17 258
rect -17 156 17 190
rect -17 88 17 122
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect -17 -184 17 -150
rect -17 -252 17 -218
rect -17 -320 17 -286
rect -17 -388 17 -354
rect -17 -456 17 -422
rect -17 -524 17 -490
rect -17 -592 17 -558
rect -17 -660 17 -626
rect -17 -728 17 -694
rect -17 -796 17 -762
rect -17 -864 17 -830
rect -17 -932 17 -898
rect -17 -1000 17 -966
rect -17 -1068 17 -1034
rect -17 -1136 17 -1102
rect -17 -1204 17 -1170
rect -17 -1272 17 -1238
rect -17 -1340 17 -1306
rect -17 -1408 17 -1374
rect 441 1312 475 1346
rect 441 1244 475 1278
rect 441 1176 475 1210
rect 441 1108 475 1142
rect 441 1040 475 1074
rect 441 972 475 1006
rect 441 904 475 938
rect 441 836 475 870
rect 441 768 475 802
rect 441 700 475 734
rect 441 632 475 666
rect 441 564 475 598
rect 441 496 475 530
rect 441 428 475 462
rect 441 360 475 394
rect 441 292 475 326
rect 441 224 475 258
rect 441 156 475 190
rect 441 88 475 122
rect 441 20 475 54
rect 441 -48 475 -14
rect 441 -116 475 -82
rect 441 -184 475 -150
rect 441 -252 475 -218
rect 441 -320 475 -286
rect 441 -388 475 -354
rect 441 -456 475 -422
rect 441 -524 475 -490
rect 441 -592 475 -558
rect 441 -660 475 -626
rect 441 -728 475 -694
rect 441 -796 475 -762
rect 441 -864 475 -830
rect 441 -932 475 -898
rect 441 -1000 475 -966
rect 441 -1068 475 -1034
rect 441 -1136 475 -1102
rect 441 -1204 475 -1170
rect 441 -1272 475 -1238
rect 441 -1340 475 -1306
rect 441 -1408 475 -1374
<< poly >>
rect -429 1441 -29 1457
rect -429 1407 -382 1441
rect -348 1407 -314 1441
rect -280 1407 -246 1441
rect -212 1407 -178 1441
rect -144 1407 -110 1441
rect -76 1407 -29 1441
rect -429 1369 -29 1407
rect 29 1441 429 1457
rect 29 1407 76 1441
rect 110 1407 144 1441
rect 178 1407 212 1441
rect 246 1407 280 1441
rect 314 1407 348 1441
rect 382 1407 429 1441
rect 29 1369 429 1407
rect -429 -1457 -29 -1431
rect 29 -1457 429 -1431
<< polycont >>
rect -382 1407 -348 1441
rect -314 1407 -280 1441
rect -246 1407 -212 1441
rect -178 1407 -144 1441
rect -110 1407 -76 1441
rect 76 1407 110 1441
rect 144 1407 178 1441
rect 212 1407 246 1441
rect 280 1407 314 1441
rect 348 1407 382 1441
<< locali >>
rect -429 1407 -390 1441
rect -348 1407 -318 1441
rect -280 1407 -246 1441
rect -212 1407 -178 1441
rect -140 1407 -110 1441
rect -68 1407 -29 1441
rect 29 1407 68 1441
rect 110 1407 140 1441
rect 178 1407 212 1441
rect 246 1407 280 1441
rect 318 1407 348 1441
rect 390 1407 429 1441
rect -475 1354 -441 1373
rect -475 1282 -441 1312
rect -475 1210 -441 1244
rect -475 1142 -441 1176
rect -475 1074 -441 1104
rect -475 1006 -441 1032
rect -475 938 -441 960
rect -475 870 -441 888
rect -475 802 -441 816
rect -475 734 -441 744
rect -475 666 -441 672
rect -475 598 -441 600
rect -475 562 -441 564
rect -475 490 -441 496
rect -475 418 -441 428
rect -475 346 -441 360
rect -475 274 -441 292
rect -475 202 -441 224
rect -475 130 -441 156
rect -475 58 -441 88
rect -475 -14 -441 20
rect -475 -82 -441 -48
rect -475 -150 -441 -120
rect -475 -218 -441 -192
rect -475 -286 -441 -264
rect -475 -354 -441 -336
rect -475 -422 -441 -408
rect -475 -490 -441 -480
rect -475 -558 -441 -552
rect -475 -626 -441 -624
rect -475 -662 -441 -660
rect -475 -734 -441 -728
rect -475 -806 -441 -796
rect -475 -878 -441 -864
rect -475 -950 -441 -932
rect -475 -1022 -441 -1000
rect -475 -1094 -441 -1068
rect -475 -1166 -441 -1136
rect -475 -1238 -441 -1204
rect -475 -1306 -441 -1272
rect -475 -1374 -441 -1344
rect -475 -1435 -441 -1416
rect -17 1354 17 1373
rect -17 1282 17 1312
rect -17 1210 17 1244
rect -17 1142 17 1176
rect -17 1074 17 1104
rect -17 1006 17 1032
rect -17 938 17 960
rect -17 870 17 888
rect -17 802 17 816
rect -17 734 17 744
rect -17 666 17 672
rect -17 598 17 600
rect -17 562 17 564
rect -17 490 17 496
rect -17 418 17 428
rect -17 346 17 360
rect -17 274 17 292
rect -17 202 17 224
rect -17 130 17 156
rect -17 58 17 88
rect -17 -14 17 20
rect -17 -82 17 -48
rect -17 -150 17 -120
rect -17 -218 17 -192
rect -17 -286 17 -264
rect -17 -354 17 -336
rect -17 -422 17 -408
rect -17 -490 17 -480
rect -17 -558 17 -552
rect -17 -626 17 -624
rect -17 -662 17 -660
rect -17 -734 17 -728
rect -17 -806 17 -796
rect -17 -878 17 -864
rect -17 -950 17 -932
rect -17 -1022 17 -1000
rect -17 -1094 17 -1068
rect -17 -1166 17 -1136
rect -17 -1238 17 -1204
rect -17 -1306 17 -1272
rect -17 -1374 17 -1344
rect -17 -1435 17 -1416
rect 441 1354 475 1373
rect 441 1282 475 1312
rect 441 1210 475 1244
rect 441 1142 475 1176
rect 441 1074 475 1104
rect 441 1006 475 1032
rect 441 938 475 960
rect 441 870 475 888
rect 441 802 475 816
rect 441 734 475 744
rect 441 666 475 672
rect 441 598 475 600
rect 441 562 475 564
rect 441 490 475 496
rect 441 418 475 428
rect 441 346 475 360
rect 441 274 475 292
rect 441 202 475 224
rect 441 130 475 156
rect 441 58 475 88
rect 441 -14 475 20
rect 441 -82 475 -48
rect 441 -150 475 -120
rect 441 -218 475 -192
rect 441 -286 475 -264
rect 441 -354 475 -336
rect 441 -422 475 -408
rect 441 -490 475 -480
rect 441 -558 475 -552
rect 441 -626 475 -624
rect 441 -662 475 -660
rect 441 -734 475 -728
rect 441 -806 475 -796
rect 441 -878 475 -864
rect 441 -950 475 -932
rect 441 -1022 475 -1000
rect 441 -1094 475 -1068
rect 441 -1166 475 -1136
rect 441 -1238 475 -1204
rect 441 -1306 475 -1272
rect 441 -1374 475 -1344
rect 441 -1435 475 -1416
<< viali >>
rect -390 1407 -382 1441
rect -382 1407 -356 1441
rect -318 1407 -314 1441
rect -314 1407 -284 1441
rect -246 1407 -212 1441
rect -174 1407 -144 1441
rect -144 1407 -140 1441
rect -102 1407 -76 1441
rect -76 1407 -68 1441
rect 68 1407 76 1441
rect 76 1407 102 1441
rect 140 1407 144 1441
rect 144 1407 174 1441
rect 212 1407 246 1441
rect 284 1407 314 1441
rect 314 1407 318 1441
rect 356 1407 382 1441
rect 382 1407 390 1441
rect -475 1346 -441 1354
rect -475 1320 -441 1346
rect -475 1278 -441 1282
rect -475 1248 -441 1278
rect -475 1176 -441 1210
rect -475 1108 -441 1138
rect -475 1104 -441 1108
rect -475 1040 -441 1066
rect -475 1032 -441 1040
rect -475 972 -441 994
rect -475 960 -441 972
rect -475 904 -441 922
rect -475 888 -441 904
rect -475 836 -441 850
rect -475 816 -441 836
rect -475 768 -441 778
rect -475 744 -441 768
rect -475 700 -441 706
rect -475 672 -441 700
rect -475 632 -441 634
rect -475 600 -441 632
rect -475 530 -441 562
rect -475 528 -441 530
rect -475 462 -441 490
rect -475 456 -441 462
rect -475 394 -441 418
rect -475 384 -441 394
rect -475 326 -441 346
rect -475 312 -441 326
rect -475 258 -441 274
rect -475 240 -441 258
rect -475 190 -441 202
rect -475 168 -441 190
rect -475 122 -441 130
rect -475 96 -441 122
rect -475 54 -441 58
rect -475 24 -441 54
rect -475 -48 -441 -14
rect -475 -116 -441 -86
rect -475 -120 -441 -116
rect -475 -184 -441 -158
rect -475 -192 -441 -184
rect -475 -252 -441 -230
rect -475 -264 -441 -252
rect -475 -320 -441 -302
rect -475 -336 -441 -320
rect -475 -388 -441 -374
rect -475 -408 -441 -388
rect -475 -456 -441 -446
rect -475 -480 -441 -456
rect -475 -524 -441 -518
rect -475 -552 -441 -524
rect -475 -592 -441 -590
rect -475 -624 -441 -592
rect -475 -694 -441 -662
rect -475 -696 -441 -694
rect -475 -762 -441 -734
rect -475 -768 -441 -762
rect -475 -830 -441 -806
rect -475 -840 -441 -830
rect -475 -898 -441 -878
rect -475 -912 -441 -898
rect -475 -966 -441 -950
rect -475 -984 -441 -966
rect -475 -1034 -441 -1022
rect -475 -1056 -441 -1034
rect -475 -1102 -441 -1094
rect -475 -1128 -441 -1102
rect -475 -1170 -441 -1166
rect -475 -1200 -441 -1170
rect -475 -1272 -441 -1238
rect -475 -1340 -441 -1310
rect -475 -1344 -441 -1340
rect -475 -1408 -441 -1382
rect -475 -1416 -441 -1408
rect -17 1346 17 1354
rect -17 1320 17 1346
rect -17 1278 17 1282
rect -17 1248 17 1278
rect -17 1176 17 1210
rect -17 1108 17 1138
rect -17 1104 17 1108
rect -17 1040 17 1066
rect -17 1032 17 1040
rect -17 972 17 994
rect -17 960 17 972
rect -17 904 17 922
rect -17 888 17 904
rect -17 836 17 850
rect -17 816 17 836
rect -17 768 17 778
rect -17 744 17 768
rect -17 700 17 706
rect -17 672 17 700
rect -17 632 17 634
rect -17 600 17 632
rect -17 530 17 562
rect -17 528 17 530
rect -17 462 17 490
rect -17 456 17 462
rect -17 394 17 418
rect -17 384 17 394
rect -17 326 17 346
rect -17 312 17 326
rect -17 258 17 274
rect -17 240 17 258
rect -17 190 17 202
rect -17 168 17 190
rect -17 122 17 130
rect -17 96 17 122
rect -17 54 17 58
rect -17 24 17 54
rect -17 -48 17 -14
rect -17 -116 17 -86
rect -17 -120 17 -116
rect -17 -184 17 -158
rect -17 -192 17 -184
rect -17 -252 17 -230
rect -17 -264 17 -252
rect -17 -320 17 -302
rect -17 -336 17 -320
rect -17 -388 17 -374
rect -17 -408 17 -388
rect -17 -456 17 -446
rect -17 -480 17 -456
rect -17 -524 17 -518
rect -17 -552 17 -524
rect -17 -592 17 -590
rect -17 -624 17 -592
rect -17 -694 17 -662
rect -17 -696 17 -694
rect -17 -762 17 -734
rect -17 -768 17 -762
rect -17 -830 17 -806
rect -17 -840 17 -830
rect -17 -898 17 -878
rect -17 -912 17 -898
rect -17 -966 17 -950
rect -17 -984 17 -966
rect -17 -1034 17 -1022
rect -17 -1056 17 -1034
rect -17 -1102 17 -1094
rect -17 -1128 17 -1102
rect -17 -1170 17 -1166
rect -17 -1200 17 -1170
rect -17 -1272 17 -1238
rect -17 -1340 17 -1310
rect -17 -1344 17 -1340
rect -17 -1408 17 -1382
rect -17 -1416 17 -1408
rect 441 1346 475 1354
rect 441 1320 475 1346
rect 441 1278 475 1282
rect 441 1248 475 1278
rect 441 1176 475 1210
rect 441 1108 475 1138
rect 441 1104 475 1108
rect 441 1040 475 1066
rect 441 1032 475 1040
rect 441 972 475 994
rect 441 960 475 972
rect 441 904 475 922
rect 441 888 475 904
rect 441 836 475 850
rect 441 816 475 836
rect 441 768 475 778
rect 441 744 475 768
rect 441 700 475 706
rect 441 672 475 700
rect 441 632 475 634
rect 441 600 475 632
rect 441 530 475 562
rect 441 528 475 530
rect 441 462 475 490
rect 441 456 475 462
rect 441 394 475 418
rect 441 384 475 394
rect 441 326 475 346
rect 441 312 475 326
rect 441 258 475 274
rect 441 240 475 258
rect 441 190 475 202
rect 441 168 475 190
rect 441 122 475 130
rect 441 96 475 122
rect 441 54 475 58
rect 441 24 475 54
rect 441 -48 475 -14
rect 441 -116 475 -86
rect 441 -120 475 -116
rect 441 -184 475 -158
rect 441 -192 475 -184
rect 441 -252 475 -230
rect 441 -264 475 -252
rect 441 -320 475 -302
rect 441 -336 475 -320
rect 441 -388 475 -374
rect 441 -408 475 -388
rect 441 -456 475 -446
rect 441 -480 475 -456
rect 441 -524 475 -518
rect 441 -552 475 -524
rect 441 -592 475 -590
rect 441 -624 475 -592
rect 441 -694 475 -662
rect 441 -696 475 -694
rect 441 -762 475 -734
rect 441 -768 475 -762
rect 441 -830 475 -806
rect 441 -840 475 -830
rect 441 -898 475 -878
rect 441 -912 475 -898
rect 441 -966 475 -950
rect 441 -984 475 -966
rect 441 -1034 475 -1022
rect 441 -1056 475 -1034
rect 441 -1102 475 -1094
rect 441 -1128 475 -1102
rect 441 -1170 475 -1166
rect 441 -1200 475 -1170
rect 441 -1272 475 -1238
rect 441 -1340 475 -1310
rect 441 -1344 475 -1340
rect 441 -1408 475 -1382
rect 441 -1416 475 -1408
<< metal1 >>
rect -425 1441 -33 1447
rect -425 1407 -390 1441
rect -356 1407 -318 1441
rect -284 1407 -246 1441
rect -212 1407 -174 1441
rect -140 1407 -102 1441
rect -68 1407 -33 1441
rect -425 1401 -33 1407
rect 33 1441 425 1447
rect 33 1407 68 1441
rect 102 1407 140 1441
rect 174 1407 212 1441
rect 246 1407 284 1441
rect 318 1407 356 1441
rect 390 1407 425 1441
rect 33 1401 425 1407
rect -481 1354 -435 1369
rect -481 1320 -475 1354
rect -441 1320 -435 1354
rect -481 1282 -435 1320
rect -481 1248 -475 1282
rect -441 1248 -435 1282
rect -481 1210 -435 1248
rect -481 1176 -475 1210
rect -441 1176 -435 1210
rect -481 1138 -435 1176
rect -481 1104 -475 1138
rect -441 1104 -435 1138
rect -481 1066 -435 1104
rect -481 1032 -475 1066
rect -441 1032 -435 1066
rect -481 994 -435 1032
rect -481 960 -475 994
rect -441 960 -435 994
rect -481 922 -435 960
rect -481 888 -475 922
rect -441 888 -435 922
rect -481 850 -435 888
rect -481 816 -475 850
rect -441 816 -435 850
rect -481 778 -435 816
rect -481 744 -475 778
rect -441 744 -435 778
rect -481 706 -435 744
rect -481 672 -475 706
rect -441 672 -435 706
rect -481 634 -435 672
rect -481 600 -475 634
rect -441 600 -435 634
rect -481 562 -435 600
rect -481 528 -475 562
rect -441 528 -435 562
rect -481 490 -435 528
rect -481 456 -475 490
rect -441 456 -435 490
rect -481 418 -435 456
rect -481 384 -475 418
rect -441 384 -435 418
rect -481 346 -435 384
rect -481 312 -475 346
rect -441 312 -435 346
rect -481 274 -435 312
rect -481 240 -475 274
rect -441 240 -435 274
rect -481 202 -435 240
rect -481 168 -475 202
rect -441 168 -435 202
rect -481 130 -435 168
rect -481 96 -475 130
rect -441 96 -435 130
rect -481 58 -435 96
rect -481 24 -475 58
rect -441 24 -435 58
rect -481 -14 -435 24
rect -481 -48 -475 -14
rect -441 -48 -435 -14
rect -481 -86 -435 -48
rect -481 -120 -475 -86
rect -441 -120 -435 -86
rect -481 -158 -435 -120
rect -481 -192 -475 -158
rect -441 -192 -435 -158
rect -481 -230 -435 -192
rect -481 -264 -475 -230
rect -441 -264 -435 -230
rect -481 -302 -435 -264
rect -481 -336 -475 -302
rect -441 -336 -435 -302
rect -481 -374 -435 -336
rect -481 -408 -475 -374
rect -441 -408 -435 -374
rect -481 -446 -435 -408
rect -481 -480 -475 -446
rect -441 -480 -435 -446
rect -481 -518 -435 -480
rect -481 -552 -475 -518
rect -441 -552 -435 -518
rect -481 -590 -435 -552
rect -481 -624 -475 -590
rect -441 -624 -435 -590
rect -481 -662 -435 -624
rect -481 -696 -475 -662
rect -441 -696 -435 -662
rect -481 -734 -435 -696
rect -481 -768 -475 -734
rect -441 -768 -435 -734
rect -481 -806 -435 -768
rect -481 -840 -475 -806
rect -441 -840 -435 -806
rect -481 -878 -435 -840
rect -481 -912 -475 -878
rect -441 -912 -435 -878
rect -481 -950 -435 -912
rect -481 -984 -475 -950
rect -441 -984 -435 -950
rect -481 -1022 -435 -984
rect -481 -1056 -475 -1022
rect -441 -1056 -435 -1022
rect -481 -1094 -435 -1056
rect -481 -1128 -475 -1094
rect -441 -1128 -435 -1094
rect -481 -1166 -435 -1128
rect -481 -1200 -475 -1166
rect -441 -1200 -435 -1166
rect -481 -1238 -435 -1200
rect -481 -1272 -475 -1238
rect -441 -1272 -435 -1238
rect -481 -1310 -435 -1272
rect -481 -1344 -475 -1310
rect -441 -1344 -435 -1310
rect -481 -1382 -435 -1344
rect -481 -1416 -475 -1382
rect -441 -1416 -435 -1382
rect -481 -1431 -435 -1416
rect -23 1354 23 1369
rect -23 1320 -17 1354
rect 17 1320 23 1354
rect -23 1282 23 1320
rect -23 1248 -17 1282
rect 17 1248 23 1282
rect -23 1210 23 1248
rect -23 1176 -17 1210
rect 17 1176 23 1210
rect -23 1138 23 1176
rect -23 1104 -17 1138
rect 17 1104 23 1138
rect -23 1066 23 1104
rect -23 1032 -17 1066
rect 17 1032 23 1066
rect -23 994 23 1032
rect -23 960 -17 994
rect 17 960 23 994
rect -23 922 23 960
rect -23 888 -17 922
rect 17 888 23 922
rect -23 850 23 888
rect -23 816 -17 850
rect 17 816 23 850
rect -23 778 23 816
rect -23 744 -17 778
rect 17 744 23 778
rect -23 706 23 744
rect -23 672 -17 706
rect 17 672 23 706
rect -23 634 23 672
rect -23 600 -17 634
rect 17 600 23 634
rect -23 562 23 600
rect -23 528 -17 562
rect 17 528 23 562
rect -23 490 23 528
rect -23 456 -17 490
rect 17 456 23 490
rect -23 418 23 456
rect -23 384 -17 418
rect 17 384 23 418
rect -23 346 23 384
rect -23 312 -17 346
rect 17 312 23 346
rect -23 274 23 312
rect -23 240 -17 274
rect 17 240 23 274
rect -23 202 23 240
rect -23 168 -17 202
rect 17 168 23 202
rect -23 130 23 168
rect -23 96 -17 130
rect 17 96 23 130
rect -23 58 23 96
rect -23 24 -17 58
rect 17 24 23 58
rect -23 -14 23 24
rect -23 -48 -17 -14
rect 17 -48 23 -14
rect -23 -86 23 -48
rect -23 -120 -17 -86
rect 17 -120 23 -86
rect -23 -158 23 -120
rect -23 -192 -17 -158
rect 17 -192 23 -158
rect -23 -230 23 -192
rect -23 -264 -17 -230
rect 17 -264 23 -230
rect -23 -302 23 -264
rect -23 -336 -17 -302
rect 17 -336 23 -302
rect -23 -374 23 -336
rect -23 -408 -17 -374
rect 17 -408 23 -374
rect -23 -446 23 -408
rect -23 -480 -17 -446
rect 17 -480 23 -446
rect -23 -518 23 -480
rect -23 -552 -17 -518
rect 17 -552 23 -518
rect -23 -590 23 -552
rect -23 -624 -17 -590
rect 17 -624 23 -590
rect -23 -662 23 -624
rect -23 -696 -17 -662
rect 17 -696 23 -662
rect -23 -734 23 -696
rect -23 -768 -17 -734
rect 17 -768 23 -734
rect -23 -806 23 -768
rect -23 -840 -17 -806
rect 17 -840 23 -806
rect -23 -878 23 -840
rect -23 -912 -17 -878
rect 17 -912 23 -878
rect -23 -950 23 -912
rect -23 -984 -17 -950
rect 17 -984 23 -950
rect -23 -1022 23 -984
rect -23 -1056 -17 -1022
rect 17 -1056 23 -1022
rect -23 -1094 23 -1056
rect -23 -1128 -17 -1094
rect 17 -1128 23 -1094
rect -23 -1166 23 -1128
rect -23 -1200 -17 -1166
rect 17 -1200 23 -1166
rect -23 -1238 23 -1200
rect -23 -1272 -17 -1238
rect 17 -1272 23 -1238
rect -23 -1310 23 -1272
rect -23 -1344 -17 -1310
rect 17 -1344 23 -1310
rect -23 -1382 23 -1344
rect -23 -1416 -17 -1382
rect 17 -1416 23 -1382
rect -23 -1431 23 -1416
rect 435 1354 481 1369
rect 435 1320 441 1354
rect 475 1320 481 1354
rect 435 1282 481 1320
rect 435 1248 441 1282
rect 475 1248 481 1282
rect 435 1210 481 1248
rect 435 1176 441 1210
rect 475 1176 481 1210
rect 435 1138 481 1176
rect 435 1104 441 1138
rect 475 1104 481 1138
rect 435 1066 481 1104
rect 435 1032 441 1066
rect 475 1032 481 1066
rect 435 994 481 1032
rect 435 960 441 994
rect 475 960 481 994
rect 435 922 481 960
rect 435 888 441 922
rect 475 888 481 922
rect 435 850 481 888
rect 435 816 441 850
rect 475 816 481 850
rect 435 778 481 816
rect 435 744 441 778
rect 475 744 481 778
rect 435 706 481 744
rect 435 672 441 706
rect 475 672 481 706
rect 435 634 481 672
rect 435 600 441 634
rect 475 600 481 634
rect 435 562 481 600
rect 435 528 441 562
rect 475 528 481 562
rect 435 490 481 528
rect 435 456 441 490
rect 475 456 481 490
rect 435 418 481 456
rect 435 384 441 418
rect 475 384 481 418
rect 435 346 481 384
rect 435 312 441 346
rect 475 312 481 346
rect 435 274 481 312
rect 435 240 441 274
rect 475 240 481 274
rect 435 202 481 240
rect 435 168 441 202
rect 475 168 481 202
rect 435 130 481 168
rect 435 96 441 130
rect 475 96 481 130
rect 435 58 481 96
rect 435 24 441 58
rect 475 24 481 58
rect 435 -14 481 24
rect 435 -48 441 -14
rect 475 -48 481 -14
rect 435 -86 481 -48
rect 435 -120 441 -86
rect 475 -120 481 -86
rect 435 -158 481 -120
rect 435 -192 441 -158
rect 475 -192 481 -158
rect 435 -230 481 -192
rect 435 -264 441 -230
rect 475 -264 481 -230
rect 435 -302 481 -264
rect 435 -336 441 -302
rect 475 -336 481 -302
rect 435 -374 481 -336
rect 435 -408 441 -374
rect 475 -408 481 -374
rect 435 -446 481 -408
rect 435 -480 441 -446
rect 475 -480 481 -446
rect 435 -518 481 -480
rect 435 -552 441 -518
rect 475 -552 481 -518
rect 435 -590 481 -552
rect 435 -624 441 -590
rect 475 -624 481 -590
rect 435 -662 481 -624
rect 435 -696 441 -662
rect 475 -696 481 -662
rect 435 -734 481 -696
rect 435 -768 441 -734
rect 475 -768 481 -734
rect 435 -806 481 -768
rect 435 -840 441 -806
rect 475 -840 481 -806
rect 435 -878 481 -840
rect 435 -912 441 -878
rect 475 -912 481 -878
rect 435 -950 481 -912
rect 435 -984 441 -950
rect 475 -984 481 -950
rect 435 -1022 481 -984
rect 435 -1056 441 -1022
rect 475 -1056 481 -1022
rect 435 -1094 481 -1056
rect 435 -1128 441 -1094
rect 475 -1128 481 -1094
rect 435 -1166 481 -1128
rect 435 -1200 441 -1166
rect 475 -1200 481 -1166
rect 435 -1238 481 -1200
rect 435 -1272 441 -1238
rect 475 -1272 481 -1238
rect 435 -1310 481 -1272
rect 435 -1344 441 -1310
rect 475 -1344 481 -1310
rect 435 -1382 481 -1344
rect 435 -1416 441 -1382
rect 475 -1416 481 -1382
rect 435 -1431 481 -1416
<< end >>
