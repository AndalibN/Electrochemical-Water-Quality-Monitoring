magic
tech sky130A
magscale 1 2
timestamp 1667400309
<< xpolycontact >>
rect -35 1265 35 1697
rect -35 -1697 35 -1265
<< xpolyres >>
rect -35 -1265 35 1265
<< viali >>
rect -19 1282 19 1679
rect -19 -1679 19 -1282
<< metal1 >>
rect -25 1679 25 1691
rect -25 1282 -19 1679
rect 19 1282 25 1679
rect -25 1270 25 1282
rect -25 -1282 25 -1270
rect -25 -1679 -19 -1282
rect 19 -1679 25 -1282
rect -25 -1691 25 -1679
<< res0p35 >>
rect -37 -1267 37 1267
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 12.65 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 73.361k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
