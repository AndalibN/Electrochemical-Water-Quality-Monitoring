magic
tech sky130A
magscale 1 2
timestamp 1667411791
<< error_p >>
rect -941 18143 -883 18149
rect -749 18143 -691 18149
rect -557 18143 -499 18149
rect -365 18143 -307 18149
rect -173 18143 -115 18149
rect 19 18143 77 18149
rect 211 18143 269 18149
rect 403 18143 461 18149
rect 595 18143 653 18149
rect 787 18143 845 18149
rect -941 18109 -929 18143
rect -749 18109 -737 18143
rect -557 18109 -545 18143
rect -365 18109 -353 18143
rect -173 18109 -161 18143
rect 19 18109 31 18143
rect 211 18109 223 18143
rect 403 18109 415 18143
rect 595 18109 607 18143
rect 787 18109 799 18143
rect -941 18103 -883 18109
rect -749 18103 -691 18109
rect -557 18103 -499 18109
rect -365 18103 -307 18109
rect -173 18103 -115 18109
rect 19 18103 77 18109
rect 211 18103 269 18109
rect 403 18103 461 18109
rect 595 18103 653 18109
rect 787 18103 845 18109
rect -1025 14600 1025 14780
rect -929 14562 1025 14600
rect -845 14507 -787 14513
rect -653 14507 -595 14513
rect -461 14507 -403 14513
rect -269 14507 -211 14513
rect -77 14507 -19 14513
rect 115 14507 173 14513
rect 307 14507 365 14513
rect 499 14507 557 14513
rect 691 14507 749 14513
rect 883 14507 941 14513
rect -845 14473 -833 14507
rect -653 14473 -641 14507
rect -461 14473 -449 14507
rect -269 14473 -257 14507
rect -77 14473 -65 14507
rect 115 14473 127 14507
rect 307 14473 319 14507
rect 499 14473 511 14507
rect 691 14473 703 14507
rect 883 14473 895 14507
rect -845 14467 -787 14473
rect -653 14467 -595 14473
rect -461 14467 -403 14473
rect -269 14467 -211 14473
rect -77 14467 -19 14473
rect 115 14467 173 14473
rect 307 14467 365 14473
rect 499 14467 557 14473
rect 691 14467 749 14473
rect 883 14467 941 14473
rect -1025 10964 1025 11144
rect -1025 10926 929 10964
rect -941 10871 -883 10877
rect -749 10871 -691 10877
rect -557 10871 -499 10877
rect -365 10871 -307 10877
rect -173 10871 -115 10877
rect 19 10871 77 10877
rect 211 10871 269 10877
rect 403 10871 461 10877
rect 595 10871 653 10877
rect 787 10871 845 10877
rect -941 10837 -929 10871
rect -749 10837 -737 10871
rect -557 10837 -545 10871
rect -365 10837 -353 10871
rect -173 10837 -161 10871
rect 19 10837 31 10871
rect 211 10837 223 10871
rect 403 10837 415 10871
rect 595 10837 607 10871
rect 787 10837 799 10871
rect -941 10831 -883 10837
rect -749 10831 -691 10837
rect -557 10831 -499 10837
rect -365 10831 -307 10837
rect -173 10831 -115 10837
rect 19 10831 77 10837
rect 211 10831 269 10837
rect 403 10831 461 10837
rect 595 10831 653 10837
rect 787 10831 845 10837
rect -1025 7328 1025 7508
rect -929 7290 1025 7328
rect -845 7235 -787 7241
rect -653 7235 -595 7241
rect -461 7235 -403 7241
rect -269 7235 -211 7241
rect -77 7235 -19 7241
rect 115 7235 173 7241
rect 307 7235 365 7241
rect 499 7235 557 7241
rect 691 7235 749 7241
rect 883 7235 941 7241
rect -845 7201 -833 7235
rect -653 7201 -641 7235
rect -461 7201 -449 7235
rect -269 7201 -257 7235
rect -77 7201 -65 7235
rect 115 7201 127 7235
rect 307 7201 319 7235
rect 499 7201 511 7235
rect 691 7201 703 7235
rect 883 7201 895 7235
rect -845 7195 -787 7201
rect -653 7195 -595 7201
rect -461 7195 -403 7201
rect -269 7195 -211 7201
rect -77 7195 -19 7201
rect 115 7195 173 7201
rect 307 7195 365 7201
rect 499 7195 557 7201
rect 691 7195 749 7201
rect 883 7195 941 7201
rect -1025 3692 1025 3872
rect -1025 3654 929 3692
rect -941 3599 -883 3605
rect -749 3599 -691 3605
rect -557 3599 -499 3605
rect -365 3599 -307 3605
rect -173 3599 -115 3605
rect 19 3599 77 3605
rect 211 3599 269 3605
rect 403 3599 461 3605
rect 595 3599 653 3605
rect 787 3599 845 3605
rect -941 3565 -929 3599
rect -749 3565 -737 3599
rect -557 3565 -545 3599
rect -365 3565 -353 3599
rect -173 3565 -161 3599
rect 19 3565 31 3599
rect 211 3565 223 3599
rect 403 3565 415 3599
rect 595 3565 607 3599
rect 787 3565 799 3599
rect -941 3559 -883 3565
rect -749 3559 -691 3565
rect -557 3559 -499 3565
rect -365 3559 -307 3565
rect -173 3559 -115 3565
rect 19 3559 77 3565
rect 211 3559 269 3565
rect 403 3559 461 3565
rect 595 3559 653 3565
rect 787 3559 845 3565
rect -1025 56 1025 236
rect -929 18 1025 56
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect -1025 -3580 1025 -3400
rect -1025 -3618 929 -3580
rect -941 -3673 -883 -3667
rect -749 -3673 -691 -3667
rect -557 -3673 -499 -3667
rect -365 -3673 -307 -3667
rect -173 -3673 -115 -3667
rect 19 -3673 77 -3667
rect 211 -3673 269 -3667
rect 403 -3673 461 -3667
rect 595 -3673 653 -3667
rect 787 -3673 845 -3667
rect -941 -3707 -929 -3673
rect -749 -3707 -737 -3673
rect -557 -3707 -545 -3673
rect -365 -3707 -353 -3673
rect -173 -3707 -161 -3673
rect 19 -3707 31 -3673
rect 211 -3707 223 -3673
rect 403 -3707 415 -3673
rect 595 -3707 607 -3673
rect 787 -3707 799 -3673
rect -941 -3713 -883 -3707
rect -749 -3713 -691 -3707
rect -557 -3713 -499 -3707
rect -365 -3713 -307 -3707
rect -173 -3713 -115 -3707
rect 19 -3713 77 -3707
rect 211 -3713 269 -3707
rect 403 -3713 461 -3707
rect 595 -3713 653 -3707
rect 787 -3713 845 -3707
rect -1025 -7216 1025 -7036
rect -929 -7254 1025 -7216
rect -845 -7309 -787 -7303
rect -653 -7309 -595 -7303
rect -461 -7309 -403 -7303
rect -269 -7309 -211 -7303
rect -77 -7309 -19 -7303
rect 115 -7309 173 -7303
rect 307 -7309 365 -7303
rect 499 -7309 557 -7303
rect 691 -7309 749 -7303
rect 883 -7309 941 -7303
rect -845 -7343 -833 -7309
rect -653 -7343 -641 -7309
rect -461 -7343 -449 -7309
rect -269 -7343 -257 -7309
rect -77 -7343 -65 -7309
rect 115 -7343 127 -7309
rect 307 -7343 319 -7309
rect 499 -7343 511 -7309
rect 691 -7343 703 -7309
rect 883 -7343 895 -7309
rect -845 -7349 -787 -7343
rect -653 -7349 -595 -7343
rect -461 -7349 -403 -7343
rect -269 -7349 -211 -7343
rect -77 -7349 -19 -7343
rect 115 -7349 173 -7343
rect 307 -7349 365 -7343
rect 499 -7349 557 -7343
rect 691 -7349 749 -7343
rect 883 -7349 941 -7343
rect -1025 -10852 1025 -10672
rect -1025 -10890 929 -10852
rect -941 -10945 -883 -10939
rect -749 -10945 -691 -10939
rect -557 -10945 -499 -10939
rect -365 -10945 -307 -10939
rect -173 -10945 -115 -10939
rect 19 -10945 77 -10939
rect 211 -10945 269 -10939
rect 403 -10945 461 -10939
rect 595 -10945 653 -10939
rect 787 -10945 845 -10939
rect -941 -10979 -929 -10945
rect -749 -10979 -737 -10945
rect -557 -10979 -545 -10945
rect -365 -10979 -353 -10945
rect -173 -10979 -161 -10945
rect 19 -10979 31 -10945
rect 211 -10979 223 -10945
rect 403 -10979 415 -10945
rect 595 -10979 607 -10945
rect 787 -10979 799 -10945
rect -941 -10985 -883 -10979
rect -749 -10985 -691 -10979
rect -557 -10985 -499 -10979
rect -365 -10985 -307 -10979
rect -173 -10985 -115 -10979
rect 19 -10985 77 -10979
rect 211 -10985 269 -10979
rect 403 -10985 461 -10979
rect 595 -10985 653 -10979
rect 787 -10985 845 -10979
rect -1025 -14488 1025 -14308
rect -929 -14526 1025 -14488
rect -845 -14581 -787 -14575
rect -653 -14581 -595 -14575
rect -461 -14581 -403 -14575
rect -269 -14581 -211 -14575
rect -77 -14581 -19 -14575
rect 115 -14581 173 -14575
rect 307 -14581 365 -14575
rect 499 -14581 557 -14575
rect 691 -14581 749 -14575
rect 883 -14581 941 -14575
rect -845 -14615 -833 -14581
rect -653 -14615 -641 -14581
rect -461 -14615 -449 -14581
rect -269 -14615 -257 -14581
rect -77 -14615 -65 -14581
rect 115 -14615 127 -14581
rect 307 -14615 319 -14581
rect 499 -14615 511 -14581
rect 691 -14615 703 -14581
rect 883 -14615 895 -14581
rect -845 -14621 -787 -14615
rect -653 -14621 -595 -14615
rect -461 -14621 -403 -14615
rect -269 -14621 -211 -14615
rect -77 -14621 -19 -14615
rect 115 -14621 173 -14615
rect 307 -14621 365 -14615
rect 499 -14621 557 -14615
rect 691 -14621 749 -14615
rect 883 -14621 941 -14615
rect -941 -18109 -883 -18103
rect -749 -18109 -691 -18103
rect -557 -18109 -499 -18103
rect -365 -18109 -307 -18103
rect -173 -18109 -115 -18103
rect 19 -18109 77 -18103
rect 211 -18109 269 -18103
rect 403 -18109 461 -18103
rect 595 -18109 653 -18103
rect 787 -18109 845 -18103
rect -941 -18143 -929 -18109
rect -749 -18143 -737 -18109
rect -557 -18143 -545 -18109
rect -365 -18143 -353 -18109
rect -173 -18143 -161 -18109
rect 19 -18143 31 -18109
rect 211 -18143 223 -18109
rect 403 -18143 415 -18109
rect 595 -18143 607 -18109
rect 787 -18143 799 -18109
rect -941 -18149 -883 -18143
rect -749 -18149 -691 -18143
rect -557 -18149 -499 -18143
rect -365 -18149 -307 -18143
rect -173 -18149 -115 -18143
rect 19 -18149 77 -18143
rect 211 -18149 269 -18143
rect 403 -18149 461 -18143
rect 595 -18149 653 -18143
rect 787 -18149 845 -18143
<< nwell >>
rect -1025 18124 929 18162
rect -1025 14600 1025 18124
rect -929 14562 1025 14600
rect -929 14488 1025 14526
rect -1025 10964 1025 14488
rect -1025 10926 929 10964
rect -1025 10852 929 10890
rect -1025 7328 1025 10852
rect -929 7290 1025 7328
rect -929 7216 1025 7254
rect -1025 3692 1025 7216
rect -1025 3654 929 3692
rect -1025 3580 929 3618
rect -1025 56 1025 3580
rect -929 18 1025 56
rect -929 -56 1025 -18
rect -1025 -3580 1025 -56
rect -1025 -3618 929 -3580
rect -1025 -3692 929 -3654
rect -1025 -7216 1025 -3692
rect -929 -7254 1025 -7216
rect -929 -7328 1025 -7290
rect -1025 -10852 1025 -7328
rect -1025 -10890 929 -10852
rect -1025 -10964 929 -10926
rect -1025 -14488 1025 -10964
rect -929 -14526 1025 -14488
rect -929 -14600 1025 -14562
rect -1025 -18124 1025 -14600
rect -1025 -18162 929 -18124
<< pmos >>
rect -927 14662 -897 18062
rect -831 14662 -801 18062
rect -735 14662 -705 18062
rect -639 14662 -609 18062
rect -543 14662 -513 18062
rect -447 14662 -417 18062
rect -351 14662 -321 18062
rect -255 14662 -225 18062
rect -159 14662 -129 18062
rect -63 14662 -33 18062
rect 33 14662 63 18062
rect 129 14662 159 18062
rect 225 14662 255 18062
rect 321 14662 351 18062
rect 417 14662 447 18062
rect 513 14662 543 18062
rect 609 14662 639 18062
rect 705 14662 735 18062
rect 801 14662 831 18062
rect 897 14662 927 18062
rect -927 11026 -897 14426
rect -831 11026 -801 14426
rect -735 11026 -705 14426
rect -639 11026 -609 14426
rect -543 11026 -513 14426
rect -447 11026 -417 14426
rect -351 11026 -321 14426
rect -255 11026 -225 14426
rect -159 11026 -129 14426
rect -63 11026 -33 14426
rect 33 11026 63 14426
rect 129 11026 159 14426
rect 225 11026 255 14426
rect 321 11026 351 14426
rect 417 11026 447 14426
rect 513 11026 543 14426
rect 609 11026 639 14426
rect 705 11026 735 14426
rect 801 11026 831 14426
rect 897 11026 927 14426
rect -927 7390 -897 10790
rect -831 7390 -801 10790
rect -735 7390 -705 10790
rect -639 7390 -609 10790
rect -543 7390 -513 10790
rect -447 7390 -417 10790
rect -351 7390 -321 10790
rect -255 7390 -225 10790
rect -159 7390 -129 10790
rect -63 7390 -33 10790
rect 33 7390 63 10790
rect 129 7390 159 10790
rect 225 7390 255 10790
rect 321 7390 351 10790
rect 417 7390 447 10790
rect 513 7390 543 10790
rect 609 7390 639 10790
rect 705 7390 735 10790
rect 801 7390 831 10790
rect 897 7390 927 10790
rect -927 3754 -897 7154
rect -831 3754 -801 7154
rect -735 3754 -705 7154
rect -639 3754 -609 7154
rect -543 3754 -513 7154
rect -447 3754 -417 7154
rect -351 3754 -321 7154
rect -255 3754 -225 7154
rect -159 3754 -129 7154
rect -63 3754 -33 7154
rect 33 3754 63 7154
rect 129 3754 159 7154
rect 225 3754 255 7154
rect 321 3754 351 7154
rect 417 3754 447 7154
rect 513 3754 543 7154
rect 609 3754 639 7154
rect 705 3754 735 7154
rect 801 3754 831 7154
rect 897 3754 927 7154
rect -927 118 -897 3518
rect -831 118 -801 3518
rect -735 118 -705 3518
rect -639 118 -609 3518
rect -543 118 -513 3518
rect -447 118 -417 3518
rect -351 118 -321 3518
rect -255 118 -225 3518
rect -159 118 -129 3518
rect -63 118 -33 3518
rect 33 118 63 3518
rect 129 118 159 3518
rect 225 118 255 3518
rect 321 118 351 3518
rect 417 118 447 3518
rect 513 118 543 3518
rect 609 118 639 3518
rect 705 118 735 3518
rect 801 118 831 3518
rect 897 118 927 3518
rect -927 -3518 -897 -118
rect -831 -3518 -801 -118
rect -735 -3518 -705 -118
rect -639 -3518 -609 -118
rect -543 -3518 -513 -118
rect -447 -3518 -417 -118
rect -351 -3518 -321 -118
rect -255 -3518 -225 -118
rect -159 -3518 -129 -118
rect -63 -3518 -33 -118
rect 33 -3518 63 -118
rect 129 -3518 159 -118
rect 225 -3518 255 -118
rect 321 -3518 351 -118
rect 417 -3518 447 -118
rect 513 -3518 543 -118
rect 609 -3518 639 -118
rect 705 -3518 735 -118
rect 801 -3518 831 -118
rect 897 -3518 927 -118
rect -927 -7154 -897 -3754
rect -831 -7154 -801 -3754
rect -735 -7154 -705 -3754
rect -639 -7154 -609 -3754
rect -543 -7154 -513 -3754
rect -447 -7154 -417 -3754
rect -351 -7154 -321 -3754
rect -255 -7154 -225 -3754
rect -159 -7154 -129 -3754
rect -63 -7154 -33 -3754
rect 33 -7154 63 -3754
rect 129 -7154 159 -3754
rect 225 -7154 255 -3754
rect 321 -7154 351 -3754
rect 417 -7154 447 -3754
rect 513 -7154 543 -3754
rect 609 -7154 639 -3754
rect 705 -7154 735 -3754
rect 801 -7154 831 -3754
rect 897 -7154 927 -3754
rect -927 -10790 -897 -7390
rect -831 -10790 -801 -7390
rect -735 -10790 -705 -7390
rect -639 -10790 -609 -7390
rect -543 -10790 -513 -7390
rect -447 -10790 -417 -7390
rect -351 -10790 -321 -7390
rect -255 -10790 -225 -7390
rect -159 -10790 -129 -7390
rect -63 -10790 -33 -7390
rect 33 -10790 63 -7390
rect 129 -10790 159 -7390
rect 225 -10790 255 -7390
rect 321 -10790 351 -7390
rect 417 -10790 447 -7390
rect 513 -10790 543 -7390
rect 609 -10790 639 -7390
rect 705 -10790 735 -7390
rect 801 -10790 831 -7390
rect 897 -10790 927 -7390
rect -927 -14426 -897 -11026
rect -831 -14426 -801 -11026
rect -735 -14426 -705 -11026
rect -639 -14426 -609 -11026
rect -543 -14426 -513 -11026
rect -447 -14426 -417 -11026
rect -351 -14426 -321 -11026
rect -255 -14426 -225 -11026
rect -159 -14426 -129 -11026
rect -63 -14426 -33 -11026
rect 33 -14426 63 -11026
rect 129 -14426 159 -11026
rect 225 -14426 255 -11026
rect 321 -14426 351 -11026
rect 417 -14426 447 -11026
rect 513 -14426 543 -11026
rect 609 -14426 639 -11026
rect 705 -14426 735 -11026
rect 801 -14426 831 -11026
rect 897 -14426 927 -11026
rect -927 -18062 -897 -14662
rect -831 -18062 -801 -14662
rect -735 -18062 -705 -14662
rect -639 -18062 -609 -14662
rect -543 -18062 -513 -14662
rect -447 -18062 -417 -14662
rect -351 -18062 -321 -14662
rect -255 -18062 -225 -14662
rect -159 -18062 -129 -14662
rect -63 -18062 -33 -14662
rect 33 -18062 63 -14662
rect 129 -18062 159 -14662
rect 225 -18062 255 -14662
rect 321 -18062 351 -14662
rect 417 -18062 447 -14662
rect 513 -18062 543 -14662
rect 609 -18062 639 -14662
rect 705 -18062 735 -14662
rect 801 -18062 831 -14662
rect 897 -18062 927 -14662
<< pdiff >>
rect -989 18050 -927 18062
rect -989 14674 -977 18050
rect -943 14674 -927 18050
rect -989 14662 -927 14674
rect -897 18050 -831 18062
rect -897 14674 -881 18050
rect -847 14674 -831 18050
rect -897 14662 -831 14674
rect -801 18050 -735 18062
rect -801 14674 -785 18050
rect -751 14674 -735 18050
rect -801 14662 -735 14674
rect -705 18050 -639 18062
rect -705 14674 -689 18050
rect -655 14674 -639 18050
rect -705 14662 -639 14674
rect -609 18050 -543 18062
rect -609 14674 -593 18050
rect -559 14674 -543 18050
rect -609 14662 -543 14674
rect -513 18050 -447 18062
rect -513 14674 -497 18050
rect -463 14674 -447 18050
rect -513 14662 -447 14674
rect -417 18050 -351 18062
rect -417 14674 -401 18050
rect -367 14674 -351 18050
rect -417 14662 -351 14674
rect -321 18050 -255 18062
rect -321 14674 -305 18050
rect -271 14674 -255 18050
rect -321 14662 -255 14674
rect -225 18050 -159 18062
rect -225 14674 -209 18050
rect -175 14674 -159 18050
rect -225 14662 -159 14674
rect -129 18050 -63 18062
rect -129 14674 -113 18050
rect -79 14674 -63 18050
rect -129 14662 -63 14674
rect -33 18050 33 18062
rect -33 14674 -17 18050
rect 17 14674 33 18050
rect -33 14662 33 14674
rect 63 18050 129 18062
rect 63 14674 79 18050
rect 113 14674 129 18050
rect 63 14662 129 14674
rect 159 18050 225 18062
rect 159 14674 175 18050
rect 209 14674 225 18050
rect 159 14662 225 14674
rect 255 18050 321 18062
rect 255 14674 271 18050
rect 305 14674 321 18050
rect 255 14662 321 14674
rect 351 18050 417 18062
rect 351 14674 367 18050
rect 401 14674 417 18050
rect 351 14662 417 14674
rect 447 18050 513 18062
rect 447 14674 463 18050
rect 497 14674 513 18050
rect 447 14662 513 14674
rect 543 18050 609 18062
rect 543 14674 559 18050
rect 593 14674 609 18050
rect 543 14662 609 14674
rect 639 18050 705 18062
rect 639 14674 655 18050
rect 689 14674 705 18050
rect 639 14662 705 14674
rect 735 18050 801 18062
rect 735 14674 751 18050
rect 785 14674 801 18050
rect 735 14662 801 14674
rect 831 18050 897 18062
rect 831 14674 847 18050
rect 881 14674 897 18050
rect 831 14662 897 14674
rect 927 18050 989 18062
rect 927 14674 943 18050
rect 977 14674 989 18050
rect 927 14662 989 14674
rect -989 14414 -927 14426
rect -989 11038 -977 14414
rect -943 11038 -927 14414
rect -989 11026 -927 11038
rect -897 14414 -831 14426
rect -897 11038 -881 14414
rect -847 11038 -831 14414
rect -897 11026 -831 11038
rect -801 14414 -735 14426
rect -801 11038 -785 14414
rect -751 11038 -735 14414
rect -801 11026 -735 11038
rect -705 14414 -639 14426
rect -705 11038 -689 14414
rect -655 11038 -639 14414
rect -705 11026 -639 11038
rect -609 14414 -543 14426
rect -609 11038 -593 14414
rect -559 11038 -543 14414
rect -609 11026 -543 11038
rect -513 14414 -447 14426
rect -513 11038 -497 14414
rect -463 11038 -447 14414
rect -513 11026 -447 11038
rect -417 14414 -351 14426
rect -417 11038 -401 14414
rect -367 11038 -351 14414
rect -417 11026 -351 11038
rect -321 14414 -255 14426
rect -321 11038 -305 14414
rect -271 11038 -255 14414
rect -321 11026 -255 11038
rect -225 14414 -159 14426
rect -225 11038 -209 14414
rect -175 11038 -159 14414
rect -225 11026 -159 11038
rect -129 14414 -63 14426
rect -129 11038 -113 14414
rect -79 11038 -63 14414
rect -129 11026 -63 11038
rect -33 14414 33 14426
rect -33 11038 -17 14414
rect 17 11038 33 14414
rect -33 11026 33 11038
rect 63 14414 129 14426
rect 63 11038 79 14414
rect 113 11038 129 14414
rect 63 11026 129 11038
rect 159 14414 225 14426
rect 159 11038 175 14414
rect 209 11038 225 14414
rect 159 11026 225 11038
rect 255 14414 321 14426
rect 255 11038 271 14414
rect 305 11038 321 14414
rect 255 11026 321 11038
rect 351 14414 417 14426
rect 351 11038 367 14414
rect 401 11038 417 14414
rect 351 11026 417 11038
rect 447 14414 513 14426
rect 447 11038 463 14414
rect 497 11038 513 14414
rect 447 11026 513 11038
rect 543 14414 609 14426
rect 543 11038 559 14414
rect 593 11038 609 14414
rect 543 11026 609 11038
rect 639 14414 705 14426
rect 639 11038 655 14414
rect 689 11038 705 14414
rect 639 11026 705 11038
rect 735 14414 801 14426
rect 735 11038 751 14414
rect 785 11038 801 14414
rect 735 11026 801 11038
rect 831 14414 897 14426
rect 831 11038 847 14414
rect 881 11038 897 14414
rect 831 11026 897 11038
rect 927 14414 989 14426
rect 927 11038 943 14414
rect 977 11038 989 14414
rect 927 11026 989 11038
rect -989 10778 -927 10790
rect -989 7402 -977 10778
rect -943 7402 -927 10778
rect -989 7390 -927 7402
rect -897 10778 -831 10790
rect -897 7402 -881 10778
rect -847 7402 -831 10778
rect -897 7390 -831 7402
rect -801 10778 -735 10790
rect -801 7402 -785 10778
rect -751 7402 -735 10778
rect -801 7390 -735 7402
rect -705 10778 -639 10790
rect -705 7402 -689 10778
rect -655 7402 -639 10778
rect -705 7390 -639 7402
rect -609 10778 -543 10790
rect -609 7402 -593 10778
rect -559 7402 -543 10778
rect -609 7390 -543 7402
rect -513 10778 -447 10790
rect -513 7402 -497 10778
rect -463 7402 -447 10778
rect -513 7390 -447 7402
rect -417 10778 -351 10790
rect -417 7402 -401 10778
rect -367 7402 -351 10778
rect -417 7390 -351 7402
rect -321 10778 -255 10790
rect -321 7402 -305 10778
rect -271 7402 -255 10778
rect -321 7390 -255 7402
rect -225 10778 -159 10790
rect -225 7402 -209 10778
rect -175 7402 -159 10778
rect -225 7390 -159 7402
rect -129 10778 -63 10790
rect -129 7402 -113 10778
rect -79 7402 -63 10778
rect -129 7390 -63 7402
rect -33 10778 33 10790
rect -33 7402 -17 10778
rect 17 7402 33 10778
rect -33 7390 33 7402
rect 63 10778 129 10790
rect 63 7402 79 10778
rect 113 7402 129 10778
rect 63 7390 129 7402
rect 159 10778 225 10790
rect 159 7402 175 10778
rect 209 7402 225 10778
rect 159 7390 225 7402
rect 255 10778 321 10790
rect 255 7402 271 10778
rect 305 7402 321 10778
rect 255 7390 321 7402
rect 351 10778 417 10790
rect 351 7402 367 10778
rect 401 7402 417 10778
rect 351 7390 417 7402
rect 447 10778 513 10790
rect 447 7402 463 10778
rect 497 7402 513 10778
rect 447 7390 513 7402
rect 543 10778 609 10790
rect 543 7402 559 10778
rect 593 7402 609 10778
rect 543 7390 609 7402
rect 639 10778 705 10790
rect 639 7402 655 10778
rect 689 7402 705 10778
rect 639 7390 705 7402
rect 735 10778 801 10790
rect 735 7402 751 10778
rect 785 7402 801 10778
rect 735 7390 801 7402
rect 831 10778 897 10790
rect 831 7402 847 10778
rect 881 7402 897 10778
rect 831 7390 897 7402
rect 927 10778 989 10790
rect 927 7402 943 10778
rect 977 7402 989 10778
rect 927 7390 989 7402
rect -989 7142 -927 7154
rect -989 3766 -977 7142
rect -943 3766 -927 7142
rect -989 3754 -927 3766
rect -897 7142 -831 7154
rect -897 3766 -881 7142
rect -847 3766 -831 7142
rect -897 3754 -831 3766
rect -801 7142 -735 7154
rect -801 3766 -785 7142
rect -751 3766 -735 7142
rect -801 3754 -735 3766
rect -705 7142 -639 7154
rect -705 3766 -689 7142
rect -655 3766 -639 7142
rect -705 3754 -639 3766
rect -609 7142 -543 7154
rect -609 3766 -593 7142
rect -559 3766 -543 7142
rect -609 3754 -543 3766
rect -513 7142 -447 7154
rect -513 3766 -497 7142
rect -463 3766 -447 7142
rect -513 3754 -447 3766
rect -417 7142 -351 7154
rect -417 3766 -401 7142
rect -367 3766 -351 7142
rect -417 3754 -351 3766
rect -321 7142 -255 7154
rect -321 3766 -305 7142
rect -271 3766 -255 7142
rect -321 3754 -255 3766
rect -225 7142 -159 7154
rect -225 3766 -209 7142
rect -175 3766 -159 7142
rect -225 3754 -159 3766
rect -129 7142 -63 7154
rect -129 3766 -113 7142
rect -79 3766 -63 7142
rect -129 3754 -63 3766
rect -33 7142 33 7154
rect -33 3766 -17 7142
rect 17 3766 33 7142
rect -33 3754 33 3766
rect 63 7142 129 7154
rect 63 3766 79 7142
rect 113 3766 129 7142
rect 63 3754 129 3766
rect 159 7142 225 7154
rect 159 3766 175 7142
rect 209 3766 225 7142
rect 159 3754 225 3766
rect 255 7142 321 7154
rect 255 3766 271 7142
rect 305 3766 321 7142
rect 255 3754 321 3766
rect 351 7142 417 7154
rect 351 3766 367 7142
rect 401 3766 417 7142
rect 351 3754 417 3766
rect 447 7142 513 7154
rect 447 3766 463 7142
rect 497 3766 513 7142
rect 447 3754 513 3766
rect 543 7142 609 7154
rect 543 3766 559 7142
rect 593 3766 609 7142
rect 543 3754 609 3766
rect 639 7142 705 7154
rect 639 3766 655 7142
rect 689 3766 705 7142
rect 639 3754 705 3766
rect 735 7142 801 7154
rect 735 3766 751 7142
rect 785 3766 801 7142
rect 735 3754 801 3766
rect 831 7142 897 7154
rect 831 3766 847 7142
rect 881 3766 897 7142
rect 831 3754 897 3766
rect 927 7142 989 7154
rect 927 3766 943 7142
rect 977 3766 989 7142
rect 927 3754 989 3766
rect -989 3506 -927 3518
rect -989 130 -977 3506
rect -943 130 -927 3506
rect -989 118 -927 130
rect -897 3506 -831 3518
rect -897 130 -881 3506
rect -847 130 -831 3506
rect -897 118 -831 130
rect -801 3506 -735 3518
rect -801 130 -785 3506
rect -751 130 -735 3506
rect -801 118 -735 130
rect -705 3506 -639 3518
rect -705 130 -689 3506
rect -655 130 -639 3506
rect -705 118 -639 130
rect -609 3506 -543 3518
rect -609 130 -593 3506
rect -559 130 -543 3506
rect -609 118 -543 130
rect -513 3506 -447 3518
rect -513 130 -497 3506
rect -463 130 -447 3506
rect -513 118 -447 130
rect -417 3506 -351 3518
rect -417 130 -401 3506
rect -367 130 -351 3506
rect -417 118 -351 130
rect -321 3506 -255 3518
rect -321 130 -305 3506
rect -271 130 -255 3506
rect -321 118 -255 130
rect -225 3506 -159 3518
rect -225 130 -209 3506
rect -175 130 -159 3506
rect -225 118 -159 130
rect -129 3506 -63 3518
rect -129 130 -113 3506
rect -79 130 -63 3506
rect -129 118 -63 130
rect -33 3506 33 3518
rect -33 130 -17 3506
rect 17 130 33 3506
rect -33 118 33 130
rect 63 3506 129 3518
rect 63 130 79 3506
rect 113 130 129 3506
rect 63 118 129 130
rect 159 3506 225 3518
rect 159 130 175 3506
rect 209 130 225 3506
rect 159 118 225 130
rect 255 3506 321 3518
rect 255 130 271 3506
rect 305 130 321 3506
rect 255 118 321 130
rect 351 3506 417 3518
rect 351 130 367 3506
rect 401 130 417 3506
rect 351 118 417 130
rect 447 3506 513 3518
rect 447 130 463 3506
rect 497 130 513 3506
rect 447 118 513 130
rect 543 3506 609 3518
rect 543 130 559 3506
rect 593 130 609 3506
rect 543 118 609 130
rect 639 3506 705 3518
rect 639 130 655 3506
rect 689 130 705 3506
rect 639 118 705 130
rect 735 3506 801 3518
rect 735 130 751 3506
rect 785 130 801 3506
rect 735 118 801 130
rect 831 3506 897 3518
rect 831 130 847 3506
rect 881 130 897 3506
rect 831 118 897 130
rect 927 3506 989 3518
rect 927 130 943 3506
rect 977 130 989 3506
rect 927 118 989 130
rect -989 -130 -927 -118
rect -989 -3506 -977 -130
rect -943 -3506 -927 -130
rect -989 -3518 -927 -3506
rect -897 -130 -831 -118
rect -897 -3506 -881 -130
rect -847 -3506 -831 -130
rect -897 -3518 -831 -3506
rect -801 -130 -735 -118
rect -801 -3506 -785 -130
rect -751 -3506 -735 -130
rect -801 -3518 -735 -3506
rect -705 -130 -639 -118
rect -705 -3506 -689 -130
rect -655 -3506 -639 -130
rect -705 -3518 -639 -3506
rect -609 -130 -543 -118
rect -609 -3506 -593 -130
rect -559 -3506 -543 -130
rect -609 -3518 -543 -3506
rect -513 -130 -447 -118
rect -513 -3506 -497 -130
rect -463 -3506 -447 -130
rect -513 -3518 -447 -3506
rect -417 -130 -351 -118
rect -417 -3506 -401 -130
rect -367 -3506 -351 -130
rect -417 -3518 -351 -3506
rect -321 -130 -255 -118
rect -321 -3506 -305 -130
rect -271 -3506 -255 -130
rect -321 -3518 -255 -3506
rect -225 -130 -159 -118
rect -225 -3506 -209 -130
rect -175 -3506 -159 -130
rect -225 -3518 -159 -3506
rect -129 -130 -63 -118
rect -129 -3506 -113 -130
rect -79 -3506 -63 -130
rect -129 -3518 -63 -3506
rect -33 -130 33 -118
rect -33 -3506 -17 -130
rect 17 -3506 33 -130
rect -33 -3518 33 -3506
rect 63 -130 129 -118
rect 63 -3506 79 -130
rect 113 -3506 129 -130
rect 63 -3518 129 -3506
rect 159 -130 225 -118
rect 159 -3506 175 -130
rect 209 -3506 225 -130
rect 159 -3518 225 -3506
rect 255 -130 321 -118
rect 255 -3506 271 -130
rect 305 -3506 321 -130
rect 255 -3518 321 -3506
rect 351 -130 417 -118
rect 351 -3506 367 -130
rect 401 -3506 417 -130
rect 351 -3518 417 -3506
rect 447 -130 513 -118
rect 447 -3506 463 -130
rect 497 -3506 513 -130
rect 447 -3518 513 -3506
rect 543 -130 609 -118
rect 543 -3506 559 -130
rect 593 -3506 609 -130
rect 543 -3518 609 -3506
rect 639 -130 705 -118
rect 639 -3506 655 -130
rect 689 -3506 705 -130
rect 639 -3518 705 -3506
rect 735 -130 801 -118
rect 735 -3506 751 -130
rect 785 -3506 801 -130
rect 735 -3518 801 -3506
rect 831 -130 897 -118
rect 831 -3506 847 -130
rect 881 -3506 897 -130
rect 831 -3518 897 -3506
rect 927 -130 989 -118
rect 927 -3506 943 -130
rect 977 -3506 989 -130
rect 927 -3518 989 -3506
rect -989 -3766 -927 -3754
rect -989 -7142 -977 -3766
rect -943 -7142 -927 -3766
rect -989 -7154 -927 -7142
rect -897 -3766 -831 -3754
rect -897 -7142 -881 -3766
rect -847 -7142 -831 -3766
rect -897 -7154 -831 -7142
rect -801 -3766 -735 -3754
rect -801 -7142 -785 -3766
rect -751 -7142 -735 -3766
rect -801 -7154 -735 -7142
rect -705 -3766 -639 -3754
rect -705 -7142 -689 -3766
rect -655 -7142 -639 -3766
rect -705 -7154 -639 -7142
rect -609 -3766 -543 -3754
rect -609 -7142 -593 -3766
rect -559 -7142 -543 -3766
rect -609 -7154 -543 -7142
rect -513 -3766 -447 -3754
rect -513 -7142 -497 -3766
rect -463 -7142 -447 -3766
rect -513 -7154 -447 -7142
rect -417 -3766 -351 -3754
rect -417 -7142 -401 -3766
rect -367 -7142 -351 -3766
rect -417 -7154 -351 -7142
rect -321 -3766 -255 -3754
rect -321 -7142 -305 -3766
rect -271 -7142 -255 -3766
rect -321 -7154 -255 -7142
rect -225 -3766 -159 -3754
rect -225 -7142 -209 -3766
rect -175 -7142 -159 -3766
rect -225 -7154 -159 -7142
rect -129 -3766 -63 -3754
rect -129 -7142 -113 -3766
rect -79 -7142 -63 -3766
rect -129 -7154 -63 -7142
rect -33 -3766 33 -3754
rect -33 -7142 -17 -3766
rect 17 -7142 33 -3766
rect -33 -7154 33 -7142
rect 63 -3766 129 -3754
rect 63 -7142 79 -3766
rect 113 -7142 129 -3766
rect 63 -7154 129 -7142
rect 159 -3766 225 -3754
rect 159 -7142 175 -3766
rect 209 -7142 225 -3766
rect 159 -7154 225 -7142
rect 255 -3766 321 -3754
rect 255 -7142 271 -3766
rect 305 -7142 321 -3766
rect 255 -7154 321 -7142
rect 351 -3766 417 -3754
rect 351 -7142 367 -3766
rect 401 -7142 417 -3766
rect 351 -7154 417 -7142
rect 447 -3766 513 -3754
rect 447 -7142 463 -3766
rect 497 -7142 513 -3766
rect 447 -7154 513 -7142
rect 543 -3766 609 -3754
rect 543 -7142 559 -3766
rect 593 -7142 609 -3766
rect 543 -7154 609 -7142
rect 639 -3766 705 -3754
rect 639 -7142 655 -3766
rect 689 -7142 705 -3766
rect 639 -7154 705 -7142
rect 735 -3766 801 -3754
rect 735 -7142 751 -3766
rect 785 -7142 801 -3766
rect 735 -7154 801 -7142
rect 831 -3766 897 -3754
rect 831 -7142 847 -3766
rect 881 -7142 897 -3766
rect 831 -7154 897 -7142
rect 927 -3766 989 -3754
rect 927 -7142 943 -3766
rect 977 -7142 989 -3766
rect 927 -7154 989 -7142
rect -989 -7402 -927 -7390
rect -989 -10778 -977 -7402
rect -943 -10778 -927 -7402
rect -989 -10790 -927 -10778
rect -897 -7402 -831 -7390
rect -897 -10778 -881 -7402
rect -847 -10778 -831 -7402
rect -897 -10790 -831 -10778
rect -801 -7402 -735 -7390
rect -801 -10778 -785 -7402
rect -751 -10778 -735 -7402
rect -801 -10790 -735 -10778
rect -705 -7402 -639 -7390
rect -705 -10778 -689 -7402
rect -655 -10778 -639 -7402
rect -705 -10790 -639 -10778
rect -609 -7402 -543 -7390
rect -609 -10778 -593 -7402
rect -559 -10778 -543 -7402
rect -609 -10790 -543 -10778
rect -513 -7402 -447 -7390
rect -513 -10778 -497 -7402
rect -463 -10778 -447 -7402
rect -513 -10790 -447 -10778
rect -417 -7402 -351 -7390
rect -417 -10778 -401 -7402
rect -367 -10778 -351 -7402
rect -417 -10790 -351 -10778
rect -321 -7402 -255 -7390
rect -321 -10778 -305 -7402
rect -271 -10778 -255 -7402
rect -321 -10790 -255 -10778
rect -225 -7402 -159 -7390
rect -225 -10778 -209 -7402
rect -175 -10778 -159 -7402
rect -225 -10790 -159 -10778
rect -129 -7402 -63 -7390
rect -129 -10778 -113 -7402
rect -79 -10778 -63 -7402
rect -129 -10790 -63 -10778
rect -33 -7402 33 -7390
rect -33 -10778 -17 -7402
rect 17 -10778 33 -7402
rect -33 -10790 33 -10778
rect 63 -7402 129 -7390
rect 63 -10778 79 -7402
rect 113 -10778 129 -7402
rect 63 -10790 129 -10778
rect 159 -7402 225 -7390
rect 159 -10778 175 -7402
rect 209 -10778 225 -7402
rect 159 -10790 225 -10778
rect 255 -7402 321 -7390
rect 255 -10778 271 -7402
rect 305 -10778 321 -7402
rect 255 -10790 321 -10778
rect 351 -7402 417 -7390
rect 351 -10778 367 -7402
rect 401 -10778 417 -7402
rect 351 -10790 417 -10778
rect 447 -7402 513 -7390
rect 447 -10778 463 -7402
rect 497 -10778 513 -7402
rect 447 -10790 513 -10778
rect 543 -7402 609 -7390
rect 543 -10778 559 -7402
rect 593 -10778 609 -7402
rect 543 -10790 609 -10778
rect 639 -7402 705 -7390
rect 639 -10778 655 -7402
rect 689 -10778 705 -7402
rect 639 -10790 705 -10778
rect 735 -7402 801 -7390
rect 735 -10778 751 -7402
rect 785 -10778 801 -7402
rect 735 -10790 801 -10778
rect 831 -7402 897 -7390
rect 831 -10778 847 -7402
rect 881 -10778 897 -7402
rect 831 -10790 897 -10778
rect 927 -7402 989 -7390
rect 927 -10778 943 -7402
rect 977 -10778 989 -7402
rect 927 -10790 989 -10778
rect -989 -11038 -927 -11026
rect -989 -14414 -977 -11038
rect -943 -14414 -927 -11038
rect -989 -14426 -927 -14414
rect -897 -11038 -831 -11026
rect -897 -14414 -881 -11038
rect -847 -14414 -831 -11038
rect -897 -14426 -831 -14414
rect -801 -11038 -735 -11026
rect -801 -14414 -785 -11038
rect -751 -14414 -735 -11038
rect -801 -14426 -735 -14414
rect -705 -11038 -639 -11026
rect -705 -14414 -689 -11038
rect -655 -14414 -639 -11038
rect -705 -14426 -639 -14414
rect -609 -11038 -543 -11026
rect -609 -14414 -593 -11038
rect -559 -14414 -543 -11038
rect -609 -14426 -543 -14414
rect -513 -11038 -447 -11026
rect -513 -14414 -497 -11038
rect -463 -14414 -447 -11038
rect -513 -14426 -447 -14414
rect -417 -11038 -351 -11026
rect -417 -14414 -401 -11038
rect -367 -14414 -351 -11038
rect -417 -14426 -351 -14414
rect -321 -11038 -255 -11026
rect -321 -14414 -305 -11038
rect -271 -14414 -255 -11038
rect -321 -14426 -255 -14414
rect -225 -11038 -159 -11026
rect -225 -14414 -209 -11038
rect -175 -14414 -159 -11038
rect -225 -14426 -159 -14414
rect -129 -11038 -63 -11026
rect -129 -14414 -113 -11038
rect -79 -14414 -63 -11038
rect -129 -14426 -63 -14414
rect -33 -11038 33 -11026
rect -33 -14414 -17 -11038
rect 17 -14414 33 -11038
rect -33 -14426 33 -14414
rect 63 -11038 129 -11026
rect 63 -14414 79 -11038
rect 113 -14414 129 -11038
rect 63 -14426 129 -14414
rect 159 -11038 225 -11026
rect 159 -14414 175 -11038
rect 209 -14414 225 -11038
rect 159 -14426 225 -14414
rect 255 -11038 321 -11026
rect 255 -14414 271 -11038
rect 305 -14414 321 -11038
rect 255 -14426 321 -14414
rect 351 -11038 417 -11026
rect 351 -14414 367 -11038
rect 401 -14414 417 -11038
rect 351 -14426 417 -14414
rect 447 -11038 513 -11026
rect 447 -14414 463 -11038
rect 497 -14414 513 -11038
rect 447 -14426 513 -14414
rect 543 -11038 609 -11026
rect 543 -14414 559 -11038
rect 593 -14414 609 -11038
rect 543 -14426 609 -14414
rect 639 -11038 705 -11026
rect 639 -14414 655 -11038
rect 689 -14414 705 -11038
rect 639 -14426 705 -14414
rect 735 -11038 801 -11026
rect 735 -14414 751 -11038
rect 785 -14414 801 -11038
rect 735 -14426 801 -14414
rect 831 -11038 897 -11026
rect 831 -14414 847 -11038
rect 881 -14414 897 -11038
rect 831 -14426 897 -14414
rect 927 -11038 989 -11026
rect 927 -14414 943 -11038
rect 977 -14414 989 -11038
rect 927 -14426 989 -14414
rect -989 -14674 -927 -14662
rect -989 -18050 -977 -14674
rect -943 -18050 -927 -14674
rect -989 -18062 -927 -18050
rect -897 -14674 -831 -14662
rect -897 -18050 -881 -14674
rect -847 -18050 -831 -14674
rect -897 -18062 -831 -18050
rect -801 -14674 -735 -14662
rect -801 -18050 -785 -14674
rect -751 -18050 -735 -14674
rect -801 -18062 -735 -18050
rect -705 -14674 -639 -14662
rect -705 -18050 -689 -14674
rect -655 -18050 -639 -14674
rect -705 -18062 -639 -18050
rect -609 -14674 -543 -14662
rect -609 -18050 -593 -14674
rect -559 -18050 -543 -14674
rect -609 -18062 -543 -18050
rect -513 -14674 -447 -14662
rect -513 -18050 -497 -14674
rect -463 -18050 -447 -14674
rect -513 -18062 -447 -18050
rect -417 -14674 -351 -14662
rect -417 -18050 -401 -14674
rect -367 -18050 -351 -14674
rect -417 -18062 -351 -18050
rect -321 -14674 -255 -14662
rect -321 -18050 -305 -14674
rect -271 -18050 -255 -14674
rect -321 -18062 -255 -18050
rect -225 -14674 -159 -14662
rect -225 -18050 -209 -14674
rect -175 -18050 -159 -14674
rect -225 -18062 -159 -18050
rect -129 -14674 -63 -14662
rect -129 -18050 -113 -14674
rect -79 -18050 -63 -14674
rect -129 -18062 -63 -18050
rect -33 -14674 33 -14662
rect -33 -18050 -17 -14674
rect 17 -18050 33 -14674
rect -33 -18062 33 -18050
rect 63 -14674 129 -14662
rect 63 -18050 79 -14674
rect 113 -18050 129 -14674
rect 63 -18062 129 -18050
rect 159 -14674 225 -14662
rect 159 -18050 175 -14674
rect 209 -18050 225 -14674
rect 159 -18062 225 -18050
rect 255 -14674 321 -14662
rect 255 -18050 271 -14674
rect 305 -18050 321 -14674
rect 255 -18062 321 -18050
rect 351 -14674 417 -14662
rect 351 -18050 367 -14674
rect 401 -18050 417 -14674
rect 351 -18062 417 -18050
rect 447 -14674 513 -14662
rect 447 -18050 463 -14674
rect 497 -18050 513 -14674
rect 447 -18062 513 -18050
rect 543 -14674 609 -14662
rect 543 -18050 559 -14674
rect 593 -18050 609 -14674
rect 543 -18062 609 -18050
rect 639 -14674 705 -14662
rect 639 -18050 655 -14674
rect 689 -18050 705 -14674
rect 639 -18062 705 -18050
rect 735 -14674 801 -14662
rect 735 -18050 751 -14674
rect 785 -18050 801 -14674
rect 735 -18062 801 -18050
rect 831 -14674 897 -14662
rect 831 -18050 847 -14674
rect 881 -18050 897 -14674
rect 831 -18062 897 -18050
rect 927 -14674 989 -14662
rect 927 -18050 943 -14674
rect 977 -18050 989 -14674
rect 927 -18062 989 -18050
<< pdiffc >>
rect -977 14674 -943 18050
rect -881 14674 -847 18050
rect -785 14674 -751 18050
rect -689 14674 -655 18050
rect -593 14674 -559 18050
rect -497 14674 -463 18050
rect -401 14674 -367 18050
rect -305 14674 -271 18050
rect -209 14674 -175 18050
rect -113 14674 -79 18050
rect -17 14674 17 18050
rect 79 14674 113 18050
rect 175 14674 209 18050
rect 271 14674 305 18050
rect 367 14674 401 18050
rect 463 14674 497 18050
rect 559 14674 593 18050
rect 655 14674 689 18050
rect 751 14674 785 18050
rect 847 14674 881 18050
rect 943 14674 977 18050
rect -977 11038 -943 14414
rect -881 11038 -847 14414
rect -785 11038 -751 14414
rect -689 11038 -655 14414
rect -593 11038 -559 14414
rect -497 11038 -463 14414
rect -401 11038 -367 14414
rect -305 11038 -271 14414
rect -209 11038 -175 14414
rect -113 11038 -79 14414
rect -17 11038 17 14414
rect 79 11038 113 14414
rect 175 11038 209 14414
rect 271 11038 305 14414
rect 367 11038 401 14414
rect 463 11038 497 14414
rect 559 11038 593 14414
rect 655 11038 689 14414
rect 751 11038 785 14414
rect 847 11038 881 14414
rect 943 11038 977 14414
rect -977 7402 -943 10778
rect -881 7402 -847 10778
rect -785 7402 -751 10778
rect -689 7402 -655 10778
rect -593 7402 -559 10778
rect -497 7402 -463 10778
rect -401 7402 -367 10778
rect -305 7402 -271 10778
rect -209 7402 -175 10778
rect -113 7402 -79 10778
rect -17 7402 17 10778
rect 79 7402 113 10778
rect 175 7402 209 10778
rect 271 7402 305 10778
rect 367 7402 401 10778
rect 463 7402 497 10778
rect 559 7402 593 10778
rect 655 7402 689 10778
rect 751 7402 785 10778
rect 847 7402 881 10778
rect 943 7402 977 10778
rect -977 3766 -943 7142
rect -881 3766 -847 7142
rect -785 3766 -751 7142
rect -689 3766 -655 7142
rect -593 3766 -559 7142
rect -497 3766 -463 7142
rect -401 3766 -367 7142
rect -305 3766 -271 7142
rect -209 3766 -175 7142
rect -113 3766 -79 7142
rect -17 3766 17 7142
rect 79 3766 113 7142
rect 175 3766 209 7142
rect 271 3766 305 7142
rect 367 3766 401 7142
rect 463 3766 497 7142
rect 559 3766 593 7142
rect 655 3766 689 7142
rect 751 3766 785 7142
rect 847 3766 881 7142
rect 943 3766 977 7142
rect -977 130 -943 3506
rect -881 130 -847 3506
rect -785 130 -751 3506
rect -689 130 -655 3506
rect -593 130 -559 3506
rect -497 130 -463 3506
rect -401 130 -367 3506
rect -305 130 -271 3506
rect -209 130 -175 3506
rect -113 130 -79 3506
rect -17 130 17 3506
rect 79 130 113 3506
rect 175 130 209 3506
rect 271 130 305 3506
rect 367 130 401 3506
rect 463 130 497 3506
rect 559 130 593 3506
rect 655 130 689 3506
rect 751 130 785 3506
rect 847 130 881 3506
rect 943 130 977 3506
rect -977 -3506 -943 -130
rect -881 -3506 -847 -130
rect -785 -3506 -751 -130
rect -689 -3506 -655 -130
rect -593 -3506 -559 -130
rect -497 -3506 -463 -130
rect -401 -3506 -367 -130
rect -305 -3506 -271 -130
rect -209 -3506 -175 -130
rect -113 -3506 -79 -130
rect -17 -3506 17 -130
rect 79 -3506 113 -130
rect 175 -3506 209 -130
rect 271 -3506 305 -130
rect 367 -3506 401 -130
rect 463 -3506 497 -130
rect 559 -3506 593 -130
rect 655 -3506 689 -130
rect 751 -3506 785 -130
rect 847 -3506 881 -130
rect 943 -3506 977 -130
rect -977 -7142 -943 -3766
rect -881 -7142 -847 -3766
rect -785 -7142 -751 -3766
rect -689 -7142 -655 -3766
rect -593 -7142 -559 -3766
rect -497 -7142 -463 -3766
rect -401 -7142 -367 -3766
rect -305 -7142 -271 -3766
rect -209 -7142 -175 -3766
rect -113 -7142 -79 -3766
rect -17 -7142 17 -3766
rect 79 -7142 113 -3766
rect 175 -7142 209 -3766
rect 271 -7142 305 -3766
rect 367 -7142 401 -3766
rect 463 -7142 497 -3766
rect 559 -7142 593 -3766
rect 655 -7142 689 -3766
rect 751 -7142 785 -3766
rect 847 -7142 881 -3766
rect 943 -7142 977 -3766
rect -977 -10778 -943 -7402
rect -881 -10778 -847 -7402
rect -785 -10778 -751 -7402
rect -689 -10778 -655 -7402
rect -593 -10778 -559 -7402
rect -497 -10778 -463 -7402
rect -401 -10778 -367 -7402
rect -305 -10778 -271 -7402
rect -209 -10778 -175 -7402
rect -113 -10778 -79 -7402
rect -17 -10778 17 -7402
rect 79 -10778 113 -7402
rect 175 -10778 209 -7402
rect 271 -10778 305 -7402
rect 367 -10778 401 -7402
rect 463 -10778 497 -7402
rect 559 -10778 593 -7402
rect 655 -10778 689 -7402
rect 751 -10778 785 -7402
rect 847 -10778 881 -7402
rect 943 -10778 977 -7402
rect -977 -14414 -943 -11038
rect -881 -14414 -847 -11038
rect -785 -14414 -751 -11038
rect -689 -14414 -655 -11038
rect -593 -14414 -559 -11038
rect -497 -14414 -463 -11038
rect -401 -14414 -367 -11038
rect -305 -14414 -271 -11038
rect -209 -14414 -175 -11038
rect -113 -14414 -79 -11038
rect -17 -14414 17 -11038
rect 79 -14414 113 -11038
rect 175 -14414 209 -11038
rect 271 -14414 305 -11038
rect 367 -14414 401 -11038
rect 463 -14414 497 -11038
rect 559 -14414 593 -11038
rect 655 -14414 689 -11038
rect 751 -14414 785 -11038
rect 847 -14414 881 -11038
rect 943 -14414 977 -11038
rect -977 -18050 -943 -14674
rect -881 -18050 -847 -14674
rect -785 -18050 -751 -14674
rect -689 -18050 -655 -14674
rect -593 -18050 -559 -14674
rect -497 -18050 -463 -14674
rect -401 -18050 -367 -14674
rect -305 -18050 -271 -14674
rect -209 -18050 -175 -14674
rect -113 -18050 -79 -14674
rect -17 -18050 17 -14674
rect 79 -18050 113 -14674
rect 175 -18050 209 -14674
rect 271 -18050 305 -14674
rect 367 -18050 401 -14674
rect 463 -18050 497 -14674
rect 559 -18050 593 -14674
rect 655 -18050 689 -14674
rect 751 -18050 785 -14674
rect 847 -18050 881 -14674
rect 943 -18050 977 -14674
<< poly >>
rect -945 18143 -879 18159
rect -945 18109 -929 18143
rect -895 18109 -879 18143
rect -945 18093 -879 18109
rect -753 18143 -687 18159
rect -753 18109 -737 18143
rect -703 18109 -687 18143
rect -753 18093 -687 18109
rect -561 18143 -495 18159
rect -561 18109 -545 18143
rect -511 18109 -495 18143
rect -561 18093 -495 18109
rect -369 18143 -303 18159
rect -369 18109 -353 18143
rect -319 18109 -303 18143
rect -369 18093 -303 18109
rect -177 18143 -111 18159
rect -177 18109 -161 18143
rect -127 18109 -111 18143
rect -177 18093 -111 18109
rect 15 18143 81 18159
rect 15 18109 31 18143
rect 65 18109 81 18143
rect 15 18093 81 18109
rect 207 18143 273 18159
rect 207 18109 223 18143
rect 257 18109 273 18143
rect 207 18093 273 18109
rect 399 18143 465 18159
rect 399 18109 415 18143
rect 449 18109 465 18143
rect 399 18093 465 18109
rect 591 18143 657 18159
rect 591 18109 607 18143
rect 641 18109 657 18143
rect 591 18093 657 18109
rect 783 18143 849 18159
rect 783 18109 799 18143
rect 833 18109 849 18143
rect 783 18093 849 18109
rect -927 18062 -897 18093
rect -831 18062 -801 18088
rect -735 18062 -705 18093
rect -639 18062 -609 18088
rect -543 18062 -513 18093
rect -447 18062 -417 18088
rect -351 18062 -321 18093
rect -255 18062 -225 18088
rect -159 18062 -129 18093
rect -63 18062 -33 18088
rect 33 18062 63 18093
rect 129 18062 159 18088
rect 225 18062 255 18093
rect 321 18062 351 18088
rect 417 18062 447 18093
rect 513 18062 543 18088
rect 609 18062 639 18093
rect 705 18062 735 18088
rect 801 18062 831 18093
rect 897 18062 927 18088
rect -927 14636 -897 14662
rect -831 14631 -801 14662
rect -735 14636 -705 14662
rect -639 14631 -609 14662
rect -543 14636 -513 14662
rect -447 14631 -417 14662
rect -351 14636 -321 14662
rect -255 14631 -225 14662
rect -159 14636 -129 14662
rect -63 14631 -33 14662
rect 33 14636 63 14662
rect 129 14631 159 14662
rect 225 14636 255 14662
rect 321 14631 351 14662
rect 417 14636 447 14662
rect 513 14631 543 14662
rect 609 14636 639 14662
rect 705 14631 735 14662
rect 801 14636 831 14662
rect 897 14631 927 14662
rect -849 14615 -783 14631
rect -849 14581 -833 14615
rect -799 14581 -783 14615
rect -849 14565 -783 14581
rect -657 14615 -591 14631
rect -657 14581 -641 14615
rect -607 14581 -591 14615
rect -657 14565 -591 14581
rect -465 14615 -399 14631
rect -465 14581 -449 14615
rect -415 14581 -399 14615
rect -465 14565 -399 14581
rect -273 14615 -207 14631
rect -273 14581 -257 14615
rect -223 14581 -207 14615
rect -273 14565 -207 14581
rect -81 14615 -15 14631
rect -81 14581 -65 14615
rect -31 14581 -15 14615
rect -81 14565 -15 14581
rect 111 14615 177 14631
rect 111 14581 127 14615
rect 161 14581 177 14615
rect 111 14565 177 14581
rect 303 14615 369 14631
rect 303 14581 319 14615
rect 353 14581 369 14615
rect 303 14565 369 14581
rect 495 14615 561 14631
rect 495 14581 511 14615
rect 545 14581 561 14615
rect 495 14565 561 14581
rect 687 14615 753 14631
rect 687 14581 703 14615
rect 737 14581 753 14615
rect 687 14565 753 14581
rect 879 14615 945 14631
rect 879 14581 895 14615
rect 929 14581 945 14615
rect 879 14565 945 14581
rect -849 14507 -783 14523
rect -849 14473 -833 14507
rect -799 14473 -783 14507
rect -849 14457 -783 14473
rect -657 14507 -591 14523
rect -657 14473 -641 14507
rect -607 14473 -591 14507
rect -657 14457 -591 14473
rect -465 14507 -399 14523
rect -465 14473 -449 14507
rect -415 14473 -399 14507
rect -465 14457 -399 14473
rect -273 14507 -207 14523
rect -273 14473 -257 14507
rect -223 14473 -207 14507
rect -273 14457 -207 14473
rect -81 14507 -15 14523
rect -81 14473 -65 14507
rect -31 14473 -15 14507
rect -81 14457 -15 14473
rect 111 14507 177 14523
rect 111 14473 127 14507
rect 161 14473 177 14507
rect 111 14457 177 14473
rect 303 14507 369 14523
rect 303 14473 319 14507
rect 353 14473 369 14507
rect 303 14457 369 14473
rect 495 14507 561 14523
rect 495 14473 511 14507
rect 545 14473 561 14507
rect 495 14457 561 14473
rect 687 14507 753 14523
rect 687 14473 703 14507
rect 737 14473 753 14507
rect 687 14457 753 14473
rect 879 14507 945 14523
rect 879 14473 895 14507
rect 929 14473 945 14507
rect 879 14457 945 14473
rect -927 14426 -897 14452
rect -831 14426 -801 14457
rect -735 14426 -705 14452
rect -639 14426 -609 14457
rect -543 14426 -513 14452
rect -447 14426 -417 14457
rect -351 14426 -321 14452
rect -255 14426 -225 14457
rect -159 14426 -129 14452
rect -63 14426 -33 14457
rect 33 14426 63 14452
rect 129 14426 159 14457
rect 225 14426 255 14452
rect 321 14426 351 14457
rect 417 14426 447 14452
rect 513 14426 543 14457
rect 609 14426 639 14452
rect 705 14426 735 14457
rect 801 14426 831 14452
rect 897 14426 927 14457
rect -927 10995 -897 11026
rect -831 11000 -801 11026
rect -735 10995 -705 11026
rect -639 11000 -609 11026
rect -543 10995 -513 11026
rect -447 11000 -417 11026
rect -351 10995 -321 11026
rect -255 11000 -225 11026
rect -159 10995 -129 11026
rect -63 11000 -33 11026
rect 33 10995 63 11026
rect 129 11000 159 11026
rect 225 10995 255 11026
rect 321 11000 351 11026
rect 417 10995 447 11026
rect 513 11000 543 11026
rect 609 10995 639 11026
rect 705 11000 735 11026
rect 801 10995 831 11026
rect 897 11000 927 11026
rect -945 10979 -879 10995
rect -945 10945 -929 10979
rect -895 10945 -879 10979
rect -945 10929 -879 10945
rect -753 10979 -687 10995
rect -753 10945 -737 10979
rect -703 10945 -687 10979
rect -753 10929 -687 10945
rect -561 10979 -495 10995
rect -561 10945 -545 10979
rect -511 10945 -495 10979
rect -561 10929 -495 10945
rect -369 10979 -303 10995
rect -369 10945 -353 10979
rect -319 10945 -303 10979
rect -369 10929 -303 10945
rect -177 10979 -111 10995
rect -177 10945 -161 10979
rect -127 10945 -111 10979
rect -177 10929 -111 10945
rect 15 10979 81 10995
rect 15 10945 31 10979
rect 65 10945 81 10979
rect 15 10929 81 10945
rect 207 10979 273 10995
rect 207 10945 223 10979
rect 257 10945 273 10979
rect 207 10929 273 10945
rect 399 10979 465 10995
rect 399 10945 415 10979
rect 449 10945 465 10979
rect 399 10929 465 10945
rect 591 10979 657 10995
rect 591 10945 607 10979
rect 641 10945 657 10979
rect 591 10929 657 10945
rect 783 10979 849 10995
rect 783 10945 799 10979
rect 833 10945 849 10979
rect 783 10929 849 10945
rect -945 10871 -879 10887
rect -945 10837 -929 10871
rect -895 10837 -879 10871
rect -945 10821 -879 10837
rect -753 10871 -687 10887
rect -753 10837 -737 10871
rect -703 10837 -687 10871
rect -753 10821 -687 10837
rect -561 10871 -495 10887
rect -561 10837 -545 10871
rect -511 10837 -495 10871
rect -561 10821 -495 10837
rect -369 10871 -303 10887
rect -369 10837 -353 10871
rect -319 10837 -303 10871
rect -369 10821 -303 10837
rect -177 10871 -111 10887
rect -177 10837 -161 10871
rect -127 10837 -111 10871
rect -177 10821 -111 10837
rect 15 10871 81 10887
rect 15 10837 31 10871
rect 65 10837 81 10871
rect 15 10821 81 10837
rect 207 10871 273 10887
rect 207 10837 223 10871
rect 257 10837 273 10871
rect 207 10821 273 10837
rect 399 10871 465 10887
rect 399 10837 415 10871
rect 449 10837 465 10871
rect 399 10821 465 10837
rect 591 10871 657 10887
rect 591 10837 607 10871
rect 641 10837 657 10871
rect 591 10821 657 10837
rect 783 10871 849 10887
rect 783 10837 799 10871
rect 833 10837 849 10871
rect 783 10821 849 10837
rect -927 10790 -897 10821
rect -831 10790 -801 10816
rect -735 10790 -705 10821
rect -639 10790 -609 10816
rect -543 10790 -513 10821
rect -447 10790 -417 10816
rect -351 10790 -321 10821
rect -255 10790 -225 10816
rect -159 10790 -129 10821
rect -63 10790 -33 10816
rect 33 10790 63 10821
rect 129 10790 159 10816
rect 225 10790 255 10821
rect 321 10790 351 10816
rect 417 10790 447 10821
rect 513 10790 543 10816
rect 609 10790 639 10821
rect 705 10790 735 10816
rect 801 10790 831 10821
rect 897 10790 927 10816
rect -927 7364 -897 7390
rect -831 7359 -801 7390
rect -735 7364 -705 7390
rect -639 7359 -609 7390
rect -543 7364 -513 7390
rect -447 7359 -417 7390
rect -351 7364 -321 7390
rect -255 7359 -225 7390
rect -159 7364 -129 7390
rect -63 7359 -33 7390
rect 33 7364 63 7390
rect 129 7359 159 7390
rect 225 7364 255 7390
rect 321 7359 351 7390
rect 417 7364 447 7390
rect 513 7359 543 7390
rect 609 7364 639 7390
rect 705 7359 735 7390
rect 801 7364 831 7390
rect 897 7359 927 7390
rect -849 7343 -783 7359
rect -849 7309 -833 7343
rect -799 7309 -783 7343
rect -849 7293 -783 7309
rect -657 7343 -591 7359
rect -657 7309 -641 7343
rect -607 7309 -591 7343
rect -657 7293 -591 7309
rect -465 7343 -399 7359
rect -465 7309 -449 7343
rect -415 7309 -399 7343
rect -465 7293 -399 7309
rect -273 7343 -207 7359
rect -273 7309 -257 7343
rect -223 7309 -207 7343
rect -273 7293 -207 7309
rect -81 7343 -15 7359
rect -81 7309 -65 7343
rect -31 7309 -15 7343
rect -81 7293 -15 7309
rect 111 7343 177 7359
rect 111 7309 127 7343
rect 161 7309 177 7343
rect 111 7293 177 7309
rect 303 7343 369 7359
rect 303 7309 319 7343
rect 353 7309 369 7343
rect 303 7293 369 7309
rect 495 7343 561 7359
rect 495 7309 511 7343
rect 545 7309 561 7343
rect 495 7293 561 7309
rect 687 7343 753 7359
rect 687 7309 703 7343
rect 737 7309 753 7343
rect 687 7293 753 7309
rect 879 7343 945 7359
rect 879 7309 895 7343
rect 929 7309 945 7343
rect 879 7293 945 7309
rect -849 7235 -783 7251
rect -849 7201 -833 7235
rect -799 7201 -783 7235
rect -849 7185 -783 7201
rect -657 7235 -591 7251
rect -657 7201 -641 7235
rect -607 7201 -591 7235
rect -657 7185 -591 7201
rect -465 7235 -399 7251
rect -465 7201 -449 7235
rect -415 7201 -399 7235
rect -465 7185 -399 7201
rect -273 7235 -207 7251
rect -273 7201 -257 7235
rect -223 7201 -207 7235
rect -273 7185 -207 7201
rect -81 7235 -15 7251
rect -81 7201 -65 7235
rect -31 7201 -15 7235
rect -81 7185 -15 7201
rect 111 7235 177 7251
rect 111 7201 127 7235
rect 161 7201 177 7235
rect 111 7185 177 7201
rect 303 7235 369 7251
rect 303 7201 319 7235
rect 353 7201 369 7235
rect 303 7185 369 7201
rect 495 7235 561 7251
rect 495 7201 511 7235
rect 545 7201 561 7235
rect 495 7185 561 7201
rect 687 7235 753 7251
rect 687 7201 703 7235
rect 737 7201 753 7235
rect 687 7185 753 7201
rect 879 7235 945 7251
rect 879 7201 895 7235
rect 929 7201 945 7235
rect 879 7185 945 7201
rect -927 7154 -897 7180
rect -831 7154 -801 7185
rect -735 7154 -705 7180
rect -639 7154 -609 7185
rect -543 7154 -513 7180
rect -447 7154 -417 7185
rect -351 7154 -321 7180
rect -255 7154 -225 7185
rect -159 7154 -129 7180
rect -63 7154 -33 7185
rect 33 7154 63 7180
rect 129 7154 159 7185
rect 225 7154 255 7180
rect 321 7154 351 7185
rect 417 7154 447 7180
rect 513 7154 543 7185
rect 609 7154 639 7180
rect 705 7154 735 7185
rect 801 7154 831 7180
rect 897 7154 927 7185
rect -927 3723 -897 3754
rect -831 3728 -801 3754
rect -735 3723 -705 3754
rect -639 3728 -609 3754
rect -543 3723 -513 3754
rect -447 3728 -417 3754
rect -351 3723 -321 3754
rect -255 3728 -225 3754
rect -159 3723 -129 3754
rect -63 3728 -33 3754
rect 33 3723 63 3754
rect 129 3728 159 3754
rect 225 3723 255 3754
rect 321 3728 351 3754
rect 417 3723 447 3754
rect 513 3728 543 3754
rect 609 3723 639 3754
rect 705 3728 735 3754
rect 801 3723 831 3754
rect 897 3728 927 3754
rect -945 3707 -879 3723
rect -945 3673 -929 3707
rect -895 3673 -879 3707
rect -945 3657 -879 3673
rect -753 3707 -687 3723
rect -753 3673 -737 3707
rect -703 3673 -687 3707
rect -753 3657 -687 3673
rect -561 3707 -495 3723
rect -561 3673 -545 3707
rect -511 3673 -495 3707
rect -561 3657 -495 3673
rect -369 3707 -303 3723
rect -369 3673 -353 3707
rect -319 3673 -303 3707
rect -369 3657 -303 3673
rect -177 3707 -111 3723
rect -177 3673 -161 3707
rect -127 3673 -111 3707
rect -177 3657 -111 3673
rect 15 3707 81 3723
rect 15 3673 31 3707
rect 65 3673 81 3707
rect 15 3657 81 3673
rect 207 3707 273 3723
rect 207 3673 223 3707
rect 257 3673 273 3707
rect 207 3657 273 3673
rect 399 3707 465 3723
rect 399 3673 415 3707
rect 449 3673 465 3707
rect 399 3657 465 3673
rect 591 3707 657 3723
rect 591 3673 607 3707
rect 641 3673 657 3707
rect 591 3657 657 3673
rect 783 3707 849 3723
rect 783 3673 799 3707
rect 833 3673 849 3707
rect 783 3657 849 3673
rect -945 3599 -879 3615
rect -945 3565 -929 3599
rect -895 3565 -879 3599
rect -945 3549 -879 3565
rect -753 3599 -687 3615
rect -753 3565 -737 3599
rect -703 3565 -687 3599
rect -753 3549 -687 3565
rect -561 3599 -495 3615
rect -561 3565 -545 3599
rect -511 3565 -495 3599
rect -561 3549 -495 3565
rect -369 3599 -303 3615
rect -369 3565 -353 3599
rect -319 3565 -303 3599
rect -369 3549 -303 3565
rect -177 3599 -111 3615
rect -177 3565 -161 3599
rect -127 3565 -111 3599
rect -177 3549 -111 3565
rect 15 3599 81 3615
rect 15 3565 31 3599
rect 65 3565 81 3599
rect 15 3549 81 3565
rect 207 3599 273 3615
rect 207 3565 223 3599
rect 257 3565 273 3599
rect 207 3549 273 3565
rect 399 3599 465 3615
rect 399 3565 415 3599
rect 449 3565 465 3599
rect 399 3549 465 3565
rect 591 3599 657 3615
rect 591 3565 607 3599
rect 641 3565 657 3599
rect 591 3549 657 3565
rect 783 3599 849 3615
rect 783 3565 799 3599
rect 833 3565 849 3599
rect 783 3549 849 3565
rect -927 3518 -897 3549
rect -831 3518 -801 3544
rect -735 3518 -705 3549
rect -639 3518 -609 3544
rect -543 3518 -513 3549
rect -447 3518 -417 3544
rect -351 3518 -321 3549
rect -255 3518 -225 3544
rect -159 3518 -129 3549
rect -63 3518 -33 3544
rect 33 3518 63 3549
rect 129 3518 159 3544
rect 225 3518 255 3549
rect 321 3518 351 3544
rect 417 3518 447 3549
rect 513 3518 543 3544
rect 609 3518 639 3549
rect 705 3518 735 3544
rect 801 3518 831 3549
rect 897 3518 927 3544
rect -927 92 -897 118
rect -831 87 -801 118
rect -735 92 -705 118
rect -639 87 -609 118
rect -543 92 -513 118
rect -447 87 -417 118
rect -351 92 -321 118
rect -255 87 -225 118
rect -159 92 -129 118
rect -63 87 -33 118
rect 33 92 63 118
rect 129 87 159 118
rect 225 92 255 118
rect 321 87 351 118
rect 417 92 447 118
rect 513 87 543 118
rect 609 92 639 118
rect 705 87 735 118
rect 801 92 831 118
rect 897 87 927 118
rect -849 71 -783 87
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 879 -87 945 -71
rect -927 -118 -897 -92
rect -831 -118 -801 -87
rect -735 -118 -705 -92
rect -639 -118 -609 -87
rect -543 -118 -513 -92
rect -447 -118 -417 -87
rect -351 -118 -321 -92
rect -255 -118 -225 -87
rect -159 -118 -129 -92
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect 129 -118 159 -87
rect 225 -118 255 -92
rect 321 -118 351 -87
rect 417 -118 447 -92
rect 513 -118 543 -87
rect 609 -118 639 -92
rect 705 -118 735 -87
rect 801 -118 831 -92
rect 897 -118 927 -87
rect -927 -3549 -897 -3518
rect -831 -3544 -801 -3518
rect -735 -3549 -705 -3518
rect -639 -3544 -609 -3518
rect -543 -3549 -513 -3518
rect -447 -3544 -417 -3518
rect -351 -3549 -321 -3518
rect -255 -3544 -225 -3518
rect -159 -3549 -129 -3518
rect -63 -3544 -33 -3518
rect 33 -3549 63 -3518
rect 129 -3544 159 -3518
rect 225 -3549 255 -3518
rect 321 -3544 351 -3518
rect 417 -3549 447 -3518
rect 513 -3544 543 -3518
rect 609 -3549 639 -3518
rect 705 -3544 735 -3518
rect 801 -3549 831 -3518
rect 897 -3544 927 -3518
rect -945 -3565 -879 -3549
rect -945 -3599 -929 -3565
rect -895 -3599 -879 -3565
rect -945 -3615 -879 -3599
rect -753 -3565 -687 -3549
rect -753 -3599 -737 -3565
rect -703 -3599 -687 -3565
rect -753 -3615 -687 -3599
rect -561 -3565 -495 -3549
rect -561 -3599 -545 -3565
rect -511 -3599 -495 -3565
rect -561 -3615 -495 -3599
rect -369 -3565 -303 -3549
rect -369 -3599 -353 -3565
rect -319 -3599 -303 -3565
rect -369 -3615 -303 -3599
rect -177 -3565 -111 -3549
rect -177 -3599 -161 -3565
rect -127 -3599 -111 -3565
rect -177 -3615 -111 -3599
rect 15 -3565 81 -3549
rect 15 -3599 31 -3565
rect 65 -3599 81 -3565
rect 15 -3615 81 -3599
rect 207 -3565 273 -3549
rect 207 -3599 223 -3565
rect 257 -3599 273 -3565
rect 207 -3615 273 -3599
rect 399 -3565 465 -3549
rect 399 -3599 415 -3565
rect 449 -3599 465 -3565
rect 399 -3615 465 -3599
rect 591 -3565 657 -3549
rect 591 -3599 607 -3565
rect 641 -3599 657 -3565
rect 591 -3615 657 -3599
rect 783 -3565 849 -3549
rect 783 -3599 799 -3565
rect 833 -3599 849 -3565
rect 783 -3615 849 -3599
rect -945 -3673 -879 -3657
rect -945 -3707 -929 -3673
rect -895 -3707 -879 -3673
rect -945 -3723 -879 -3707
rect -753 -3673 -687 -3657
rect -753 -3707 -737 -3673
rect -703 -3707 -687 -3673
rect -753 -3723 -687 -3707
rect -561 -3673 -495 -3657
rect -561 -3707 -545 -3673
rect -511 -3707 -495 -3673
rect -561 -3723 -495 -3707
rect -369 -3673 -303 -3657
rect -369 -3707 -353 -3673
rect -319 -3707 -303 -3673
rect -369 -3723 -303 -3707
rect -177 -3673 -111 -3657
rect -177 -3707 -161 -3673
rect -127 -3707 -111 -3673
rect -177 -3723 -111 -3707
rect 15 -3673 81 -3657
rect 15 -3707 31 -3673
rect 65 -3707 81 -3673
rect 15 -3723 81 -3707
rect 207 -3673 273 -3657
rect 207 -3707 223 -3673
rect 257 -3707 273 -3673
rect 207 -3723 273 -3707
rect 399 -3673 465 -3657
rect 399 -3707 415 -3673
rect 449 -3707 465 -3673
rect 399 -3723 465 -3707
rect 591 -3673 657 -3657
rect 591 -3707 607 -3673
rect 641 -3707 657 -3673
rect 591 -3723 657 -3707
rect 783 -3673 849 -3657
rect 783 -3707 799 -3673
rect 833 -3707 849 -3673
rect 783 -3723 849 -3707
rect -927 -3754 -897 -3723
rect -831 -3754 -801 -3728
rect -735 -3754 -705 -3723
rect -639 -3754 -609 -3728
rect -543 -3754 -513 -3723
rect -447 -3754 -417 -3728
rect -351 -3754 -321 -3723
rect -255 -3754 -225 -3728
rect -159 -3754 -129 -3723
rect -63 -3754 -33 -3728
rect 33 -3754 63 -3723
rect 129 -3754 159 -3728
rect 225 -3754 255 -3723
rect 321 -3754 351 -3728
rect 417 -3754 447 -3723
rect 513 -3754 543 -3728
rect 609 -3754 639 -3723
rect 705 -3754 735 -3728
rect 801 -3754 831 -3723
rect 897 -3754 927 -3728
rect -927 -7180 -897 -7154
rect -831 -7185 -801 -7154
rect -735 -7180 -705 -7154
rect -639 -7185 -609 -7154
rect -543 -7180 -513 -7154
rect -447 -7185 -417 -7154
rect -351 -7180 -321 -7154
rect -255 -7185 -225 -7154
rect -159 -7180 -129 -7154
rect -63 -7185 -33 -7154
rect 33 -7180 63 -7154
rect 129 -7185 159 -7154
rect 225 -7180 255 -7154
rect 321 -7185 351 -7154
rect 417 -7180 447 -7154
rect 513 -7185 543 -7154
rect 609 -7180 639 -7154
rect 705 -7185 735 -7154
rect 801 -7180 831 -7154
rect 897 -7185 927 -7154
rect -849 -7201 -783 -7185
rect -849 -7235 -833 -7201
rect -799 -7235 -783 -7201
rect -849 -7251 -783 -7235
rect -657 -7201 -591 -7185
rect -657 -7235 -641 -7201
rect -607 -7235 -591 -7201
rect -657 -7251 -591 -7235
rect -465 -7201 -399 -7185
rect -465 -7235 -449 -7201
rect -415 -7235 -399 -7201
rect -465 -7251 -399 -7235
rect -273 -7201 -207 -7185
rect -273 -7235 -257 -7201
rect -223 -7235 -207 -7201
rect -273 -7251 -207 -7235
rect -81 -7201 -15 -7185
rect -81 -7235 -65 -7201
rect -31 -7235 -15 -7201
rect -81 -7251 -15 -7235
rect 111 -7201 177 -7185
rect 111 -7235 127 -7201
rect 161 -7235 177 -7201
rect 111 -7251 177 -7235
rect 303 -7201 369 -7185
rect 303 -7235 319 -7201
rect 353 -7235 369 -7201
rect 303 -7251 369 -7235
rect 495 -7201 561 -7185
rect 495 -7235 511 -7201
rect 545 -7235 561 -7201
rect 495 -7251 561 -7235
rect 687 -7201 753 -7185
rect 687 -7235 703 -7201
rect 737 -7235 753 -7201
rect 687 -7251 753 -7235
rect 879 -7201 945 -7185
rect 879 -7235 895 -7201
rect 929 -7235 945 -7201
rect 879 -7251 945 -7235
rect -849 -7309 -783 -7293
rect -849 -7343 -833 -7309
rect -799 -7343 -783 -7309
rect -849 -7359 -783 -7343
rect -657 -7309 -591 -7293
rect -657 -7343 -641 -7309
rect -607 -7343 -591 -7309
rect -657 -7359 -591 -7343
rect -465 -7309 -399 -7293
rect -465 -7343 -449 -7309
rect -415 -7343 -399 -7309
rect -465 -7359 -399 -7343
rect -273 -7309 -207 -7293
rect -273 -7343 -257 -7309
rect -223 -7343 -207 -7309
rect -273 -7359 -207 -7343
rect -81 -7309 -15 -7293
rect -81 -7343 -65 -7309
rect -31 -7343 -15 -7309
rect -81 -7359 -15 -7343
rect 111 -7309 177 -7293
rect 111 -7343 127 -7309
rect 161 -7343 177 -7309
rect 111 -7359 177 -7343
rect 303 -7309 369 -7293
rect 303 -7343 319 -7309
rect 353 -7343 369 -7309
rect 303 -7359 369 -7343
rect 495 -7309 561 -7293
rect 495 -7343 511 -7309
rect 545 -7343 561 -7309
rect 495 -7359 561 -7343
rect 687 -7309 753 -7293
rect 687 -7343 703 -7309
rect 737 -7343 753 -7309
rect 687 -7359 753 -7343
rect 879 -7309 945 -7293
rect 879 -7343 895 -7309
rect 929 -7343 945 -7309
rect 879 -7359 945 -7343
rect -927 -7390 -897 -7364
rect -831 -7390 -801 -7359
rect -735 -7390 -705 -7364
rect -639 -7390 -609 -7359
rect -543 -7390 -513 -7364
rect -447 -7390 -417 -7359
rect -351 -7390 -321 -7364
rect -255 -7390 -225 -7359
rect -159 -7390 -129 -7364
rect -63 -7390 -33 -7359
rect 33 -7390 63 -7364
rect 129 -7390 159 -7359
rect 225 -7390 255 -7364
rect 321 -7390 351 -7359
rect 417 -7390 447 -7364
rect 513 -7390 543 -7359
rect 609 -7390 639 -7364
rect 705 -7390 735 -7359
rect 801 -7390 831 -7364
rect 897 -7390 927 -7359
rect -927 -10821 -897 -10790
rect -831 -10816 -801 -10790
rect -735 -10821 -705 -10790
rect -639 -10816 -609 -10790
rect -543 -10821 -513 -10790
rect -447 -10816 -417 -10790
rect -351 -10821 -321 -10790
rect -255 -10816 -225 -10790
rect -159 -10821 -129 -10790
rect -63 -10816 -33 -10790
rect 33 -10821 63 -10790
rect 129 -10816 159 -10790
rect 225 -10821 255 -10790
rect 321 -10816 351 -10790
rect 417 -10821 447 -10790
rect 513 -10816 543 -10790
rect 609 -10821 639 -10790
rect 705 -10816 735 -10790
rect 801 -10821 831 -10790
rect 897 -10816 927 -10790
rect -945 -10837 -879 -10821
rect -945 -10871 -929 -10837
rect -895 -10871 -879 -10837
rect -945 -10887 -879 -10871
rect -753 -10837 -687 -10821
rect -753 -10871 -737 -10837
rect -703 -10871 -687 -10837
rect -753 -10887 -687 -10871
rect -561 -10837 -495 -10821
rect -561 -10871 -545 -10837
rect -511 -10871 -495 -10837
rect -561 -10887 -495 -10871
rect -369 -10837 -303 -10821
rect -369 -10871 -353 -10837
rect -319 -10871 -303 -10837
rect -369 -10887 -303 -10871
rect -177 -10837 -111 -10821
rect -177 -10871 -161 -10837
rect -127 -10871 -111 -10837
rect -177 -10887 -111 -10871
rect 15 -10837 81 -10821
rect 15 -10871 31 -10837
rect 65 -10871 81 -10837
rect 15 -10887 81 -10871
rect 207 -10837 273 -10821
rect 207 -10871 223 -10837
rect 257 -10871 273 -10837
rect 207 -10887 273 -10871
rect 399 -10837 465 -10821
rect 399 -10871 415 -10837
rect 449 -10871 465 -10837
rect 399 -10887 465 -10871
rect 591 -10837 657 -10821
rect 591 -10871 607 -10837
rect 641 -10871 657 -10837
rect 591 -10887 657 -10871
rect 783 -10837 849 -10821
rect 783 -10871 799 -10837
rect 833 -10871 849 -10837
rect 783 -10887 849 -10871
rect -945 -10945 -879 -10929
rect -945 -10979 -929 -10945
rect -895 -10979 -879 -10945
rect -945 -10995 -879 -10979
rect -753 -10945 -687 -10929
rect -753 -10979 -737 -10945
rect -703 -10979 -687 -10945
rect -753 -10995 -687 -10979
rect -561 -10945 -495 -10929
rect -561 -10979 -545 -10945
rect -511 -10979 -495 -10945
rect -561 -10995 -495 -10979
rect -369 -10945 -303 -10929
rect -369 -10979 -353 -10945
rect -319 -10979 -303 -10945
rect -369 -10995 -303 -10979
rect -177 -10945 -111 -10929
rect -177 -10979 -161 -10945
rect -127 -10979 -111 -10945
rect -177 -10995 -111 -10979
rect 15 -10945 81 -10929
rect 15 -10979 31 -10945
rect 65 -10979 81 -10945
rect 15 -10995 81 -10979
rect 207 -10945 273 -10929
rect 207 -10979 223 -10945
rect 257 -10979 273 -10945
rect 207 -10995 273 -10979
rect 399 -10945 465 -10929
rect 399 -10979 415 -10945
rect 449 -10979 465 -10945
rect 399 -10995 465 -10979
rect 591 -10945 657 -10929
rect 591 -10979 607 -10945
rect 641 -10979 657 -10945
rect 591 -10995 657 -10979
rect 783 -10945 849 -10929
rect 783 -10979 799 -10945
rect 833 -10979 849 -10945
rect 783 -10995 849 -10979
rect -927 -11026 -897 -10995
rect -831 -11026 -801 -11000
rect -735 -11026 -705 -10995
rect -639 -11026 -609 -11000
rect -543 -11026 -513 -10995
rect -447 -11026 -417 -11000
rect -351 -11026 -321 -10995
rect -255 -11026 -225 -11000
rect -159 -11026 -129 -10995
rect -63 -11026 -33 -11000
rect 33 -11026 63 -10995
rect 129 -11026 159 -11000
rect 225 -11026 255 -10995
rect 321 -11026 351 -11000
rect 417 -11026 447 -10995
rect 513 -11026 543 -11000
rect 609 -11026 639 -10995
rect 705 -11026 735 -11000
rect 801 -11026 831 -10995
rect 897 -11026 927 -11000
rect -927 -14452 -897 -14426
rect -831 -14457 -801 -14426
rect -735 -14452 -705 -14426
rect -639 -14457 -609 -14426
rect -543 -14452 -513 -14426
rect -447 -14457 -417 -14426
rect -351 -14452 -321 -14426
rect -255 -14457 -225 -14426
rect -159 -14452 -129 -14426
rect -63 -14457 -33 -14426
rect 33 -14452 63 -14426
rect 129 -14457 159 -14426
rect 225 -14452 255 -14426
rect 321 -14457 351 -14426
rect 417 -14452 447 -14426
rect 513 -14457 543 -14426
rect 609 -14452 639 -14426
rect 705 -14457 735 -14426
rect 801 -14452 831 -14426
rect 897 -14457 927 -14426
rect -849 -14473 -783 -14457
rect -849 -14507 -833 -14473
rect -799 -14507 -783 -14473
rect -849 -14523 -783 -14507
rect -657 -14473 -591 -14457
rect -657 -14507 -641 -14473
rect -607 -14507 -591 -14473
rect -657 -14523 -591 -14507
rect -465 -14473 -399 -14457
rect -465 -14507 -449 -14473
rect -415 -14507 -399 -14473
rect -465 -14523 -399 -14507
rect -273 -14473 -207 -14457
rect -273 -14507 -257 -14473
rect -223 -14507 -207 -14473
rect -273 -14523 -207 -14507
rect -81 -14473 -15 -14457
rect -81 -14507 -65 -14473
rect -31 -14507 -15 -14473
rect -81 -14523 -15 -14507
rect 111 -14473 177 -14457
rect 111 -14507 127 -14473
rect 161 -14507 177 -14473
rect 111 -14523 177 -14507
rect 303 -14473 369 -14457
rect 303 -14507 319 -14473
rect 353 -14507 369 -14473
rect 303 -14523 369 -14507
rect 495 -14473 561 -14457
rect 495 -14507 511 -14473
rect 545 -14507 561 -14473
rect 495 -14523 561 -14507
rect 687 -14473 753 -14457
rect 687 -14507 703 -14473
rect 737 -14507 753 -14473
rect 687 -14523 753 -14507
rect 879 -14473 945 -14457
rect 879 -14507 895 -14473
rect 929 -14507 945 -14473
rect 879 -14523 945 -14507
rect -849 -14581 -783 -14565
rect -849 -14615 -833 -14581
rect -799 -14615 -783 -14581
rect -849 -14631 -783 -14615
rect -657 -14581 -591 -14565
rect -657 -14615 -641 -14581
rect -607 -14615 -591 -14581
rect -657 -14631 -591 -14615
rect -465 -14581 -399 -14565
rect -465 -14615 -449 -14581
rect -415 -14615 -399 -14581
rect -465 -14631 -399 -14615
rect -273 -14581 -207 -14565
rect -273 -14615 -257 -14581
rect -223 -14615 -207 -14581
rect -273 -14631 -207 -14615
rect -81 -14581 -15 -14565
rect -81 -14615 -65 -14581
rect -31 -14615 -15 -14581
rect -81 -14631 -15 -14615
rect 111 -14581 177 -14565
rect 111 -14615 127 -14581
rect 161 -14615 177 -14581
rect 111 -14631 177 -14615
rect 303 -14581 369 -14565
rect 303 -14615 319 -14581
rect 353 -14615 369 -14581
rect 303 -14631 369 -14615
rect 495 -14581 561 -14565
rect 495 -14615 511 -14581
rect 545 -14615 561 -14581
rect 495 -14631 561 -14615
rect 687 -14581 753 -14565
rect 687 -14615 703 -14581
rect 737 -14615 753 -14581
rect 687 -14631 753 -14615
rect 879 -14581 945 -14565
rect 879 -14615 895 -14581
rect 929 -14615 945 -14581
rect 879 -14631 945 -14615
rect -927 -14662 -897 -14636
rect -831 -14662 -801 -14631
rect -735 -14662 -705 -14636
rect -639 -14662 -609 -14631
rect -543 -14662 -513 -14636
rect -447 -14662 -417 -14631
rect -351 -14662 -321 -14636
rect -255 -14662 -225 -14631
rect -159 -14662 -129 -14636
rect -63 -14662 -33 -14631
rect 33 -14662 63 -14636
rect 129 -14662 159 -14631
rect 225 -14662 255 -14636
rect 321 -14662 351 -14631
rect 417 -14662 447 -14636
rect 513 -14662 543 -14631
rect 609 -14662 639 -14636
rect 705 -14662 735 -14631
rect 801 -14662 831 -14636
rect 897 -14662 927 -14631
rect -927 -18093 -897 -18062
rect -831 -18088 -801 -18062
rect -735 -18093 -705 -18062
rect -639 -18088 -609 -18062
rect -543 -18093 -513 -18062
rect -447 -18088 -417 -18062
rect -351 -18093 -321 -18062
rect -255 -18088 -225 -18062
rect -159 -18093 -129 -18062
rect -63 -18088 -33 -18062
rect 33 -18093 63 -18062
rect 129 -18088 159 -18062
rect 225 -18093 255 -18062
rect 321 -18088 351 -18062
rect 417 -18093 447 -18062
rect 513 -18088 543 -18062
rect 609 -18093 639 -18062
rect 705 -18088 735 -18062
rect 801 -18093 831 -18062
rect 897 -18088 927 -18062
rect -945 -18109 -879 -18093
rect -945 -18143 -929 -18109
rect -895 -18143 -879 -18109
rect -945 -18159 -879 -18143
rect -753 -18109 -687 -18093
rect -753 -18143 -737 -18109
rect -703 -18143 -687 -18109
rect -753 -18159 -687 -18143
rect -561 -18109 -495 -18093
rect -561 -18143 -545 -18109
rect -511 -18143 -495 -18109
rect -561 -18159 -495 -18143
rect -369 -18109 -303 -18093
rect -369 -18143 -353 -18109
rect -319 -18143 -303 -18109
rect -369 -18159 -303 -18143
rect -177 -18109 -111 -18093
rect -177 -18143 -161 -18109
rect -127 -18143 -111 -18109
rect -177 -18159 -111 -18143
rect 15 -18109 81 -18093
rect 15 -18143 31 -18109
rect 65 -18143 81 -18109
rect 15 -18159 81 -18143
rect 207 -18109 273 -18093
rect 207 -18143 223 -18109
rect 257 -18143 273 -18109
rect 207 -18159 273 -18143
rect 399 -18109 465 -18093
rect 399 -18143 415 -18109
rect 449 -18143 465 -18109
rect 399 -18159 465 -18143
rect 591 -18109 657 -18093
rect 591 -18143 607 -18109
rect 641 -18143 657 -18109
rect 591 -18159 657 -18143
rect 783 -18109 849 -18093
rect 783 -18143 799 -18109
rect 833 -18143 849 -18109
rect 783 -18159 849 -18143
<< polycont >>
rect -929 18109 -895 18143
rect -737 18109 -703 18143
rect -545 18109 -511 18143
rect -353 18109 -319 18143
rect -161 18109 -127 18143
rect 31 18109 65 18143
rect 223 18109 257 18143
rect 415 18109 449 18143
rect 607 18109 641 18143
rect 799 18109 833 18143
rect -833 14581 -799 14615
rect -641 14581 -607 14615
rect -449 14581 -415 14615
rect -257 14581 -223 14615
rect -65 14581 -31 14615
rect 127 14581 161 14615
rect 319 14581 353 14615
rect 511 14581 545 14615
rect 703 14581 737 14615
rect 895 14581 929 14615
rect -833 14473 -799 14507
rect -641 14473 -607 14507
rect -449 14473 -415 14507
rect -257 14473 -223 14507
rect -65 14473 -31 14507
rect 127 14473 161 14507
rect 319 14473 353 14507
rect 511 14473 545 14507
rect 703 14473 737 14507
rect 895 14473 929 14507
rect -929 10945 -895 10979
rect -737 10945 -703 10979
rect -545 10945 -511 10979
rect -353 10945 -319 10979
rect -161 10945 -127 10979
rect 31 10945 65 10979
rect 223 10945 257 10979
rect 415 10945 449 10979
rect 607 10945 641 10979
rect 799 10945 833 10979
rect -929 10837 -895 10871
rect -737 10837 -703 10871
rect -545 10837 -511 10871
rect -353 10837 -319 10871
rect -161 10837 -127 10871
rect 31 10837 65 10871
rect 223 10837 257 10871
rect 415 10837 449 10871
rect 607 10837 641 10871
rect 799 10837 833 10871
rect -833 7309 -799 7343
rect -641 7309 -607 7343
rect -449 7309 -415 7343
rect -257 7309 -223 7343
rect -65 7309 -31 7343
rect 127 7309 161 7343
rect 319 7309 353 7343
rect 511 7309 545 7343
rect 703 7309 737 7343
rect 895 7309 929 7343
rect -833 7201 -799 7235
rect -641 7201 -607 7235
rect -449 7201 -415 7235
rect -257 7201 -223 7235
rect -65 7201 -31 7235
rect 127 7201 161 7235
rect 319 7201 353 7235
rect 511 7201 545 7235
rect 703 7201 737 7235
rect 895 7201 929 7235
rect -929 3673 -895 3707
rect -737 3673 -703 3707
rect -545 3673 -511 3707
rect -353 3673 -319 3707
rect -161 3673 -127 3707
rect 31 3673 65 3707
rect 223 3673 257 3707
rect 415 3673 449 3707
rect 607 3673 641 3707
rect 799 3673 833 3707
rect -929 3565 -895 3599
rect -737 3565 -703 3599
rect -545 3565 -511 3599
rect -353 3565 -319 3599
rect -161 3565 -127 3599
rect 31 3565 65 3599
rect 223 3565 257 3599
rect 415 3565 449 3599
rect 607 3565 641 3599
rect 799 3565 833 3599
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -929 -3599 -895 -3565
rect -737 -3599 -703 -3565
rect -545 -3599 -511 -3565
rect -353 -3599 -319 -3565
rect -161 -3599 -127 -3565
rect 31 -3599 65 -3565
rect 223 -3599 257 -3565
rect 415 -3599 449 -3565
rect 607 -3599 641 -3565
rect 799 -3599 833 -3565
rect -929 -3707 -895 -3673
rect -737 -3707 -703 -3673
rect -545 -3707 -511 -3673
rect -353 -3707 -319 -3673
rect -161 -3707 -127 -3673
rect 31 -3707 65 -3673
rect 223 -3707 257 -3673
rect 415 -3707 449 -3673
rect 607 -3707 641 -3673
rect 799 -3707 833 -3673
rect -833 -7235 -799 -7201
rect -641 -7235 -607 -7201
rect -449 -7235 -415 -7201
rect -257 -7235 -223 -7201
rect -65 -7235 -31 -7201
rect 127 -7235 161 -7201
rect 319 -7235 353 -7201
rect 511 -7235 545 -7201
rect 703 -7235 737 -7201
rect 895 -7235 929 -7201
rect -833 -7343 -799 -7309
rect -641 -7343 -607 -7309
rect -449 -7343 -415 -7309
rect -257 -7343 -223 -7309
rect -65 -7343 -31 -7309
rect 127 -7343 161 -7309
rect 319 -7343 353 -7309
rect 511 -7343 545 -7309
rect 703 -7343 737 -7309
rect 895 -7343 929 -7309
rect -929 -10871 -895 -10837
rect -737 -10871 -703 -10837
rect -545 -10871 -511 -10837
rect -353 -10871 -319 -10837
rect -161 -10871 -127 -10837
rect 31 -10871 65 -10837
rect 223 -10871 257 -10837
rect 415 -10871 449 -10837
rect 607 -10871 641 -10837
rect 799 -10871 833 -10837
rect -929 -10979 -895 -10945
rect -737 -10979 -703 -10945
rect -545 -10979 -511 -10945
rect -353 -10979 -319 -10945
rect -161 -10979 -127 -10945
rect 31 -10979 65 -10945
rect 223 -10979 257 -10945
rect 415 -10979 449 -10945
rect 607 -10979 641 -10945
rect 799 -10979 833 -10945
rect -833 -14507 -799 -14473
rect -641 -14507 -607 -14473
rect -449 -14507 -415 -14473
rect -257 -14507 -223 -14473
rect -65 -14507 -31 -14473
rect 127 -14507 161 -14473
rect 319 -14507 353 -14473
rect 511 -14507 545 -14473
rect 703 -14507 737 -14473
rect 895 -14507 929 -14473
rect -833 -14615 -799 -14581
rect -641 -14615 -607 -14581
rect -449 -14615 -415 -14581
rect -257 -14615 -223 -14581
rect -65 -14615 -31 -14581
rect 127 -14615 161 -14581
rect 319 -14615 353 -14581
rect 511 -14615 545 -14581
rect 703 -14615 737 -14581
rect 895 -14615 929 -14581
rect -929 -18143 -895 -18109
rect -737 -18143 -703 -18109
rect -545 -18143 -511 -18109
rect -353 -18143 -319 -18109
rect -161 -18143 -127 -18109
rect 31 -18143 65 -18109
rect 223 -18143 257 -18109
rect 415 -18143 449 -18109
rect 607 -18143 641 -18109
rect 799 -18143 833 -18109
<< locali >>
rect -945 18109 -929 18143
rect -895 18109 -879 18143
rect -753 18109 -737 18143
rect -703 18109 -687 18143
rect -561 18109 -545 18143
rect -511 18109 -495 18143
rect -369 18109 -353 18143
rect -319 18109 -303 18143
rect -177 18109 -161 18143
rect -127 18109 -111 18143
rect 15 18109 31 18143
rect 65 18109 81 18143
rect 207 18109 223 18143
rect 257 18109 273 18143
rect 399 18109 415 18143
rect 449 18109 465 18143
rect 591 18109 607 18143
rect 641 18109 657 18143
rect 783 18109 799 18143
rect 833 18109 849 18143
rect -977 18050 -943 18066
rect -977 14658 -943 14674
rect -881 18050 -847 18066
rect -881 14658 -847 14674
rect -785 18050 -751 18066
rect -785 14658 -751 14674
rect -689 18050 -655 18066
rect -689 14658 -655 14674
rect -593 18050 -559 18066
rect -593 14658 -559 14674
rect -497 18050 -463 18066
rect -497 14658 -463 14674
rect -401 18050 -367 18066
rect -401 14658 -367 14674
rect -305 18050 -271 18066
rect -305 14658 -271 14674
rect -209 18050 -175 18066
rect -209 14658 -175 14674
rect -113 18050 -79 18066
rect -113 14658 -79 14674
rect -17 18050 17 18066
rect -17 14658 17 14674
rect 79 18050 113 18066
rect 79 14658 113 14674
rect 175 18050 209 18066
rect 175 14658 209 14674
rect 271 18050 305 18066
rect 271 14658 305 14674
rect 367 18050 401 18066
rect 367 14658 401 14674
rect 463 18050 497 18066
rect 463 14658 497 14674
rect 559 18050 593 18066
rect 559 14658 593 14674
rect 655 18050 689 18066
rect 655 14658 689 14674
rect 751 18050 785 18066
rect 751 14658 785 14674
rect 847 18050 881 18066
rect 847 14658 881 14674
rect 943 18050 977 18066
rect 943 14658 977 14674
rect -849 14581 -833 14615
rect -799 14581 -783 14615
rect -657 14581 -641 14615
rect -607 14581 -591 14615
rect -465 14581 -449 14615
rect -415 14581 -399 14615
rect -273 14581 -257 14615
rect -223 14581 -207 14615
rect -81 14581 -65 14615
rect -31 14581 -15 14615
rect 111 14581 127 14615
rect 161 14581 177 14615
rect 303 14581 319 14615
rect 353 14581 369 14615
rect 495 14581 511 14615
rect 545 14581 561 14615
rect 687 14581 703 14615
rect 737 14581 753 14615
rect 879 14581 895 14615
rect 929 14581 945 14615
rect -849 14473 -833 14507
rect -799 14473 -783 14507
rect -657 14473 -641 14507
rect -607 14473 -591 14507
rect -465 14473 -449 14507
rect -415 14473 -399 14507
rect -273 14473 -257 14507
rect -223 14473 -207 14507
rect -81 14473 -65 14507
rect -31 14473 -15 14507
rect 111 14473 127 14507
rect 161 14473 177 14507
rect 303 14473 319 14507
rect 353 14473 369 14507
rect 495 14473 511 14507
rect 545 14473 561 14507
rect 687 14473 703 14507
rect 737 14473 753 14507
rect 879 14473 895 14507
rect 929 14473 945 14507
rect -977 14414 -943 14430
rect -977 11022 -943 11038
rect -881 14414 -847 14430
rect -881 11022 -847 11038
rect -785 14414 -751 14430
rect -785 11022 -751 11038
rect -689 14414 -655 14430
rect -689 11022 -655 11038
rect -593 14414 -559 14430
rect -593 11022 -559 11038
rect -497 14414 -463 14430
rect -497 11022 -463 11038
rect -401 14414 -367 14430
rect -401 11022 -367 11038
rect -305 14414 -271 14430
rect -305 11022 -271 11038
rect -209 14414 -175 14430
rect -209 11022 -175 11038
rect -113 14414 -79 14430
rect -113 11022 -79 11038
rect -17 14414 17 14430
rect -17 11022 17 11038
rect 79 14414 113 14430
rect 79 11022 113 11038
rect 175 14414 209 14430
rect 175 11022 209 11038
rect 271 14414 305 14430
rect 271 11022 305 11038
rect 367 14414 401 14430
rect 367 11022 401 11038
rect 463 14414 497 14430
rect 463 11022 497 11038
rect 559 14414 593 14430
rect 559 11022 593 11038
rect 655 14414 689 14430
rect 655 11022 689 11038
rect 751 14414 785 14430
rect 751 11022 785 11038
rect 847 14414 881 14430
rect 847 11022 881 11038
rect 943 14414 977 14430
rect 943 11022 977 11038
rect -945 10945 -929 10979
rect -895 10945 -879 10979
rect -753 10945 -737 10979
rect -703 10945 -687 10979
rect -561 10945 -545 10979
rect -511 10945 -495 10979
rect -369 10945 -353 10979
rect -319 10945 -303 10979
rect -177 10945 -161 10979
rect -127 10945 -111 10979
rect 15 10945 31 10979
rect 65 10945 81 10979
rect 207 10945 223 10979
rect 257 10945 273 10979
rect 399 10945 415 10979
rect 449 10945 465 10979
rect 591 10945 607 10979
rect 641 10945 657 10979
rect 783 10945 799 10979
rect 833 10945 849 10979
rect -945 10837 -929 10871
rect -895 10837 -879 10871
rect -753 10837 -737 10871
rect -703 10837 -687 10871
rect -561 10837 -545 10871
rect -511 10837 -495 10871
rect -369 10837 -353 10871
rect -319 10837 -303 10871
rect -177 10837 -161 10871
rect -127 10837 -111 10871
rect 15 10837 31 10871
rect 65 10837 81 10871
rect 207 10837 223 10871
rect 257 10837 273 10871
rect 399 10837 415 10871
rect 449 10837 465 10871
rect 591 10837 607 10871
rect 641 10837 657 10871
rect 783 10837 799 10871
rect 833 10837 849 10871
rect -977 10778 -943 10794
rect -977 7386 -943 7402
rect -881 10778 -847 10794
rect -881 7386 -847 7402
rect -785 10778 -751 10794
rect -785 7386 -751 7402
rect -689 10778 -655 10794
rect -689 7386 -655 7402
rect -593 10778 -559 10794
rect -593 7386 -559 7402
rect -497 10778 -463 10794
rect -497 7386 -463 7402
rect -401 10778 -367 10794
rect -401 7386 -367 7402
rect -305 10778 -271 10794
rect -305 7386 -271 7402
rect -209 10778 -175 10794
rect -209 7386 -175 7402
rect -113 10778 -79 10794
rect -113 7386 -79 7402
rect -17 10778 17 10794
rect -17 7386 17 7402
rect 79 10778 113 10794
rect 79 7386 113 7402
rect 175 10778 209 10794
rect 175 7386 209 7402
rect 271 10778 305 10794
rect 271 7386 305 7402
rect 367 10778 401 10794
rect 367 7386 401 7402
rect 463 10778 497 10794
rect 463 7386 497 7402
rect 559 10778 593 10794
rect 559 7386 593 7402
rect 655 10778 689 10794
rect 655 7386 689 7402
rect 751 10778 785 10794
rect 751 7386 785 7402
rect 847 10778 881 10794
rect 847 7386 881 7402
rect 943 10778 977 10794
rect 943 7386 977 7402
rect -849 7309 -833 7343
rect -799 7309 -783 7343
rect -657 7309 -641 7343
rect -607 7309 -591 7343
rect -465 7309 -449 7343
rect -415 7309 -399 7343
rect -273 7309 -257 7343
rect -223 7309 -207 7343
rect -81 7309 -65 7343
rect -31 7309 -15 7343
rect 111 7309 127 7343
rect 161 7309 177 7343
rect 303 7309 319 7343
rect 353 7309 369 7343
rect 495 7309 511 7343
rect 545 7309 561 7343
rect 687 7309 703 7343
rect 737 7309 753 7343
rect 879 7309 895 7343
rect 929 7309 945 7343
rect -849 7201 -833 7235
rect -799 7201 -783 7235
rect -657 7201 -641 7235
rect -607 7201 -591 7235
rect -465 7201 -449 7235
rect -415 7201 -399 7235
rect -273 7201 -257 7235
rect -223 7201 -207 7235
rect -81 7201 -65 7235
rect -31 7201 -15 7235
rect 111 7201 127 7235
rect 161 7201 177 7235
rect 303 7201 319 7235
rect 353 7201 369 7235
rect 495 7201 511 7235
rect 545 7201 561 7235
rect 687 7201 703 7235
rect 737 7201 753 7235
rect 879 7201 895 7235
rect 929 7201 945 7235
rect -977 7142 -943 7158
rect -977 3750 -943 3766
rect -881 7142 -847 7158
rect -881 3750 -847 3766
rect -785 7142 -751 7158
rect -785 3750 -751 3766
rect -689 7142 -655 7158
rect -689 3750 -655 3766
rect -593 7142 -559 7158
rect -593 3750 -559 3766
rect -497 7142 -463 7158
rect -497 3750 -463 3766
rect -401 7142 -367 7158
rect -401 3750 -367 3766
rect -305 7142 -271 7158
rect -305 3750 -271 3766
rect -209 7142 -175 7158
rect -209 3750 -175 3766
rect -113 7142 -79 7158
rect -113 3750 -79 3766
rect -17 7142 17 7158
rect -17 3750 17 3766
rect 79 7142 113 7158
rect 79 3750 113 3766
rect 175 7142 209 7158
rect 175 3750 209 3766
rect 271 7142 305 7158
rect 271 3750 305 3766
rect 367 7142 401 7158
rect 367 3750 401 3766
rect 463 7142 497 7158
rect 463 3750 497 3766
rect 559 7142 593 7158
rect 559 3750 593 3766
rect 655 7142 689 7158
rect 655 3750 689 3766
rect 751 7142 785 7158
rect 751 3750 785 3766
rect 847 7142 881 7158
rect 847 3750 881 3766
rect 943 7142 977 7158
rect 943 3750 977 3766
rect -945 3673 -929 3707
rect -895 3673 -879 3707
rect -753 3673 -737 3707
rect -703 3673 -687 3707
rect -561 3673 -545 3707
rect -511 3673 -495 3707
rect -369 3673 -353 3707
rect -319 3673 -303 3707
rect -177 3673 -161 3707
rect -127 3673 -111 3707
rect 15 3673 31 3707
rect 65 3673 81 3707
rect 207 3673 223 3707
rect 257 3673 273 3707
rect 399 3673 415 3707
rect 449 3673 465 3707
rect 591 3673 607 3707
rect 641 3673 657 3707
rect 783 3673 799 3707
rect 833 3673 849 3707
rect -945 3565 -929 3599
rect -895 3565 -879 3599
rect -753 3565 -737 3599
rect -703 3565 -687 3599
rect -561 3565 -545 3599
rect -511 3565 -495 3599
rect -369 3565 -353 3599
rect -319 3565 -303 3599
rect -177 3565 -161 3599
rect -127 3565 -111 3599
rect 15 3565 31 3599
rect 65 3565 81 3599
rect 207 3565 223 3599
rect 257 3565 273 3599
rect 399 3565 415 3599
rect 449 3565 465 3599
rect 591 3565 607 3599
rect 641 3565 657 3599
rect 783 3565 799 3599
rect 833 3565 849 3599
rect -977 3506 -943 3522
rect -977 114 -943 130
rect -881 3506 -847 3522
rect -881 114 -847 130
rect -785 3506 -751 3522
rect -785 114 -751 130
rect -689 3506 -655 3522
rect -689 114 -655 130
rect -593 3506 -559 3522
rect -593 114 -559 130
rect -497 3506 -463 3522
rect -497 114 -463 130
rect -401 3506 -367 3522
rect -401 114 -367 130
rect -305 3506 -271 3522
rect -305 114 -271 130
rect -209 3506 -175 3522
rect -209 114 -175 130
rect -113 3506 -79 3522
rect -113 114 -79 130
rect -17 3506 17 3522
rect -17 114 17 130
rect 79 3506 113 3522
rect 79 114 113 130
rect 175 3506 209 3522
rect 175 114 209 130
rect 271 3506 305 3522
rect 271 114 305 130
rect 367 3506 401 3522
rect 367 114 401 130
rect 463 3506 497 3522
rect 463 114 497 130
rect 559 3506 593 3522
rect 559 114 593 130
rect 655 3506 689 3522
rect 655 114 689 130
rect 751 3506 785 3522
rect 751 114 785 130
rect 847 3506 881 3522
rect 847 114 881 130
rect 943 3506 977 3522
rect 943 114 977 130
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect -977 -130 -943 -114
rect -977 -3522 -943 -3506
rect -881 -130 -847 -114
rect -881 -3522 -847 -3506
rect -785 -130 -751 -114
rect -785 -3522 -751 -3506
rect -689 -130 -655 -114
rect -689 -3522 -655 -3506
rect -593 -130 -559 -114
rect -593 -3522 -559 -3506
rect -497 -130 -463 -114
rect -497 -3522 -463 -3506
rect -401 -130 -367 -114
rect -401 -3522 -367 -3506
rect -305 -130 -271 -114
rect -305 -3522 -271 -3506
rect -209 -130 -175 -114
rect -209 -3522 -175 -3506
rect -113 -130 -79 -114
rect -113 -3522 -79 -3506
rect -17 -130 17 -114
rect -17 -3522 17 -3506
rect 79 -130 113 -114
rect 79 -3522 113 -3506
rect 175 -130 209 -114
rect 175 -3522 209 -3506
rect 271 -130 305 -114
rect 271 -3522 305 -3506
rect 367 -130 401 -114
rect 367 -3522 401 -3506
rect 463 -130 497 -114
rect 463 -3522 497 -3506
rect 559 -130 593 -114
rect 559 -3522 593 -3506
rect 655 -130 689 -114
rect 655 -3522 689 -3506
rect 751 -130 785 -114
rect 751 -3522 785 -3506
rect 847 -130 881 -114
rect 847 -3522 881 -3506
rect 943 -130 977 -114
rect 943 -3522 977 -3506
rect -945 -3599 -929 -3565
rect -895 -3599 -879 -3565
rect -753 -3599 -737 -3565
rect -703 -3599 -687 -3565
rect -561 -3599 -545 -3565
rect -511 -3599 -495 -3565
rect -369 -3599 -353 -3565
rect -319 -3599 -303 -3565
rect -177 -3599 -161 -3565
rect -127 -3599 -111 -3565
rect 15 -3599 31 -3565
rect 65 -3599 81 -3565
rect 207 -3599 223 -3565
rect 257 -3599 273 -3565
rect 399 -3599 415 -3565
rect 449 -3599 465 -3565
rect 591 -3599 607 -3565
rect 641 -3599 657 -3565
rect 783 -3599 799 -3565
rect 833 -3599 849 -3565
rect -945 -3707 -929 -3673
rect -895 -3707 -879 -3673
rect -753 -3707 -737 -3673
rect -703 -3707 -687 -3673
rect -561 -3707 -545 -3673
rect -511 -3707 -495 -3673
rect -369 -3707 -353 -3673
rect -319 -3707 -303 -3673
rect -177 -3707 -161 -3673
rect -127 -3707 -111 -3673
rect 15 -3707 31 -3673
rect 65 -3707 81 -3673
rect 207 -3707 223 -3673
rect 257 -3707 273 -3673
rect 399 -3707 415 -3673
rect 449 -3707 465 -3673
rect 591 -3707 607 -3673
rect 641 -3707 657 -3673
rect 783 -3707 799 -3673
rect 833 -3707 849 -3673
rect -977 -3766 -943 -3750
rect -977 -7158 -943 -7142
rect -881 -3766 -847 -3750
rect -881 -7158 -847 -7142
rect -785 -3766 -751 -3750
rect -785 -7158 -751 -7142
rect -689 -3766 -655 -3750
rect -689 -7158 -655 -7142
rect -593 -3766 -559 -3750
rect -593 -7158 -559 -7142
rect -497 -3766 -463 -3750
rect -497 -7158 -463 -7142
rect -401 -3766 -367 -3750
rect -401 -7158 -367 -7142
rect -305 -3766 -271 -3750
rect -305 -7158 -271 -7142
rect -209 -3766 -175 -3750
rect -209 -7158 -175 -7142
rect -113 -3766 -79 -3750
rect -113 -7158 -79 -7142
rect -17 -3766 17 -3750
rect -17 -7158 17 -7142
rect 79 -3766 113 -3750
rect 79 -7158 113 -7142
rect 175 -3766 209 -3750
rect 175 -7158 209 -7142
rect 271 -3766 305 -3750
rect 271 -7158 305 -7142
rect 367 -3766 401 -3750
rect 367 -7158 401 -7142
rect 463 -3766 497 -3750
rect 463 -7158 497 -7142
rect 559 -3766 593 -3750
rect 559 -7158 593 -7142
rect 655 -3766 689 -3750
rect 655 -7158 689 -7142
rect 751 -3766 785 -3750
rect 751 -7158 785 -7142
rect 847 -3766 881 -3750
rect 847 -7158 881 -7142
rect 943 -3766 977 -3750
rect 943 -7158 977 -7142
rect -849 -7235 -833 -7201
rect -799 -7235 -783 -7201
rect -657 -7235 -641 -7201
rect -607 -7235 -591 -7201
rect -465 -7235 -449 -7201
rect -415 -7235 -399 -7201
rect -273 -7235 -257 -7201
rect -223 -7235 -207 -7201
rect -81 -7235 -65 -7201
rect -31 -7235 -15 -7201
rect 111 -7235 127 -7201
rect 161 -7235 177 -7201
rect 303 -7235 319 -7201
rect 353 -7235 369 -7201
rect 495 -7235 511 -7201
rect 545 -7235 561 -7201
rect 687 -7235 703 -7201
rect 737 -7235 753 -7201
rect 879 -7235 895 -7201
rect 929 -7235 945 -7201
rect -849 -7343 -833 -7309
rect -799 -7343 -783 -7309
rect -657 -7343 -641 -7309
rect -607 -7343 -591 -7309
rect -465 -7343 -449 -7309
rect -415 -7343 -399 -7309
rect -273 -7343 -257 -7309
rect -223 -7343 -207 -7309
rect -81 -7343 -65 -7309
rect -31 -7343 -15 -7309
rect 111 -7343 127 -7309
rect 161 -7343 177 -7309
rect 303 -7343 319 -7309
rect 353 -7343 369 -7309
rect 495 -7343 511 -7309
rect 545 -7343 561 -7309
rect 687 -7343 703 -7309
rect 737 -7343 753 -7309
rect 879 -7343 895 -7309
rect 929 -7343 945 -7309
rect -977 -7402 -943 -7386
rect -977 -10794 -943 -10778
rect -881 -7402 -847 -7386
rect -881 -10794 -847 -10778
rect -785 -7402 -751 -7386
rect -785 -10794 -751 -10778
rect -689 -7402 -655 -7386
rect -689 -10794 -655 -10778
rect -593 -7402 -559 -7386
rect -593 -10794 -559 -10778
rect -497 -7402 -463 -7386
rect -497 -10794 -463 -10778
rect -401 -7402 -367 -7386
rect -401 -10794 -367 -10778
rect -305 -7402 -271 -7386
rect -305 -10794 -271 -10778
rect -209 -7402 -175 -7386
rect -209 -10794 -175 -10778
rect -113 -7402 -79 -7386
rect -113 -10794 -79 -10778
rect -17 -7402 17 -7386
rect -17 -10794 17 -10778
rect 79 -7402 113 -7386
rect 79 -10794 113 -10778
rect 175 -7402 209 -7386
rect 175 -10794 209 -10778
rect 271 -7402 305 -7386
rect 271 -10794 305 -10778
rect 367 -7402 401 -7386
rect 367 -10794 401 -10778
rect 463 -7402 497 -7386
rect 463 -10794 497 -10778
rect 559 -7402 593 -7386
rect 559 -10794 593 -10778
rect 655 -7402 689 -7386
rect 655 -10794 689 -10778
rect 751 -7402 785 -7386
rect 751 -10794 785 -10778
rect 847 -7402 881 -7386
rect 847 -10794 881 -10778
rect 943 -7402 977 -7386
rect 943 -10794 977 -10778
rect -945 -10871 -929 -10837
rect -895 -10871 -879 -10837
rect -753 -10871 -737 -10837
rect -703 -10871 -687 -10837
rect -561 -10871 -545 -10837
rect -511 -10871 -495 -10837
rect -369 -10871 -353 -10837
rect -319 -10871 -303 -10837
rect -177 -10871 -161 -10837
rect -127 -10871 -111 -10837
rect 15 -10871 31 -10837
rect 65 -10871 81 -10837
rect 207 -10871 223 -10837
rect 257 -10871 273 -10837
rect 399 -10871 415 -10837
rect 449 -10871 465 -10837
rect 591 -10871 607 -10837
rect 641 -10871 657 -10837
rect 783 -10871 799 -10837
rect 833 -10871 849 -10837
rect -945 -10979 -929 -10945
rect -895 -10979 -879 -10945
rect -753 -10979 -737 -10945
rect -703 -10979 -687 -10945
rect -561 -10979 -545 -10945
rect -511 -10979 -495 -10945
rect -369 -10979 -353 -10945
rect -319 -10979 -303 -10945
rect -177 -10979 -161 -10945
rect -127 -10979 -111 -10945
rect 15 -10979 31 -10945
rect 65 -10979 81 -10945
rect 207 -10979 223 -10945
rect 257 -10979 273 -10945
rect 399 -10979 415 -10945
rect 449 -10979 465 -10945
rect 591 -10979 607 -10945
rect 641 -10979 657 -10945
rect 783 -10979 799 -10945
rect 833 -10979 849 -10945
rect -977 -11038 -943 -11022
rect -977 -14430 -943 -14414
rect -881 -11038 -847 -11022
rect -881 -14430 -847 -14414
rect -785 -11038 -751 -11022
rect -785 -14430 -751 -14414
rect -689 -11038 -655 -11022
rect -689 -14430 -655 -14414
rect -593 -11038 -559 -11022
rect -593 -14430 -559 -14414
rect -497 -11038 -463 -11022
rect -497 -14430 -463 -14414
rect -401 -11038 -367 -11022
rect -401 -14430 -367 -14414
rect -305 -11038 -271 -11022
rect -305 -14430 -271 -14414
rect -209 -11038 -175 -11022
rect -209 -14430 -175 -14414
rect -113 -11038 -79 -11022
rect -113 -14430 -79 -14414
rect -17 -11038 17 -11022
rect -17 -14430 17 -14414
rect 79 -11038 113 -11022
rect 79 -14430 113 -14414
rect 175 -11038 209 -11022
rect 175 -14430 209 -14414
rect 271 -11038 305 -11022
rect 271 -14430 305 -14414
rect 367 -11038 401 -11022
rect 367 -14430 401 -14414
rect 463 -11038 497 -11022
rect 463 -14430 497 -14414
rect 559 -11038 593 -11022
rect 559 -14430 593 -14414
rect 655 -11038 689 -11022
rect 655 -14430 689 -14414
rect 751 -11038 785 -11022
rect 751 -14430 785 -14414
rect 847 -11038 881 -11022
rect 847 -14430 881 -14414
rect 943 -11038 977 -11022
rect 943 -14430 977 -14414
rect -849 -14507 -833 -14473
rect -799 -14507 -783 -14473
rect -657 -14507 -641 -14473
rect -607 -14507 -591 -14473
rect -465 -14507 -449 -14473
rect -415 -14507 -399 -14473
rect -273 -14507 -257 -14473
rect -223 -14507 -207 -14473
rect -81 -14507 -65 -14473
rect -31 -14507 -15 -14473
rect 111 -14507 127 -14473
rect 161 -14507 177 -14473
rect 303 -14507 319 -14473
rect 353 -14507 369 -14473
rect 495 -14507 511 -14473
rect 545 -14507 561 -14473
rect 687 -14507 703 -14473
rect 737 -14507 753 -14473
rect 879 -14507 895 -14473
rect 929 -14507 945 -14473
rect -849 -14615 -833 -14581
rect -799 -14615 -783 -14581
rect -657 -14615 -641 -14581
rect -607 -14615 -591 -14581
rect -465 -14615 -449 -14581
rect -415 -14615 -399 -14581
rect -273 -14615 -257 -14581
rect -223 -14615 -207 -14581
rect -81 -14615 -65 -14581
rect -31 -14615 -15 -14581
rect 111 -14615 127 -14581
rect 161 -14615 177 -14581
rect 303 -14615 319 -14581
rect 353 -14615 369 -14581
rect 495 -14615 511 -14581
rect 545 -14615 561 -14581
rect 687 -14615 703 -14581
rect 737 -14615 753 -14581
rect 879 -14615 895 -14581
rect 929 -14615 945 -14581
rect -977 -14674 -943 -14658
rect -977 -18066 -943 -18050
rect -881 -14674 -847 -14658
rect -881 -18066 -847 -18050
rect -785 -14674 -751 -14658
rect -785 -18066 -751 -18050
rect -689 -14674 -655 -14658
rect -689 -18066 -655 -18050
rect -593 -14674 -559 -14658
rect -593 -18066 -559 -18050
rect -497 -14674 -463 -14658
rect -497 -18066 -463 -18050
rect -401 -14674 -367 -14658
rect -401 -18066 -367 -18050
rect -305 -14674 -271 -14658
rect -305 -18066 -271 -18050
rect -209 -14674 -175 -14658
rect -209 -18066 -175 -18050
rect -113 -14674 -79 -14658
rect -113 -18066 -79 -18050
rect -17 -14674 17 -14658
rect -17 -18066 17 -18050
rect 79 -14674 113 -14658
rect 79 -18066 113 -18050
rect 175 -14674 209 -14658
rect 175 -18066 209 -18050
rect 271 -14674 305 -14658
rect 271 -18066 305 -18050
rect 367 -14674 401 -14658
rect 367 -18066 401 -18050
rect 463 -14674 497 -14658
rect 463 -18066 497 -18050
rect 559 -14674 593 -14658
rect 559 -18066 593 -18050
rect 655 -14674 689 -14658
rect 655 -18066 689 -18050
rect 751 -14674 785 -14658
rect 751 -18066 785 -18050
rect 847 -14674 881 -14658
rect 847 -18066 881 -18050
rect 943 -14674 977 -14658
rect 943 -18066 977 -18050
rect -945 -18143 -929 -18109
rect -895 -18143 -879 -18109
rect -753 -18143 -737 -18109
rect -703 -18143 -687 -18109
rect -561 -18143 -545 -18109
rect -511 -18143 -495 -18109
rect -369 -18143 -353 -18109
rect -319 -18143 -303 -18109
rect -177 -18143 -161 -18109
rect -127 -18143 -111 -18109
rect 15 -18143 31 -18109
rect 65 -18143 81 -18109
rect 207 -18143 223 -18109
rect 257 -18143 273 -18109
rect 399 -18143 415 -18109
rect 449 -18143 465 -18109
rect 591 -18143 607 -18109
rect 641 -18143 657 -18109
rect 783 -18143 799 -18109
rect 833 -18143 849 -18109
<< viali >>
rect -929 18109 -895 18143
rect -737 18109 -703 18143
rect -545 18109 -511 18143
rect -353 18109 -319 18143
rect -161 18109 -127 18143
rect 31 18109 65 18143
rect 223 18109 257 18143
rect 415 18109 449 18143
rect 607 18109 641 18143
rect 799 18109 833 18143
rect -977 14674 -943 18050
rect -881 14674 -847 18050
rect -785 14674 -751 18050
rect -689 14674 -655 18050
rect -593 14674 -559 18050
rect -497 14674 -463 18050
rect -401 14674 -367 18050
rect -305 14674 -271 18050
rect -209 14674 -175 18050
rect -113 14674 -79 18050
rect -17 14674 17 18050
rect 79 14674 113 18050
rect 175 14674 209 18050
rect 271 14674 305 18050
rect 367 14674 401 18050
rect 463 14674 497 18050
rect 559 14674 593 18050
rect 655 14674 689 18050
rect 751 14674 785 18050
rect 847 14674 881 18050
rect 943 14674 977 18050
rect -833 14581 -799 14615
rect -641 14581 -607 14615
rect -449 14581 -415 14615
rect -257 14581 -223 14615
rect -65 14581 -31 14615
rect 127 14581 161 14615
rect 319 14581 353 14615
rect 511 14581 545 14615
rect 703 14581 737 14615
rect 895 14581 929 14615
rect -833 14473 -799 14507
rect -641 14473 -607 14507
rect -449 14473 -415 14507
rect -257 14473 -223 14507
rect -65 14473 -31 14507
rect 127 14473 161 14507
rect 319 14473 353 14507
rect 511 14473 545 14507
rect 703 14473 737 14507
rect 895 14473 929 14507
rect -977 11038 -943 14414
rect -881 11038 -847 14414
rect -785 11038 -751 14414
rect -689 11038 -655 14414
rect -593 11038 -559 14414
rect -497 11038 -463 14414
rect -401 11038 -367 14414
rect -305 11038 -271 14414
rect -209 11038 -175 14414
rect -113 11038 -79 14414
rect -17 11038 17 14414
rect 79 11038 113 14414
rect 175 11038 209 14414
rect 271 11038 305 14414
rect 367 11038 401 14414
rect 463 11038 497 14414
rect 559 11038 593 14414
rect 655 11038 689 14414
rect 751 11038 785 14414
rect 847 11038 881 14414
rect 943 11038 977 14414
rect -929 10945 -895 10979
rect -737 10945 -703 10979
rect -545 10945 -511 10979
rect -353 10945 -319 10979
rect -161 10945 -127 10979
rect 31 10945 65 10979
rect 223 10945 257 10979
rect 415 10945 449 10979
rect 607 10945 641 10979
rect 799 10945 833 10979
rect -929 10837 -895 10871
rect -737 10837 -703 10871
rect -545 10837 -511 10871
rect -353 10837 -319 10871
rect -161 10837 -127 10871
rect 31 10837 65 10871
rect 223 10837 257 10871
rect 415 10837 449 10871
rect 607 10837 641 10871
rect 799 10837 833 10871
rect -977 7402 -943 10778
rect -881 7402 -847 10778
rect -785 7402 -751 10778
rect -689 7402 -655 10778
rect -593 7402 -559 10778
rect -497 7402 -463 10778
rect -401 7402 -367 10778
rect -305 7402 -271 10778
rect -209 7402 -175 10778
rect -113 7402 -79 10778
rect -17 7402 17 10778
rect 79 7402 113 10778
rect 175 7402 209 10778
rect 271 7402 305 10778
rect 367 7402 401 10778
rect 463 7402 497 10778
rect 559 7402 593 10778
rect 655 7402 689 10778
rect 751 7402 785 10778
rect 847 7402 881 10778
rect 943 7402 977 10778
rect -833 7309 -799 7343
rect -641 7309 -607 7343
rect -449 7309 -415 7343
rect -257 7309 -223 7343
rect -65 7309 -31 7343
rect 127 7309 161 7343
rect 319 7309 353 7343
rect 511 7309 545 7343
rect 703 7309 737 7343
rect 895 7309 929 7343
rect -833 7201 -799 7235
rect -641 7201 -607 7235
rect -449 7201 -415 7235
rect -257 7201 -223 7235
rect -65 7201 -31 7235
rect 127 7201 161 7235
rect 319 7201 353 7235
rect 511 7201 545 7235
rect 703 7201 737 7235
rect 895 7201 929 7235
rect -977 3766 -943 7142
rect -881 3766 -847 7142
rect -785 3766 -751 7142
rect -689 3766 -655 7142
rect -593 3766 -559 7142
rect -497 3766 -463 7142
rect -401 3766 -367 7142
rect -305 3766 -271 7142
rect -209 3766 -175 7142
rect -113 3766 -79 7142
rect -17 3766 17 7142
rect 79 3766 113 7142
rect 175 3766 209 7142
rect 271 3766 305 7142
rect 367 3766 401 7142
rect 463 3766 497 7142
rect 559 3766 593 7142
rect 655 3766 689 7142
rect 751 3766 785 7142
rect 847 3766 881 7142
rect 943 3766 977 7142
rect -929 3673 -895 3707
rect -737 3673 -703 3707
rect -545 3673 -511 3707
rect -353 3673 -319 3707
rect -161 3673 -127 3707
rect 31 3673 65 3707
rect 223 3673 257 3707
rect 415 3673 449 3707
rect 607 3673 641 3707
rect 799 3673 833 3707
rect -929 3565 -895 3599
rect -737 3565 -703 3599
rect -545 3565 -511 3599
rect -353 3565 -319 3599
rect -161 3565 -127 3599
rect 31 3565 65 3599
rect 223 3565 257 3599
rect 415 3565 449 3599
rect 607 3565 641 3599
rect 799 3565 833 3599
rect -977 130 -943 3506
rect -881 130 -847 3506
rect -785 130 -751 3506
rect -689 130 -655 3506
rect -593 130 -559 3506
rect -497 130 -463 3506
rect -401 130 -367 3506
rect -305 130 -271 3506
rect -209 130 -175 3506
rect -113 130 -79 3506
rect -17 130 17 3506
rect 79 130 113 3506
rect 175 130 209 3506
rect 271 130 305 3506
rect 367 130 401 3506
rect 463 130 497 3506
rect 559 130 593 3506
rect 655 130 689 3506
rect 751 130 785 3506
rect 847 130 881 3506
rect 943 130 977 3506
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -977 -3506 -943 -130
rect -881 -3506 -847 -130
rect -785 -3506 -751 -130
rect -689 -3506 -655 -130
rect -593 -3506 -559 -130
rect -497 -3506 -463 -130
rect -401 -3506 -367 -130
rect -305 -3506 -271 -130
rect -209 -3506 -175 -130
rect -113 -3506 -79 -130
rect -17 -3506 17 -130
rect 79 -3506 113 -130
rect 175 -3506 209 -130
rect 271 -3506 305 -130
rect 367 -3506 401 -130
rect 463 -3506 497 -130
rect 559 -3506 593 -130
rect 655 -3506 689 -130
rect 751 -3506 785 -130
rect 847 -3506 881 -130
rect 943 -3506 977 -130
rect -929 -3599 -895 -3565
rect -737 -3599 -703 -3565
rect -545 -3599 -511 -3565
rect -353 -3599 -319 -3565
rect -161 -3599 -127 -3565
rect 31 -3599 65 -3565
rect 223 -3599 257 -3565
rect 415 -3599 449 -3565
rect 607 -3599 641 -3565
rect 799 -3599 833 -3565
rect -929 -3707 -895 -3673
rect -737 -3707 -703 -3673
rect -545 -3707 -511 -3673
rect -353 -3707 -319 -3673
rect -161 -3707 -127 -3673
rect 31 -3707 65 -3673
rect 223 -3707 257 -3673
rect 415 -3707 449 -3673
rect 607 -3707 641 -3673
rect 799 -3707 833 -3673
rect -977 -7142 -943 -3766
rect -881 -7142 -847 -3766
rect -785 -7142 -751 -3766
rect -689 -7142 -655 -3766
rect -593 -7142 -559 -3766
rect -497 -7142 -463 -3766
rect -401 -7142 -367 -3766
rect -305 -7142 -271 -3766
rect -209 -7142 -175 -3766
rect -113 -7142 -79 -3766
rect -17 -7142 17 -3766
rect 79 -7142 113 -3766
rect 175 -7142 209 -3766
rect 271 -7142 305 -3766
rect 367 -7142 401 -3766
rect 463 -7142 497 -3766
rect 559 -7142 593 -3766
rect 655 -7142 689 -3766
rect 751 -7142 785 -3766
rect 847 -7142 881 -3766
rect 943 -7142 977 -3766
rect -833 -7235 -799 -7201
rect -641 -7235 -607 -7201
rect -449 -7235 -415 -7201
rect -257 -7235 -223 -7201
rect -65 -7235 -31 -7201
rect 127 -7235 161 -7201
rect 319 -7235 353 -7201
rect 511 -7235 545 -7201
rect 703 -7235 737 -7201
rect 895 -7235 929 -7201
rect -833 -7343 -799 -7309
rect -641 -7343 -607 -7309
rect -449 -7343 -415 -7309
rect -257 -7343 -223 -7309
rect -65 -7343 -31 -7309
rect 127 -7343 161 -7309
rect 319 -7343 353 -7309
rect 511 -7343 545 -7309
rect 703 -7343 737 -7309
rect 895 -7343 929 -7309
rect -977 -10778 -943 -7402
rect -881 -10778 -847 -7402
rect -785 -10778 -751 -7402
rect -689 -10778 -655 -7402
rect -593 -10778 -559 -7402
rect -497 -10778 -463 -7402
rect -401 -10778 -367 -7402
rect -305 -10778 -271 -7402
rect -209 -10778 -175 -7402
rect -113 -10778 -79 -7402
rect -17 -10778 17 -7402
rect 79 -10778 113 -7402
rect 175 -10778 209 -7402
rect 271 -10778 305 -7402
rect 367 -10778 401 -7402
rect 463 -10778 497 -7402
rect 559 -10778 593 -7402
rect 655 -10778 689 -7402
rect 751 -10778 785 -7402
rect 847 -10778 881 -7402
rect 943 -10778 977 -7402
rect -929 -10871 -895 -10837
rect -737 -10871 -703 -10837
rect -545 -10871 -511 -10837
rect -353 -10871 -319 -10837
rect -161 -10871 -127 -10837
rect 31 -10871 65 -10837
rect 223 -10871 257 -10837
rect 415 -10871 449 -10837
rect 607 -10871 641 -10837
rect 799 -10871 833 -10837
rect -929 -10979 -895 -10945
rect -737 -10979 -703 -10945
rect -545 -10979 -511 -10945
rect -353 -10979 -319 -10945
rect -161 -10979 -127 -10945
rect 31 -10979 65 -10945
rect 223 -10979 257 -10945
rect 415 -10979 449 -10945
rect 607 -10979 641 -10945
rect 799 -10979 833 -10945
rect -977 -14414 -943 -11038
rect -881 -14414 -847 -11038
rect -785 -14414 -751 -11038
rect -689 -14414 -655 -11038
rect -593 -14414 -559 -11038
rect -497 -14414 -463 -11038
rect -401 -14414 -367 -11038
rect -305 -14414 -271 -11038
rect -209 -14414 -175 -11038
rect -113 -14414 -79 -11038
rect -17 -14414 17 -11038
rect 79 -14414 113 -11038
rect 175 -14414 209 -11038
rect 271 -14414 305 -11038
rect 367 -14414 401 -11038
rect 463 -14414 497 -11038
rect 559 -14414 593 -11038
rect 655 -14414 689 -11038
rect 751 -14414 785 -11038
rect 847 -14414 881 -11038
rect 943 -14414 977 -11038
rect -833 -14507 -799 -14473
rect -641 -14507 -607 -14473
rect -449 -14507 -415 -14473
rect -257 -14507 -223 -14473
rect -65 -14507 -31 -14473
rect 127 -14507 161 -14473
rect 319 -14507 353 -14473
rect 511 -14507 545 -14473
rect 703 -14507 737 -14473
rect 895 -14507 929 -14473
rect -833 -14615 -799 -14581
rect -641 -14615 -607 -14581
rect -449 -14615 -415 -14581
rect -257 -14615 -223 -14581
rect -65 -14615 -31 -14581
rect 127 -14615 161 -14581
rect 319 -14615 353 -14581
rect 511 -14615 545 -14581
rect 703 -14615 737 -14581
rect 895 -14615 929 -14581
rect -977 -18050 -943 -14674
rect -881 -18050 -847 -14674
rect -785 -18050 -751 -14674
rect -689 -18050 -655 -14674
rect -593 -18050 -559 -14674
rect -497 -18050 -463 -14674
rect -401 -18050 -367 -14674
rect -305 -18050 -271 -14674
rect -209 -18050 -175 -14674
rect -113 -18050 -79 -14674
rect -17 -18050 17 -14674
rect 79 -18050 113 -14674
rect 175 -18050 209 -14674
rect 271 -18050 305 -14674
rect 367 -18050 401 -14674
rect 463 -18050 497 -14674
rect 559 -18050 593 -14674
rect 655 -18050 689 -14674
rect 751 -18050 785 -14674
rect 847 -18050 881 -14674
rect 943 -18050 977 -14674
rect -929 -18143 -895 -18109
rect -737 -18143 -703 -18109
rect -545 -18143 -511 -18109
rect -353 -18143 -319 -18109
rect -161 -18143 -127 -18109
rect 31 -18143 65 -18109
rect 223 -18143 257 -18109
rect 415 -18143 449 -18109
rect 607 -18143 641 -18109
rect 799 -18143 833 -18109
<< metal1 >>
rect -941 18143 -883 18149
rect -941 18109 -929 18143
rect -895 18109 -883 18143
rect -941 18103 -883 18109
rect -749 18143 -691 18149
rect -749 18109 -737 18143
rect -703 18109 -691 18143
rect -749 18103 -691 18109
rect -557 18143 -499 18149
rect -557 18109 -545 18143
rect -511 18109 -499 18143
rect -557 18103 -499 18109
rect -365 18143 -307 18149
rect -365 18109 -353 18143
rect -319 18109 -307 18143
rect -365 18103 -307 18109
rect -173 18143 -115 18149
rect -173 18109 -161 18143
rect -127 18109 -115 18143
rect -173 18103 -115 18109
rect 19 18143 77 18149
rect 19 18109 31 18143
rect 65 18109 77 18143
rect 19 18103 77 18109
rect 211 18143 269 18149
rect 211 18109 223 18143
rect 257 18109 269 18143
rect 211 18103 269 18109
rect 403 18143 461 18149
rect 403 18109 415 18143
rect 449 18109 461 18143
rect 403 18103 461 18109
rect 595 18143 653 18149
rect 595 18109 607 18143
rect 641 18109 653 18143
rect 595 18103 653 18109
rect 787 18143 845 18149
rect 787 18109 799 18143
rect 833 18109 845 18143
rect 787 18103 845 18109
rect -983 18050 -937 18062
rect -983 14674 -977 18050
rect -943 14674 -937 18050
rect -983 14662 -937 14674
rect -887 18050 -841 18062
rect -887 14674 -881 18050
rect -847 14674 -841 18050
rect -887 14662 -841 14674
rect -791 18050 -745 18062
rect -791 14674 -785 18050
rect -751 14674 -745 18050
rect -791 14662 -745 14674
rect -695 18050 -649 18062
rect -695 14674 -689 18050
rect -655 14674 -649 18050
rect -695 14662 -649 14674
rect -599 18050 -553 18062
rect -599 14674 -593 18050
rect -559 14674 -553 18050
rect -599 14662 -553 14674
rect -503 18050 -457 18062
rect -503 14674 -497 18050
rect -463 14674 -457 18050
rect -503 14662 -457 14674
rect -407 18050 -361 18062
rect -407 14674 -401 18050
rect -367 14674 -361 18050
rect -407 14662 -361 14674
rect -311 18050 -265 18062
rect -311 14674 -305 18050
rect -271 14674 -265 18050
rect -311 14662 -265 14674
rect -215 18050 -169 18062
rect -215 14674 -209 18050
rect -175 14674 -169 18050
rect -215 14662 -169 14674
rect -119 18050 -73 18062
rect -119 14674 -113 18050
rect -79 14674 -73 18050
rect -119 14662 -73 14674
rect -23 18050 23 18062
rect -23 14674 -17 18050
rect 17 14674 23 18050
rect -23 14662 23 14674
rect 73 18050 119 18062
rect 73 14674 79 18050
rect 113 14674 119 18050
rect 73 14662 119 14674
rect 169 18050 215 18062
rect 169 14674 175 18050
rect 209 14674 215 18050
rect 169 14662 215 14674
rect 265 18050 311 18062
rect 265 14674 271 18050
rect 305 14674 311 18050
rect 265 14662 311 14674
rect 361 18050 407 18062
rect 361 14674 367 18050
rect 401 14674 407 18050
rect 361 14662 407 14674
rect 457 18050 503 18062
rect 457 14674 463 18050
rect 497 14674 503 18050
rect 457 14662 503 14674
rect 553 18050 599 18062
rect 553 14674 559 18050
rect 593 14674 599 18050
rect 553 14662 599 14674
rect 649 18050 695 18062
rect 649 14674 655 18050
rect 689 14674 695 18050
rect 649 14662 695 14674
rect 745 18050 791 18062
rect 745 14674 751 18050
rect 785 14674 791 18050
rect 745 14662 791 14674
rect 841 18050 887 18062
rect 841 14674 847 18050
rect 881 14674 887 18050
rect 841 14662 887 14674
rect 937 18050 983 18062
rect 937 14674 943 18050
rect 977 14674 983 18050
rect 937 14662 983 14674
rect -845 14615 -787 14621
rect -845 14581 -833 14615
rect -799 14581 -787 14615
rect -845 14575 -787 14581
rect -653 14615 -595 14621
rect -653 14581 -641 14615
rect -607 14581 -595 14615
rect -653 14575 -595 14581
rect -461 14615 -403 14621
rect -461 14581 -449 14615
rect -415 14581 -403 14615
rect -461 14575 -403 14581
rect -269 14615 -211 14621
rect -269 14581 -257 14615
rect -223 14581 -211 14615
rect -269 14575 -211 14581
rect -77 14615 -19 14621
rect -77 14581 -65 14615
rect -31 14581 -19 14615
rect -77 14575 -19 14581
rect 115 14615 173 14621
rect 115 14581 127 14615
rect 161 14581 173 14615
rect 115 14575 173 14581
rect 307 14615 365 14621
rect 307 14581 319 14615
rect 353 14581 365 14615
rect 307 14575 365 14581
rect 499 14615 557 14621
rect 499 14581 511 14615
rect 545 14581 557 14615
rect 499 14575 557 14581
rect 691 14615 749 14621
rect 691 14581 703 14615
rect 737 14581 749 14615
rect 691 14575 749 14581
rect 883 14615 941 14621
rect 883 14581 895 14615
rect 929 14581 941 14615
rect 883 14575 941 14581
rect -845 14507 -787 14513
rect -845 14473 -833 14507
rect -799 14473 -787 14507
rect -845 14467 -787 14473
rect -653 14507 -595 14513
rect -653 14473 -641 14507
rect -607 14473 -595 14507
rect -653 14467 -595 14473
rect -461 14507 -403 14513
rect -461 14473 -449 14507
rect -415 14473 -403 14507
rect -461 14467 -403 14473
rect -269 14507 -211 14513
rect -269 14473 -257 14507
rect -223 14473 -211 14507
rect -269 14467 -211 14473
rect -77 14507 -19 14513
rect -77 14473 -65 14507
rect -31 14473 -19 14507
rect -77 14467 -19 14473
rect 115 14507 173 14513
rect 115 14473 127 14507
rect 161 14473 173 14507
rect 115 14467 173 14473
rect 307 14507 365 14513
rect 307 14473 319 14507
rect 353 14473 365 14507
rect 307 14467 365 14473
rect 499 14507 557 14513
rect 499 14473 511 14507
rect 545 14473 557 14507
rect 499 14467 557 14473
rect 691 14507 749 14513
rect 691 14473 703 14507
rect 737 14473 749 14507
rect 691 14467 749 14473
rect 883 14507 941 14513
rect 883 14473 895 14507
rect 929 14473 941 14507
rect 883 14467 941 14473
rect -983 14414 -937 14426
rect -983 11038 -977 14414
rect -943 11038 -937 14414
rect -983 11026 -937 11038
rect -887 14414 -841 14426
rect -887 11038 -881 14414
rect -847 11038 -841 14414
rect -887 11026 -841 11038
rect -791 14414 -745 14426
rect -791 11038 -785 14414
rect -751 11038 -745 14414
rect -791 11026 -745 11038
rect -695 14414 -649 14426
rect -695 11038 -689 14414
rect -655 11038 -649 14414
rect -695 11026 -649 11038
rect -599 14414 -553 14426
rect -599 11038 -593 14414
rect -559 11038 -553 14414
rect -599 11026 -553 11038
rect -503 14414 -457 14426
rect -503 11038 -497 14414
rect -463 11038 -457 14414
rect -503 11026 -457 11038
rect -407 14414 -361 14426
rect -407 11038 -401 14414
rect -367 11038 -361 14414
rect -407 11026 -361 11038
rect -311 14414 -265 14426
rect -311 11038 -305 14414
rect -271 11038 -265 14414
rect -311 11026 -265 11038
rect -215 14414 -169 14426
rect -215 11038 -209 14414
rect -175 11038 -169 14414
rect -215 11026 -169 11038
rect -119 14414 -73 14426
rect -119 11038 -113 14414
rect -79 11038 -73 14414
rect -119 11026 -73 11038
rect -23 14414 23 14426
rect -23 11038 -17 14414
rect 17 11038 23 14414
rect -23 11026 23 11038
rect 73 14414 119 14426
rect 73 11038 79 14414
rect 113 11038 119 14414
rect 73 11026 119 11038
rect 169 14414 215 14426
rect 169 11038 175 14414
rect 209 11038 215 14414
rect 169 11026 215 11038
rect 265 14414 311 14426
rect 265 11038 271 14414
rect 305 11038 311 14414
rect 265 11026 311 11038
rect 361 14414 407 14426
rect 361 11038 367 14414
rect 401 11038 407 14414
rect 361 11026 407 11038
rect 457 14414 503 14426
rect 457 11038 463 14414
rect 497 11038 503 14414
rect 457 11026 503 11038
rect 553 14414 599 14426
rect 553 11038 559 14414
rect 593 11038 599 14414
rect 553 11026 599 11038
rect 649 14414 695 14426
rect 649 11038 655 14414
rect 689 11038 695 14414
rect 649 11026 695 11038
rect 745 14414 791 14426
rect 745 11038 751 14414
rect 785 11038 791 14414
rect 745 11026 791 11038
rect 841 14414 887 14426
rect 841 11038 847 14414
rect 881 11038 887 14414
rect 841 11026 887 11038
rect 937 14414 983 14426
rect 937 11038 943 14414
rect 977 11038 983 14414
rect 937 11026 983 11038
rect -941 10979 -883 10985
rect -941 10945 -929 10979
rect -895 10945 -883 10979
rect -941 10939 -883 10945
rect -749 10979 -691 10985
rect -749 10945 -737 10979
rect -703 10945 -691 10979
rect -749 10939 -691 10945
rect -557 10979 -499 10985
rect -557 10945 -545 10979
rect -511 10945 -499 10979
rect -557 10939 -499 10945
rect -365 10979 -307 10985
rect -365 10945 -353 10979
rect -319 10945 -307 10979
rect -365 10939 -307 10945
rect -173 10979 -115 10985
rect -173 10945 -161 10979
rect -127 10945 -115 10979
rect -173 10939 -115 10945
rect 19 10979 77 10985
rect 19 10945 31 10979
rect 65 10945 77 10979
rect 19 10939 77 10945
rect 211 10979 269 10985
rect 211 10945 223 10979
rect 257 10945 269 10979
rect 211 10939 269 10945
rect 403 10979 461 10985
rect 403 10945 415 10979
rect 449 10945 461 10979
rect 403 10939 461 10945
rect 595 10979 653 10985
rect 595 10945 607 10979
rect 641 10945 653 10979
rect 595 10939 653 10945
rect 787 10979 845 10985
rect 787 10945 799 10979
rect 833 10945 845 10979
rect 787 10939 845 10945
rect -941 10871 -883 10877
rect -941 10837 -929 10871
rect -895 10837 -883 10871
rect -941 10831 -883 10837
rect -749 10871 -691 10877
rect -749 10837 -737 10871
rect -703 10837 -691 10871
rect -749 10831 -691 10837
rect -557 10871 -499 10877
rect -557 10837 -545 10871
rect -511 10837 -499 10871
rect -557 10831 -499 10837
rect -365 10871 -307 10877
rect -365 10837 -353 10871
rect -319 10837 -307 10871
rect -365 10831 -307 10837
rect -173 10871 -115 10877
rect -173 10837 -161 10871
rect -127 10837 -115 10871
rect -173 10831 -115 10837
rect 19 10871 77 10877
rect 19 10837 31 10871
rect 65 10837 77 10871
rect 19 10831 77 10837
rect 211 10871 269 10877
rect 211 10837 223 10871
rect 257 10837 269 10871
rect 211 10831 269 10837
rect 403 10871 461 10877
rect 403 10837 415 10871
rect 449 10837 461 10871
rect 403 10831 461 10837
rect 595 10871 653 10877
rect 595 10837 607 10871
rect 641 10837 653 10871
rect 595 10831 653 10837
rect 787 10871 845 10877
rect 787 10837 799 10871
rect 833 10837 845 10871
rect 787 10831 845 10837
rect -983 10778 -937 10790
rect -983 7402 -977 10778
rect -943 7402 -937 10778
rect -983 7390 -937 7402
rect -887 10778 -841 10790
rect -887 7402 -881 10778
rect -847 7402 -841 10778
rect -887 7390 -841 7402
rect -791 10778 -745 10790
rect -791 7402 -785 10778
rect -751 7402 -745 10778
rect -791 7390 -745 7402
rect -695 10778 -649 10790
rect -695 7402 -689 10778
rect -655 7402 -649 10778
rect -695 7390 -649 7402
rect -599 10778 -553 10790
rect -599 7402 -593 10778
rect -559 7402 -553 10778
rect -599 7390 -553 7402
rect -503 10778 -457 10790
rect -503 7402 -497 10778
rect -463 7402 -457 10778
rect -503 7390 -457 7402
rect -407 10778 -361 10790
rect -407 7402 -401 10778
rect -367 7402 -361 10778
rect -407 7390 -361 7402
rect -311 10778 -265 10790
rect -311 7402 -305 10778
rect -271 7402 -265 10778
rect -311 7390 -265 7402
rect -215 10778 -169 10790
rect -215 7402 -209 10778
rect -175 7402 -169 10778
rect -215 7390 -169 7402
rect -119 10778 -73 10790
rect -119 7402 -113 10778
rect -79 7402 -73 10778
rect -119 7390 -73 7402
rect -23 10778 23 10790
rect -23 7402 -17 10778
rect 17 7402 23 10778
rect -23 7390 23 7402
rect 73 10778 119 10790
rect 73 7402 79 10778
rect 113 7402 119 10778
rect 73 7390 119 7402
rect 169 10778 215 10790
rect 169 7402 175 10778
rect 209 7402 215 10778
rect 169 7390 215 7402
rect 265 10778 311 10790
rect 265 7402 271 10778
rect 305 7402 311 10778
rect 265 7390 311 7402
rect 361 10778 407 10790
rect 361 7402 367 10778
rect 401 7402 407 10778
rect 361 7390 407 7402
rect 457 10778 503 10790
rect 457 7402 463 10778
rect 497 7402 503 10778
rect 457 7390 503 7402
rect 553 10778 599 10790
rect 553 7402 559 10778
rect 593 7402 599 10778
rect 553 7390 599 7402
rect 649 10778 695 10790
rect 649 7402 655 10778
rect 689 7402 695 10778
rect 649 7390 695 7402
rect 745 10778 791 10790
rect 745 7402 751 10778
rect 785 7402 791 10778
rect 745 7390 791 7402
rect 841 10778 887 10790
rect 841 7402 847 10778
rect 881 7402 887 10778
rect 841 7390 887 7402
rect 937 10778 983 10790
rect 937 7402 943 10778
rect 977 7402 983 10778
rect 937 7390 983 7402
rect -845 7343 -787 7349
rect -845 7309 -833 7343
rect -799 7309 -787 7343
rect -845 7303 -787 7309
rect -653 7343 -595 7349
rect -653 7309 -641 7343
rect -607 7309 -595 7343
rect -653 7303 -595 7309
rect -461 7343 -403 7349
rect -461 7309 -449 7343
rect -415 7309 -403 7343
rect -461 7303 -403 7309
rect -269 7343 -211 7349
rect -269 7309 -257 7343
rect -223 7309 -211 7343
rect -269 7303 -211 7309
rect -77 7343 -19 7349
rect -77 7309 -65 7343
rect -31 7309 -19 7343
rect -77 7303 -19 7309
rect 115 7343 173 7349
rect 115 7309 127 7343
rect 161 7309 173 7343
rect 115 7303 173 7309
rect 307 7343 365 7349
rect 307 7309 319 7343
rect 353 7309 365 7343
rect 307 7303 365 7309
rect 499 7343 557 7349
rect 499 7309 511 7343
rect 545 7309 557 7343
rect 499 7303 557 7309
rect 691 7343 749 7349
rect 691 7309 703 7343
rect 737 7309 749 7343
rect 691 7303 749 7309
rect 883 7343 941 7349
rect 883 7309 895 7343
rect 929 7309 941 7343
rect 883 7303 941 7309
rect -845 7235 -787 7241
rect -845 7201 -833 7235
rect -799 7201 -787 7235
rect -845 7195 -787 7201
rect -653 7235 -595 7241
rect -653 7201 -641 7235
rect -607 7201 -595 7235
rect -653 7195 -595 7201
rect -461 7235 -403 7241
rect -461 7201 -449 7235
rect -415 7201 -403 7235
rect -461 7195 -403 7201
rect -269 7235 -211 7241
rect -269 7201 -257 7235
rect -223 7201 -211 7235
rect -269 7195 -211 7201
rect -77 7235 -19 7241
rect -77 7201 -65 7235
rect -31 7201 -19 7235
rect -77 7195 -19 7201
rect 115 7235 173 7241
rect 115 7201 127 7235
rect 161 7201 173 7235
rect 115 7195 173 7201
rect 307 7235 365 7241
rect 307 7201 319 7235
rect 353 7201 365 7235
rect 307 7195 365 7201
rect 499 7235 557 7241
rect 499 7201 511 7235
rect 545 7201 557 7235
rect 499 7195 557 7201
rect 691 7235 749 7241
rect 691 7201 703 7235
rect 737 7201 749 7235
rect 691 7195 749 7201
rect 883 7235 941 7241
rect 883 7201 895 7235
rect 929 7201 941 7235
rect 883 7195 941 7201
rect -983 7142 -937 7154
rect -983 3766 -977 7142
rect -943 3766 -937 7142
rect -983 3754 -937 3766
rect -887 7142 -841 7154
rect -887 3766 -881 7142
rect -847 3766 -841 7142
rect -887 3754 -841 3766
rect -791 7142 -745 7154
rect -791 3766 -785 7142
rect -751 3766 -745 7142
rect -791 3754 -745 3766
rect -695 7142 -649 7154
rect -695 3766 -689 7142
rect -655 3766 -649 7142
rect -695 3754 -649 3766
rect -599 7142 -553 7154
rect -599 3766 -593 7142
rect -559 3766 -553 7142
rect -599 3754 -553 3766
rect -503 7142 -457 7154
rect -503 3766 -497 7142
rect -463 3766 -457 7142
rect -503 3754 -457 3766
rect -407 7142 -361 7154
rect -407 3766 -401 7142
rect -367 3766 -361 7142
rect -407 3754 -361 3766
rect -311 7142 -265 7154
rect -311 3766 -305 7142
rect -271 3766 -265 7142
rect -311 3754 -265 3766
rect -215 7142 -169 7154
rect -215 3766 -209 7142
rect -175 3766 -169 7142
rect -215 3754 -169 3766
rect -119 7142 -73 7154
rect -119 3766 -113 7142
rect -79 3766 -73 7142
rect -119 3754 -73 3766
rect -23 7142 23 7154
rect -23 3766 -17 7142
rect 17 3766 23 7142
rect -23 3754 23 3766
rect 73 7142 119 7154
rect 73 3766 79 7142
rect 113 3766 119 7142
rect 73 3754 119 3766
rect 169 7142 215 7154
rect 169 3766 175 7142
rect 209 3766 215 7142
rect 169 3754 215 3766
rect 265 7142 311 7154
rect 265 3766 271 7142
rect 305 3766 311 7142
rect 265 3754 311 3766
rect 361 7142 407 7154
rect 361 3766 367 7142
rect 401 3766 407 7142
rect 361 3754 407 3766
rect 457 7142 503 7154
rect 457 3766 463 7142
rect 497 3766 503 7142
rect 457 3754 503 3766
rect 553 7142 599 7154
rect 553 3766 559 7142
rect 593 3766 599 7142
rect 553 3754 599 3766
rect 649 7142 695 7154
rect 649 3766 655 7142
rect 689 3766 695 7142
rect 649 3754 695 3766
rect 745 7142 791 7154
rect 745 3766 751 7142
rect 785 3766 791 7142
rect 745 3754 791 3766
rect 841 7142 887 7154
rect 841 3766 847 7142
rect 881 3766 887 7142
rect 841 3754 887 3766
rect 937 7142 983 7154
rect 937 3766 943 7142
rect 977 3766 983 7142
rect 937 3754 983 3766
rect -941 3707 -883 3713
rect -941 3673 -929 3707
rect -895 3673 -883 3707
rect -941 3667 -883 3673
rect -749 3707 -691 3713
rect -749 3673 -737 3707
rect -703 3673 -691 3707
rect -749 3667 -691 3673
rect -557 3707 -499 3713
rect -557 3673 -545 3707
rect -511 3673 -499 3707
rect -557 3667 -499 3673
rect -365 3707 -307 3713
rect -365 3673 -353 3707
rect -319 3673 -307 3707
rect -365 3667 -307 3673
rect -173 3707 -115 3713
rect -173 3673 -161 3707
rect -127 3673 -115 3707
rect -173 3667 -115 3673
rect 19 3707 77 3713
rect 19 3673 31 3707
rect 65 3673 77 3707
rect 19 3667 77 3673
rect 211 3707 269 3713
rect 211 3673 223 3707
rect 257 3673 269 3707
rect 211 3667 269 3673
rect 403 3707 461 3713
rect 403 3673 415 3707
rect 449 3673 461 3707
rect 403 3667 461 3673
rect 595 3707 653 3713
rect 595 3673 607 3707
rect 641 3673 653 3707
rect 595 3667 653 3673
rect 787 3707 845 3713
rect 787 3673 799 3707
rect 833 3673 845 3707
rect 787 3667 845 3673
rect -941 3599 -883 3605
rect -941 3565 -929 3599
rect -895 3565 -883 3599
rect -941 3559 -883 3565
rect -749 3599 -691 3605
rect -749 3565 -737 3599
rect -703 3565 -691 3599
rect -749 3559 -691 3565
rect -557 3599 -499 3605
rect -557 3565 -545 3599
rect -511 3565 -499 3599
rect -557 3559 -499 3565
rect -365 3599 -307 3605
rect -365 3565 -353 3599
rect -319 3565 -307 3599
rect -365 3559 -307 3565
rect -173 3599 -115 3605
rect -173 3565 -161 3599
rect -127 3565 -115 3599
rect -173 3559 -115 3565
rect 19 3599 77 3605
rect 19 3565 31 3599
rect 65 3565 77 3599
rect 19 3559 77 3565
rect 211 3599 269 3605
rect 211 3565 223 3599
rect 257 3565 269 3599
rect 211 3559 269 3565
rect 403 3599 461 3605
rect 403 3565 415 3599
rect 449 3565 461 3599
rect 403 3559 461 3565
rect 595 3599 653 3605
rect 595 3565 607 3599
rect 641 3565 653 3599
rect 595 3559 653 3565
rect 787 3599 845 3605
rect 787 3565 799 3599
rect 833 3565 845 3599
rect 787 3559 845 3565
rect -983 3506 -937 3518
rect -983 130 -977 3506
rect -943 130 -937 3506
rect -983 118 -937 130
rect -887 3506 -841 3518
rect -887 130 -881 3506
rect -847 130 -841 3506
rect -887 118 -841 130
rect -791 3506 -745 3518
rect -791 130 -785 3506
rect -751 130 -745 3506
rect -791 118 -745 130
rect -695 3506 -649 3518
rect -695 130 -689 3506
rect -655 130 -649 3506
rect -695 118 -649 130
rect -599 3506 -553 3518
rect -599 130 -593 3506
rect -559 130 -553 3506
rect -599 118 -553 130
rect -503 3506 -457 3518
rect -503 130 -497 3506
rect -463 130 -457 3506
rect -503 118 -457 130
rect -407 3506 -361 3518
rect -407 130 -401 3506
rect -367 130 -361 3506
rect -407 118 -361 130
rect -311 3506 -265 3518
rect -311 130 -305 3506
rect -271 130 -265 3506
rect -311 118 -265 130
rect -215 3506 -169 3518
rect -215 130 -209 3506
rect -175 130 -169 3506
rect -215 118 -169 130
rect -119 3506 -73 3518
rect -119 130 -113 3506
rect -79 130 -73 3506
rect -119 118 -73 130
rect -23 3506 23 3518
rect -23 130 -17 3506
rect 17 130 23 3506
rect -23 118 23 130
rect 73 3506 119 3518
rect 73 130 79 3506
rect 113 130 119 3506
rect 73 118 119 130
rect 169 3506 215 3518
rect 169 130 175 3506
rect 209 130 215 3506
rect 169 118 215 130
rect 265 3506 311 3518
rect 265 130 271 3506
rect 305 130 311 3506
rect 265 118 311 130
rect 361 3506 407 3518
rect 361 130 367 3506
rect 401 130 407 3506
rect 361 118 407 130
rect 457 3506 503 3518
rect 457 130 463 3506
rect 497 130 503 3506
rect 457 118 503 130
rect 553 3506 599 3518
rect 553 130 559 3506
rect 593 130 599 3506
rect 553 118 599 130
rect 649 3506 695 3518
rect 649 130 655 3506
rect 689 130 695 3506
rect 649 118 695 130
rect 745 3506 791 3518
rect 745 130 751 3506
rect 785 130 791 3506
rect 745 118 791 130
rect 841 3506 887 3518
rect 841 130 847 3506
rect 881 130 887 3506
rect 841 118 887 130
rect 937 3506 983 3518
rect 937 130 943 3506
rect 977 130 983 3506
rect 937 118 983 130
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect -983 -130 -937 -118
rect -983 -3506 -977 -130
rect -943 -3506 -937 -130
rect -983 -3518 -937 -3506
rect -887 -130 -841 -118
rect -887 -3506 -881 -130
rect -847 -3506 -841 -130
rect -887 -3518 -841 -3506
rect -791 -130 -745 -118
rect -791 -3506 -785 -130
rect -751 -3506 -745 -130
rect -791 -3518 -745 -3506
rect -695 -130 -649 -118
rect -695 -3506 -689 -130
rect -655 -3506 -649 -130
rect -695 -3518 -649 -3506
rect -599 -130 -553 -118
rect -599 -3506 -593 -130
rect -559 -3506 -553 -130
rect -599 -3518 -553 -3506
rect -503 -130 -457 -118
rect -503 -3506 -497 -130
rect -463 -3506 -457 -130
rect -503 -3518 -457 -3506
rect -407 -130 -361 -118
rect -407 -3506 -401 -130
rect -367 -3506 -361 -130
rect -407 -3518 -361 -3506
rect -311 -130 -265 -118
rect -311 -3506 -305 -130
rect -271 -3506 -265 -130
rect -311 -3518 -265 -3506
rect -215 -130 -169 -118
rect -215 -3506 -209 -130
rect -175 -3506 -169 -130
rect -215 -3518 -169 -3506
rect -119 -130 -73 -118
rect -119 -3506 -113 -130
rect -79 -3506 -73 -130
rect -119 -3518 -73 -3506
rect -23 -130 23 -118
rect -23 -3506 -17 -130
rect 17 -3506 23 -130
rect -23 -3518 23 -3506
rect 73 -130 119 -118
rect 73 -3506 79 -130
rect 113 -3506 119 -130
rect 73 -3518 119 -3506
rect 169 -130 215 -118
rect 169 -3506 175 -130
rect 209 -3506 215 -130
rect 169 -3518 215 -3506
rect 265 -130 311 -118
rect 265 -3506 271 -130
rect 305 -3506 311 -130
rect 265 -3518 311 -3506
rect 361 -130 407 -118
rect 361 -3506 367 -130
rect 401 -3506 407 -130
rect 361 -3518 407 -3506
rect 457 -130 503 -118
rect 457 -3506 463 -130
rect 497 -3506 503 -130
rect 457 -3518 503 -3506
rect 553 -130 599 -118
rect 553 -3506 559 -130
rect 593 -3506 599 -130
rect 553 -3518 599 -3506
rect 649 -130 695 -118
rect 649 -3506 655 -130
rect 689 -3506 695 -130
rect 649 -3518 695 -3506
rect 745 -130 791 -118
rect 745 -3506 751 -130
rect 785 -3506 791 -130
rect 745 -3518 791 -3506
rect 841 -130 887 -118
rect 841 -3506 847 -130
rect 881 -3506 887 -130
rect 841 -3518 887 -3506
rect 937 -130 983 -118
rect 937 -3506 943 -130
rect 977 -3506 983 -130
rect 937 -3518 983 -3506
rect -941 -3565 -883 -3559
rect -941 -3599 -929 -3565
rect -895 -3599 -883 -3565
rect -941 -3605 -883 -3599
rect -749 -3565 -691 -3559
rect -749 -3599 -737 -3565
rect -703 -3599 -691 -3565
rect -749 -3605 -691 -3599
rect -557 -3565 -499 -3559
rect -557 -3599 -545 -3565
rect -511 -3599 -499 -3565
rect -557 -3605 -499 -3599
rect -365 -3565 -307 -3559
rect -365 -3599 -353 -3565
rect -319 -3599 -307 -3565
rect -365 -3605 -307 -3599
rect -173 -3565 -115 -3559
rect -173 -3599 -161 -3565
rect -127 -3599 -115 -3565
rect -173 -3605 -115 -3599
rect 19 -3565 77 -3559
rect 19 -3599 31 -3565
rect 65 -3599 77 -3565
rect 19 -3605 77 -3599
rect 211 -3565 269 -3559
rect 211 -3599 223 -3565
rect 257 -3599 269 -3565
rect 211 -3605 269 -3599
rect 403 -3565 461 -3559
rect 403 -3599 415 -3565
rect 449 -3599 461 -3565
rect 403 -3605 461 -3599
rect 595 -3565 653 -3559
rect 595 -3599 607 -3565
rect 641 -3599 653 -3565
rect 595 -3605 653 -3599
rect 787 -3565 845 -3559
rect 787 -3599 799 -3565
rect 833 -3599 845 -3565
rect 787 -3605 845 -3599
rect -941 -3673 -883 -3667
rect -941 -3707 -929 -3673
rect -895 -3707 -883 -3673
rect -941 -3713 -883 -3707
rect -749 -3673 -691 -3667
rect -749 -3707 -737 -3673
rect -703 -3707 -691 -3673
rect -749 -3713 -691 -3707
rect -557 -3673 -499 -3667
rect -557 -3707 -545 -3673
rect -511 -3707 -499 -3673
rect -557 -3713 -499 -3707
rect -365 -3673 -307 -3667
rect -365 -3707 -353 -3673
rect -319 -3707 -307 -3673
rect -365 -3713 -307 -3707
rect -173 -3673 -115 -3667
rect -173 -3707 -161 -3673
rect -127 -3707 -115 -3673
rect -173 -3713 -115 -3707
rect 19 -3673 77 -3667
rect 19 -3707 31 -3673
rect 65 -3707 77 -3673
rect 19 -3713 77 -3707
rect 211 -3673 269 -3667
rect 211 -3707 223 -3673
rect 257 -3707 269 -3673
rect 211 -3713 269 -3707
rect 403 -3673 461 -3667
rect 403 -3707 415 -3673
rect 449 -3707 461 -3673
rect 403 -3713 461 -3707
rect 595 -3673 653 -3667
rect 595 -3707 607 -3673
rect 641 -3707 653 -3673
rect 595 -3713 653 -3707
rect 787 -3673 845 -3667
rect 787 -3707 799 -3673
rect 833 -3707 845 -3673
rect 787 -3713 845 -3707
rect -983 -3766 -937 -3754
rect -983 -7142 -977 -3766
rect -943 -7142 -937 -3766
rect -983 -7154 -937 -7142
rect -887 -3766 -841 -3754
rect -887 -7142 -881 -3766
rect -847 -7142 -841 -3766
rect -887 -7154 -841 -7142
rect -791 -3766 -745 -3754
rect -791 -7142 -785 -3766
rect -751 -7142 -745 -3766
rect -791 -7154 -745 -7142
rect -695 -3766 -649 -3754
rect -695 -7142 -689 -3766
rect -655 -7142 -649 -3766
rect -695 -7154 -649 -7142
rect -599 -3766 -553 -3754
rect -599 -7142 -593 -3766
rect -559 -7142 -553 -3766
rect -599 -7154 -553 -7142
rect -503 -3766 -457 -3754
rect -503 -7142 -497 -3766
rect -463 -7142 -457 -3766
rect -503 -7154 -457 -7142
rect -407 -3766 -361 -3754
rect -407 -7142 -401 -3766
rect -367 -7142 -361 -3766
rect -407 -7154 -361 -7142
rect -311 -3766 -265 -3754
rect -311 -7142 -305 -3766
rect -271 -7142 -265 -3766
rect -311 -7154 -265 -7142
rect -215 -3766 -169 -3754
rect -215 -7142 -209 -3766
rect -175 -7142 -169 -3766
rect -215 -7154 -169 -7142
rect -119 -3766 -73 -3754
rect -119 -7142 -113 -3766
rect -79 -7142 -73 -3766
rect -119 -7154 -73 -7142
rect -23 -3766 23 -3754
rect -23 -7142 -17 -3766
rect 17 -7142 23 -3766
rect -23 -7154 23 -7142
rect 73 -3766 119 -3754
rect 73 -7142 79 -3766
rect 113 -7142 119 -3766
rect 73 -7154 119 -7142
rect 169 -3766 215 -3754
rect 169 -7142 175 -3766
rect 209 -7142 215 -3766
rect 169 -7154 215 -7142
rect 265 -3766 311 -3754
rect 265 -7142 271 -3766
rect 305 -7142 311 -3766
rect 265 -7154 311 -7142
rect 361 -3766 407 -3754
rect 361 -7142 367 -3766
rect 401 -7142 407 -3766
rect 361 -7154 407 -7142
rect 457 -3766 503 -3754
rect 457 -7142 463 -3766
rect 497 -7142 503 -3766
rect 457 -7154 503 -7142
rect 553 -3766 599 -3754
rect 553 -7142 559 -3766
rect 593 -7142 599 -3766
rect 553 -7154 599 -7142
rect 649 -3766 695 -3754
rect 649 -7142 655 -3766
rect 689 -7142 695 -3766
rect 649 -7154 695 -7142
rect 745 -3766 791 -3754
rect 745 -7142 751 -3766
rect 785 -7142 791 -3766
rect 745 -7154 791 -7142
rect 841 -3766 887 -3754
rect 841 -7142 847 -3766
rect 881 -7142 887 -3766
rect 841 -7154 887 -7142
rect 937 -3766 983 -3754
rect 937 -7142 943 -3766
rect 977 -7142 983 -3766
rect 937 -7154 983 -7142
rect -845 -7201 -787 -7195
rect -845 -7235 -833 -7201
rect -799 -7235 -787 -7201
rect -845 -7241 -787 -7235
rect -653 -7201 -595 -7195
rect -653 -7235 -641 -7201
rect -607 -7235 -595 -7201
rect -653 -7241 -595 -7235
rect -461 -7201 -403 -7195
rect -461 -7235 -449 -7201
rect -415 -7235 -403 -7201
rect -461 -7241 -403 -7235
rect -269 -7201 -211 -7195
rect -269 -7235 -257 -7201
rect -223 -7235 -211 -7201
rect -269 -7241 -211 -7235
rect -77 -7201 -19 -7195
rect -77 -7235 -65 -7201
rect -31 -7235 -19 -7201
rect -77 -7241 -19 -7235
rect 115 -7201 173 -7195
rect 115 -7235 127 -7201
rect 161 -7235 173 -7201
rect 115 -7241 173 -7235
rect 307 -7201 365 -7195
rect 307 -7235 319 -7201
rect 353 -7235 365 -7201
rect 307 -7241 365 -7235
rect 499 -7201 557 -7195
rect 499 -7235 511 -7201
rect 545 -7235 557 -7201
rect 499 -7241 557 -7235
rect 691 -7201 749 -7195
rect 691 -7235 703 -7201
rect 737 -7235 749 -7201
rect 691 -7241 749 -7235
rect 883 -7201 941 -7195
rect 883 -7235 895 -7201
rect 929 -7235 941 -7201
rect 883 -7241 941 -7235
rect -845 -7309 -787 -7303
rect -845 -7343 -833 -7309
rect -799 -7343 -787 -7309
rect -845 -7349 -787 -7343
rect -653 -7309 -595 -7303
rect -653 -7343 -641 -7309
rect -607 -7343 -595 -7309
rect -653 -7349 -595 -7343
rect -461 -7309 -403 -7303
rect -461 -7343 -449 -7309
rect -415 -7343 -403 -7309
rect -461 -7349 -403 -7343
rect -269 -7309 -211 -7303
rect -269 -7343 -257 -7309
rect -223 -7343 -211 -7309
rect -269 -7349 -211 -7343
rect -77 -7309 -19 -7303
rect -77 -7343 -65 -7309
rect -31 -7343 -19 -7309
rect -77 -7349 -19 -7343
rect 115 -7309 173 -7303
rect 115 -7343 127 -7309
rect 161 -7343 173 -7309
rect 115 -7349 173 -7343
rect 307 -7309 365 -7303
rect 307 -7343 319 -7309
rect 353 -7343 365 -7309
rect 307 -7349 365 -7343
rect 499 -7309 557 -7303
rect 499 -7343 511 -7309
rect 545 -7343 557 -7309
rect 499 -7349 557 -7343
rect 691 -7309 749 -7303
rect 691 -7343 703 -7309
rect 737 -7343 749 -7309
rect 691 -7349 749 -7343
rect 883 -7309 941 -7303
rect 883 -7343 895 -7309
rect 929 -7343 941 -7309
rect 883 -7349 941 -7343
rect -983 -7402 -937 -7390
rect -983 -10778 -977 -7402
rect -943 -10778 -937 -7402
rect -983 -10790 -937 -10778
rect -887 -7402 -841 -7390
rect -887 -10778 -881 -7402
rect -847 -10778 -841 -7402
rect -887 -10790 -841 -10778
rect -791 -7402 -745 -7390
rect -791 -10778 -785 -7402
rect -751 -10778 -745 -7402
rect -791 -10790 -745 -10778
rect -695 -7402 -649 -7390
rect -695 -10778 -689 -7402
rect -655 -10778 -649 -7402
rect -695 -10790 -649 -10778
rect -599 -7402 -553 -7390
rect -599 -10778 -593 -7402
rect -559 -10778 -553 -7402
rect -599 -10790 -553 -10778
rect -503 -7402 -457 -7390
rect -503 -10778 -497 -7402
rect -463 -10778 -457 -7402
rect -503 -10790 -457 -10778
rect -407 -7402 -361 -7390
rect -407 -10778 -401 -7402
rect -367 -10778 -361 -7402
rect -407 -10790 -361 -10778
rect -311 -7402 -265 -7390
rect -311 -10778 -305 -7402
rect -271 -10778 -265 -7402
rect -311 -10790 -265 -10778
rect -215 -7402 -169 -7390
rect -215 -10778 -209 -7402
rect -175 -10778 -169 -7402
rect -215 -10790 -169 -10778
rect -119 -7402 -73 -7390
rect -119 -10778 -113 -7402
rect -79 -10778 -73 -7402
rect -119 -10790 -73 -10778
rect -23 -7402 23 -7390
rect -23 -10778 -17 -7402
rect 17 -10778 23 -7402
rect -23 -10790 23 -10778
rect 73 -7402 119 -7390
rect 73 -10778 79 -7402
rect 113 -10778 119 -7402
rect 73 -10790 119 -10778
rect 169 -7402 215 -7390
rect 169 -10778 175 -7402
rect 209 -10778 215 -7402
rect 169 -10790 215 -10778
rect 265 -7402 311 -7390
rect 265 -10778 271 -7402
rect 305 -10778 311 -7402
rect 265 -10790 311 -10778
rect 361 -7402 407 -7390
rect 361 -10778 367 -7402
rect 401 -10778 407 -7402
rect 361 -10790 407 -10778
rect 457 -7402 503 -7390
rect 457 -10778 463 -7402
rect 497 -10778 503 -7402
rect 457 -10790 503 -10778
rect 553 -7402 599 -7390
rect 553 -10778 559 -7402
rect 593 -10778 599 -7402
rect 553 -10790 599 -10778
rect 649 -7402 695 -7390
rect 649 -10778 655 -7402
rect 689 -10778 695 -7402
rect 649 -10790 695 -10778
rect 745 -7402 791 -7390
rect 745 -10778 751 -7402
rect 785 -10778 791 -7402
rect 745 -10790 791 -10778
rect 841 -7402 887 -7390
rect 841 -10778 847 -7402
rect 881 -10778 887 -7402
rect 841 -10790 887 -10778
rect 937 -7402 983 -7390
rect 937 -10778 943 -7402
rect 977 -10778 983 -7402
rect 937 -10790 983 -10778
rect -941 -10837 -883 -10831
rect -941 -10871 -929 -10837
rect -895 -10871 -883 -10837
rect -941 -10877 -883 -10871
rect -749 -10837 -691 -10831
rect -749 -10871 -737 -10837
rect -703 -10871 -691 -10837
rect -749 -10877 -691 -10871
rect -557 -10837 -499 -10831
rect -557 -10871 -545 -10837
rect -511 -10871 -499 -10837
rect -557 -10877 -499 -10871
rect -365 -10837 -307 -10831
rect -365 -10871 -353 -10837
rect -319 -10871 -307 -10837
rect -365 -10877 -307 -10871
rect -173 -10837 -115 -10831
rect -173 -10871 -161 -10837
rect -127 -10871 -115 -10837
rect -173 -10877 -115 -10871
rect 19 -10837 77 -10831
rect 19 -10871 31 -10837
rect 65 -10871 77 -10837
rect 19 -10877 77 -10871
rect 211 -10837 269 -10831
rect 211 -10871 223 -10837
rect 257 -10871 269 -10837
rect 211 -10877 269 -10871
rect 403 -10837 461 -10831
rect 403 -10871 415 -10837
rect 449 -10871 461 -10837
rect 403 -10877 461 -10871
rect 595 -10837 653 -10831
rect 595 -10871 607 -10837
rect 641 -10871 653 -10837
rect 595 -10877 653 -10871
rect 787 -10837 845 -10831
rect 787 -10871 799 -10837
rect 833 -10871 845 -10837
rect 787 -10877 845 -10871
rect -941 -10945 -883 -10939
rect -941 -10979 -929 -10945
rect -895 -10979 -883 -10945
rect -941 -10985 -883 -10979
rect -749 -10945 -691 -10939
rect -749 -10979 -737 -10945
rect -703 -10979 -691 -10945
rect -749 -10985 -691 -10979
rect -557 -10945 -499 -10939
rect -557 -10979 -545 -10945
rect -511 -10979 -499 -10945
rect -557 -10985 -499 -10979
rect -365 -10945 -307 -10939
rect -365 -10979 -353 -10945
rect -319 -10979 -307 -10945
rect -365 -10985 -307 -10979
rect -173 -10945 -115 -10939
rect -173 -10979 -161 -10945
rect -127 -10979 -115 -10945
rect -173 -10985 -115 -10979
rect 19 -10945 77 -10939
rect 19 -10979 31 -10945
rect 65 -10979 77 -10945
rect 19 -10985 77 -10979
rect 211 -10945 269 -10939
rect 211 -10979 223 -10945
rect 257 -10979 269 -10945
rect 211 -10985 269 -10979
rect 403 -10945 461 -10939
rect 403 -10979 415 -10945
rect 449 -10979 461 -10945
rect 403 -10985 461 -10979
rect 595 -10945 653 -10939
rect 595 -10979 607 -10945
rect 641 -10979 653 -10945
rect 595 -10985 653 -10979
rect 787 -10945 845 -10939
rect 787 -10979 799 -10945
rect 833 -10979 845 -10945
rect 787 -10985 845 -10979
rect -983 -11038 -937 -11026
rect -983 -14414 -977 -11038
rect -943 -14414 -937 -11038
rect -983 -14426 -937 -14414
rect -887 -11038 -841 -11026
rect -887 -14414 -881 -11038
rect -847 -14414 -841 -11038
rect -887 -14426 -841 -14414
rect -791 -11038 -745 -11026
rect -791 -14414 -785 -11038
rect -751 -14414 -745 -11038
rect -791 -14426 -745 -14414
rect -695 -11038 -649 -11026
rect -695 -14414 -689 -11038
rect -655 -14414 -649 -11038
rect -695 -14426 -649 -14414
rect -599 -11038 -553 -11026
rect -599 -14414 -593 -11038
rect -559 -14414 -553 -11038
rect -599 -14426 -553 -14414
rect -503 -11038 -457 -11026
rect -503 -14414 -497 -11038
rect -463 -14414 -457 -11038
rect -503 -14426 -457 -14414
rect -407 -11038 -361 -11026
rect -407 -14414 -401 -11038
rect -367 -14414 -361 -11038
rect -407 -14426 -361 -14414
rect -311 -11038 -265 -11026
rect -311 -14414 -305 -11038
rect -271 -14414 -265 -11038
rect -311 -14426 -265 -14414
rect -215 -11038 -169 -11026
rect -215 -14414 -209 -11038
rect -175 -14414 -169 -11038
rect -215 -14426 -169 -14414
rect -119 -11038 -73 -11026
rect -119 -14414 -113 -11038
rect -79 -14414 -73 -11038
rect -119 -14426 -73 -14414
rect -23 -11038 23 -11026
rect -23 -14414 -17 -11038
rect 17 -14414 23 -11038
rect -23 -14426 23 -14414
rect 73 -11038 119 -11026
rect 73 -14414 79 -11038
rect 113 -14414 119 -11038
rect 73 -14426 119 -14414
rect 169 -11038 215 -11026
rect 169 -14414 175 -11038
rect 209 -14414 215 -11038
rect 169 -14426 215 -14414
rect 265 -11038 311 -11026
rect 265 -14414 271 -11038
rect 305 -14414 311 -11038
rect 265 -14426 311 -14414
rect 361 -11038 407 -11026
rect 361 -14414 367 -11038
rect 401 -14414 407 -11038
rect 361 -14426 407 -14414
rect 457 -11038 503 -11026
rect 457 -14414 463 -11038
rect 497 -14414 503 -11038
rect 457 -14426 503 -14414
rect 553 -11038 599 -11026
rect 553 -14414 559 -11038
rect 593 -14414 599 -11038
rect 553 -14426 599 -14414
rect 649 -11038 695 -11026
rect 649 -14414 655 -11038
rect 689 -14414 695 -11038
rect 649 -14426 695 -14414
rect 745 -11038 791 -11026
rect 745 -14414 751 -11038
rect 785 -14414 791 -11038
rect 745 -14426 791 -14414
rect 841 -11038 887 -11026
rect 841 -14414 847 -11038
rect 881 -14414 887 -11038
rect 841 -14426 887 -14414
rect 937 -11038 983 -11026
rect 937 -14414 943 -11038
rect 977 -14414 983 -11038
rect 937 -14426 983 -14414
rect -845 -14473 -787 -14467
rect -845 -14507 -833 -14473
rect -799 -14507 -787 -14473
rect -845 -14513 -787 -14507
rect -653 -14473 -595 -14467
rect -653 -14507 -641 -14473
rect -607 -14507 -595 -14473
rect -653 -14513 -595 -14507
rect -461 -14473 -403 -14467
rect -461 -14507 -449 -14473
rect -415 -14507 -403 -14473
rect -461 -14513 -403 -14507
rect -269 -14473 -211 -14467
rect -269 -14507 -257 -14473
rect -223 -14507 -211 -14473
rect -269 -14513 -211 -14507
rect -77 -14473 -19 -14467
rect -77 -14507 -65 -14473
rect -31 -14507 -19 -14473
rect -77 -14513 -19 -14507
rect 115 -14473 173 -14467
rect 115 -14507 127 -14473
rect 161 -14507 173 -14473
rect 115 -14513 173 -14507
rect 307 -14473 365 -14467
rect 307 -14507 319 -14473
rect 353 -14507 365 -14473
rect 307 -14513 365 -14507
rect 499 -14473 557 -14467
rect 499 -14507 511 -14473
rect 545 -14507 557 -14473
rect 499 -14513 557 -14507
rect 691 -14473 749 -14467
rect 691 -14507 703 -14473
rect 737 -14507 749 -14473
rect 691 -14513 749 -14507
rect 883 -14473 941 -14467
rect 883 -14507 895 -14473
rect 929 -14507 941 -14473
rect 883 -14513 941 -14507
rect -845 -14581 -787 -14575
rect -845 -14615 -833 -14581
rect -799 -14615 -787 -14581
rect -845 -14621 -787 -14615
rect -653 -14581 -595 -14575
rect -653 -14615 -641 -14581
rect -607 -14615 -595 -14581
rect -653 -14621 -595 -14615
rect -461 -14581 -403 -14575
rect -461 -14615 -449 -14581
rect -415 -14615 -403 -14581
rect -461 -14621 -403 -14615
rect -269 -14581 -211 -14575
rect -269 -14615 -257 -14581
rect -223 -14615 -211 -14581
rect -269 -14621 -211 -14615
rect -77 -14581 -19 -14575
rect -77 -14615 -65 -14581
rect -31 -14615 -19 -14581
rect -77 -14621 -19 -14615
rect 115 -14581 173 -14575
rect 115 -14615 127 -14581
rect 161 -14615 173 -14581
rect 115 -14621 173 -14615
rect 307 -14581 365 -14575
rect 307 -14615 319 -14581
rect 353 -14615 365 -14581
rect 307 -14621 365 -14615
rect 499 -14581 557 -14575
rect 499 -14615 511 -14581
rect 545 -14615 557 -14581
rect 499 -14621 557 -14615
rect 691 -14581 749 -14575
rect 691 -14615 703 -14581
rect 737 -14615 749 -14581
rect 691 -14621 749 -14615
rect 883 -14581 941 -14575
rect 883 -14615 895 -14581
rect 929 -14615 941 -14581
rect 883 -14621 941 -14615
rect -983 -14674 -937 -14662
rect -983 -18050 -977 -14674
rect -943 -18050 -937 -14674
rect -983 -18062 -937 -18050
rect -887 -14674 -841 -14662
rect -887 -18050 -881 -14674
rect -847 -18050 -841 -14674
rect -887 -18062 -841 -18050
rect -791 -14674 -745 -14662
rect -791 -18050 -785 -14674
rect -751 -18050 -745 -14674
rect -791 -18062 -745 -18050
rect -695 -14674 -649 -14662
rect -695 -18050 -689 -14674
rect -655 -18050 -649 -14674
rect -695 -18062 -649 -18050
rect -599 -14674 -553 -14662
rect -599 -18050 -593 -14674
rect -559 -18050 -553 -14674
rect -599 -18062 -553 -18050
rect -503 -14674 -457 -14662
rect -503 -18050 -497 -14674
rect -463 -18050 -457 -14674
rect -503 -18062 -457 -18050
rect -407 -14674 -361 -14662
rect -407 -18050 -401 -14674
rect -367 -18050 -361 -14674
rect -407 -18062 -361 -18050
rect -311 -14674 -265 -14662
rect -311 -18050 -305 -14674
rect -271 -18050 -265 -14674
rect -311 -18062 -265 -18050
rect -215 -14674 -169 -14662
rect -215 -18050 -209 -14674
rect -175 -18050 -169 -14674
rect -215 -18062 -169 -18050
rect -119 -14674 -73 -14662
rect -119 -18050 -113 -14674
rect -79 -18050 -73 -14674
rect -119 -18062 -73 -18050
rect -23 -14674 23 -14662
rect -23 -18050 -17 -14674
rect 17 -18050 23 -14674
rect -23 -18062 23 -18050
rect 73 -14674 119 -14662
rect 73 -18050 79 -14674
rect 113 -18050 119 -14674
rect 73 -18062 119 -18050
rect 169 -14674 215 -14662
rect 169 -18050 175 -14674
rect 209 -18050 215 -14674
rect 169 -18062 215 -18050
rect 265 -14674 311 -14662
rect 265 -18050 271 -14674
rect 305 -18050 311 -14674
rect 265 -18062 311 -18050
rect 361 -14674 407 -14662
rect 361 -18050 367 -14674
rect 401 -18050 407 -14674
rect 361 -18062 407 -18050
rect 457 -14674 503 -14662
rect 457 -18050 463 -14674
rect 497 -18050 503 -14674
rect 457 -18062 503 -18050
rect 553 -14674 599 -14662
rect 553 -18050 559 -14674
rect 593 -18050 599 -14674
rect 553 -18062 599 -18050
rect 649 -14674 695 -14662
rect 649 -18050 655 -14674
rect 689 -18050 695 -14674
rect 649 -18062 695 -18050
rect 745 -14674 791 -14662
rect 745 -18050 751 -14674
rect 785 -18050 791 -14674
rect 745 -18062 791 -18050
rect 841 -14674 887 -14662
rect 841 -18050 847 -14674
rect 881 -18050 887 -14674
rect 841 -18062 887 -18050
rect 937 -14674 983 -14662
rect 937 -18050 943 -14674
rect 977 -18050 983 -14674
rect 937 -18062 983 -18050
rect -941 -18109 -883 -18103
rect -941 -18143 -929 -18109
rect -895 -18143 -883 -18109
rect -941 -18149 -883 -18143
rect -749 -18109 -691 -18103
rect -749 -18143 -737 -18109
rect -703 -18143 -691 -18109
rect -749 -18149 -691 -18143
rect -557 -18109 -499 -18103
rect -557 -18143 -545 -18109
rect -511 -18143 -499 -18109
rect -557 -18149 -499 -18143
rect -365 -18109 -307 -18103
rect -365 -18143 -353 -18109
rect -319 -18143 -307 -18109
rect -365 -18149 -307 -18143
rect -173 -18109 -115 -18103
rect -173 -18143 -161 -18109
rect -127 -18143 -115 -18109
rect -173 -18149 -115 -18143
rect 19 -18109 77 -18103
rect 19 -18143 31 -18109
rect 65 -18143 77 -18109
rect 19 -18149 77 -18143
rect 211 -18109 269 -18103
rect 211 -18143 223 -18109
rect 257 -18143 269 -18109
rect 211 -18149 269 -18143
rect 403 -18109 461 -18103
rect 403 -18143 415 -18109
rect 449 -18143 461 -18109
rect 403 -18149 461 -18143
rect 595 -18109 653 -18103
rect 595 -18143 607 -18109
rect 641 -18143 653 -18109
rect 595 -18149 653 -18143
rect 787 -18109 845 -18103
rect 787 -18143 799 -18109
rect 833 -18143 845 -18109
rect 787 -18149 845 -18143
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 17 l 0.15 m 10 nf 20 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
