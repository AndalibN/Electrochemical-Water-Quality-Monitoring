magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_s >>
rect 2390 3987 2478 4125
rect 4185 4009 4273 4147
rect 2094 2360 2182 2498
rect 3889 2382 3977 2520
<< pwell >>
rect 1181 334 1408 733
rect 2949 333 3179 1009
<< psubdiff >>
rect 2975 929 3153 983
rect 1207 661 1382 707
rect 1207 627 1278 661
rect 1312 627 1382 661
rect 1207 593 1382 627
rect 1207 559 1278 593
rect 1312 559 1382 593
rect 1207 525 1382 559
rect 1207 491 1278 525
rect 1312 491 1382 525
rect 1207 457 1382 491
rect 1207 423 1278 457
rect 1312 423 1382 457
rect 1207 360 1382 423
rect 2975 419 3010 929
rect 3112 419 3153 929
rect 2975 359 3153 419
<< psubdiffcont >>
rect 1278 627 1312 661
rect 1278 559 1312 593
rect 1278 491 1312 525
rect 1278 423 1312 457
rect 3010 419 3112 929
<< poly >>
rect 726 3926 766 3954
<< locali >>
rect 2989 929 3134 967
rect 1237 661 1356 688
rect 1237 627 1278 661
rect 1312 627 1356 661
rect 1237 593 1356 627
rect 1237 559 1278 593
rect 1312 559 1356 593
rect 1237 525 1356 559
rect 1237 491 1278 525
rect 1312 491 1356 525
rect 1237 457 1356 491
rect 1237 423 1278 457
rect 1312 423 1356 457
rect 1237 383 1356 423
rect 2989 419 3010 929
rect 3112 419 3134 929
rect 2989 378 3134 419
<< metal1 >>
rect 710 4039 964 4048
rect 710 3987 741 4039
rect 793 3987 889 4039
rect 941 3987 964 4039
rect 710 3977 964 3987
rect 675 3909 1009 3940
rect 675 3854 710 3909
rect 971 3872 1009 3909
rect 1222 3874 1319 4325
rect 2999 4255 3099 4324
rect 1894 4090 1977 4094
rect 1894 4078 1910 4090
rect 1698 4042 1910 4078
rect 1698 3914 1732 4042
rect 1894 4038 1910 4042
rect 1962 4038 1977 4090
rect 1894 4036 1977 4038
rect 2044 4090 2127 4095
rect 2044 4038 2059 4090
rect 2111 4038 2127 4090
rect 2492 4086 2575 4090
rect 2492 4076 2505 4086
rect 2044 4037 2127 4038
rect 2290 4042 2505 4076
rect 1846 3953 2177 3987
rect 1846 3914 1880 3953
rect 2142 3914 2177 3953
rect 2290 3914 2324 4042
rect 2492 4034 2505 4042
rect 2557 4034 2575 4086
rect 2492 4032 2575 4034
rect 2634 4086 2717 4090
rect 2634 4034 2651 4086
rect 2703 4034 2717 4086
rect 2634 4032 2717 4034
rect 2438 3953 2768 3987
rect 2438 3921 2472 3953
rect 1216 3872 1319 3874
rect 676 3294 710 3854
rect 822 3827 858 3870
rect 822 3304 859 3827
rect 373 2553 710 3294
rect 823 3261 859 3304
rect 971 3675 1319 3872
rect 373 2230 469 2553
rect 823 2364 858 3261
rect 971 2552 1318 3675
rect 972 2527 1318 2552
rect 1216 2428 1318 2527
rect 1549 2527 1584 3913
rect 1697 2572 1732 3914
rect 1845 2582 1880 3914
rect 1845 2572 1881 2582
rect 1846 2527 1881 2572
rect 1549 2492 1881 2527
rect 1600 2453 1683 2456
rect 1600 2401 1615 2453
rect 1667 2401 1683 2453
rect 1600 2398 1683 2401
rect 1747 2452 1830 2456
rect 1747 2400 1762 2452
rect 1814 2400 1830 2452
rect 1747 2398 1830 2400
rect 1612 2364 1670 2398
rect 823 2331 1671 2364
rect 1993 2230 2028 3914
rect 2141 2621 2177 3914
rect 2141 2595 2176 2621
rect 2141 2572 2177 2595
rect 2289 2572 2324 3914
rect 2142 2524 2177 2572
rect 2437 2524 2472 3921
rect 2734 3914 2768 3953
rect 2142 2489 2472 2524
rect 2194 2451 2277 2455
rect 2194 2399 2207 2451
rect 2259 2399 2277 2451
rect 2194 2397 2277 2399
rect 2338 2452 2421 2456
rect 2338 2400 2354 2452
rect 2406 2400 2421 2452
rect 2338 2398 2421 2400
rect 2585 2230 2620 3914
rect 2733 2572 2768 3914
rect 2998 3710 3099 4255
rect 3697 4102 3771 4106
rect 3837 4103 3920 4106
rect 3697 4099 3781 4102
rect 3697 4098 3709 4099
rect 3492 4064 3709 4098
rect 2999 2230 3099 2654
rect 3344 2640 3379 3935
rect 3492 2641 3527 4064
rect 3697 4047 3709 4064
rect 3761 4047 3781 4099
rect 3837 4051 3854 4103
rect 3906 4051 3920 4103
rect 4284 4103 4367 4106
rect 4284 4098 4297 4103
rect 3837 4048 3920 4051
rect 4084 4064 4297 4098
rect 3697 4044 3781 4047
rect 3697 4040 3771 4044
rect 3640 3979 3971 4009
rect 3344 2594 3380 2640
rect 3492 2594 3528 2641
rect 3640 2625 3675 3979
rect 3937 3942 3971 3979
rect 3344 2537 3379 2594
rect 3640 2579 3676 2625
rect 3640 2537 3675 2579
rect 3344 2503 3675 2537
rect 3395 2470 3478 2474
rect 3395 2418 3409 2470
rect 3461 2418 3478 2470
rect 3395 2416 3478 2418
rect 3544 2471 3627 2474
rect 3544 2419 3557 2471
rect 3609 2419 3627 2471
rect 3544 2416 3627 2419
rect 3788 2240 3823 3941
rect 3936 2548 3971 3942
rect 4084 2594 4119 4064
rect 4284 4051 4297 4064
rect 4349 4051 4367 4103
rect 4284 4048 4367 4051
rect 4428 4103 4511 4106
rect 4428 4051 4445 4103
rect 4497 4051 4511 4103
rect 4428 4048 4511 4051
rect 4233 3979 4563 4009
rect 4233 3936 4268 3979
rect 4232 3930 4268 3936
rect 4379 3936 4413 3950
rect 4232 2548 4267 3930
rect 4379 3327 4415 3936
rect 4380 2629 4415 3327
rect 4379 2594 4415 2629
rect 3936 2514 4267 2548
rect 3985 2472 4068 2475
rect 3985 2420 4000 2472
rect 4052 2420 4068 2472
rect 3985 2417 4068 2420
rect 4132 2472 4215 2475
rect 4132 2420 4149 2472
rect 4201 2420 4215 2472
rect 4132 2417 4215 2420
rect 3787 2230 3823 2240
rect 4380 2230 4415 2594
rect 4528 3935 4563 3979
rect 4528 2593 4562 3935
rect 373 2104 4887 2230
rect 1893 1933 3634 1951
rect 1893 1881 1908 1933
rect 1960 1932 3634 1933
rect 1960 1881 3546 1932
rect 1893 1880 3546 1881
rect 3598 1880 3634 1932
rect 1893 1869 3634 1880
rect 1893 1817 1908 1869
rect 1960 1868 3634 1869
rect 1960 1817 3546 1868
rect 1893 1816 3546 1817
rect 3598 1816 3634 1868
rect 1893 1799 3634 1816
rect 708 1655 2430 1692
rect 708 1654 2343 1655
rect 708 1538 746 1654
rect 926 1603 2343 1654
rect 2395 1603 2430 1655
rect 926 1591 2430 1603
rect 926 1539 2343 1591
rect 2395 1539 2430 1591
rect 926 1538 2430 1539
rect 708 1503 2430 1538
rect 953 1502 2430 1503
rect 2490 1425 4229 1442
rect 2490 1373 2506 1425
rect 2558 1424 4229 1425
rect 2558 1373 4143 1424
rect 2490 1372 4143 1373
rect 4195 1372 4229 1424
rect 2490 1361 4229 1372
rect 2490 1309 2506 1361
rect 2558 1360 4229 1361
rect 2558 1309 4143 1360
rect 2490 1308 4143 1309
rect 4195 1308 4229 1360
rect 2490 1291 4229 1308
rect 800 877 883 880
rect 1895 879 1978 882
rect 800 825 815 877
rect 867 825 883 877
rect 1749 875 1832 879
rect 1749 868 1762 875
rect 800 822 883 825
rect 1624 833 1762 868
rect 1624 797 1667 833
rect 1749 823 1762 833
rect 1814 823 1832 875
rect 1895 827 1911 879
rect 1963 827 1978 879
rect 2344 881 2427 883
rect 2344 829 2358 881
rect 2410 829 2427 881
rect 2344 827 2427 829
rect 2491 879 2574 883
rect 2491 827 2506 879
rect 2558 827 2574 879
rect 1895 824 1978 827
rect 2491 825 2574 827
rect 1749 821 1832 823
rect 898 756 1667 797
rect 1907 786 1966 824
rect 2503 791 2562 825
rect 3008 791 3113 1223
rect 3549 876 3632 879
rect 3549 824 3564 876
rect 3616 824 3632 876
rect 3549 821 3632 824
rect 3702 872 3777 878
rect 3702 820 3712 872
rect 3764 820 3777 872
rect 4137 876 4220 880
rect 4137 824 4151 876
rect 4203 824 4220 876
rect 4137 822 4220 824
rect 4286 873 4367 880
rect 3702 791 3777 820
rect 4286 821 4300 873
rect 4352 821 4367 873
rect 4286 815 4367 821
rect 356 511 784 713
rect 898 511 932 756
rect 1698 754 1966 786
rect 2294 759 2562 791
rect 356 205 477 511
rect 1260 205 1329 546
rect 1698 511 1732 754
rect 1842 449 1882 715
rect 1838 444 1905 449
rect 1838 392 1845 444
rect 1897 392 1905 444
rect 1838 385 1905 392
rect 1993 205 2028 713
rect 2294 511 2328 759
rect 3499 754 3777 791
rect 4287 786 4362 815
rect 4085 756 4362 786
rect 2439 449 2479 713
rect 2417 445 2485 449
rect 2417 393 2426 445
rect 2478 393 2485 445
rect 2417 388 2485 393
rect 2589 205 2624 725
rect 3008 205 3113 649
rect 3499 511 3535 754
rect 3648 429 3682 713
rect 3647 421 3722 429
rect 3647 369 3657 421
rect 3709 369 3722 421
rect 3647 361 3722 369
rect 3795 205 3830 726
rect 4085 510 4121 756
rect 4234 431 4268 714
rect 4192 423 4268 431
rect 4192 371 4204 423
rect 4256 393 4268 423
rect 4256 371 4267 393
rect 4192 363 4267 371
rect 4381 205 4416 726
rect 356 74 4427 205
<< via1 >>
rect 741 3987 793 4039
rect 889 3987 941 4039
rect 1910 4038 1962 4090
rect 2059 4038 2111 4090
rect 2505 4034 2557 4086
rect 2651 4034 2703 4086
rect 1615 2401 1667 2453
rect 1762 2400 1814 2452
rect 2207 2399 2259 2451
rect 2354 2400 2406 2452
rect 3709 4047 3761 4099
rect 3854 4051 3906 4103
rect 3409 2418 3461 2470
rect 3557 2419 3609 2471
rect 4297 4051 4349 4103
rect 4445 4051 4497 4103
rect 4000 2420 4052 2472
rect 4149 2420 4201 2472
rect 1908 1881 1960 1933
rect 3546 1880 3598 1932
rect 1908 1817 1960 1869
rect 3546 1816 3598 1868
rect 746 1538 926 1654
rect 2343 1603 2395 1655
rect 2343 1539 2395 1591
rect 2506 1373 2558 1425
rect 4143 1372 4195 1424
rect 2506 1309 2558 1361
rect 4143 1308 4195 1360
rect 815 825 867 877
rect 1762 823 1814 875
rect 1911 827 1963 879
rect 2358 829 2410 881
rect 2506 827 2558 879
rect 3564 824 3616 876
rect 3712 820 3764 872
rect 4151 824 4203 876
rect 4300 821 4352 873
rect 1845 392 1897 444
rect 2426 393 2478 445
rect 3657 369 3709 421
rect 4204 371 4256 423
<< metal2 >>
rect 3696 4103 3925 4110
rect 3696 4099 3854 4103
rect 1894 4090 2127 4097
rect 710 4039 965 4048
rect 710 3993 741 4039
rect 709 3987 741 3993
rect 793 3987 889 4039
rect 941 3987 965 4039
rect 1894 4038 1910 4090
rect 1962 4038 2059 4090
rect 2111 4038 2127 4090
rect 1894 4026 2127 4038
rect 2491 4086 2724 4093
rect 2491 4034 2505 4086
rect 2557 4034 2651 4086
rect 2703 4034 2724 4086
rect 2491 4026 2724 4034
rect 3696 4047 3709 4099
rect 3761 4051 3854 4099
rect 3906 4051 3925 4103
rect 3761 4047 3925 4051
rect 3696 4040 3925 4047
rect 4284 4103 4517 4112
rect 4284 4051 4297 4103
rect 4349 4051 4445 4103
rect 4497 4051 4517 4103
rect 4284 4045 4517 4051
rect 709 1756 812 3987
rect 1894 2712 1977 4026
rect 1594 2453 1836 2460
rect 1594 2401 1615 2453
rect 1667 2452 1836 2453
rect 1667 2401 1762 2452
rect 1594 2400 1762 2401
rect 1814 2400 1836 2452
rect 1594 2383 1836 2400
rect 709 1683 964 1756
rect 710 1681 964 1683
rect 710 1654 965 1681
rect 710 1538 746 1654
rect 926 1538 965 1654
rect 710 877 965 1538
rect 710 825 815 877
rect 867 825 965 877
rect 710 818 965 825
rect 1717 875 1836 2383
rect 1717 823 1762 875
rect 1814 823 1836 875
rect 1717 814 1836 823
rect 1893 1933 1977 2712
rect 2187 2452 2431 2459
rect 2187 2451 2354 2452
rect 2187 2399 2207 2451
rect 2259 2400 2354 2451
rect 2406 2400 2431 2452
rect 2259 2399 2431 2400
rect 2187 2384 2431 2399
rect 1893 1881 1908 1933
rect 1960 1881 1977 1933
rect 1893 1869 1977 1881
rect 1893 1817 1908 1869
rect 1960 1817 1977 1869
rect 1893 879 1977 1817
rect 1893 827 1911 879
rect 1963 827 1977 879
rect 1893 819 1977 827
rect 2312 1655 2431 2384
rect 2312 1603 2343 1655
rect 2395 1603 2431 1655
rect 2312 1591 2431 1603
rect 2312 1539 2343 1591
rect 2395 1539 2431 1591
rect 2312 881 2431 1539
rect 2312 829 2358 881
rect 2410 829 2431 881
rect 2312 821 2431 829
rect 2491 1425 2574 4026
rect 3390 2471 3634 2481
rect 3390 2470 3557 2471
rect 3390 2418 3409 2470
rect 3461 2419 3557 2470
rect 3609 2419 3634 2471
rect 3461 2418 3634 2419
rect 3390 2406 3634 2418
rect 2491 1373 2506 1425
rect 2558 1373 2574 1425
rect 2491 1361 2574 1373
rect 2491 1309 2506 1361
rect 2558 1309 2574 1361
rect 2491 879 2574 1309
rect 2491 827 2506 879
rect 2558 827 2574 879
rect 2491 805 2574 827
rect 3515 1932 3634 2406
rect 3515 1880 3546 1932
rect 3598 1880 3634 1932
rect 3515 1868 3634 1880
rect 3515 1816 3546 1868
rect 3598 1816 3634 1868
rect 3515 876 3634 1816
rect 3515 824 3564 876
rect 3616 824 3634 876
rect 3515 816 3634 824
rect 3696 872 3774 4040
rect 3983 2472 4229 2482
rect 3983 2420 4000 2472
rect 4052 2420 4149 2472
rect 4201 2420 4229 2472
rect 3983 2400 4229 2420
rect 3696 820 3712 872
rect 3764 820 3774 872
rect 3696 814 3774 820
rect 4110 1424 4229 2400
rect 4110 1372 4143 1424
rect 4195 1372 4229 1424
rect 4110 1360 4229 1372
rect 4110 1308 4143 1360
rect 4195 1308 4229 1360
rect 4110 876 4229 1308
rect 4110 824 4151 876
rect 4203 824 4229 876
rect 4110 802 4229 824
rect 4284 873 4370 4045
rect 4284 821 4300 873
rect 4352 821 4370 873
rect 4284 814 4370 821
rect 1838 455 1888 720
rect 2436 455 2486 719
rect 1838 445 2486 455
rect 1838 444 2426 445
rect 1838 392 1845 444
rect 1897 393 2426 444
rect 2478 393 2486 445
rect 1897 392 2486 393
rect 1838 383 2486 392
rect 1898 382 2486 383
rect 3641 436 3688 727
rect 4227 436 4277 724
rect 3641 423 4277 436
rect 3641 421 4204 423
rect 3641 369 3657 421
rect 3709 371 4204 421
rect 4256 371 4277 423
rect 3709 369 4277 371
rect 3641 356 4277 369
rect 3641 355 4275 356
use sky130_fd_pr__pfet_01v8_BKDUYV  XM3
timestamp 1669522153
transform -1 0 2307 0 -1 3207
box -213 -780 213 847
use sky130_fd_pr__nfet_01v8_RFHF3H  XM4
timestamp 1669522153
transform 1 0 2384 0 1 643
box -129 -170 129 240
use sky130_fd_pr__pfet_01v8_BKDUYV  XM5
timestamp 1669522153
transform 1 0 2603 0 1 3278
box -213 -780 213 847
use sky130_fd_pr__nfet_01v8_RFHF3H  XM6
timestamp 1669522153
transform -1 0 2532 0 1 643
box -129 -170 129 240
use sky130_fd_pr__pfet_01v8_BKDUYV  XM7
timestamp 1669522153
transform -1 0 1715 0 -1 3207
box -213 -780 213 847
use sky130_fd_pr__pfet_01v8_BKDUYV  XM8
timestamp 1669522153
transform -1 0 4102 0 -1 3229
box -213 -780 213 847
use sky130_fd_pr__pfet_01v8_BKDUYV  XM9
timestamp 1669522153
transform -1 0 3510 0 -1 3229
box -213 -780 213 847
use sky130_fd_pr__pfet_01v8_BKDUYV  XM10
timestamp 1669522153
transform 1 0 2011 0 1 3278
box -213 -780 213 847
use sky130_fd_pr__pfet_01v8_BKDUYV  XM11
timestamp 1669522153
transform 1 0 4398 0 1 3300
box -213 -780 213 847
use sky130_fd_pr__pfet_01v8_BKDUYV  XM12
timestamp 1669522153
transform 1 0 3806 0 1 3300
box -213 -780 213 847
use sky130_fd_pr__nfet_01v8_RFHF3H  XM13
timestamp 1669522153
transform 1 0 1790 0 1 643
box -129 -170 129 240
use sky130_fd_pr__nfet_01v8_RFHF3H  XM14
timestamp 1669522153
transform 1 0 4178 0 1 643
box -129 -170 129 240
use sky130_fd_pr__nfet_01v8_RFHF3H  XM15
timestamp 1669522153
transform 1 0 3590 0 1 643
box -129 -170 129 240
use sky130_fd_pr__nfet_01v8_RFHF3H  XM16
timestamp 1669522153
transform 1 0 1938 0 1 643
box -129 -170 129 240
use sky130_fd_pr__nfet_01v8_RFHF3H  XM17
timestamp 1669522153
transform 1 0 4326 0 1 643
box -129 -170 129 240
use sky130_fd_pr__nfet_01v8_RFHF3H  sky130_fd_pr__nfet_01v8_RFHF3H_0
timestamp 1669522153
transform 1 0 841 0 1 643
box -129 -170 129 240
use sky130_fd_pr__nfet_01v8_RFHF3H  sky130_fd_pr__nfet_01v8_RFHF3H_1
timestamp 1669522153
transform -1 0 3738 0 1 643
box -129 -170 129 240
use sky130_fd_pr__pfet_01v8_BKDUYV  sky130_fd_pr__pfet_01v8_BKDUYV_0
timestamp 1669522153
transform 1 0 841 0 1 3233
box -213 -780 213 847
<< labels >>
rlabel metal1 s 1050 1624 1050 1624 4 Vin
port 1 nsew
rlabel metal1 s 4584 2156 4584 2156 4 Vdd
port 2 nsew
rlabel metal1 s 4254 3052 4254 3052 4 Vs11
port 3 nsew
rlabel metal1 s 2452 2640 2452 2640 4 Vs5
port 4 nsew
rlabel metal2 s 3738 916 3738 916 4 Voutinverted
port 5 nsew
rlabel metal2 s 4328 906 4328 906 4 Voutfinal
port 6 nsew
rlabel metal2 s 1930 930 1930 930 4 Vout3
port 7 nsew
rlabel metal2 s 1750 942 1750 942 4 Vout1
port 8 nsew
rlabel metal2 s 4246 626 4246 626 4 Vs14
port 9 nsew
rlabel metal2 s 2546 916 2546 916 4 Vout2
port 10 nsew
rlabel metal2 s 2456 526 2456 526 4 Vs4
port 11 nsew
<< end >>
