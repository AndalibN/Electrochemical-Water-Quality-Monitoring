magic
tech sky130A
magscale 1 2
timestamp 1667331940
<< pwell >>
rect -201 -793 201 793
<< psubdiff >>
rect -165 723 -69 757
rect 69 723 165 757
rect -165 661 -131 723
rect 131 661 165 723
rect -165 -723 -131 -661
rect 131 -723 165 -661
rect -165 -757 -69 -723
rect 69 -757 165 -723
<< psubdiffcont >>
rect -69 723 69 757
rect -165 -661 -131 661
rect 131 -661 165 661
rect -69 -757 69 -723
<< xpolycontact >>
rect -35 195 35 627
rect -35 -627 35 -195
<< ppolyres >>
rect -35 -195 35 195
<< locali >>
rect -165 723 -69 757
rect 69 723 165 757
rect -165 661 -131 723
rect 131 661 165 723
rect -165 -723 -131 -661
rect 131 -723 165 -661
rect -165 -757 -69 -723
rect 69 -757 165 -723
<< viali >>
rect -19 212 19 609
rect -19 -609 19 -212
<< metal1 >>
rect -25 609 25 621
rect -25 212 -19 609
rect 19 212 25 609
rect -25 200 25 212
rect -25 -212 25 -200
rect -25 -609 -19 -212
rect 19 -609 25 -212
rect -25 -621 25 -609
<< res0p35 >>
rect -37 -197 37 197
<< properties >>
string FIXED_BBOX -148 -740 148 740
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 1.95 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.895k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
