magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 372 29 378
rect -29 338 -17 372
rect -29 332 29 338
rect -29 -338 29 -332
rect -29 -372 -17 -338
rect -29 -378 29 -372
<< pwell >>
rect -114 -326 114 326
<< nmos >>
rect -30 -300 30 300
<< ndiff >>
rect -88 255 -30 300
rect -88 221 -76 255
rect -42 221 -30 255
rect -88 187 -30 221
rect -88 153 -76 187
rect -42 153 -30 187
rect -88 119 -30 153
rect -88 85 -76 119
rect -42 85 -30 119
rect -88 51 -30 85
rect -88 17 -76 51
rect -42 17 -30 51
rect -88 -17 -30 17
rect -88 -51 -76 -17
rect -42 -51 -30 -17
rect -88 -85 -30 -51
rect -88 -119 -76 -85
rect -42 -119 -30 -85
rect -88 -153 -30 -119
rect -88 -187 -76 -153
rect -42 -187 -30 -153
rect -88 -221 -30 -187
rect -88 -255 -76 -221
rect -42 -255 -30 -221
rect -88 -300 -30 -255
rect 30 255 88 300
rect 30 221 42 255
rect 76 221 88 255
rect 30 187 88 221
rect 30 153 42 187
rect 76 153 88 187
rect 30 119 88 153
rect 30 85 42 119
rect 76 85 88 119
rect 30 51 88 85
rect 30 17 42 51
rect 76 17 88 51
rect 30 -17 88 17
rect 30 -51 42 -17
rect 76 -51 88 -17
rect 30 -85 88 -51
rect 30 -119 42 -85
rect 76 -119 88 -85
rect 30 -153 88 -119
rect 30 -187 42 -153
rect 76 -187 88 -153
rect 30 -221 88 -187
rect 30 -255 42 -221
rect 76 -255 88 -221
rect 30 -300 88 -255
<< ndiffc >>
rect -76 221 -42 255
rect -76 153 -42 187
rect -76 85 -42 119
rect -76 17 -42 51
rect -76 -51 -42 -17
rect -76 -119 -42 -85
rect -76 -187 -42 -153
rect -76 -255 -42 -221
rect 42 221 76 255
rect 42 153 76 187
rect 42 85 76 119
rect 42 17 76 51
rect 42 -51 76 -17
rect 42 -119 76 -85
rect 42 -187 76 -153
rect 42 -255 76 -221
<< poly >>
rect -33 372 33 388
rect -33 338 -17 372
rect 17 338 33 372
rect -33 322 33 338
rect -30 300 30 322
rect -30 -322 30 -300
rect -33 -338 33 -322
rect -33 -372 -17 -338
rect 17 -372 33 -338
rect -33 -388 33 -372
<< polycont >>
rect -17 338 17 372
rect -17 -372 17 -338
<< locali >>
rect -33 338 -17 372
rect 17 338 33 372
rect -76 269 -42 304
rect -76 197 -42 221
rect -76 125 -42 153
rect -76 53 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -53
rect -76 -153 -42 -125
rect -76 -221 -42 -197
rect -76 -304 -42 -269
rect 42 269 76 304
rect 42 197 76 221
rect 42 125 76 153
rect 42 53 76 85
rect 42 -17 76 17
rect 42 -85 76 -53
rect 42 -153 76 -125
rect 42 -221 76 -197
rect 42 -304 76 -269
rect -33 -372 -17 -338
rect 17 -372 33 -338
<< viali >>
rect -17 338 17 372
rect -76 255 -42 269
rect -76 235 -42 255
rect -76 187 -42 197
rect -76 163 -42 187
rect -76 119 -42 125
rect -76 91 -42 119
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect -76 -119 -42 -91
rect -76 -125 -42 -119
rect -76 -187 -42 -163
rect -76 -197 -42 -187
rect -76 -255 -42 -235
rect -76 -269 -42 -255
rect 42 255 76 269
rect 42 235 76 255
rect 42 187 76 197
rect 42 163 76 187
rect 42 119 76 125
rect 42 91 76 119
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect 42 -119 76 -91
rect 42 -125 76 -119
rect 42 -187 76 -163
rect 42 -197 76 -187
rect 42 -255 76 -235
rect 42 -269 76 -255
rect -17 -372 17 -338
<< metal1 >>
rect -29 372 29 378
rect -29 338 -17 372
rect 17 338 29 372
rect -29 332 29 338
rect -82 269 -36 300
rect -82 235 -76 269
rect -42 235 -36 269
rect -82 197 -36 235
rect -82 163 -76 197
rect -42 163 -36 197
rect -82 125 -36 163
rect -82 91 -76 125
rect -42 91 -36 125
rect -82 53 -36 91
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -91 -36 -53
rect -82 -125 -76 -91
rect -42 -125 -36 -91
rect -82 -163 -36 -125
rect -82 -197 -76 -163
rect -42 -197 -36 -163
rect -82 -235 -36 -197
rect -82 -269 -76 -235
rect -42 -269 -36 -235
rect -82 -300 -36 -269
rect 36 269 82 300
rect 36 235 42 269
rect 76 235 82 269
rect 36 197 82 235
rect 36 163 42 197
rect 76 163 82 197
rect 36 125 82 163
rect 36 91 42 125
rect 76 91 82 125
rect 36 53 82 91
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -91 82 -53
rect 36 -125 42 -91
rect 76 -125 82 -91
rect 36 -163 82 -125
rect 36 -197 42 -163
rect 76 -197 82 -163
rect 36 -235 82 -197
rect 36 -269 42 -235
rect 76 -269 82 -235
rect 36 -300 82 -269
rect -29 -338 29 -332
rect -29 -372 -17 -338
rect 17 -372 29 -338
rect -29 -378 29 -372
<< end >>
