magic
tech sky130B
timestamp 1658697764
<< metal4 >>
rect 2300 -2850 2800 700
rect 2300 -3000 2350 -2850
rect 2500 -3000 2550 -2850
rect 2700 -3000 2800 -2850
rect 2300 -3050 2800 -3000
rect 2300 -3200 2400 -3050
rect 2550 -3200 2600 -3050
rect 2750 -3200 2800 -3050
rect 2300 -3300 2800 -3200
<< via4 >>
rect 2350 -3000 2500 -2850
rect 2550 -3000 2700 -2850
rect 2400 -3200 2550 -3050
rect 2600 -3200 2750 -3050
<< metal5 >>
rect -100 -100 9900 400
rect -100 -900 9100 -400
rect -100 -9100 400 -900
rect 700 -1700 8300 -1200
rect 700 -8300 1200 -1700
rect 1500 -2500 7500 -2000
rect 1500 -7500 2000 -2500
rect 2300 -2850 2800 -2800
rect 2300 -3000 2350 -2850
rect 2500 -3000 2550 -2850
rect 2700 -3000 2800 -2850
rect 2300 -3050 2800 -3000
rect 2300 -3200 2400 -3050
rect 2550 -3200 2600 -3050
rect 2750 -3200 2800 -3050
rect 2300 -6700 2800 -3200
rect 7000 -6700 7500 -2500
rect 2300 -7200 7500 -6700
rect 7800 -7500 8300 -1700
rect 1500 -8000 8300 -7500
rect 8600 -8300 9100 -900
rect 700 -8800 9100 -8300
rect 9400 -9100 9900 -100
rect -100 -9600 9900 -9100
<< end >>
