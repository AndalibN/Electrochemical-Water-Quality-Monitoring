magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 405 29 411
rect -29 371 -17 405
rect -29 365 29 371
<< nwell >>
rect -112 -458 112 424
<< pmos >>
rect -18 -396 18 324
<< pdiff >>
rect -76 287 -18 324
rect -76 253 -64 287
rect -30 253 -18 287
rect -76 219 -18 253
rect -76 185 -64 219
rect -30 185 -18 219
rect -76 151 -18 185
rect -76 117 -64 151
rect -30 117 -18 151
rect -76 83 -18 117
rect -76 49 -64 83
rect -30 49 -18 83
rect -76 15 -18 49
rect -76 -19 -64 15
rect -30 -19 -18 15
rect -76 -53 -18 -19
rect -76 -87 -64 -53
rect -30 -87 -18 -53
rect -76 -121 -18 -87
rect -76 -155 -64 -121
rect -30 -155 -18 -121
rect -76 -189 -18 -155
rect -76 -223 -64 -189
rect -30 -223 -18 -189
rect -76 -257 -18 -223
rect -76 -291 -64 -257
rect -30 -291 -18 -257
rect -76 -325 -18 -291
rect -76 -359 -64 -325
rect -30 -359 -18 -325
rect -76 -396 -18 -359
rect 18 287 76 324
rect 18 253 30 287
rect 64 253 76 287
rect 18 219 76 253
rect 18 185 30 219
rect 64 185 76 219
rect 18 151 76 185
rect 18 117 30 151
rect 64 117 76 151
rect 18 83 76 117
rect 18 49 30 83
rect 64 49 76 83
rect 18 15 76 49
rect 18 -19 30 15
rect 64 -19 76 15
rect 18 -53 76 -19
rect 18 -87 30 -53
rect 64 -87 76 -53
rect 18 -121 76 -87
rect 18 -155 30 -121
rect 64 -155 76 -121
rect 18 -189 76 -155
rect 18 -223 30 -189
rect 64 -223 76 -189
rect 18 -257 76 -223
rect 18 -291 30 -257
rect 64 -291 76 -257
rect 18 -325 76 -291
rect 18 -359 30 -325
rect 64 -359 76 -325
rect 18 -396 76 -359
<< pdiffc >>
rect -64 253 -30 287
rect -64 185 -30 219
rect -64 117 -30 151
rect -64 49 -30 83
rect -64 -19 -30 15
rect -64 -87 -30 -53
rect -64 -155 -30 -121
rect -64 -223 -30 -189
rect -64 -291 -30 -257
rect -64 -359 -30 -325
rect 30 253 64 287
rect 30 185 64 219
rect 30 117 64 151
rect 30 49 64 83
rect 30 -19 64 15
rect 30 -87 64 -53
rect 30 -155 64 -121
rect 30 -223 64 -189
rect 30 -291 64 -257
rect 30 -359 64 -325
<< poly >>
rect -33 405 33 421
rect -33 371 -17 405
rect 17 371 33 405
rect -33 355 33 371
rect -18 324 18 355
rect -18 -422 18 -396
<< polycont >>
rect -17 371 17 405
<< locali >>
rect -33 371 -17 405
rect 17 371 33 405
rect -64 305 -30 328
rect -64 233 -30 253
rect -64 161 -30 185
rect -64 89 -30 117
rect -64 17 -30 49
rect -64 -53 -30 -19
rect -64 -121 -30 -89
rect -64 -189 -30 -161
rect -64 -257 -30 -233
rect -64 -325 -30 -305
rect -64 -400 -30 -377
rect 30 305 64 328
rect 30 233 64 253
rect 30 161 64 185
rect 30 89 64 117
rect 30 17 64 49
rect 30 -53 64 -19
rect 30 -121 64 -89
rect 30 -189 64 -161
rect 30 -257 64 -233
rect 30 -325 64 -305
rect 30 -400 64 -377
<< viali >>
rect -17 371 17 405
rect -64 287 -30 305
rect -64 271 -30 287
rect -64 219 -30 233
rect -64 199 -30 219
rect -64 151 -30 161
rect -64 127 -30 151
rect -64 83 -30 89
rect -64 55 -30 83
rect -64 15 -30 17
rect -64 -17 -30 15
rect -64 -87 -30 -55
rect -64 -89 -30 -87
rect -64 -155 -30 -127
rect -64 -161 -30 -155
rect -64 -223 -30 -199
rect -64 -233 -30 -223
rect -64 -291 -30 -271
rect -64 -305 -30 -291
rect -64 -359 -30 -343
rect -64 -377 -30 -359
rect 30 287 64 305
rect 30 271 64 287
rect 30 219 64 233
rect 30 199 64 219
rect 30 151 64 161
rect 30 127 64 151
rect 30 83 64 89
rect 30 55 64 83
rect 30 15 64 17
rect 30 -17 64 15
rect 30 -87 64 -55
rect 30 -89 64 -87
rect 30 -155 64 -127
rect 30 -161 64 -155
rect 30 -223 64 -199
rect 30 -233 64 -223
rect 30 -291 64 -271
rect 30 -305 64 -291
rect 30 -359 64 -343
rect 30 -377 64 -359
<< metal1 >>
rect -29 405 29 411
rect -29 371 -17 405
rect 17 371 29 405
rect -29 365 29 371
rect -70 305 -24 324
rect -70 271 -64 305
rect -30 271 -24 305
rect -70 233 -24 271
rect -70 199 -64 233
rect -30 199 -24 233
rect -70 161 -24 199
rect -70 127 -64 161
rect -30 127 -24 161
rect -70 89 -24 127
rect -70 55 -64 89
rect -30 55 -24 89
rect -70 17 -24 55
rect -70 -17 -64 17
rect -30 -17 -24 17
rect -70 -55 -24 -17
rect -70 -89 -64 -55
rect -30 -89 -24 -55
rect -70 -127 -24 -89
rect -70 -161 -64 -127
rect -30 -161 -24 -127
rect -70 -199 -24 -161
rect -70 -233 -64 -199
rect -30 -233 -24 -199
rect -70 -271 -24 -233
rect -70 -305 -64 -271
rect -30 -305 -24 -271
rect -70 -343 -24 -305
rect -70 -377 -64 -343
rect -30 -377 -24 -343
rect -70 -396 -24 -377
rect 24 305 70 324
rect 24 271 30 305
rect 64 271 70 305
rect 24 233 70 271
rect 24 199 30 233
rect 64 199 70 233
rect 24 161 70 199
rect 24 127 30 161
rect 64 127 70 161
rect 24 89 70 127
rect 24 55 30 89
rect 64 55 70 89
rect 24 17 70 55
rect 24 -17 30 17
rect 64 -17 70 17
rect 24 -55 70 -17
rect 24 -89 30 -55
rect 64 -89 70 -55
rect 24 -127 70 -89
rect 24 -161 30 -127
rect 64 -161 70 -127
rect 24 -199 70 -161
rect 24 -233 30 -199
rect 64 -233 70 -199
rect 24 -271 70 -233
rect 24 -305 30 -271
rect 64 -305 70 -271
rect 24 -343 70 -305
rect 24 -377 30 -343
rect 64 -377 70 -343
rect 24 -396 70 -377
<< end >>
