magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -294 -2100 294 2100
<< pmos >>
rect -200 -2000 200 2000
<< pdiff >>
rect -258 1955 -200 2000
rect -258 1921 -246 1955
rect -212 1921 -200 1955
rect -258 1887 -200 1921
rect -258 1853 -246 1887
rect -212 1853 -200 1887
rect -258 1819 -200 1853
rect -258 1785 -246 1819
rect -212 1785 -200 1819
rect -258 1751 -200 1785
rect -258 1717 -246 1751
rect -212 1717 -200 1751
rect -258 1683 -200 1717
rect -258 1649 -246 1683
rect -212 1649 -200 1683
rect -258 1615 -200 1649
rect -258 1581 -246 1615
rect -212 1581 -200 1615
rect -258 1547 -200 1581
rect -258 1513 -246 1547
rect -212 1513 -200 1547
rect -258 1479 -200 1513
rect -258 1445 -246 1479
rect -212 1445 -200 1479
rect -258 1411 -200 1445
rect -258 1377 -246 1411
rect -212 1377 -200 1411
rect -258 1343 -200 1377
rect -258 1309 -246 1343
rect -212 1309 -200 1343
rect -258 1275 -200 1309
rect -258 1241 -246 1275
rect -212 1241 -200 1275
rect -258 1207 -200 1241
rect -258 1173 -246 1207
rect -212 1173 -200 1207
rect -258 1139 -200 1173
rect -258 1105 -246 1139
rect -212 1105 -200 1139
rect -258 1071 -200 1105
rect -258 1037 -246 1071
rect -212 1037 -200 1071
rect -258 1003 -200 1037
rect -258 969 -246 1003
rect -212 969 -200 1003
rect -258 935 -200 969
rect -258 901 -246 935
rect -212 901 -200 935
rect -258 867 -200 901
rect -258 833 -246 867
rect -212 833 -200 867
rect -258 799 -200 833
rect -258 765 -246 799
rect -212 765 -200 799
rect -258 731 -200 765
rect -258 697 -246 731
rect -212 697 -200 731
rect -258 663 -200 697
rect -258 629 -246 663
rect -212 629 -200 663
rect -258 595 -200 629
rect -258 561 -246 595
rect -212 561 -200 595
rect -258 527 -200 561
rect -258 493 -246 527
rect -212 493 -200 527
rect -258 459 -200 493
rect -258 425 -246 459
rect -212 425 -200 459
rect -258 391 -200 425
rect -258 357 -246 391
rect -212 357 -200 391
rect -258 323 -200 357
rect -258 289 -246 323
rect -212 289 -200 323
rect -258 255 -200 289
rect -258 221 -246 255
rect -212 221 -200 255
rect -258 187 -200 221
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -221 -200 -187
rect -258 -255 -246 -221
rect -212 -255 -200 -221
rect -258 -289 -200 -255
rect -258 -323 -246 -289
rect -212 -323 -200 -289
rect -258 -357 -200 -323
rect -258 -391 -246 -357
rect -212 -391 -200 -357
rect -258 -425 -200 -391
rect -258 -459 -246 -425
rect -212 -459 -200 -425
rect -258 -493 -200 -459
rect -258 -527 -246 -493
rect -212 -527 -200 -493
rect -258 -561 -200 -527
rect -258 -595 -246 -561
rect -212 -595 -200 -561
rect -258 -629 -200 -595
rect -258 -663 -246 -629
rect -212 -663 -200 -629
rect -258 -697 -200 -663
rect -258 -731 -246 -697
rect -212 -731 -200 -697
rect -258 -765 -200 -731
rect -258 -799 -246 -765
rect -212 -799 -200 -765
rect -258 -833 -200 -799
rect -258 -867 -246 -833
rect -212 -867 -200 -833
rect -258 -901 -200 -867
rect -258 -935 -246 -901
rect -212 -935 -200 -901
rect -258 -969 -200 -935
rect -258 -1003 -246 -969
rect -212 -1003 -200 -969
rect -258 -1037 -200 -1003
rect -258 -1071 -246 -1037
rect -212 -1071 -200 -1037
rect -258 -1105 -200 -1071
rect -258 -1139 -246 -1105
rect -212 -1139 -200 -1105
rect -258 -1173 -200 -1139
rect -258 -1207 -246 -1173
rect -212 -1207 -200 -1173
rect -258 -1241 -200 -1207
rect -258 -1275 -246 -1241
rect -212 -1275 -200 -1241
rect -258 -1309 -200 -1275
rect -258 -1343 -246 -1309
rect -212 -1343 -200 -1309
rect -258 -1377 -200 -1343
rect -258 -1411 -246 -1377
rect -212 -1411 -200 -1377
rect -258 -1445 -200 -1411
rect -258 -1479 -246 -1445
rect -212 -1479 -200 -1445
rect -258 -1513 -200 -1479
rect -258 -1547 -246 -1513
rect -212 -1547 -200 -1513
rect -258 -1581 -200 -1547
rect -258 -1615 -246 -1581
rect -212 -1615 -200 -1581
rect -258 -1649 -200 -1615
rect -258 -1683 -246 -1649
rect -212 -1683 -200 -1649
rect -258 -1717 -200 -1683
rect -258 -1751 -246 -1717
rect -212 -1751 -200 -1717
rect -258 -1785 -200 -1751
rect -258 -1819 -246 -1785
rect -212 -1819 -200 -1785
rect -258 -1853 -200 -1819
rect -258 -1887 -246 -1853
rect -212 -1887 -200 -1853
rect -258 -1921 -200 -1887
rect -258 -1955 -246 -1921
rect -212 -1955 -200 -1921
rect -258 -2000 -200 -1955
rect 200 1955 258 2000
rect 200 1921 212 1955
rect 246 1921 258 1955
rect 200 1887 258 1921
rect 200 1853 212 1887
rect 246 1853 258 1887
rect 200 1819 258 1853
rect 200 1785 212 1819
rect 246 1785 258 1819
rect 200 1751 258 1785
rect 200 1717 212 1751
rect 246 1717 258 1751
rect 200 1683 258 1717
rect 200 1649 212 1683
rect 246 1649 258 1683
rect 200 1615 258 1649
rect 200 1581 212 1615
rect 246 1581 258 1615
rect 200 1547 258 1581
rect 200 1513 212 1547
rect 246 1513 258 1547
rect 200 1479 258 1513
rect 200 1445 212 1479
rect 246 1445 258 1479
rect 200 1411 258 1445
rect 200 1377 212 1411
rect 246 1377 258 1411
rect 200 1343 258 1377
rect 200 1309 212 1343
rect 246 1309 258 1343
rect 200 1275 258 1309
rect 200 1241 212 1275
rect 246 1241 258 1275
rect 200 1207 258 1241
rect 200 1173 212 1207
rect 246 1173 258 1207
rect 200 1139 258 1173
rect 200 1105 212 1139
rect 246 1105 258 1139
rect 200 1071 258 1105
rect 200 1037 212 1071
rect 246 1037 258 1071
rect 200 1003 258 1037
rect 200 969 212 1003
rect 246 969 258 1003
rect 200 935 258 969
rect 200 901 212 935
rect 246 901 258 935
rect 200 867 258 901
rect 200 833 212 867
rect 246 833 258 867
rect 200 799 258 833
rect 200 765 212 799
rect 246 765 258 799
rect 200 731 258 765
rect 200 697 212 731
rect 246 697 258 731
rect 200 663 258 697
rect 200 629 212 663
rect 246 629 258 663
rect 200 595 258 629
rect 200 561 212 595
rect 246 561 258 595
rect 200 527 258 561
rect 200 493 212 527
rect 246 493 258 527
rect 200 459 258 493
rect 200 425 212 459
rect 246 425 258 459
rect 200 391 258 425
rect 200 357 212 391
rect 246 357 258 391
rect 200 323 258 357
rect 200 289 212 323
rect 246 289 258 323
rect 200 255 258 289
rect 200 221 212 255
rect 246 221 258 255
rect 200 187 258 221
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -221 258 -187
rect 200 -255 212 -221
rect 246 -255 258 -221
rect 200 -289 258 -255
rect 200 -323 212 -289
rect 246 -323 258 -289
rect 200 -357 258 -323
rect 200 -391 212 -357
rect 246 -391 258 -357
rect 200 -425 258 -391
rect 200 -459 212 -425
rect 246 -459 258 -425
rect 200 -493 258 -459
rect 200 -527 212 -493
rect 246 -527 258 -493
rect 200 -561 258 -527
rect 200 -595 212 -561
rect 246 -595 258 -561
rect 200 -629 258 -595
rect 200 -663 212 -629
rect 246 -663 258 -629
rect 200 -697 258 -663
rect 200 -731 212 -697
rect 246 -731 258 -697
rect 200 -765 258 -731
rect 200 -799 212 -765
rect 246 -799 258 -765
rect 200 -833 258 -799
rect 200 -867 212 -833
rect 246 -867 258 -833
rect 200 -901 258 -867
rect 200 -935 212 -901
rect 246 -935 258 -901
rect 200 -969 258 -935
rect 200 -1003 212 -969
rect 246 -1003 258 -969
rect 200 -1037 258 -1003
rect 200 -1071 212 -1037
rect 246 -1071 258 -1037
rect 200 -1105 258 -1071
rect 200 -1139 212 -1105
rect 246 -1139 258 -1105
rect 200 -1173 258 -1139
rect 200 -1207 212 -1173
rect 246 -1207 258 -1173
rect 200 -1241 258 -1207
rect 200 -1275 212 -1241
rect 246 -1275 258 -1241
rect 200 -1309 258 -1275
rect 200 -1343 212 -1309
rect 246 -1343 258 -1309
rect 200 -1377 258 -1343
rect 200 -1411 212 -1377
rect 246 -1411 258 -1377
rect 200 -1445 258 -1411
rect 200 -1479 212 -1445
rect 246 -1479 258 -1445
rect 200 -1513 258 -1479
rect 200 -1547 212 -1513
rect 246 -1547 258 -1513
rect 200 -1581 258 -1547
rect 200 -1615 212 -1581
rect 246 -1615 258 -1581
rect 200 -1649 258 -1615
rect 200 -1683 212 -1649
rect 246 -1683 258 -1649
rect 200 -1717 258 -1683
rect 200 -1751 212 -1717
rect 246 -1751 258 -1717
rect 200 -1785 258 -1751
rect 200 -1819 212 -1785
rect 246 -1819 258 -1785
rect 200 -1853 258 -1819
rect 200 -1887 212 -1853
rect 246 -1887 258 -1853
rect 200 -1921 258 -1887
rect 200 -1955 212 -1921
rect 246 -1955 258 -1921
rect 200 -2000 258 -1955
<< pdiffc >>
rect -246 1921 -212 1955
rect -246 1853 -212 1887
rect -246 1785 -212 1819
rect -246 1717 -212 1751
rect -246 1649 -212 1683
rect -246 1581 -212 1615
rect -246 1513 -212 1547
rect -246 1445 -212 1479
rect -246 1377 -212 1411
rect -246 1309 -212 1343
rect -246 1241 -212 1275
rect -246 1173 -212 1207
rect -246 1105 -212 1139
rect -246 1037 -212 1071
rect -246 969 -212 1003
rect -246 901 -212 935
rect -246 833 -212 867
rect -246 765 -212 799
rect -246 697 -212 731
rect -246 629 -212 663
rect -246 561 -212 595
rect -246 493 -212 527
rect -246 425 -212 459
rect -246 357 -212 391
rect -246 289 -212 323
rect -246 221 -212 255
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect -246 -255 -212 -221
rect -246 -323 -212 -289
rect -246 -391 -212 -357
rect -246 -459 -212 -425
rect -246 -527 -212 -493
rect -246 -595 -212 -561
rect -246 -663 -212 -629
rect -246 -731 -212 -697
rect -246 -799 -212 -765
rect -246 -867 -212 -833
rect -246 -935 -212 -901
rect -246 -1003 -212 -969
rect -246 -1071 -212 -1037
rect -246 -1139 -212 -1105
rect -246 -1207 -212 -1173
rect -246 -1275 -212 -1241
rect -246 -1343 -212 -1309
rect -246 -1411 -212 -1377
rect -246 -1479 -212 -1445
rect -246 -1547 -212 -1513
rect -246 -1615 -212 -1581
rect -246 -1683 -212 -1649
rect -246 -1751 -212 -1717
rect -246 -1819 -212 -1785
rect -246 -1887 -212 -1853
rect -246 -1955 -212 -1921
rect 212 1921 246 1955
rect 212 1853 246 1887
rect 212 1785 246 1819
rect 212 1717 246 1751
rect 212 1649 246 1683
rect 212 1581 246 1615
rect 212 1513 246 1547
rect 212 1445 246 1479
rect 212 1377 246 1411
rect 212 1309 246 1343
rect 212 1241 246 1275
rect 212 1173 246 1207
rect 212 1105 246 1139
rect 212 1037 246 1071
rect 212 969 246 1003
rect 212 901 246 935
rect 212 833 246 867
rect 212 765 246 799
rect 212 697 246 731
rect 212 629 246 663
rect 212 561 246 595
rect 212 493 246 527
rect 212 425 246 459
rect 212 357 246 391
rect 212 289 246 323
rect 212 221 246 255
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
rect 212 -255 246 -221
rect 212 -323 246 -289
rect 212 -391 246 -357
rect 212 -459 246 -425
rect 212 -527 246 -493
rect 212 -595 246 -561
rect 212 -663 246 -629
rect 212 -731 246 -697
rect 212 -799 246 -765
rect 212 -867 246 -833
rect 212 -935 246 -901
rect 212 -1003 246 -969
rect 212 -1071 246 -1037
rect 212 -1139 246 -1105
rect 212 -1207 246 -1173
rect 212 -1275 246 -1241
rect 212 -1343 246 -1309
rect 212 -1411 246 -1377
rect 212 -1479 246 -1445
rect 212 -1547 246 -1513
rect 212 -1615 246 -1581
rect 212 -1683 246 -1649
rect 212 -1751 246 -1717
rect 212 -1819 246 -1785
rect 212 -1887 246 -1853
rect 212 -1955 246 -1921
<< poly >>
rect -200 2081 200 2097
rect -200 2047 -153 2081
rect -119 2047 -85 2081
rect -51 2047 -17 2081
rect 17 2047 51 2081
rect 85 2047 119 2081
rect 153 2047 200 2081
rect -200 2000 200 2047
rect -200 -2047 200 -2000
rect -200 -2081 -153 -2047
rect -119 -2081 -85 -2047
rect -51 -2081 -17 -2047
rect 17 -2081 51 -2047
rect 85 -2081 119 -2047
rect 153 -2081 200 -2047
rect -200 -2097 200 -2081
<< polycont >>
rect -153 2047 -119 2081
rect -85 2047 -51 2081
rect -17 2047 17 2081
rect 51 2047 85 2081
rect 119 2047 153 2081
rect -153 -2081 -119 -2047
rect -85 -2081 -51 -2047
rect -17 -2081 17 -2047
rect 51 -2081 85 -2047
rect 119 -2081 153 -2047
<< locali >>
rect -200 2047 -161 2081
rect -119 2047 -89 2081
rect -51 2047 -17 2081
rect 17 2047 51 2081
rect 89 2047 119 2081
rect 161 2047 200 2081
rect -246 1961 -212 2004
rect -246 1889 -212 1921
rect -246 1819 -212 1853
rect -246 1751 -212 1783
rect -246 1683 -212 1711
rect -246 1615 -212 1639
rect -246 1547 -212 1567
rect -246 1479 -212 1495
rect -246 1411 -212 1423
rect -246 1343 -212 1351
rect -246 1275 -212 1279
rect -246 1169 -212 1173
rect -246 1097 -212 1105
rect -246 1025 -212 1037
rect -246 953 -212 969
rect -246 881 -212 901
rect -246 809 -212 833
rect -246 737 -212 765
rect -246 665 -212 697
rect -246 595 -212 629
rect -246 527 -212 559
rect -246 459 -212 487
rect -246 391 -212 415
rect -246 323 -212 343
rect -246 255 -212 271
rect -246 187 -212 199
rect -246 119 -212 127
rect -246 51 -212 55
rect -246 -55 -212 -51
rect -246 -127 -212 -119
rect -246 -199 -212 -187
rect -246 -271 -212 -255
rect -246 -343 -212 -323
rect -246 -415 -212 -391
rect -246 -487 -212 -459
rect -246 -559 -212 -527
rect -246 -629 -212 -595
rect -246 -697 -212 -665
rect -246 -765 -212 -737
rect -246 -833 -212 -809
rect -246 -901 -212 -881
rect -246 -969 -212 -953
rect -246 -1037 -212 -1025
rect -246 -1105 -212 -1097
rect -246 -1173 -212 -1169
rect -246 -1279 -212 -1275
rect -246 -1351 -212 -1343
rect -246 -1423 -212 -1411
rect -246 -1495 -212 -1479
rect -246 -1567 -212 -1547
rect -246 -1639 -212 -1615
rect -246 -1711 -212 -1683
rect -246 -1783 -212 -1751
rect -246 -1853 -212 -1819
rect -246 -1921 -212 -1889
rect -246 -2004 -212 -1961
rect 212 1961 246 2004
rect 212 1889 246 1921
rect 212 1819 246 1853
rect 212 1751 246 1783
rect 212 1683 246 1711
rect 212 1615 246 1639
rect 212 1547 246 1567
rect 212 1479 246 1495
rect 212 1411 246 1423
rect 212 1343 246 1351
rect 212 1275 246 1279
rect 212 1169 246 1173
rect 212 1097 246 1105
rect 212 1025 246 1037
rect 212 953 246 969
rect 212 881 246 901
rect 212 809 246 833
rect 212 737 246 765
rect 212 665 246 697
rect 212 595 246 629
rect 212 527 246 559
rect 212 459 246 487
rect 212 391 246 415
rect 212 323 246 343
rect 212 255 246 271
rect 212 187 246 199
rect 212 119 246 127
rect 212 51 246 55
rect 212 -55 246 -51
rect 212 -127 246 -119
rect 212 -199 246 -187
rect 212 -271 246 -255
rect 212 -343 246 -323
rect 212 -415 246 -391
rect 212 -487 246 -459
rect 212 -559 246 -527
rect 212 -629 246 -595
rect 212 -697 246 -665
rect 212 -765 246 -737
rect 212 -833 246 -809
rect 212 -901 246 -881
rect 212 -969 246 -953
rect 212 -1037 246 -1025
rect 212 -1105 246 -1097
rect 212 -1173 246 -1169
rect 212 -1279 246 -1275
rect 212 -1351 246 -1343
rect 212 -1423 246 -1411
rect 212 -1495 246 -1479
rect 212 -1567 246 -1547
rect 212 -1639 246 -1615
rect 212 -1711 246 -1683
rect 212 -1783 246 -1751
rect 212 -1853 246 -1819
rect 212 -1921 246 -1889
rect 212 -2004 246 -1961
rect -200 -2081 -161 -2047
rect -119 -2081 -89 -2047
rect -51 -2081 -17 -2047
rect 17 -2081 51 -2047
rect 89 -2081 119 -2047
rect 161 -2081 200 -2047
<< viali >>
rect -161 2047 -153 2081
rect -153 2047 -127 2081
rect -89 2047 -85 2081
rect -85 2047 -55 2081
rect -17 2047 17 2081
rect 55 2047 85 2081
rect 85 2047 89 2081
rect 127 2047 153 2081
rect 153 2047 161 2081
rect -246 1955 -212 1961
rect -246 1927 -212 1955
rect -246 1887 -212 1889
rect -246 1855 -212 1887
rect -246 1785 -212 1817
rect -246 1783 -212 1785
rect -246 1717 -212 1745
rect -246 1711 -212 1717
rect -246 1649 -212 1673
rect -246 1639 -212 1649
rect -246 1581 -212 1601
rect -246 1567 -212 1581
rect -246 1513 -212 1529
rect -246 1495 -212 1513
rect -246 1445 -212 1457
rect -246 1423 -212 1445
rect -246 1377 -212 1385
rect -246 1351 -212 1377
rect -246 1309 -212 1313
rect -246 1279 -212 1309
rect -246 1207 -212 1241
rect -246 1139 -212 1169
rect -246 1135 -212 1139
rect -246 1071 -212 1097
rect -246 1063 -212 1071
rect -246 1003 -212 1025
rect -246 991 -212 1003
rect -246 935 -212 953
rect -246 919 -212 935
rect -246 867 -212 881
rect -246 847 -212 867
rect -246 799 -212 809
rect -246 775 -212 799
rect -246 731 -212 737
rect -246 703 -212 731
rect -246 663 -212 665
rect -246 631 -212 663
rect -246 561 -212 593
rect -246 559 -212 561
rect -246 493 -212 521
rect -246 487 -212 493
rect -246 425 -212 449
rect -246 415 -212 425
rect -246 357 -212 377
rect -246 343 -212 357
rect -246 289 -212 305
rect -246 271 -212 289
rect -246 221 -212 233
rect -246 199 -212 221
rect -246 153 -212 161
rect -246 127 -212 153
rect -246 85 -212 89
rect -246 55 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -55
rect -246 -89 -212 -85
rect -246 -153 -212 -127
rect -246 -161 -212 -153
rect -246 -221 -212 -199
rect -246 -233 -212 -221
rect -246 -289 -212 -271
rect -246 -305 -212 -289
rect -246 -357 -212 -343
rect -246 -377 -212 -357
rect -246 -425 -212 -415
rect -246 -449 -212 -425
rect -246 -493 -212 -487
rect -246 -521 -212 -493
rect -246 -561 -212 -559
rect -246 -593 -212 -561
rect -246 -663 -212 -631
rect -246 -665 -212 -663
rect -246 -731 -212 -703
rect -246 -737 -212 -731
rect -246 -799 -212 -775
rect -246 -809 -212 -799
rect -246 -867 -212 -847
rect -246 -881 -212 -867
rect -246 -935 -212 -919
rect -246 -953 -212 -935
rect -246 -1003 -212 -991
rect -246 -1025 -212 -1003
rect -246 -1071 -212 -1063
rect -246 -1097 -212 -1071
rect -246 -1139 -212 -1135
rect -246 -1169 -212 -1139
rect -246 -1241 -212 -1207
rect -246 -1309 -212 -1279
rect -246 -1313 -212 -1309
rect -246 -1377 -212 -1351
rect -246 -1385 -212 -1377
rect -246 -1445 -212 -1423
rect -246 -1457 -212 -1445
rect -246 -1513 -212 -1495
rect -246 -1529 -212 -1513
rect -246 -1581 -212 -1567
rect -246 -1601 -212 -1581
rect -246 -1649 -212 -1639
rect -246 -1673 -212 -1649
rect -246 -1717 -212 -1711
rect -246 -1745 -212 -1717
rect -246 -1785 -212 -1783
rect -246 -1817 -212 -1785
rect -246 -1887 -212 -1855
rect -246 -1889 -212 -1887
rect -246 -1955 -212 -1927
rect -246 -1961 -212 -1955
rect 212 1955 246 1961
rect 212 1927 246 1955
rect 212 1887 246 1889
rect 212 1855 246 1887
rect 212 1785 246 1817
rect 212 1783 246 1785
rect 212 1717 246 1745
rect 212 1711 246 1717
rect 212 1649 246 1673
rect 212 1639 246 1649
rect 212 1581 246 1601
rect 212 1567 246 1581
rect 212 1513 246 1529
rect 212 1495 246 1513
rect 212 1445 246 1457
rect 212 1423 246 1445
rect 212 1377 246 1385
rect 212 1351 246 1377
rect 212 1309 246 1313
rect 212 1279 246 1309
rect 212 1207 246 1241
rect 212 1139 246 1169
rect 212 1135 246 1139
rect 212 1071 246 1097
rect 212 1063 246 1071
rect 212 1003 246 1025
rect 212 991 246 1003
rect 212 935 246 953
rect 212 919 246 935
rect 212 867 246 881
rect 212 847 246 867
rect 212 799 246 809
rect 212 775 246 799
rect 212 731 246 737
rect 212 703 246 731
rect 212 663 246 665
rect 212 631 246 663
rect 212 561 246 593
rect 212 559 246 561
rect 212 493 246 521
rect 212 487 246 493
rect 212 425 246 449
rect 212 415 246 425
rect 212 357 246 377
rect 212 343 246 357
rect 212 289 246 305
rect 212 271 246 289
rect 212 221 246 233
rect 212 199 246 221
rect 212 153 246 161
rect 212 127 246 153
rect 212 85 246 89
rect 212 55 246 85
rect 212 -17 246 17
rect 212 -85 246 -55
rect 212 -89 246 -85
rect 212 -153 246 -127
rect 212 -161 246 -153
rect 212 -221 246 -199
rect 212 -233 246 -221
rect 212 -289 246 -271
rect 212 -305 246 -289
rect 212 -357 246 -343
rect 212 -377 246 -357
rect 212 -425 246 -415
rect 212 -449 246 -425
rect 212 -493 246 -487
rect 212 -521 246 -493
rect 212 -561 246 -559
rect 212 -593 246 -561
rect 212 -663 246 -631
rect 212 -665 246 -663
rect 212 -731 246 -703
rect 212 -737 246 -731
rect 212 -799 246 -775
rect 212 -809 246 -799
rect 212 -867 246 -847
rect 212 -881 246 -867
rect 212 -935 246 -919
rect 212 -953 246 -935
rect 212 -1003 246 -991
rect 212 -1025 246 -1003
rect 212 -1071 246 -1063
rect 212 -1097 246 -1071
rect 212 -1139 246 -1135
rect 212 -1169 246 -1139
rect 212 -1241 246 -1207
rect 212 -1309 246 -1279
rect 212 -1313 246 -1309
rect 212 -1377 246 -1351
rect 212 -1385 246 -1377
rect 212 -1445 246 -1423
rect 212 -1457 246 -1445
rect 212 -1513 246 -1495
rect 212 -1529 246 -1513
rect 212 -1581 246 -1567
rect 212 -1601 246 -1581
rect 212 -1649 246 -1639
rect 212 -1673 246 -1649
rect 212 -1717 246 -1711
rect 212 -1745 246 -1717
rect 212 -1785 246 -1783
rect 212 -1817 246 -1785
rect 212 -1887 246 -1855
rect 212 -1889 246 -1887
rect 212 -1955 246 -1927
rect 212 -1961 246 -1955
rect -161 -2081 -153 -2047
rect -153 -2081 -127 -2047
rect -89 -2081 -85 -2047
rect -85 -2081 -55 -2047
rect -17 -2081 17 -2047
rect 55 -2081 85 -2047
rect 85 -2081 89 -2047
rect 127 -2081 153 -2047
rect 153 -2081 161 -2047
<< metal1 >>
rect -196 2081 196 2087
rect -196 2047 -161 2081
rect -127 2047 -89 2081
rect -55 2047 -17 2081
rect 17 2047 55 2081
rect 89 2047 127 2081
rect 161 2047 196 2081
rect -196 2041 196 2047
rect -252 1961 -206 2000
rect -252 1927 -246 1961
rect -212 1927 -206 1961
rect -252 1889 -206 1927
rect -252 1855 -246 1889
rect -212 1855 -206 1889
rect -252 1817 -206 1855
rect -252 1783 -246 1817
rect -212 1783 -206 1817
rect -252 1745 -206 1783
rect -252 1711 -246 1745
rect -212 1711 -206 1745
rect -252 1673 -206 1711
rect -252 1639 -246 1673
rect -212 1639 -206 1673
rect -252 1601 -206 1639
rect -252 1567 -246 1601
rect -212 1567 -206 1601
rect -252 1529 -206 1567
rect -252 1495 -246 1529
rect -212 1495 -206 1529
rect -252 1457 -206 1495
rect -252 1423 -246 1457
rect -212 1423 -206 1457
rect -252 1385 -206 1423
rect -252 1351 -246 1385
rect -212 1351 -206 1385
rect -252 1313 -206 1351
rect -252 1279 -246 1313
rect -212 1279 -206 1313
rect -252 1241 -206 1279
rect -252 1207 -246 1241
rect -212 1207 -206 1241
rect -252 1169 -206 1207
rect -252 1135 -246 1169
rect -212 1135 -206 1169
rect -252 1097 -206 1135
rect -252 1063 -246 1097
rect -212 1063 -206 1097
rect -252 1025 -206 1063
rect -252 991 -246 1025
rect -212 991 -206 1025
rect -252 953 -206 991
rect -252 919 -246 953
rect -212 919 -206 953
rect -252 881 -206 919
rect -252 847 -246 881
rect -212 847 -206 881
rect -252 809 -206 847
rect -252 775 -246 809
rect -212 775 -206 809
rect -252 737 -206 775
rect -252 703 -246 737
rect -212 703 -206 737
rect -252 665 -206 703
rect -252 631 -246 665
rect -212 631 -206 665
rect -252 593 -206 631
rect -252 559 -246 593
rect -212 559 -206 593
rect -252 521 -206 559
rect -252 487 -246 521
rect -212 487 -206 521
rect -252 449 -206 487
rect -252 415 -246 449
rect -212 415 -206 449
rect -252 377 -206 415
rect -252 343 -246 377
rect -212 343 -206 377
rect -252 305 -206 343
rect -252 271 -246 305
rect -212 271 -206 305
rect -252 233 -206 271
rect -252 199 -246 233
rect -212 199 -206 233
rect -252 161 -206 199
rect -252 127 -246 161
rect -212 127 -206 161
rect -252 89 -206 127
rect -252 55 -246 89
rect -212 55 -206 89
rect -252 17 -206 55
rect -252 -17 -246 17
rect -212 -17 -206 17
rect -252 -55 -206 -17
rect -252 -89 -246 -55
rect -212 -89 -206 -55
rect -252 -127 -206 -89
rect -252 -161 -246 -127
rect -212 -161 -206 -127
rect -252 -199 -206 -161
rect -252 -233 -246 -199
rect -212 -233 -206 -199
rect -252 -271 -206 -233
rect -252 -305 -246 -271
rect -212 -305 -206 -271
rect -252 -343 -206 -305
rect -252 -377 -246 -343
rect -212 -377 -206 -343
rect -252 -415 -206 -377
rect -252 -449 -246 -415
rect -212 -449 -206 -415
rect -252 -487 -206 -449
rect -252 -521 -246 -487
rect -212 -521 -206 -487
rect -252 -559 -206 -521
rect -252 -593 -246 -559
rect -212 -593 -206 -559
rect -252 -631 -206 -593
rect -252 -665 -246 -631
rect -212 -665 -206 -631
rect -252 -703 -206 -665
rect -252 -737 -246 -703
rect -212 -737 -206 -703
rect -252 -775 -206 -737
rect -252 -809 -246 -775
rect -212 -809 -206 -775
rect -252 -847 -206 -809
rect -252 -881 -246 -847
rect -212 -881 -206 -847
rect -252 -919 -206 -881
rect -252 -953 -246 -919
rect -212 -953 -206 -919
rect -252 -991 -206 -953
rect -252 -1025 -246 -991
rect -212 -1025 -206 -991
rect -252 -1063 -206 -1025
rect -252 -1097 -246 -1063
rect -212 -1097 -206 -1063
rect -252 -1135 -206 -1097
rect -252 -1169 -246 -1135
rect -212 -1169 -206 -1135
rect -252 -1207 -206 -1169
rect -252 -1241 -246 -1207
rect -212 -1241 -206 -1207
rect -252 -1279 -206 -1241
rect -252 -1313 -246 -1279
rect -212 -1313 -206 -1279
rect -252 -1351 -206 -1313
rect -252 -1385 -246 -1351
rect -212 -1385 -206 -1351
rect -252 -1423 -206 -1385
rect -252 -1457 -246 -1423
rect -212 -1457 -206 -1423
rect -252 -1495 -206 -1457
rect -252 -1529 -246 -1495
rect -212 -1529 -206 -1495
rect -252 -1567 -206 -1529
rect -252 -1601 -246 -1567
rect -212 -1601 -206 -1567
rect -252 -1639 -206 -1601
rect -252 -1673 -246 -1639
rect -212 -1673 -206 -1639
rect -252 -1711 -206 -1673
rect -252 -1745 -246 -1711
rect -212 -1745 -206 -1711
rect -252 -1783 -206 -1745
rect -252 -1817 -246 -1783
rect -212 -1817 -206 -1783
rect -252 -1855 -206 -1817
rect -252 -1889 -246 -1855
rect -212 -1889 -206 -1855
rect -252 -1927 -206 -1889
rect -252 -1961 -246 -1927
rect -212 -1961 -206 -1927
rect -252 -2000 -206 -1961
rect 206 1961 252 2000
rect 206 1927 212 1961
rect 246 1927 252 1961
rect 206 1889 252 1927
rect 206 1855 212 1889
rect 246 1855 252 1889
rect 206 1817 252 1855
rect 206 1783 212 1817
rect 246 1783 252 1817
rect 206 1745 252 1783
rect 206 1711 212 1745
rect 246 1711 252 1745
rect 206 1673 252 1711
rect 206 1639 212 1673
rect 246 1639 252 1673
rect 206 1601 252 1639
rect 206 1567 212 1601
rect 246 1567 252 1601
rect 206 1529 252 1567
rect 206 1495 212 1529
rect 246 1495 252 1529
rect 206 1457 252 1495
rect 206 1423 212 1457
rect 246 1423 252 1457
rect 206 1385 252 1423
rect 206 1351 212 1385
rect 246 1351 252 1385
rect 206 1313 252 1351
rect 206 1279 212 1313
rect 246 1279 252 1313
rect 206 1241 252 1279
rect 206 1207 212 1241
rect 246 1207 252 1241
rect 206 1169 252 1207
rect 206 1135 212 1169
rect 246 1135 252 1169
rect 206 1097 252 1135
rect 206 1063 212 1097
rect 246 1063 252 1097
rect 206 1025 252 1063
rect 206 991 212 1025
rect 246 991 252 1025
rect 206 953 252 991
rect 206 919 212 953
rect 246 919 252 953
rect 206 881 252 919
rect 206 847 212 881
rect 246 847 252 881
rect 206 809 252 847
rect 206 775 212 809
rect 246 775 252 809
rect 206 737 252 775
rect 206 703 212 737
rect 246 703 252 737
rect 206 665 252 703
rect 206 631 212 665
rect 246 631 252 665
rect 206 593 252 631
rect 206 559 212 593
rect 246 559 252 593
rect 206 521 252 559
rect 206 487 212 521
rect 246 487 252 521
rect 206 449 252 487
rect 206 415 212 449
rect 246 415 252 449
rect 206 377 252 415
rect 206 343 212 377
rect 246 343 252 377
rect 206 305 252 343
rect 206 271 212 305
rect 246 271 252 305
rect 206 233 252 271
rect 206 199 212 233
rect 246 199 252 233
rect 206 161 252 199
rect 206 127 212 161
rect 246 127 252 161
rect 206 89 252 127
rect 206 55 212 89
rect 246 55 252 89
rect 206 17 252 55
rect 206 -17 212 17
rect 246 -17 252 17
rect 206 -55 252 -17
rect 206 -89 212 -55
rect 246 -89 252 -55
rect 206 -127 252 -89
rect 206 -161 212 -127
rect 246 -161 252 -127
rect 206 -199 252 -161
rect 206 -233 212 -199
rect 246 -233 252 -199
rect 206 -271 252 -233
rect 206 -305 212 -271
rect 246 -305 252 -271
rect 206 -343 252 -305
rect 206 -377 212 -343
rect 246 -377 252 -343
rect 206 -415 252 -377
rect 206 -449 212 -415
rect 246 -449 252 -415
rect 206 -487 252 -449
rect 206 -521 212 -487
rect 246 -521 252 -487
rect 206 -559 252 -521
rect 206 -593 212 -559
rect 246 -593 252 -559
rect 206 -631 252 -593
rect 206 -665 212 -631
rect 246 -665 252 -631
rect 206 -703 252 -665
rect 206 -737 212 -703
rect 246 -737 252 -703
rect 206 -775 252 -737
rect 206 -809 212 -775
rect 246 -809 252 -775
rect 206 -847 252 -809
rect 206 -881 212 -847
rect 246 -881 252 -847
rect 206 -919 252 -881
rect 206 -953 212 -919
rect 246 -953 252 -919
rect 206 -991 252 -953
rect 206 -1025 212 -991
rect 246 -1025 252 -991
rect 206 -1063 252 -1025
rect 206 -1097 212 -1063
rect 246 -1097 252 -1063
rect 206 -1135 252 -1097
rect 206 -1169 212 -1135
rect 246 -1169 252 -1135
rect 206 -1207 252 -1169
rect 206 -1241 212 -1207
rect 246 -1241 252 -1207
rect 206 -1279 252 -1241
rect 206 -1313 212 -1279
rect 246 -1313 252 -1279
rect 206 -1351 252 -1313
rect 206 -1385 212 -1351
rect 246 -1385 252 -1351
rect 206 -1423 252 -1385
rect 206 -1457 212 -1423
rect 246 -1457 252 -1423
rect 206 -1495 252 -1457
rect 206 -1529 212 -1495
rect 246 -1529 252 -1495
rect 206 -1567 252 -1529
rect 206 -1601 212 -1567
rect 246 -1601 252 -1567
rect 206 -1639 252 -1601
rect 206 -1673 212 -1639
rect 246 -1673 252 -1639
rect 206 -1711 252 -1673
rect 206 -1745 212 -1711
rect 246 -1745 252 -1711
rect 206 -1783 252 -1745
rect 206 -1817 212 -1783
rect 246 -1817 252 -1783
rect 206 -1855 252 -1817
rect 206 -1889 212 -1855
rect 246 -1889 252 -1855
rect 206 -1927 252 -1889
rect 206 -1961 212 -1927
rect 246 -1961 252 -1927
rect 206 -2000 252 -1961
rect -196 -2047 196 -2041
rect -196 -2081 -161 -2047
rect -127 -2081 -89 -2047
rect -55 -2081 -17 -2047
rect 17 -2081 55 -2047
rect 89 -2081 127 -2047
rect 161 -2081 196 -2047
rect -196 -2087 196 -2081
<< end >>
