magic
tech sky130A
magscale 1 2
timestamp 1666407696
<< poly >>
rect 137 2693 437 2738
rect 377 2655 437 2693
<< locali >>
rect 230 3850 264 4003
rect 466 3850 500 4003
rect 702 3853 736 4006
rect 348 2921 382 3073
rect 348 2887 483 2921
rect 449 2641 483 2887
rect 642 2686 678 2972
rect -56 2599 126 2638
rect 449 2607 618 2641
rect 92 2520 126 2599
rect 331 1412 365 1637
rect 331 1378 694 1412
rect 210 1185 244 1281
rect 210 1146 1112 1185
rect -27 1078 201 1112
<< metal1 >>
rect 348 2921 382 3073
rect 348 2887 483 2921
rect 449 2641 483 2887
rect 642 2686 678 2972
rect -56 2599 126 2638
rect 449 2607 618 2641
rect 92 2520 126 2599
rect 331 1412 365 1637
rect 331 1378 694 1412
rect 210 1185 244 1281
rect 210 1146 1112 1185
rect -27 1078 201 1112
use sky130_fd_pr__cap_mim_m3_1_C9NYDN  XC1
timestamp 1666402782
transform 1 0 16043 0 1 1188
box -1150 -800 1149 800
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  XC2
timestamp 1666402782
transform 1 0 12744 0 1 2488
box -2150 -2100 2149 2100
use sky130_fd_pr__cap_mim_m3_1_MWYMHE  XC3
timestamp 1666402782
transform 1 0 7945 0 1 2488
box -2650 -2100 2649 2100
use sky130_fd_pr__cap_mim_m3_1_BTMG45  XC4
timestamp 1666402782
transform 1 0 3446 0 1 988
box -1850 -600 1849 600
use sky130_fd_pr__nfet_01v8_K6VZSH  XM1
timestamp 1666407406
transform 1 0 407 0 1 2078
box -88 -596 88 596
use sky130_fd_pr__nfet_01v8_Z3HWK5  XM2
timestamp 1666407491
transform 1 0 660 0 1 2050
box -88 -688 88 688
use sky130_fd_pr__pfet_01v8_BRZSWZ  XM6
timestamp 1666404115
transform 1 0 424 0 1 3414
box -360 -494 360 556
use sky130_fd_pr__nfet_01v8_9ZFLEJ  XM8
timestamp 1666406900
transform 1 0 168 0 1 1900
box -88 -838 88 838
<< end >>
