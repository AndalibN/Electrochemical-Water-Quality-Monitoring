magic
tech sky130A
magscale 1 2
timestamp 1666829797
<< error_p >>
rect -740 1127 -682 1133
rect -582 1127 -524 1133
rect -424 1127 -366 1133
rect -266 1127 -208 1133
rect -108 1127 -50 1133
rect 50 1127 108 1133
rect 208 1127 266 1133
rect 366 1127 424 1133
rect 524 1127 582 1133
rect 682 1127 740 1133
rect -740 1093 -728 1127
rect -582 1093 -570 1127
rect -424 1093 -412 1127
rect -266 1093 -254 1127
rect -108 1093 -96 1127
rect 50 1093 62 1127
rect 208 1093 220 1127
rect 366 1093 378 1127
rect 524 1093 536 1127
rect 682 1093 694 1127
rect -740 1087 -682 1093
rect -582 1087 -524 1093
rect -424 1087 -366 1093
rect -266 1087 -208 1093
rect -108 1087 -50 1093
rect 50 1087 108 1093
rect 208 1087 266 1093
rect 366 1087 424 1093
rect 524 1087 582 1093
rect 682 1087 740 1093
rect -740 17 -682 23
rect -582 17 -524 23
rect -424 17 -366 23
rect -266 17 -208 23
rect -108 17 -50 23
rect 50 17 108 23
rect 208 17 266 23
rect 366 17 424 23
rect 524 17 582 23
rect 682 17 740 23
rect -740 -17 -728 17
rect -582 -17 -570 17
rect -424 -17 -412 17
rect -266 -17 -254 17
rect -108 -17 -96 17
rect 50 -17 62 17
rect 208 -17 220 17
rect 366 -17 378 17
rect 524 -17 536 17
rect 682 -17 694 17
rect -740 -23 -682 -17
rect -582 -23 -524 -17
rect -424 -23 -366 -17
rect -266 -23 -208 -17
rect -108 -23 -50 -17
rect 50 -23 108 -17
rect 208 -23 266 -17
rect 366 -23 424 -17
rect 524 -23 582 -17
rect 682 -23 740 -17
rect -740 -1093 -682 -1087
rect -582 -1093 -524 -1087
rect -424 -1093 -366 -1087
rect -266 -1093 -208 -1087
rect -108 -1093 -50 -1087
rect 50 -1093 108 -1087
rect 208 -1093 266 -1087
rect 366 -1093 424 -1087
rect 524 -1093 582 -1087
rect 682 -1093 740 -1087
rect -740 -1127 -728 -1093
rect -582 -1127 -570 -1093
rect -424 -1127 -412 -1093
rect -266 -1127 -254 -1093
rect -108 -1127 -96 -1093
rect 50 -1127 62 -1093
rect 208 -1127 220 -1093
rect 366 -1127 378 -1093
rect 524 -1127 536 -1093
rect 682 -1127 694 -1093
rect -740 -1133 -682 -1127
rect -582 -1133 -524 -1127
rect -424 -1133 -366 -1127
rect -266 -1133 -208 -1127
rect -108 -1133 -50 -1127
rect 50 -1133 108 -1127
rect 208 -1133 266 -1127
rect 366 -1133 424 -1127
rect 524 -1133 582 -1127
rect 682 -1133 740 -1127
<< nmos >>
rect -761 55 -661 1055
rect -603 55 -503 1055
rect -445 55 -345 1055
rect -287 55 -187 1055
rect -129 55 -29 1055
rect 29 55 129 1055
rect 187 55 287 1055
rect 345 55 445 1055
rect 503 55 603 1055
rect 661 55 761 1055
rect -761 -1055 -661 -55
rect -603 -1055 -503 -55
rect -445 -1055 -345 -55
rect -287 -1055 -187 -55
rect -129 -1055 -29 -55
rect 29 -1055 129 -55
rect 187 -1055 287 -55
rect 345 -1055 445 -55
rect 503 -1055 603 -55
rect 661 -1055 761 -55
<< ndiff >>
rect -819 1043 -761 1055
rect -819 67 -807 1043
rect -773 67 -761 1043
rect -819 55 -761 67
rect -661 1043 -603 1055
rect -661 67 -649 1043
rect -615 67 -603 1043
rect -661 55 -603 67
rect -503 1043 -445 1055
rect -503 67 -491 1043
rect -457 67 -445 1043
rect -503 55 -445 67
rect -345 1043 -287 1055
rect -345 67 -333 1043
rect -299 67 -287 1043
rect -345 55 -287 67
rect -187 1043 -129 1055
rect -187 67 -175 1043
rect -141 67 -129 1043
rect -187 55 -129 67
rect -29 1043 29 1055
rect -29 67 -17 1043
rect 17 67 29 1043
rect -29 55 29 67
rect 129 1043 187 1055
rect 129 67 141 1043
rect 175 67 187 1043
rect 129 55 187 67
rect 287 1043 345 1055
rect 287 67 299 1043
rect 333 67 345 1043
rect 287 55 345 67
rect 445 1043 503 1055
rect 445 67 457 1043
rect 491 67 503 1043
rect 445 55 503 67
rect 603 1043 661 1055
rect 603 67 615 1043
rect 649 67 661 1043
rect 603 55 661 67
rect 761 1043 819 1055
rect 761 67 773 1043
rect 807 67 819 1043
rect 761 55 819 67
rect -819 -67 -761 -55
rect -819 -1043 -807 -67
rect -773 -1043 -761 -67
rect -819 -1055 -761 -1043
rect -661 -67 -603 -55
rect -661 -1043 -649 -67
rect -615 -1043 -603 -67
rect -661 -1055 -603 -1043
rect -503 -67 -445 -55
rect -503 -1043 -491 -67
rect -457 -1043 -445 -67
rect -503 -1055 -445 -1043
rect -345 -67 -287 -55
rect -345 -1043 -333 -67
rect -299 -1043 -287 -67
rect -345 -1055 -287 -1043
rect -187 -67 -129 -55
rect -187 -1043 -175 -67
rect -141 -1043 -129 -67
rect -187 -1055 -129 -1043
rect -29 -67 29 -55
rect -29 -1043 -17 -67
rect 17 -1043 29 -67
rect -29 -1055 29 -1043
rect 129 -67 187 -55
rect 129 -1043 141 -67
rect 175 -1043 187 -67
rect 129 -1055 187 -1043
rect 287 -67 345 -55
rect 287 -1043 299 -67
rect 333 -1043 345 -67
rect 287 -1055 345 -1043
rect 445 -67 503 -55
rect 445 -1043 457 -67
rect 491 -1043 503 -67
rect 445 -1055 503 -1043
rect 603 -67 661 -55
rect 603 -1043 615 -67
rect 649 -1043 661 -67
rect 603 -1055 661 -1043
rect 761 -67 819 -55
rect 761 -1043 773 -67
rect 807 -1043 819 -67
rect 761 -1055 819 -1043
<< ndiffc >>
rect -807 67 -773 1043
rect -649 67 -615 1043
rect -491 67 -457 1043
rect -333 67 -299 1043
rect -175 67 -141 1043
rect -17 67 17 1043
rect 141 67 175 1043
rect 299 67 333 1043
rect 457 67 491 1043
rect 615 67 649 1043
rect 773 67 807 1043
rect -807 -1043 -773 -67
rect -649 -1043 -615 -67
rect -491 -1043 -457 -67
rect -333 -1043 -299 -67
rect -175 -1043 -141 -67
rect -17 -1043 17 -67
rect 141 -1043 175 -67
rect 299 -1043 333 -67
rect 457 -1043 491 -67
rect 615 -1043 649 -67
rect 773 -1043 807 -67
<< poly >>
rect -761 1127 -661 1143
rect -761 1093 -745 1127
rect -677 1093 -661 1127
rect -761 1055 -661 1093
rect -603 1127 -503 1143
rect -603 1093 -587 1127
rect -519 1093 -503 1127
rect -603 1055 -503 1093
rect -445 1127 -345 1143
rect -445 1093 -429 1127
rect -361 1093 -345 1127
rect -445 1055 -345 1093
rect -287 1127 -187 1143
rect -287 1093 -271 1127
rect -203 1093 -187 1127
rect -287 1055 -187 1093
rect -129 1127 -29 1143
rect -129 1093 -113 1127
rect -45 1093 -29 1127
rect -129 1055 -29 1093
rect 29 1127 129 1143
rect 29 1093 45 1127
rect 113 1093 129 1127
rect 29 1055 129 1093
rect 187 1127 287 1143
rect 187 1093 203 1127
rect 271 1093 287 1127
rect 187 1055 287 1093
rect 345 1127 445 1143
rect 345 1093 361 1127
rect 429 1093 445 1127
rect 345 1055 445 1093
rect 503 1127 603 1143
rect 503 1093 519 1127
rect 587 1093 603 1127
rect 503 1055 603 1093
rect 661 1127 761 1143
rect 661 1093 677 1127
rect 745 1093 761 1127
rect 661 1055 761 1093
rect -761 17 -661 55
rect -761 -17 -745 17
rect -677 -17 -661 17
rect -761 -55 -661 -17
rect -603 17 -503 55
rect -603 -17 -587 17
rect -519 -17 -503 17
rect -603 -55 -503 -17
rect -445 17 -345 55
rect -445 -17 -429 17
rect -361 -17 -345 17
rect -445 -55 -345 -17
rect -287 17 -187 55
rect -287 -17 -271 17
rect -203 -17 -187 17
rect -287 -55 -187 -17
rect -129 17 -29 55
rect -129 -17 -113 17
rect -45 -17 -29 17
rect -129 -55 -29 -17
rect 29 17 129 55
rect 29 -17 45 17
rect 113 -17 129 17
rect 29 -55 129 -17
rect 187 17 287 55
rect 187 -17 203 17
rect 271 -17 287 17
rect 187 -55 287 -17
rect 345 17 445 55
rect 345 -17 361 17
rect 429 -17 445 17
rect 345 -55 445 -17
rect 503 17 603 55
rect 503 -17 519 17
rect 587 -17 603 17
rect 503 -55 603 -17
rect 661 17 761 55
rect 661 -17 677 17
rect 745 -17 761 17
rect 661 -55 761 -17
rect -761 -1093 -661 -1055
rect -761 -1127 -745 -1093
rect -677 -1127 -661 -1093
rect -761 -1143 -661 -1127
rect -603 -1093 -503 -1055
rect -603 -1127 -587 -1093
rect -519 -1127 -503 -1093
rect -603 -1143 -503 -1127
rect -445 -1093 -345 -1055
rect -445 -1127 -429 -1093
rect -361 -1127 -345 -1093
rect -445 -1143 -345 -1127
rect -287 -1093 -187 -1055
rect -287 -1127 -271 -1093
rect -203 -1127 -187 -1093
rect -287 -1143 -187 -1127
rect -129 -1093 -29 -1055
rect -129 -1127 -113 -1093
rect -45 -1127 -29 -1093
rect -129 -1143 -29 -1127
rect 29 -1093 129 -1055
rect 29 -1127 45 -1093
rect 113 -1127 129 -1093
rect 29 -1143 129 -1127
rect 187 -1093 287 -1055
rect 187 -1127 203 -1093
rect 271 -1127 287 -1093
rect 187 -1143 287 -1127
rect 345 -1093 445 -1055
rect 345 -1127 361 -1093
rect 429 -1127 445 -1093
rect 345 -1143 445 -1127
rect 503 -1093 603 -1055
rect 503 -1127 519 -1093
rect 587 -1127 603 -1093
rect 503 -1143 603 -1127
rect 661 -1093 761 -1055
rect 661 -1127 677 -1093
rect 745 -1127 761 -1093
rect 661 -1143 761 -1127
<< polycont >>
rect -745 1093 -677 1127
rect -587 1093 -519 1127
rect -429 1093 -361 1127
rect -271 1093 -203 1127
rect -113 1093 -45 1127
rect 45 1093 113 1127
rect 203 1093 271 1127
rect 361 1093 429 1127
rect 519 1093 587 1127
rect 677 1093 745 1127
rect -745 -17 -677 17
rect -587 -17 -519 17
rect -429 -17 -361 17
rect -271 -17 -203 17
rect -113 -17 -45 17
rect 45 -17 113 17
rect 203 -17 271 17
rect 361 -17 429 17
rect 519 -17 587 17
rect 677 -17 745 17
rect -745 -1127 -677 -1093
rect -587 -1127 -519 -1093
rect -429 -1127 -361 -1093
rect -271 -1127 -203 -1093
rect -113 -1127 -45 -1093
rect 45 -1127 113 -1093
rect 203 -1127 271 -1093
rect 361 -1127 429 -1093
rect 519 -1127 587 -1093
rect 677 -1127 745 -1093
<< locali >>
rect -761 1093 -745 1127
rect -677 1093 -661 1127
rect -603 1093 -587 1127
rect -519 1093 -503 1127
rect -445 1093 -429 1127
rect -361 1093 -345 1127
rect -287 1093 -271 1127
rect -203 1093 -187 1127
rect -129 1093 -113 1127
rect -45 1093 -29 1127
rect 29 1093 45 1127
rect 113 1093 129 1127
rect 187 1093 203 1127
rect 271 1093 287 1127
rect 345 1093 361 1127
rect 429 1093 445 1127
rect 503 1093 519 1127
rect 587 1093 603 1127
rect 661 1093 677 1127
rect 745 1093 761 1127
rect -807 1043 -773 1059
rect -807 51 -773 67
rect -649 1043 -615 1059
rect -649 51 -615 67
rect -491 1043 -457 1059
rect -491 51 -457 67
rect -333 1043 -299 1059
rect -333 51 -299 67
rect -175 1043 -141 1059
rect -175 51 -141 67
rect -17 1043 17 1059
rect -17 51 17 67
rect 141 1043 175 1059
rect 141 51 175 67
rect 299 1043 333 1059
rect 299 51 333 67
rect 457 1043 491 1059
rect 457 51 491 67
rect 615 1043 649 1059
rect 615 51 649 67
rect 773 1043 807 1059
rect 773 51 807 67
rect -761 -17 -745 17
rect -677 -17 -661 17
rect -603 -17 -587 17
rect -519 -17 -503 17
rect -445 -17 -429 17
rect -361 -17 -345 17
rect -287 -17 -271 17
rect -203 -17 -187 17
rect -129 -17 -113 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 113 -17 129 17
rect 187 -17 203 17
rect 271 -17 287 17
rect 345 -17 361 17
rect 429 -17 445 17
rect 503 -17 519 17
rect 587 -17 603 17
rect 661 -17 677 17
rect 745 -17 761 17
rect -807 -67 -773 -51
rect -807 -1059 -773 -1043
rect -649 -67 -615 -51
rect -649 -1059 -615 -1043
rect -491 -67 -457 -51
rect -491 -1059 -457 -1043
rect -333 -67 -299 -51
rect -333 -1059 -299 -1043
rect -175 -67 -141 -51
rect -175 -1059 -141 -1043
rect -17 -67 17 -51
rect -17 -1059 17 -1043
rect 141 -67 175 -51
rect 141 -1059 175 -1043
rect 299 -67 333 -51
rect 299 -1059 333 -1043
rect 457 -67 491 -51
rect 457 -1059 491 -1043
rect 615 -67 649 -51
rect 615 -1059 649 -1043
rect 773 -67 807 -51
rect 773 -1059 807 -1043
rect -761 -1127 -745 -1093
rect -677 -1127 -661 -1093
rect -603 -1127 -587 -1093
rect -519 -1127 -503 -1093
rect -445 -1127 -429 -1093
rect -361 -1127 -345 -1093
rect -287 -1127 -271 -1093
rect -203 -1127 -187 -1093
rect -129 -1127 -113 -1093
rect -45 -1127 -29 -1093
rect 29 -1127 45 -1093
rect 113 -1127 129 -1093
rect 187 -1127 203 -1093
rect 271 -1127 287 -1093
rect 345 -1127 361 -1093
rect 429 -1127 445 -1093
rect 503 -1127 519 -1093
rect 587 -1127 603 -1093
rect 661 -1127 677 -1093
rect 745 -1127 761 -1093
<< viali >>
rect -728 1093 -694 1127
rect -570 1093 -536 1127
rect -412 1093 -378 1127
rect -254 1093 -220 1127
rect -96 1093 -62 1127
rect 62 1093 96 1127
rect 220 1093 254 1127
rect 378 1093 412 1127
rect 536 1093 570 1127
rect 694 1093 728 1127
rect -807 67 -773 1043
rect -649 67 -615 1043
rect -491 67 -457 1043
rect -333 67 -299 1043
rect -175 67 -141 1043
rect -17 67 17 1043
rect 141 67 175 1043
rect 299 67 333 1043
rect 457 67 491 1043
rect 615 67 649 1043
rect 773 67 807 1043
rect -728 -17 -694 17
rect -570 -17 -536 17
rect -412 -17 -378 17
rect -254 -17 -220 17
rect -96 -17 -62 17
rect 62 -17 96 17
rect 220 -17 254 17
rect 378 -17 412 17
rect 536 -17 570 17
rect 694 -17 728 17
rect -807 -1043 -773 -67
rect -649 -1043 -615 -67
rect -491 -1043 -457 -67
rect -333 -1043 -299 -67
rect -175 -1043 -141 -67
rect -17 -1043 17 -67
rect 141 -1043 175 -67
rect 299 -1043 333 -67
rect 457 -1043 491 -67
rect 615 -1043 649 -67
rect 773 -1043 807 -67
rect -728 -1127 -694 -1093
rect -570 -1127 -536 -1093
rect -412 -1127 -378 -1093
rect -254 -1127 -220 -1093
rect -96 -1127 -62 -1093
rect 62 -1127 96 -1093
rect 220 -1127 254 -1093
rect 378 -1127 412 -1093
rect 536 -1127 570 -1093
rect 694 -1127 728 -1093
<< metal1 >>
rect -740 1127 -682 1133
rect -740 1093 -728 1127
rect -694 1093 -682 1127
rect -740 1087 -682 1093
rect -582 1127 -524 1133
rect -582 1093 -570 1127
rect -536 1093 -524 1127
rect -582 1087 -524 1093
rect -424 1127 -366 1133
rect -424 1093 -412 1127
rect -378 1093 -366 1127
rect -424 1087 -366 1093
rect -266 1127 -208 1133
rect -266 1093 -254 1127
rect -220 1093 -208 1127
rect -266 1087 -208 1093
rect -108 1127 -50 1133
rect -108 1093 -96 1127
rect -62 1093 -50 1127
rect -108 1087 -50 1093
rect 50 1127 108 1133
rect 50 1093 62 1127
rect 96 1093 108 1127
rect 50 1087 108 1093
rect 208 1127 266 1133
rect 208 1093 220 1127
rect 254 1093 266 1127
rect 208 1087 266 1093
rect 366 1127 424 1133
rect 366 1093 378 1127
rect 412 1093 424 1127
rect 366 1087 424 1093
rect 524 1127 582 1133
rect 524 1093 536 1127
rect 570 1093 582 1127
rect 524 1087 582 1093
rect 682 1127 740 1133
rect 682 1093 694 1127
rect 728 1093 740 1127
rect 682 1087 740 1093
rect -813 1043 -767 1055
rect -813 67 -807 1043
rect -773 67 -767 1043
rect -813 55 -767 67
rect -655 1043 -609 1055
rect -655 67 -649 1043
rect -615 67 -609 1043
rect -655 55 -609 67
rect -497 1043 -451 1055
rect -497 67 -491 1043
rect -457 67 -451 1043
rect -497 55 -451 67
rect -339 1043 -293 1055
rect -339 67 -333 1043
rect -299 67 -293 1043
rect -339 55 -293 67
rect -181 1043 -135 1055
rect -181 67 -175 1043
rect -141 67 -135 1043
rect -181 55 -135 67
rect -23 1043 23 1055
rect -23 67 -17 1043
rect 17 67 23 1043
rect -23 55 23 67
rect 135 1043 181 1055
rect 135 67 141 1043
rect 175 67 181 1043
rect 135 55 181 67
rect 293 1043 339 1055
rect 293 67 299 1043
rect 333 67 339 1043
rect 293 55 339 67
rect 451 1043 497 1055
rect 451 67 457 1043
rect 491 67 497 1043
rect 451 55 497 67
rect 609 1043 655 1055
rect 609 67 615 1043
rect 649 67 655 1043
rect 609 55 655 67
rect 767 1043 813 1055
rect 767 67 773 1043
rect 807 67 813 1043
rect 767 55 813 67
rect -740 17 -682 23
rect -740 -17 -728 17
rect -694 -17 -682 17
rect -740 -23 -682 -17
rect -582 17 -524 23
rect -582 -17 -570 17
rect -536 -17 -524 17
rect -582 -23 -524 -17
rect -424 17 -366 23
rect -424 -17 -412 17
rect -378 -17 -366 17
rect -424 -23 -366 -17
rect -266 17 -208 23
rect -266 -17 -254 17
rect -220 -17 -208 17
rect -266 -23 -208 -17
rect -108 17 -50 23
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -23 -50 -17
rect 50 17 108 23
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -23 108 -17
rect 208 17 266 23
rect 208 -17 220 17
rect 254 -17 266 17
rect 208 -23 266 -17
rect 366 17 424 23
rect 366 -17 378 17
rect 412 -17 424 17
rect 366 -23 424 -17
rect 524 17 582 23
rect 524 -17 536 17
rect 570 -17 582 17
rect 524 -23 582 -17
rect 682 17 740 23
rect 682 -17 694 17
rect 728 -17 740 17
rect 682 -23 740 -17
rect -813 -67 -767 -55
rect -813 -1043 -807 -67
rect -773 -1043 -767 -67
rect -813 -1055 -767 -1043
rect -655 -67 -609 -55
rect -655 -1043 -649 -67
rect -615 -1043 -609 -67
rect -655 -1055 -609 -1043
rect -497 -67 -451 -55
rect -497 -1043 -491 -67
rect -457 -1043 -451 -67
rect -497 -1055 -451 -1043
rect -339 -67 -293 -55
rect -339 -1043 -333 -67
rect -299 -1043 -293 -67
rect -339 -1055 -293 -1043
rect -181 -67 -135 -55
rect -181 -1043 -175 -67
rect -141 -1043 -135 -67
rect -181 -1055 -135 -1043
rect -23 -67 23 -55
rect -23 -1043 -17 -67
rect 17 -1043 23 -67
rect -23 -1055 23 -1043
rect 135 -67 181 -55
rect 135 -1043 141 -67
rect 175 -1043 181 -67
rect 135 -1055 181 -1043
rect 293 -67 339 -55
rect 293 -1043 299 -67
rect 333 -1043 339 -67
rect 293 -1055 339 -1043
rect 451 -67 497 -55
rect 451 -1043 457 -67
rect 491 -1043 497 -67
rect 451 -1055 497 -1043
rect 609 -67 655 -55
rect 609 -1043 615 -67
rect 649 -1043 655 -67
rect 609 -1055 655 -1043
rect 767 -67 813 -55
rect 767 -1043 773 -67
rect 807 -1043 813 -67
rect 767 -1055 813 -1043
rect -740 -1093 -682 -1087
rect -740 -1127 -728 -1093
rect -694 -1127 -682 -1093
rect -740 -1133 -682 -1127
rect -582 -1093 -524 -1087
rect -582 -1127 -570 -1093
rect -536 -1127 -524 -1093
rect -582 -1133 -524 -1127
rect -424 -1093 -366 -1087
rect -424 -1127 -412 -1093
rect -378 -1127 -366 -1093
rect -424 -1133 -366 -1127
rect -266 -1093 -208 -1087
rect -266 -1127 -254 -1093
rect -220 -1127 -208 -1093
rect -266 -1133 -208 -1127
rect -108 -1093 -50 -1087
rect -108 -1127 -96 -1093
rect -62 -1127 -50 -1093
rect -108 -1133 -50 -1127
rect 50 -1093 108 -1087
rect 50 -1127 62 -1093
rect 96 -1127 108 -1093
rect 50 -1133 108 -1127
rect 208 -1093 266 -1087
rect 208 -1127 220 -1093
rect 254 -1127 266 -1093
rect 208 -1133 266 -1127
rect 366 -1093 424 -1087
rect 366 -1127 378 -1093
rect 412 -1127 424 -1093
rect 366 -1133 424 -1127
rect 524 -1093 582 -1087
rect 524 -1127 536 -1093
rect 570 -1127 582 -1093
rect 524 -1133 582 -1127
rect 682 -1093 740 -1087
rect 682 -1127 694 -1093
rect 728 -1127 740 -1093
rect 682 -1133 740 -1127
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
