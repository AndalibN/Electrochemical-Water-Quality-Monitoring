magic
tech sky130A
magscale 1 2
timestamp 1667404707
<< nwell >>
rect -194 -2100 194 2100
<< pmos >>
rect -100 -2000 100 2000
<< pdiff >>
rect -158 1988 -100 2000
rect -158 -1988 -146 1988
rect -112 -1988 -100 1988
rect -158 -2000 -100 -1988
rect 100 1988 158 2000
rect 100 -1988 112 1988
rect 146 -1988 158 1988
rect 100 -2000 158 -1988
<< pdiffc >>
rect -146 -1988 -112 1988
rect 112 -1988 146 1988
<< poly >>
rect -100 2081 100 2097
rect -100 2047 -84 2081
rect 84 2047 100 2081
rect -100 2000 100 2047
rect -100 -2047 100 -2000
rect -100 -2081 -84 -2047
rect 84 -2081 100 -2047
rect -100 -2097 100 -2081
<< polycont >>
rect -84 2047 84 2081
rect -84 -2081 84 -2047
<< locali >>
rect -100 2047 -84 2081
rect 84 2047 100 2081
rect -146 1988 -112 2004
rect -146 -2004 -112 -1988
rect 112 1988 146 2004
rect 112 -2004 146 -1988
rect -100 -2081 -84 -2047
rect 84 -2081 100 -2047
<< viali >>
rect -84 2047 84 2081
rect -146 -1988 -112 1988
rect 112 -1988 146 1988
rect -84 -2081 84 -2047
<< metal1 >>
rect -96 2081 96 2087
rect -96 2047 -84 2081
rect 84 2047 96 2081
rect -96 2041 96 2047
rect -152 1988 -106 2000
rect -152 -1988 -146 1988
rect -112 -1988 -106 1988
rect -152 -2000 -106 -1988
rect 106 1988 152 2000
rect 106 -1988 112 1988
rect 146 -1988 152 1988
rect 106 -2000 152 -1988
rect -96 -2047 96 -2041
rect -96 -2081 -84 -2047
rect 84 -2081 96 -2047
rect -96 -2087 96 -2081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
