magic
tech sky130A
magscale 1 2
timestamp 1666707788
<< nwell >>
rect -296 -909 296 909
<< pmos >>
rect -100 -690 100 690
<< pdiff >>
rect -158 678 -100 690
rect -158 -678 -146 678
rect -112 -678 -100 678
rect -158 -690 -100 -678
rect 100 678 158 690
rect 100 -678 112 678
rect 146 -678 158 678
rect 100 -690 158 -678
<< pdiffc >>
rect -146 -678 -112 678
rect 112 -678 146 678
<< nsubdiff >>
rect -260 839 -164 873
rect 164 839 260 873
rect -260 777 -226 839
rect 226 777 260 839
rect -260 -839 -226 -777
rect 226 -839 260 -777
rect -260 -873 -164 -839
rect 164 -873 260 -839
<< nsubdiffcont >>
rect -164 839 164 873
rect -260 -777 -226 777
rect 226 -777 260 777
rect -164 -873 164 -839
<< poly >>
rect -100 771 100 787
rect -100 737 -84 771
rect 84 737 100 771
rect -100 690 100 737
rect -100 -737 100 -690
rect -100 -771 -84 -737
rect 84 -771 100 -737
rect -100 -787 100 -771
<< polycont >>
rect -84 737 84 771
rect -84 -771 84 -737
<< locali >>
rect -260 839 -164 873
rect 164 839 260 873
rect -260 777 -226 839
rect 226 777 260 839
rect -100 737 -84 771
rect 84 737 100 771
rect -146 678 -112 694
rect -146 -694 -112 -678
rect 112 678 146 694
rect 112 -694 146 -678
rect -100 -771 -84 -737
rect 84 -771 100 -737
rect -260 -839 -226 -777
rect 226 -839 260 -777
rect -260 -873 -164 -839
rect 164 -873 260 -839
<< viali >>
rect -84 737 84 771
rect -146 -678 -112 678
rect 112 -678 146 678
rect -84 -771 84 -737
<< metal1 >>
rect -96 771 96 777
rect -96 737 -84 771
rect 84 737 96 771
rect -96 731 96 737
rect -152 678 -106 690
rect -152 -678 -146 678
rect -112 -678 -106 678
rect -152 -690 -106 -678
rect 106 678 152 690
rect 106 -678 112 678
rect 146 -678 152 678
rect 106 -690 152 -678
rect -96 -737 96 -731
rect -96 -771 -84 -737
rect 84 -771 96 -737
rect -96 -777 96 -771
<< properties >>
string FIXED_BBOX -243 -856 243 856
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.9 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
