magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_s >>
rect 6997 1084 7003 1090
rect 7043 1084 7049 1090
rect 6991 1078 6997 1084
rect 7049 1078 7055 1084
rect 6991 1032 6997 1038
rect 7049 1032 7055 1038
rect 6997 1026 7003 1032
rect 7043 1026 7049 1032
rect 7004 578 7010 584
rect 7050 578 7056 584
rect 6998 572 7004 578
rect 7056 572 7062 578
rect 6998 526 7004 532
rect 7056 526 7062 532
rect 7004 520 7010 526
rect 7050 520 7056 526
rect 7001 -272 7007 -266
rect 7047 -272 7053 -266
rect 6995 -278 7001 -272
rect 7053 -278 7059 -272
rect 6995 -324 7001 -318
rect 7053 -324 7059 -318
rect 7001 -330 7007 -324
rect 7047 -330 7053 -324
rect 7002 -786 7008 -780
rect 7048 -786 7054 -780
rect 6996 -792 7002 -786
rect 7054 -792 7060 -786
rect 6996 -838 7002 -832
rect 7054 -838 7060 -832
rect 7002 -844 7008 -838
rect 7048 -844 7054 -838
rect 6997 -1636 7003 -1630
rect 7043 -1636 7049 -1630
rect 6991 -1642 6997 -1636
rect 7049 -1642 7055 -1636
rect 6991 -1688 6997 -1682
rect 7049 -1688 7055 -1682
rect 6997 -1694 7003 -1688
rect 7043 -1694 7049 -1688
rect 7000 -2154 7006 -2148
rect 7046 -2154 7052 -2148
rect 6994 -2160 7000 -2154
rect 7052 -2160 7058 -2154
rect 6994 -2206 7000 -2200
rect 7052 -2206 7058 -2200
rect 7000 -2212 7006 -2206
rect 7046 -2212 7052 -2206
rect 6999 -2994 7005 -2988
rect 7045 -2994 7051 -2988
rect 6993 -3000 6999 -2994
rect 7051 -3000 7057 -2994
rect 6993 -3046 6999 -3040
rect 7051 -3046 7057 -3040
rect 6999 -3052 7005 -3046
rect 7045 -3052 7051 -3046
rect 7011 -3508 7017 -3502
rect 7057 -3508 7063 -3502
rect 7005 -3514 7011 -3508
rect 7063 -3514 7069 -3508
rect 7005 -3560 7011 -3554
rect 7063 -3560 7069 -3554
rect 7011 -3566 7017 -3560
rect 7057 -3566 7063 -3560
<< nwell >>
rect 202 8696 484 8698
rect 5412 8696 7638 8698
rect 202 8058 10380 8696
rect 202 7158 10370 8058
rect 202 5194 10376 7158
rect 202 5116 1708 5194
rect 1966 5168 10376 5194
rect 1966 5166 3012 5168
rect 3314 5166 10376 5168
rect 4360 5148 10376 5166
rect 6864 5134 10370 5148
rect 202 5062 590 5116
rect 202 994 484 5062
rect 520 5034 560 5062
rect 860 2370 1708 5116
rect 8270 5112 8544 5134
rect 8540 4738 8544 5112
rect 860 1068 1352 2370
rect 1452 2368 1708 2370
rect 1454 2364 1708 2368
rect 1458 2248 1708 2364
rect 1630 2174 1708 2248
rect 860 986 1216 1068
<< pwell >>
rect 8180 -4928 9438 -4926
rect 9776 -4928 9912 -4926
rect 13022 -4928 13474 -4926
rect -2150 -4930 -2068 -4928
rect -1162 -4930 -892 -4928
rect 5662 -4930 10314 -4928
rect 11234 -4930 14048 -4928
rect -2150 -5242 14048 -4930
rect -2128 -5244 -1066 -5242
<< psubdiff >>
rect 8206 -4954 9412 -4952
rect 9802 -4954 9886 -4952
rect 13048 -4954 13448 -4952
rect -2124 -4956 -2094 -4954
rect -1136 -4956 -918 -4954
rect 5688 -4956 10288 -4954
rect 11260 -4956 14022 -4954
rect -2124 -5005 14022 -4956
rect -2124 -5008 11122 -5005
rect -2124 -5009 9452 -5008
rect -2124 -5010 8385 -5009
rect -2124 -5180 -2079 -5010
rect -1841 -5011 1803 -5010
rect -1841 -5020 -1174 -5011
rect -1841 -5180 -1635 -5020
rect -2124 -5190 -1635 -5180
rect -1261 -5181 -1174 -5020
rect -868 -5180 1803 -5011
rect 2109 -5011 6663 -5010
rect 2109 -5015 5301 -5011
rect 2109 -5180 2193 -5015
rect -868 -5181 2193 -5180
rect -1261 -5185 2193 -5181
rect 2499 -5038 5301 -5015
rect 2499 -5140 4546 -5038
rect 5056 -5140 5301 -5038
rect 2499 -5181 5301 -5140
rect 5879 -5180 6663 -5011
rect 7241 -5179 8385 -5010
rect 9235 -5178 9452 -5009
rect 10166 -5175 11122 -5008
rect 11496 -5009 14022 -5005
rect 11496 -5175 12224 -5009
rect 10166 -5178 12224 -5175
rect 9235 -5179 12224 -5178
rect 12666 -5011 13632 -5009
rect 12666 -5179 12833 -5011
rect 7241 -5180 12833 -5179
rect 5879 -5181 12833 -5180
rect 13207 -5179 13632 -5011
rect 13938 -5179 14022 -5009
rect 13207 -5181 14022 -5179
rect 2499 -5185 14022 -5181
rect -1261 -5190 14022 -5185
rect -2124 -5216 14022 -5190
rect -2102 -5218 -1092 -5216
<< nsubdiff >>
rect 6878 8608 7236 8614
rect 2942 8606 10338 8608
rect 516 8561 10338 8606
rect 516 8558 6897 8561
rect 516 8530 5881 8558
rect 516 8526 5340 8530
rect 516 8356 530 8526
rect 972 8525 5340 8526
rect 972 8356 2269 8525
rect 516 8355 2269 8356
rect 2711 8522 5340 8525
rect 2711 8355 3609 8522
rect 516 8352 3609 8355
rect 4051 8360 5340 8522
rect 5714 8360 5881 8530
rect 4051 8352 5881 8360
rect 516 8320 5881 8352
rect 6119 8323 6897 8558
rect 7203 8558 10338 8561
rect 7203 8323 7870 8558
rect 6119 8320 7870 8323
rect 8176 8320 8786 8558
rect 9092 8556 10338 8558
rect 9092 8320 9650 8556
rect 516 8318 9650 8320
rect 9956 8318 10338 8556
rect 516 8276 10338 8318
rect 2942 8274 4306 8276
rect 7586 8274 10338 8276
rect 3860 8272 3892 8274
<< psubdiffcont >>
rect -2079 -5180 -1841 -5010
rect -1635 -5190 -1261 -5020
rect -1174 -5181 -868 -5011
rect 1803 -5180 2109 -5010
rect 2193 -5185 2499 -5015
rect 4546 -5140 5056 -5038
rect 5301 -5181 5879 -5011
rect 6663 -5180 7241 -5010
rect 8385 -5179 9235 -5009
rect 9452 -5178 10166 -5008
rect 11122 -5175 11496 -5005
rect 12224 -5179 12666 -5009
rect 12833 -5181 13207 -5011
rect 13632 -5179 13938 -5009
<< nsubdiffcont >>
rect 530 8356 972 8526
rect 2269 8355 2711 8525
rect 3609 8352 4051 8522
rect 5340 8360 5714 8530
rect 5881 8320 6119 8558
rect 6897 8323 7203 8561
rect 7870 8320 8176 8558
rect 8786 8320 9092 8558
rect 9650 8318 9956 8556
<< locali >>
rect 6878 8576 7236 8582
rect 526 8561 10322 8576
rect 526 8558 6897 8561
rect 526 8530 5881 8558
rect 526 8526 5340 8530
rect 526 8356 530 8526
rect 972 8525 5340 8526
rect 972 8356 2269 8525
rect 526 8355 2269 8356
rect 2711 8522 5340 8525
rect 2711 8355 3609 8522
rect 526 8352 3609 8355
rect 4051 8360 5340 8522
rect 5714 8360 5881 8530
rect 4051 8352 5881 8360
rect 526 8320 5881 8352
rect 6119 8323 6897 8558
rect 7203 8558 10322 8561
rect 7203 8323 7870 8558
rect 6119 8320 7870 8323
rect 8176 8320 8786 8558
rect 9092 8556 10322 8558
rect 9092 8320 9650 8556
rect 526 8318 9650 8320
rect 9956 8318 10322 8556
rect 526 8306 10322 8318
rect 526 8276 566 8306
rect 524 8206 566 8276
rect 2476 8260 2514 8306
rect 3826 8260 3860 8306
rect 2472 8214 2512 8260
rect 3822 8214 3860 8260
rect 5458 8260 5496 8306
rect 5682 8304 7570 8306
rect 5458 8214 5492 8260
rect 5916 8214 5950 8304
rect 522 7158 566 8206
rect 2470 7158 2512 8214
rect 3820 7158 3862 8214
rect 522 5444 564 7158
rect 2470 5444 2510 7158
rect 522 5308 560 5444
rect 332 5270 562 5308
rect 332 5064 376 5270
rect 2470 5220 2508 5444
rect 2472 5086 2506 5220
rect 3820 5214 3858 7158
rect 5456 7154 5492 8214
rect 5914 7154 5950 8214
rect 6946 8278 6986 8304
rect 6946 8266 6984 8278
rect 6946 8198 6982 8266
rect 8004 8202 8038 8306
rect 8868 8208 8902 8306
rect 6946 7954 6980 8198
rect 8004 8050 8040 8202
rect 8866 8056 8902 8208
rect 9716 8202 9754 8306
rect 9716 8198 9752 8202
rect 9718 8060 9752 8198
rect 5456 7048 5490 7154
rect 5914 7064 5948 7154
rect 5946 7056 5948 7064
rect 3818 5090 3858 5214
rect -1166 4712 -1086 4796
rect 10290 4280 10506 4322
rect 10290 4278 10342 4280
rect 798 4138 1362 4194
rect 4280 3252 5096 3328
rect 4280 3250 4362 3252
rect 4468 3100 4790 3144
rect 3390 1190 3392 1200
rect 800 1132 944 1188
rect 1660 1146 2014 1182
rect 686 994 774 1054
rect 686 992 720 994
rect -1848 -1660 -1784 682
rect 896 -84 942 1132
rect 1142 992 1222 1056
rect 1136 844 1220 950
rect 1920 730 1960 1146
rect 2922 1106 2982 1178
rect 3220 1116 3362 1190
rect 3364 1120 3392 1190
rect 2710 1056 3460 1058
rect 2710 1024 3408 1056
rect 2240 950 2310 1024
rect 3562 1008 3676 1082
rect 3980 950 4040 1036
rect 4150 1004 4240 1070
rect 2240 880 4040 950
rect 4468 844 4544 3100
rect 4736 3044 4790 3100
rect 5026 2750 5096 3252
rect 10196 3116 10220 3156
rect 9340 3044 9798 3046
rect 8636 3040 8960 3044
rect 5876 3034 7472 3036
rect 8420 3034 8960 3040
rect 5876 2998 8120 3034
rect 5876 2996 7472 2998
rect 7994 2996 8120 2998
rect 8330 2996 8960 3034
rect 9272 3032 9798 3044
rect 9030 3000 9798 3032
rect 9030 2998 9498 3000
rect 8400 2994 8960 2996
rect 8420 2988 8960 2994
rect 5026 2692 8190 2750
rect 5026 2690 5286 2692
rect 5026 2594 5096 2690
rect 4926 2590 5228 2594
rect 4926 2534 5890 2590
rect 5834 1545 5890 2534
rect 8140 2586 8190 2692
rect 8698 2588 9676 2590
rect 8698 2586 9736 2588
rect 10290 2586 10340 4278
rect 8140 2518 10340 2586
rect 8140 2516 9736 2518
rect 8140 2514 9676 2516
rect 6330 2414 6412 2488
rect 6820 2156 6916 2170
rect 6820 2103 8118 2156
rect 6820 2069 6876 2103
rect 6910 2069 6948 2103
rect 6982 2069 7020 2103
rect 7054 2069 7092 2103
rect 7126 2069 7164 2103
rect 7198 2069 7236 2103
rect 7270 2069 7308 2103
rect 7342 2069 7380 2103
rect 7414 2069 7452 2103
rect 7486 2069 7524 2103
rect 7558 2069 7596 2103
rect 7630 2069 7668 2103
rect 7702 2069 7740 2103
rect 7774 2069 7812 2103
rect 7846 2069 7884 2103
rect 7918 2069 7956 2103
rect 7990 2069 8028 2103
rect 8062 2069 8118 2103
rect 6820 2050 8118 2069
rect 6820 1984 6922 2050
rect 6820 1950 6859 1984
rect 6893 1950 6922 1984
rect 6820 1912 6922 1950
rect 6986 1969 7952 1986
rect 6986 1935 7019 1969
rect 7053 1935 7091 1969
rect 7125 1935 7163 1969
rect 7197 1935 7235 1969
rect 7269 1935 7307 1969
rect 7341 1935 7379 1969
rect 7413 1935 7451 1969
rect 7485 1935 7523 1969
rect 7557 1935 7595 1969
rect 7629 1935 7667 1969
rect 7701 1935 7739 1969
rect 7773 1935 7811 1969
rect 7845 1935 7952 1969
rect 6986 1926 7952 1935
rect 6820 1878 6859 1912
rect 6893 1878 6922 1912
rect 6522 1736 6558 1864
rect 6820 1840 6922 1878
rect 6984 1918 7952 1926
rect 8014 1984 8116 2050
rect 8014 1950 8045 1984
rect 8079 1950 8116 1984
rect 6984 1883 7062 1918
rect 6984 1849 7009 1883
rect 7043 1849 7062 1883
rect 7874 1883 7948 1918
rect 6984 1846 7062 1849
rect 6820 1806 6859 1840
rect 6893 1806 6922 1840
rect 6820 1768 6922 1806
rect 5834 1124 6370 1545
rect 6520 1432 6562 1736
rect 6820 1734 6859 1768
rect 6893 1734 6922 1768
rect 6820 1696 6922 1734
rect 6820 1662 6859 1696
rect 6893 1662 6922 1696
rect 6820 1624 6922 1662
rect 6820 1590 6859 1624
rect 6893 1590 6922 1624
rect 6820 1552 6922 1590
rect 6820 1518 6859 1552
rect 6893 1518 6922 1552
rect 6820 1480 6922 1518
rect 6820 1446 6859 1480
rect 6893 1446 6922 1480
rect 3220 766 4544 844
rect 4700 972 4744 1006
rect 1660 650 1684 720
rect 1920 690 3510 730
rect 1890 522 3150 528
rect 892 -196 942 -84
rect 1862 482 3150 522
rect 1862 448 1911 482
rect 1945 448 1983 482
rect 2017 448 2055 482
rect 2089 448 2127 482
rect 2161 448 2199 482
rect 2233 448 2271 482
rect 2305 448 2343 482
rect 2377 448 2415 482
rect 2449 448 2487 482
rect 2521 448 2559 482
rect 2593 448 2631 482
rect 2665 448 2703 482
rect 2737 448 2775 482
rect 2809 448 2847 482
rect 2881 448 2919 482
rect 2953 448 2991 482
rect 3025 448 3063 482
rect 3097 448 3150 482
rect 3300 480 3368 552
rect 1862 428 3150 448
rect 1862 363 1954 428
rect 1862 329 1892 363
rect 1926 329 1954 363
rect 1862 291 1954 329
rect 2022 349 2986 368
rect 2022 315 2053 349
rect 2087 315 2125 349
rect 2159 315 2197 349
rect 2231 315 2269 349
rect 2303 315 2341 349
rect 2375 315 2413 349
rect 2447 315 2485 349
rect 2519 315 2557 349
rect 2591 315 2629 349
rect 2663 315 2701 349
rect 2735 315 2773 349
rect 2807 315 2845 349
rect 2879 315 2917 349
rect 2951 315 2986 349
rect 2022 312 2986 315
rect 1862 257 1892 291
rect 1926 257 1954 291
rect 1862 219 1954 257
rect 1862 185 1892 219
rect 1926 185 1954 219
rect 1862 147 1954 185
rect 1862 113 1892 147
rect 1926 113 1954 147
rect 1862 75 1954 113
rect 1862 41 1892 75
rect 1926 41 1954 75
rect 1862 3 1954 41
rect 1862 -31 1892 3
rect 1926 -31 1954 3
rect 1862 -69 1954 -31
rect 1862 -103 1892 -69
rect 1926 -103 1954 -69
rect 1862 -141 1954 -103
rect 1862 -175 1892 -141
rect 1926 -175 1954 -141
rect 892 -244 1266 -196
rect 1862 -213 1954 -175
rect 892 -446 940 -244
rect -910 -498 -860 -488
rect -910 -666 -836 -498
rect 1216 -582 1264 -244
rect 1862 -247 1892 -213
rect 1926 -247 1954 -213
rect 1862 -285 1954 -247
rect 1862 -319 1892 -285
rect 1926 -319 1954 -285
rect 1862 -357 1954 -319
rect 1862 -391 1892 -357
rect 1926 -391 1954 -357
rect 1862 -429 1954 -391
rect 1862 -463 1892 -429
rect 1926 -463 1954 -429
rect 1862 -501 1954 -463
rect 1862 -535 1892 -501
rect 1926 -535 1954 -501
rect 2020 298 2986 312
rect 2020 263 2090 298
rect 2020 229 2042 263
rect 2076 229 2090 263
rect 2916 263 2986 298
rect 2020 191 2090 229
rect 2020 157 2042 191
rect 2076 157 2090 191
rect 2020 119 2090 157
rect 2020 85 2042 119
rect 2076 85 2090 119
rect 2020 47 2090 85
rect 2020 13 2042 47
rect 2076 13 2090 47
rect 2020 -25 2090 13
rect 2020 -59 2042 -25
rect 2076 -59 2090 -25
rect 2020 -97 2090 -59
rect 2020 -131 2042 -97
rect 2076 -131 2090 -97
rect 2020 -169 2090 -131
rect 2020 -203 2042 -169
rect 2076 -203 2090 -169
rect 2020 -241 2090 -203
rect 2020 -275 2042 -241
rect 2076 -275 2090 -241
rect 2020 -313 2090 -275
rect 2020 -347 2042 -313
rect 2076 -347 2090 -313
rect 2020 -385 2090 -347
rect 2020 -419 2042 -385
rect 2076 -419 2090 -385
rect 2020 -457 2090 -419
rect 2020 -491 2042 -457
rect 2076 -491 2090 -457
rect 2154 -462 2844 230
rect 2916 229 2932 263
rect 2966 229 2986 263
rect 2916 191 2986 229
rect 2916 157 2932 191
rect 2966 157 2986 191
rect 2916 119 2986 157
rect 2916 85 2932 119
rect 2966 85 2986 119
rect 2916 47 2986 85
rect 2916 13 2932 47
rect 2966 13 2986 47
rect 2916 -25 2986 13
rect 2916 -59 2932 -25
rect 2966 -59 2986 -25
rect 2916 -97 2986 -59
rect 2916 -131 2932 -97
rect 2966 -131 2986 -97
rect 2916 -169 2986 -131
rect 2916 -203 2932 -169
rect 2966 -203 2986 -169
rect 2916 -241 2986 -203
rect 2916 -275 2932 -241
rect 2966 -275 2986 -241
rect 2916 -313 2986 -275
rect 2916 -347 2932 -313
rect 2966 -347 2986 -313
rect 2916 -385 2986 -347
rect 2916 -419 2932 -385
rect 2966 -419 2986 -385
rect 2916 -457 2986 -419
rect 2020 -526 2090 -491
rect 2916 -491 2932 -457
rect 2966 -491 2986 -457
rect 2916 -526 2986 -491
rect 1862 -573 1954 -535
rect 1862 -607 1892 -573
rect 1926 -607 1954 -573
rect 2018 -543 2986 -526
rect 2018 -577 2042 -543
rect 2076 -577 2127 -543
rect 2161 -577 2199 -543
rect 2233 -577 2271 -543
rect 2305 -577 2343 -543
rect 2377 -577 2415 -543
rect 2449 -577 2487 -543
rect 2521 -577 2559 -543
rect 2593 -577 2631 -543
rect 2665 -577 2703 -543
rect 2737 -577 2775 -543
rect 2809 -577 2847 -543
rect 2881 -577 2932 -543
rect 2966 -577 2986 -543
rect 2018 -596 2986 -577
rect 3052 363 3144 428
rect 3052 329 3082 363
rect 3116 329 3144 363
rect 3052 291 3144 329
rect 3052 257 3082 291
rect 3116 257 3144 291
rect 3052 219 3144 257
rect 3052 185 3082 219
rect 3116 185 3144 219
rect 3052 147 3144 185
rect 3052 113 3082 147
rect 3116 113 3144 147
rect 3052 75 3144 113
rect 3052 41 3082 75
rect 3116 41 3144 75
rect 3052 3 3144 41
rect 3052 -31 3082 3
rect 3116 -31 3144 3
rect 3052 -69 3144 -31
rect 3052 -103 3082 -69
rect 3116 -103 3144 -69
rect 3052 -141 3144 -103
rect 3052 -175 3082 -141
rect 3116 -175 3144 -141
rect 3052 -213 3144 -175
rect 3052 -247 3082 -213
rect 3116 -247 3144 -213
rect 3052 -285 3144 -247
rect 3052 -319 3082 -285
rect 3116 -319 3144 -285
rect 3052 -357 3144 -319
rect 3052 -391 3082 -357
rect 3116 -391 3144 -357
rect 3052 -429 3144 -391
rect 3052 -463 3082 -429
rect 3116 -463 3144 -429
rect 3052 -501 3144 -463
rect 3052 -535 3082 -501
rect 3116 -535 3144 -501
rect 3052 -573 3144 -535
rect 2018 -598 2100 -596
rect 1862 -660 1954 -607
rect 3052 -607 3082 -573
rect 3116 -607 3144 -573
rect 3052 -660 3144 -607
rect -2022 -1736 -1782 -1660
rect -2020 -3420 -1950 -1736
rect -1166 -2236 -1090 -1820
rect -1378 -3136 -1328 -2946
rect -2018 -4950 -1950 -3420
rect -1588 -3186 -1328 -3136
rect -1588 -4950 -1532 -3186
rect -1158 -3540 -1090 -3286
rect -1374 -3594 -1090 -3540
rect -910 -3566 -860 -666
rect 1860 -692 3144 -660
rect 1860 -726 1911 -692
rect 1945 -726 1983 -692
rect 2017 -726 2055 -692
rect 2089 -726 2127 -692
rect 2161 -726 2199 -692
rect 2233 -726 2271 -692
rect 2305 -726 2343 -692
rect 2377 -726 2415 -692
rect 2449 -726 2487 -692
rect 2521 -726 2559 -692
rect 2593 -726 2631 -692
rect 2665 -726 2703 -692
rect 2737 -726 2775 -692
rect 2809 -726 2847 -692
rect 2881 -726 2919 -692
rect 2953 -726 2991 -692
rect 3025 -726 3063 -692
rect 3097 -726 3144 -692
rect 1860 -754 3144 -726
rect 1860 -760 3120 -754
rect 1888 -1358 1952 -760
rect 3304 -826 3368 480
rect 2392 -884 3368 -826
rect 2392 -1096 2430 -884
rect 3460 -988 3510 690
rect 4700 660 4742 972
rect 3930 630 4742 660
rect 3930 608 4740 630
rect 3930 400 3980 608
rect 3928 352 4094 400
rect 3928 350 4066 352
rect 3932 -818 3976 350
rect 4580 156 5092 158
rect 6120 156 6154 274
rect 4580 122 6154 156
rect 4580 120 5096 122
rect 6120 120 6154 122
rect 3932 -864 4536 -818
rect 3932 -866 3976 -864
rect 3460 -1012 3508 -988
rect 4502 -1074 4536 -864
rect 2392 -1144 2452 -1096
rect 4482 -1110 4536 -1074
rect -912 -3570 -860 -3566
rect -1374 -4922 -1298 -3594
rect -912 -3748 -858 -3570
rect -1126 -3792 -858 -3748
rect -2018 -4978 -1948 -4950
rect -1590 -4978 -1530 -4950
rect -1374 -4978 -1296 -4922
rect -1126 -4950 -1078 -3792
rect 1890 -4950 1950 -1358
rect -1126 -4978 -1076 -4950
rect -2110 -4980 -914 -4978
rect 1890 -4980 1954 -4950
rect 4582 -4980 4644 120
rect 6520 0 6560 1432
rect 6820 1408 6922 1446
rect 6820 1374 6859 1408
rect 6893 1374 6922 1408
rect 6820 1336 6922 1374
rect 6820 1302 6859 1336
rect 6893 1302 6922 1336
rect 6820 1264 6922 1302
rect 6820 1230 6859 1264
rect 6893 1230 6922 1264
rect 6820 1192 6922 1230
rect 6820 1158 6859 1192
rect 6893 1158 6922 1192
rect 6820 1120 6922 1158
rect 6820 1086 6859 1120
rect 6893 1086 6922 1120
rect 6986 1811 7060 1846
rect 6986 1777 7009 1811
rect 7043 1777 7060 1811
rect 6986 1739 7060 1777
rect 6986 1705 7009 1739
rect 7043 1705 7060 1739
rect 6986 1667 7060 1705
rect 6986 1633 7009 1667
rect 7043 1633 7060 1667
rect 6986 1595 7060 1633
rect 6986 1561 7009 1595
rect 7043 1561 7060 1595
rect 6986 1523 7060 1561
rect 6986 1489 7009 1523
rect 7043 1489 7060 1523
rect 6986 1451 7060 1489
rect 6986 1417 7009 1451
rect 7043 1417 7060 1451
rect 6986 1379 7060 1417
rect 6986 1345 7009 1379
rect 7043 1345 7060 1379
rect 6986 1307 7060 1345
rect 6986 1273 7009 1307
rect 7043 1273 7060 1307
rect 6986 1235 7060 1273
rect 6986 1201 7009 1235
rect 7043 1201 7060 1235
rect 6986 1163 7060 1201
rect 7126 1168 7808 1858
rect 7874 1849 7899 1883
rect 7933 1849 7948 1883
rect 7874 1811 7948 1849
rect 7874 1777 7899 1811
rect 7933 1777 7948 1811
rect 7874 1739 7948 1777
rect 7874 1705 7899 1739
rect 7933 1705 7948 1739
rect 7874 1667 7948 1705
rect 7874 1633 7899 1667
rect 7933 1633 7948 1667
rect 7874 1595 7948 1633
rect 7874 1561 7899 1595
rect 7933 1561 7948 1595
rect 7874 1523 7948 1561
rect 7874 1489 7899 1523
rect 7933 1489 7948 1523
rect 7874 1451 7948 1489
rect 7874 1417 7899 1451
rect 7933 1417 7948 1451
rect 7874 1379 7948 1417
rect 7874 1345 7899 1379
rect 7933 1345 7948 1379
rect 7874 1307 7948 1345
rect 7874 1273 7899 1307
rect 7933 1273 7948 1307
rect 7874 1235 7948 1273
rect 7874 1201 7899 1235
rect 7933 1201 7948 1235
rect 6986 1129 7009 1163
rect 7043 1129 7060 1163
rect 6986 1098 7060 1129
rect 7874 1163 7948 1201
rect 7874 1129 7899 1163
rect 7933 1129 7948 1163
rect 6820 1048 6922 1086
rect 6820 1014 6859 1048
rect 6893 1014 6922 1048
rect 6980 1094 7066 1098
rect 7874 1094 7948 1129
rect 8014 1912 8116 1950
rect 8014 1878 8045 1912
rect 8079 1878 8116 1912
rect 8014 1840 8116 1878
rect 8014 1806 8045 1840
rect 8079 1806 8116 1840
rect 8014 1768 8116 1806
rect 8014 1734 8045 1768
rect 8079 1734 8116 1768
rect 8014 1696 8116 1734
rect 8014 1662 8045 1696
rect 8079 1662 8116 1696
rect 8014 1624 8116 1662
rect 8014 1590 8045 1624
rect 8079 1590 8116 1624
rect 8014 1552 8116 1590
rect 8014 1518 8045 1552
rect 8079 1518 8116 1552
rect 8014 1480 8116 1518
rect 8014 1446 8045 1480
rect 8079 1446 8116 1480
rect 8014 1408 8116 1446
rect 8014 1374 8045 1408
rect 8079 1374 8116 1408
rect 8014 1336 8116 1374
rect 8014 1302 8045 1336
rect 8079 1302 8116 1336
rect 8014 1264 8116 1302
rect 8014 1230 8045 1264
rect 8079 1230 8116 1264
rect 8014 1192 8116 1230
rect 8014 1158 8045 1192
rect 8079 1158 8116 1192
rect 8014 1120 8116 1158
rect 6980 1077 7950 1094
rect 6980 1043 7009 1077
rect 7043 1043 7094 1077
rect 7128 1043 7166 1077
rect 7200 1043 7238 1077
rect 7272 1043 7310 1077
rect 7344 1043 7382 1077
rect 7416 1043 7454 1077
rect 7488 1043 7526 1077
rect 7560 1043 7598 1077
rect 7632 1043 7670 1077
rect 7704 1043 7742 1077
rect 7776 1043 7814 1077
rect 7848 1076 7950 1077
rect 7848 1043 7899 1076
rect 6980 1042 7899 1043
rect 7933 1042 7950 1076
rect 6980 1026 7950 1042
rect 8014 1086 8045 1120
rect 8079 1086 8116 1120
rect 8014 1048 8116 1086
rect 6980 1024 7066 1026
rect 7874 1022 7948 1026
rect 6820 966 6922 1014
rect 8014 1014 8045 1048
rect 8079 1014 8116 1048
rect 8014 966 8116 1014
rect 6820 929 8118 966
rect 6820 895 6876 929
rect 6910 895 6948 929
rect 6982 895 7020 929
rect 7054 895 7092 929
rect 7126 895 7164 929
rect 7198 895 7236 929
rect 7270 895 7308 929
rect 7342 895 7380 929
rect 7414 895 7452 929
rect 7486 895 7524 929
rect 7558 895 7596 929
rect 7630 895 7668 929
rect 7702 895 7740 929
rect 7774 895 7812 929
rect 7846 895 7884 929
rect 7918 895 7956 929
rect 7990 895 8028 929
rect 8062 895 8118 929
rect 6820 886 8118 895
rect 6818 860 8118 886
rect 6818 852 6920 860
rect 6820 812 6920 852
rect 4928 -42 6560 0
rect 4930 -66 6560 -42
rect 4930 -4980 5002 -66
rect 6520 -72 6560 -66
rect 6824 800 6920 812
rect 6824 747 8122 800
rect 6824 713 6880 747
rect 6914 713 6952 747
rect 6986 713 7024 747
rect 7058 713 7096 747
rect 7130 713 7168 747
rect 7202 713 7240 747
rect 7274 713 7312 747
rect 7346 713 7384 747
rect 7418 713 7456 747
rect 7490 713 7528 747
rect 7562 713 7600 747
rect 7634 713 7672 747
rect 7706 713 7744 747
rect 7778 713 7816 747
rect 7850 713 7888 747
rect 7922 713 7960 747
rect 7994 713 8032 747
rect 8066 713 8122 747
rect 6824 694 8122 713
rect 6824 628 6926 694
rect 6824 594 6863 628
rect 6897 594 6926 628
rect 6824 556 6926 594
rect 6990 613 7956 630
rect 6990 579 7023 613
rect 7057 579 7095 613
rect 7129 579 7167 613
rect 7201 579 7239 613
rect 7273 579 7311 613
rect 7345 579 7383 613
rect 7417 579 7455 613
rect 7489 579 7527 613
rect 7561 579 7599 613
rect 7633 579 7671 613
rect 7705 579 7743 613
rect 7777 579 7815 613
rect 7849 579 7956 613
rect 6990 570 7956 579
rect 6824 522 6863 556
rect 6897 522 6926 556
rect 6824 484 6926 522
rect 6988 562 7956 570
rect 8018 628 8120 694
rect 8018 594 8049 628
rect 8083 594 8120 628
rect 6988 527 7066 562
rect 6988 493 7013 527
rect 7047 493 7066 527
rect 7878 527 7952 562
rect 6988 490 7066 493
rect 6824 450 6863 484
rect 6897 450 6926 484
rect 6824 412 6926 450
rect 6824 378 6863 412
rect 6897 378 6926 412
rect 6824 340 6926 378
rect 6824 306 6863 340
rect 6897 306 6926 340
rect 6824 268 6926 306
rect 6824 234 6863 268
rect 6897 234 6926 268
rect 6824 196 6926 234
rect 6824 162 6863 196
rect 6897 162 6926 196
rect 6824 124 6926 162
rect 6824 90 6863 124
rect 6897 90 6926 124
rect 6824 52 6926 90
rect 6824 18 6863 52
rect 6897 18 6926 52
rect 6824 -20 6926 18
rect 6824 -54 6863 -20
rect 6897 -54 6926 -20
rect 6824 -92 6926 -54
rect 6824 -126 6863 -92
rect 6897 -126 6926 -92
rect 6824 -164 6926 -126
rect 6824 -198 6863 -164
rect 6897 -198 6926 -164
rect 6824 -236 6926 -198
rect 6824 -270 6863 -236
rect 6897 -270 6926 -236
rect 6990 455 7064 490
rect 6990 421 7013 455
rect 7047 421 7064 455
rect 6990 383 7064 421
rect 6990 349 7013 383
rect 7047 349 7064 383
rect 6990 311 7064 349
rect 6990 277 7013 311
rect 7047 277 7064 311
rect 6990 239 7064 277
rect 6990 205 7013 239
rect 7047 205 7064 239
rect 6990 167 7064 205
rect 6990 133 7013 167
rect 7047 133 7064 167
rect 6990 95 7064 133
rect 6990 61 7013 95
rect 7047 61 7064 95
rect 6990 23 7064 61
rect 6990 -11 7013 23
rect 7047 -11 7064 23
rect 6990 -49 7064 -11
rect 6990 -83 7013 -49
rect 7047 -83 7064 -49
rect 6990 -121 7064 -83
rect 6990 -155 7013 -121
rect 7047 -155 7064 -121
rect 6990 -193 7064 -155
rect 7130 -188 7812 502
rect 7878 493 7903 527
rect 7937 493 7952 527
rect 7878 455 7952 493
rect 7878 421 7903 455
rect 7937 421 7952 455
rect 7878 383 7952 421
rect 7878 349 7903 383
rect 7937 349 7952 383
rect 7878 311 7952 349
rect 7878 277 7903 311
rect 7937 277 7952 311
rect 7878 239 7952 277
rect 7878 205 7903 239
rect 7937 205 7952 239
rect 7878 167 7952 205
rect 7878 133 7903 167
rect 7937 133 7952 167
rect 7878 95 7952 133
rect 7878 61 7903 95
rect 7937 61 7952 95
rect 7878 23 7952 61
rect 7878 -11 7903 23
rect 7937 -11 7952 23
rect 7878 -49 7952 -11
rect 7878 -83 7903 -49
rect 7937 -83 7952 -49
rect 7878 -121 7952 -83
rect 7878 -155 7903 -121
rect 7937 -155 7952 -121
rect 6990 -227 7013 -193
rect 7047 -227 7064 -193
rect 6990 -258 7064 -227
rect 7878 -193 7952 -155
rect 7878 -227 7903 -193
rect 7937 -227 7952 -193
rect 6824 -308 6926 -270
rect 6824 -342 6863 -308
rect 6897 -342 6926 -308
rect 6984 -262 7070 -258
rect 7878 -262 7952 -227
rect 8018 556 8120 594
rect 8018 522 8049 556
rect 8083 522 8120 556
rect 8018 484 8120 522
rect 8018 450 8049 484
rect 8083 450 8120 484
rect 8018 412 8120 450
rect 8018 378 8049 412
rect 8083 378 8120 412
rect 8018 340 8120 378
rect 8018 306 8049 340
rect 8083 306 8120 340
rect 8018 268 8120 306
rect 8018 234 8049 268
rect 8083 234 8120 268
rect 8018 196 8120 234
rect 8018 162 8049 196
rect 8083 162 8120 196
rect 8018 124 8120 162
rect 8018 90 8049 124
rect 8083 90 8120 124
rect 8018 52 8120 90
rect 8018 18 8049 52
rect 8083 18 8120 52
rect 8018 -20 8120 18
rect 8018 -54 8049 -20
rect 8083 -54 8120 -20
rect 8018 -92 8120 -54
rect 8018 -126 8049 -92
rect 8083 -126 8120 -92
rect 8018 -164 8120 -126
rect 8018 -198 8049 -164
rect 8083 -198 8120 -164
rect 8018 -236 8120 -198
rect 6984 -279 7954 -262
rect 6984 -313 7013 -279
rect 7047 -313 7098 -279
rect 7132 -313 7170 -279
rect 7204 -313 7242 -279
rect 7276 -313 7314 -279
rect 7348 -313 7386 -279
rect 7420 -313 7458 -279
rect 7492 -313 7530 -279
rect 7564 -313 7602 -279
rect 7636 -313 7674 -279
rect 7708 -313 7746 -279
rect 7780 -313 7818 -279
rect 7852 -280 7954 -279
rect 7852 -313 7903 -280
rect 6984 -314 7903 -313
rect 7937 -314 7954 -280
rect 6984 -330 7954 -314
rect 8018 -270 8049 -236
rect 8083 -270 8120 -236
rect 8018 -308 8120 -270
rect 6984 -332 7070 -330
rect 7878 -334 7952 -330
rect 6824 -390 6926 -342
rect 8018 -342 8049 -308
rect 8083 -342 8120 -308
rect 8018 -390 8120 -342
rect 6824 -427 8122 -390
rect 6824 -461 6880 -427
rect 6914 -461 6952 -427
rect 6986 -461 7024 -427
rect 7058 -461 7096 -427
rect 7130 -461 7168 -427
rect 7202 -461 7240 -427
rect 7274 -461 7312 -427
rect 7346 -461 7384 -427
rect 7418 -461 7456 -427
rect 7490 -461 7528 -427
rect 7562 -461 7600 -427
rect 7634 -461 7672 -427
rect 7706 -461 7744 -427
rect 7778 -461 7816 -427
rect 7850 -461 7888 -427
rect 7922 -461 7960 -427
rect 7994 -461 8032 -427
rect 8066 -461 8122 -427
rect 6824 -470 8122 -461
rect 6822 -494 8122 -470
rect 6820 -496 8122 -494
rect 6820 -550 6914 -496
rect 5410 -568 5506 -554
rect 6820 -564 6916 -550
rect 5410 -621 6708 -568
rect 5410 -655 5466 -621
rect 5500 -655 5538 -621
rect 5572 -655 5610 -621
rect 5644 -655 5682 -621
rect 5716 -655 5754 -621
rect 5788 -655 5826 -621
rect 5860 -655 5898 -621
rect 5932 -655 5970 -621
rect 6004 -655 6042 -621
rect 6076 -655 6114 -621
rect 6148 -655 6186 -621
rect 6220 -655 6258 -621
rect 6292 -655 6330 -621
rect 6364 -655 6402 -621
rect 6436 -655 6474 -621
rect 6508 -655 6546 -621
rect 6580 -655 6618 -621
rect 6652 -655 6708 -621
rect 5410 -674 6708 -655
rect 6820 -617 8118 -564
rect 6820 -651 6876 -617
rect 6910 -651 6948 -617
rect 6982 -651 7020 -617
rect 7054 -651 7092 -617
rect 7126 -651 7164 -617
rect 7198 -651 7236 -617
rect 7270 -651 7308 -617
rect 7342 -651 7380 -617
rect 7414 -651 7452 -617
rect 7486 -651 7524 -617
rect 7558 -651 7596 -617
rect 7630 -651 7668 -617
rect 7702 -651 7740 -617
rect 7774 -651 7812 -617
rect 7846 -651 7884 -617
rect 7918 -651 7956 -617
rect 7990 -651 8028 -617
rect 8062 -651 8118 -617
rect 6820 -670 8118 -651
rect 5410 -740 5512 -674
rect 5410 -774 5449 -740
rect 5483 -774 5512 -740
rect 5410 -812 5512 -774
rect 5576 -755 6542 -738
rect 5576 -789 5609 -755
rect 5643 -789 5681 -755
rect 5715 -789 5753 -755
rect 5787 -789 5825 -755
rect 5859 -789 5897 -755
rect 5931 -789 5969 -755
rect 6003 -789 6041 -755
rect 6075 -789 6113 -755
rect 6147 -789 6185 -755
rect 6219 -789 6257 -755
rect 6291 -789 6329 -755
rect 6363 -789 6401 -755
rect 6435 -789 6542 -755
rect 5576 -798 6542 -789
rect 5410 -846 5449 -812
rect 5483 -846 5512 -812
rect 5410 -884 5512 -846
rect 5574 -806 6542 -798
rect 6604 -740 6706 -674
rect 6604 -774 6635 -740
rect 6669 -774 6706 -740
rect 5574 -841 5652 -806
rect 5574 -875 5599 -841
rect 5633 -875 5652 -841
rect 6464 -841 6538 -806
rect 5574 -878 5652 -875
rect 5410 -918 5449 -884
rect 5483 -918 5512 -884
rect 5410 -956 5512 -918
rect 5410 -990 5449 -956
rect 5483 -990 5512 -956
rect 5410 -1028 5512 -990
rect 5410 -1062 5449 -1028
rect 5483 -1062 5512 -1028
rect 5410 -1100 5512 -1062
rect 5410 -1134 5449 -1100
rect 5483 -1134 5512 -1100
rect 5410 -1172 5512 -1134
rect 5410 -1206 5449 -1172
rect 5483 -1206 5512 -1172
rect 5410 -1244 5512 -1206
rect 5410 -1278 5449 -1244
rect 5483 -1278 5512 -1244
rect 5410 -1316 5512 -1278
rect 5410 -1350 5449 -1316
rect 5483 -1350 5512 -1316
rect 5410 -1388 5512 -1350
rect 5410 -1422 5449 -1388
rect 5483 -1422 5512 -1388
rect 5410 -1460 5512 -1422
rect 5410 -1494 5449 -1460
rect 5483 -1494 5512 -1460
rect 5410 -1532 5512 -1494
rect 5410 -1566 5449 -1532
rect 5483 -1566 5512 -1532
rect 5410 -1604 5512 -1566
rect 5410 -1638 5449 -1604
rect 5483 -1638 5512 -1604
rect 5576 -913 5650 -878
rect 5576 -947 5599 -913
rect 5633 -947 5650 -913
rect 5576 -985 5650 -947
rect 5576 -1019 5599 -985
rect 5633 -1019 5650 -985
rect 5576 -1057 5650 -1019
rect 5576 -1091 5599 -1057
rect 5633 -1091 5650 -1057
rect 5576 -1129 5650 -1091
rect 5576 -1163 5599 -1129
rect 5633 -1163 5650 -1129
rect 5576 -1201 5650 -1163
rect 5576 -1235 5599 -1201
rect 5633 -1235 5650 -1201
rect 5576 -1273 5650 -1235
rect 5576 -1307 5599 -1273
rect 5633 -1307 5650 -1273
rect 5576 -1345 5650 -1307
rect 5576 -1379 5599 -1345
rect 5633 -1379 5650 -1345
rect 5576 -1417 5650 -1379
rect 5576 -1451 5599 -1417
rect 5633 -1451 5650 -1417
rect 5576 -1489 5650 -1451
rect 5576 -1523 5599 -1489
rect 5633 -1523 5650 -1489
rect 5576 -1561 5650 -1523
rect 5716 -1556 6398 -866
rect 6464 -875 6489 -841
rect 6523 -875 6538 -841
rect 6464 -913 6538 -875
rect 6464 -947 6489 -913
rect 6523 -947 6538 -913
rect 6464 -985 6538 -947
rect 6464 -1019 6489 -985
rect 6523 -1019 6538 -985
rect 6464 -1057 6538 -1019
rect 6464 -1091 6489 -1057
rect 6523 -1091 6538 -1057
rect 6464 -1129 6538 -1091
rect 6464 -1163 6489 -1129
rect 6523 -1163 6538 -1129
rect 6464 -1201 6538 -1163
rect 6464 -1235 6489 -1201
rect 6523 -1235 6538 -1201
rect 6464 -1273 6538 -1235
rect 6464 -1307 6489 -1273
rect 6523 -1307 6538 -1273
rect 6464 -1345 6538 -1307
rect 6464 -1379 6489 -1345
rect 6523 -1379 6538 -1345
rect 6464 -1417 6538 -1379
rect 6464 -1451 6489 -1417
rect 6523 -1451 6538 -1417
rect 6464 -1489 6538 -1451
rect 6464 -1523 6489 -1489
rect 6523 -1523 6538 -1489
rect 5576 -1595 5599 -1561
rect 5633 -1595 5650 -1561
rect 5576 -1626 5650 -1595
rect 6464 -1561 6538 -1523
rect 6464 -1595 6489 -1561
rect 6523 -1595 6538 -1561
rect 5410 -1676 5512 -1638
rect 5410 -1710 5449 -1676
rect 5483 -1710 5512 -1676
rect 5570 -1630 5656 -1626
rect 6464 -1630 6538 -1595
rect 6604 -812 6706 -774
rect 6604 -846 6635 -812
rect 6669 -846 6706 -812
rect 6604 -884 6706 -846
rect 6604 -918 6635 -884
rect 6669 -918 6706 -884
rect 6604 -956 6706 -918
rect 6604 -990 6635 -956
rect 6669 -990 6706 -956
rect 6604 -1028 6706 -990
rect 6604 -1062 6635 -1028
rect 6669 -1062 6706 -1028
rect 6604 -1100 6706 -1062
rect 6604 -1134 6635 -1100
rect 6669 -1134 6706 -1100
rect 6604 -1172 6706 -1134
rect 6604 -1206 6635 -1172
rect 6669 -1206 6706 -1172
rect 6604 -1244 6706 -1206
rect 6604 -1278 6635 -1244
rect 6669 -1278 6706 -1244
rect 6604 -1316 6706 -1278
rect 6604 -1350 6635 -1316
rect 6669 -1350 6706 -1316
rect 6604 -1388 6706 -1350
rect 6604 -1422 6635 -1388
rect 6669 -1422 6706 -1388
rect 6604 -1460 6706 -1422
rect 6604 -1494 6635 -1460
rect 6669 -1494 6706 -1460
rect 6604 -1532 6706 -1494
rect 6604 -1566 6635 -1532
rect 6669 -1566 6706 -1532
rect 6604 -1604 6706 -1566
rect 5570 -1647 6540 -1630
rect 5570 -1681 5599 -1647
rect 5633 -1681 5684 -1647
rect 5718 -1681 5756 -1647
rect 5790 -1681 5828 -1647
rect 5862 -1681 5900 -1647
rect 5934 -1681 5972 -1647
rect 6006 -1681 6044 -1647
rect 6078 -1681 6116 -1647
rect 6150 -1681 6188 -1647
rect 6222 -1681 6260 -1647
rect 6294 -1681 6332 -1647
rect 6366 -1681 6404 -1647
rect 6438 -1648 6540 -1647
rect 6438 -1681 6489 -1648
rect 5570 -1682 6489 -1681
rect 6523 -1682 6540 -1648
rect 5570 -1698 6540 -1682
rect 6604 -1638 6635 -1604
rect 6669 -1638 6706 -1604
rect 6604 -1676 6706 -1638
rect 5570 -1700 5656 -1698
rect 6464 -1702 6538 -1698
rect 5410 -1758 5512 -1710
rect 6604 -1710 6635 -1676
rect 6669 -1710 6706 -1676
rect 6604 -1758 6706 -1710
rect 6820 -736 6922 -670
rect 6820 -770 6859 -736
rect 6893 -770 6922 -736
rect 6820 -808 6922 -770
rect 6986 -751 7952 -734
rect 6986 -785 7019 -751
rect 7053 -785 7091 -751
rect 7125 -785 7163 -751
rect 7197 -785 7235 -751
rect 7269 -785 7307 -751
rect 7341 -785 7379 -751
rect 7413 -785 7451 -751
rect 7485 -785 7523 -751
rect 7557 -785 7595 -751
rect 7629 -785 7667 -751
rect 7701 -785 7739 -751
rect 7773 -785 7811 -751
rect 7845 -785 7952 -751
rect 6986 -794 7952 -785
rect 6820 -842 6859 -808
rect 6893 -842 6922 -808
rect 6820 -880 6922 -842
rect 6984 -802 7952 -794
rect 8014 -736 8116 -670
rect 8014 -770 8045 -736
rect 8079 -770 8116 -736
rect 6984 -837 7062 -802
rect 6984 -871 7009 -837
rect 7043 -871 7062 -837
rect 7874 -837 7948 -802
rect 6984 -874 7062 -871
rect 6820 -914 6859 -880
rect 6893 -914 6922 -880
rect 6820 -952 6922 -914
rect 6820 -986 6859 -952
rect 6893 -986 6922 -952
rect 6820 -1024 6922 -986
rect 6820 -1058 6859 -1024
rect 6893 -1058 6922 -1024
rect 6820 -1096 6922 -1058
rect 6820 -1130 6859 -1096
rect 6893 -1130 6922 -1096
rect 6820 -1168 6922 -1130
rect 6820 -1202 6859 -1168
rect 6893 -1202 6922 -1168
rect 6820 -1240 6922 -1202
rect 6820 -1274 6859 -1240
rect 6893 -1274 6922 -1240
rect 6820 -1312 6922 -1274
rect 6820 -1346 6859 -1312
rect 6893 -1346 6922 -1312
rect 6820 -1384 6922 -1346
rect 6820 -1418 6859 -1384
rect 6893 -1418 6922 -1384
rect 6820 -1456 6922 -1418
rect 6820 -1490 6859 -1456
rect 6893 -1490 6922 -1456
rect 6820 -1528 6922 -1490
rect 6820 -1562 6859 -1528
rect 6893 -1562 6922 -1528
rect 6820 -1600 6922 -1562
rect 6820 -1634 6859 -1600
rect 6893 -1634 6922 -1600
rect 6986 -909 7060 -874
rect 6986 -943 7009 -909
rect 7043 -943 7060 -909
rect 6986 -981 7060 -943
rect 6986 -1015 7009 -981
rect 7043 -1015 7060 -981
rect 6986 -1053 7060 -1015
rect 6986 -1087 7009 -1053
rect 7043 -1087 7060 -1053
rect 6986 -1125 7060 -1087
rect 6986 -1159 7009 -1125
rect 7043 -1159 7060 -1125
rect 6986 -1197 7060 -1159
rect 6986 -1231 7009 -1197
rect 7043 -1231 7060 -1197
rect 6986 -1269 7060 -1231
rect 6986 -1303 7009 -1269
rect 7043 -1303 7060 -1269
rect 6986 -1341 7060 -1303
rect 6986 -1375 7009 -1341
rect 7043 -1375 7060 -1341
rect 6986 -1413 7060 -1375
rect 6986 -1447 7009 -1413
rect 7043 -1447 7060 -1413
rect 6986 -1485 7060 -1447
rect 6986 -1519 7009 -1485
rect 7043 -1519 7060 -1485
rect 6986 -1557 7060 -1519
rect 7126 -1552 7808 -862
rect 7874 -871 7899 -837
rect 7933 -871 7948 -837
rect 7874 -909 7948 -871
rect 7874 -943 7899 -909
rect 7933 -943 7948 -909
rect 7874 -981 7948 -943
rect 7874 -1015 7899 -981
rect 7933 -1015 7948 -981
rect 7874 -1053 7948 -1015
rect 7874 -1087 7899 -1053
rect 7933 -1087 7948 -1053
rect 7874 -1125 7948 -1087
rect 7874 -1159 7899 -1125
rect 7933 -1159 7948 -1125
rect 7874 -1197 7948 -1159
rect 7874 -1231 7899 -1197
rect 7933 -1231 7948 -1197
rect 7874 -1269 7948 -1231
rect 7874 -1303 7899 -1269
rect 7933 -1303 7948 -1269
rect 7874 -1341 7948 -1303
rect 7874 -1375 7899 -1341
rect 7933 -1375 7948 -1341
rect 7874 -1413 7948 -1375
rect 7874 -1447 7899 -1413
rect 7933 -1447 7948 -1413
rect 7874 -1485 7948 -1447
rect 7874 -1519 7899 -1485
rect 7933 -1519 7948 -1485
rect 6986 -1591 7009 -1557
rect 7043 -1591 7060 -1557
rect 6986 -1622 7060 -1591
rect 7874 -1557 7948 -1519
rect 7874 -1591 7899 -1557
rect 7933 -1591 7948 -1557
rect 6820 -1672 6922 -1634
rect 6820 -1706 6859 -1672
rect 6893 -1706 6922 -1672
rect 6980 -1626 7066 -1622
rect 7874 -1626 7948 -1591
rect 8014 -808 8116 -770
rect 8014 -842 8045 -808
rect 8079 -842 8116 -808
rect 8014 -880 8116 -842
rect 8014 -914 8045 -880
rect 8079 -914 8116 -880
rect 8014 -952 8116 -914
rect 8014 -986 8045 -952
rect 8079 -986 8116 -952
rect 8014 -1024 8116 -986
rect 8014 -1058 8045 -1024
rect 8079 -1058 8116 -1024
rect 8014 -1096 8116 -1058
rect 8014 -1130 8045 -1096
rect 8079 -1130 8116 -1096
rect 8014 -1168 8116 -1130
rect 8014 -1202 8045 -1168
rect 8079 -1202 8116 -1168
rect 8014 -1240 8116 -1202
rect 8014 -1274 8045 -1240
rect 8079 -1274 8116 -1240
rect 8014 -1312 8116 -1274
rect 8014 -1346 8045 -1312
rect 8079 -1346 8116 -1312
rect 8014 -1384 8116 -1346
rect 8014 -1418 8045 -1384
rect 8079 -1418 8116 -1384
rect 8014 -1456 8116 -1418
rect 8014 -1490 8045 -1456
rect 8079 -1490 8116 -1456
rect 8014 -1528 8116 -1490
rect 8014 -1562 8045 -1528
rect 8079 -1562 8116 -1528
rect 8014 -1600 8116 -1562
rect 6980 -1643 7950 -1626
rect 6980 -1677 7009 -1643
rect 7043 -1677 7094 -1643
rect 7128 -1677 7166 -1643
rect 7200 -1677 7238 -1643
rect 7272 -1677 7310 -1643
rect 7344 -1677 7382 -1643
rect 7416 -1677 7454 -1643
rect 7488 -1677 7526 -1643
rect 7560 -1677 7598 -1643
rect 7632 -1677 7670 -1643
rect 7704 -1677 7742 -1643
rect 7776 -1677 7814 -1643
rect 7848 -1644 7950 -1643
rect 7848 -1677 7899 -1644
rect 6980 -1678 7899 -1677
rect 7933 -1678 7950 -1644
rect 6980 -1694 7950 -1678
rect 8014 -1634 8045 -1600
rect 8079 -1634 8116 -1600
rect 8014 -1672 8116 -1634
rect 6980 -1696 7066 -1694
rect 7874 -1698 7948 -1694
rect 6820 -1754 6922 -1706
rect 8014 -1706 8045 -1672
rect 8079 -1706 8116 -1672
rect 8014 -1754 8116 -1706
rect 5410 -1795 6708 -1758
rect 5410 -1829 5466 -1795
rect 5500 -1829 5538 -1795
rect 5572 -1829 5610 -1795
rect 5644 -1829 5682 -1795
rect 5716 -1829 5754 -1795
rect 5788 -1829 5826 -1795
rect 5860 -1829 5898 -1795
rect 5932 -1829 5970 -1795
rect 6004 -1829 6042 -1795
rect 6076 -1829 6114 -1795
rect 6148 -1829 6186 -1795
rect 6220 -1829 6258 -1795
rect 6292 -1829 6330 -1795
rect 6364 -1829 6402 -1795
rect 6436 -1829 6474 -1795
rect 6508 -1829 6546 -1795
rect 6580 -1829 6618 -1795
rect 6652 -1829 6708 -1795
rect 5410 -1838 6708 -1829
rect 6820 -1791 8118 -1754
rect 6820 -1825 6876 -1791
rect 6910 -1825 6948 -1791
rect 6982 -1825 7020 -1791
rect 7054 -1825 7092 -1791
rect 7126 -1825 7164 -1791
rect 7198 -1825 7236 -1791
rect 7270 -1825 7308 -1791
rect 7342 -1825 7380 -1791
rect 7414 -1825 7452 -1791
rect 7486 -1825 7524 -1791
rect 7558 -1825 7596 -1791
rect 7630 -1825 7668 -1791
rect 7702 -1825 7740 -1791
rect 7774 -1825 7812 -1791
rect 7846 -1825 7884 -1791
rect 7918 -1825 7956 -1791
rect 7990 -1825 8028 -1791
rect 8062 -1825 8118 -1791
rect 6820 -1834 8118 -1825
rect 5408 -1864 6708 -1838
rect 6818 -1860 8118 -1834
rect 5408 -1872 5500 -1864
rect 6818 -1868 6916 -1860
rect 5410 -1910 5500 -1872
rect 6820 -1908 6916 -1868
rect 6820 -1910 6918 -1908
rect 5408 -1924 5504 -1910
rect 6822 -1922 6918 -1910
rect 5408 -1977 6706 -1924
rect 5408 -2011 5464 -1977
rect 5498 -2011 5536 -1977
rect 5570 -2011 5608 -1977
rect 5642 -2011 5680 -1977
rect 5714 -2011 5752 -1977
rect 5786 -2011 5824 -1977
rect 5858 -2011 5896 -1977
rect 5930 -2011 5968 -1977
rect 6002 -2011 6040 -1977
rect 6074 -2011 6112 -1977
rect 6146 -2011 6184 -1977
rect 6218 -2011 6256 -1977
rect 6290 -2011 6328 -1977
rect 6362 -2011 6400 -1977
rect 6434 -2011 6472 -1977
rect 6506 -2011 6544 -1977
rect 6578 -2011 6616 -1977
rect 6650 -2011 6706 -1977
rect 5408 -2030 6706 -2011
rect 6822 -1975 8120 -1922
rect 6822 -2009 6878 -1975
rect 6912 -2009 6950 -1975
rect 6984 -2009 7022 -1975
rect 7056 -2009 7094 -1975
rect 7128 -2009 7166 -1975
rect 7200 -2009 7238 -1975
rect 7272 -2009 7310 -1975
rect 7344 -2009 7382 -1975
rect 7416 -2009 7454 -1975
rect 7488 -2009 7526 -1975
rect 7560 -2009 7598 -1975
rect 7632 -2009 7670 -1975
rect 7704 -2009 7742 -1975
rect 7776 -2009 7814 -1975
rect 7848 -2009 7886 -1975
rect 7920 -2009 7958 -1975
rect 7992 -2009 8030 -1975
rect 8064 -2009 8120 -1975
rect 6822 -2028 8120 -2009
rect 5408 -2096 5510 -2030
rect 5408 -2130 5447 -2096
rect 5481 -2130 5510 -2096
rect 5408 -2168 5510 -2130
rect 5574 -2111 6540 -2094
rect 5574 -2145 5607 -2111
rect 5641 -2145 5679 -2111
rect 5713 -2145 5751 -2111
rect 5785 -2145 5823 -2111
rect 5857 -2145 5895 -2111
rect 5929 -2145 5967 -2111
rect 6001 -2145 6039 -2111
rect 6073 -2145 6111 -2111
rect 6145 -2145 6183 -2111
rect 6217 -2145 6255 -2111
rect 6289 -2145 6327 -2111
rect 6361 -2145 6399 -2111
rect 6433 -2145 6540 -2111
rect 5574 -2154 6540 -2145
rect 5408 -2202 5447 -2168
rect 5481 -2202 5510 -2168
rect 5408 -2240 5510 -2202
rect 5572 -2162 6540 -2154
rect 6602 -2096 6704 -2030
rect 6602 -2130 6633 -2096
rect 6667 -2130 6704 -2096
rect 5572 -2197 5650 -2162
rect 5572 -2231 5597 -2197
rect 5631 -2231 5650 -2197
rect 6462 -2197 6536 -2162
rect 5572 -2234 5650 -2231
rect 5408 -2274 5447 -2240
rect 5481 -2274 5510 -2240
rect 5408 -2312 5510 -2274
rect 5408 -2346 5447 -2312
rect 5481 -2346 5510 -2312
rect 5408 -2384 5510 -2346
rect 5408 -2418 5447 -2384
rect 5481 -2418 5510 -2384
rect 5408 -2456 5510 -2418
rect 5408 -2490 5447 -2456
rect 5481 -2490 5510 -2456
rect 5408 -2528 5510 -2490
rect 5408 -2562 5447 -2528
rect 5481 -2562 5510 -2528
rect 5408 -2600 5510 -2562
rect 5408 -2634 5447 -2600
rect 5481 -2634 5510 -2600
rect 5408 -2672 5510 -2634
rect 5408 -2706 5447 -2672
rect 5481 -2706 5510 -2672
rect 5408 -2744 5510 -2706
rect 5408 -2778 5447 -2744
rect 5481 -2778 5510 -2744
rect 5408 -2816 5510 -2778
rect 5408 -2850 5447 -2816
rect 5481 -2850 5510 -2816
rect 5408 -2888 5510 -2850
rect 5408 -2922 5447 -2888
rect 5481 -2922 5510 -2888
rect 5408 -2960 5510 -2922
rect 5408 -2994 5447 -2960
rect 5481 -2994 5510 -2960
rect 5574 -2269 5648 -2234
rect 5574 -2303 5597 -2269
rect 5631 -2303 5648 -2269
rect 5574 -2341 5648 -2303
rect 5574 -2375 5597 -2341
rect 5631 -2375 5648 -2341
rect 5574 -2413 5648 -2375
rect 5574 -2447 5597 -2413
rect 5631 -2447 5648 -2413
rect 5574 -2485 5648 -2447
rect 5574 -2519 5597 -2485
rect 5631 -2519 5648 -2485
rect 5574 -2557 5648 -2519
rect 5574 -2591 5597 -2557
rect 5631 -2591 5648 -2557
rect 5574 -2629 5648 -2591
rect 5574 -2663 5597 -2629
rect 5631 -2663 5648 -2629
rect 5574 -2701 5648 -2663
rect 5574 -2735 5597 -2701
rect 5631 -2735 5648 -2701
rect 5574 -2773 5648 -2735
rect 5574 -2807 5597 -2773
rect 5631 -2807 5648 -2773
rect 5574 -2845 5648 -2807
rect 5574 -2879 5597 -2845
rect 5631 -2879 5648 -2845
rect 5574 -2917 5648 -2879
rect 5714 -2912 6396 -2222
rect 6462 -2231 6487 -2197
rect 6521 -2231 6536 -2197
rect 6462 -2269 6536 -2231
rect 6462 -2303 6487 -2269
rect 6521 -2303 6536 -2269
rect 6462 -2341 6536 -2303
rect 6462 -2375 6487 -2341
rect 6521 -2375 6536 -2341
rect 6462 -2413 6536 -2375
rect 6462 -2447 6487 -2413
rect 6521 -2447 6536 -2413
rect 6462 -2485 6536 -2447
rect 6462 -2519 6487 -2485
rect 6521 -2519 6536 -2485
rect 6462 -2557 6536 -2519
rect 6462 -2591 6487 -2557
rect 6521 -2591 6536 -2557
rect 6462 -2629 6536 -2591
rect 6462 -2663 6487 -2629
rect 6521 -2663 6536 -2629
rect 6462 -2701 6536 -2663
rect 6462 -2735 6487 -2701
rect 6521 -2735 6536 -2701
rect 6462 -2773 6536 -2735
rect 6462 -2807 6487 -2773
rect 6521 -2807 6536 -2773
rect 6462 -2845 6536 -2807
rect 6462 -2879 6487 -2845
rect 6521 -2879 6536 -2845
rect 5574 -2951 5597 -2917
rect 5631 -2951 5648 -2917
rect 5574 -2982 5648 -2951
rect 6462 -2917 6536 -2879
rect 6462 -2951 6487 -2917
rect 6521 -2951 6536 -2917
rect 5408 -3032 5510 -2994
rect 5408 -3066 5447 -3032
rect 5481 -3066 5510 -3032
rect 5568 -2986 5654 -2982
rect 6462 -2986 6536 -2951
rect 6602 -2168 6704 -2130
rect 6602 -2202 6633 -2168
rect 6667 -2202 6704 -2168
rect 6602 -2240 6704 -2202
rect 6602 -2274 6633 -2240
rect 6667 -2274 6704 -2240
rect 6602 -2312 6704 -2274
rect 6602 -2346 6633 -2312
rect 6667 -2346 6704 -2312
rect 6602 -2384 6704 -2346
rect 6602 -2418 6633 -2384
rect 6667 -2418 6704 -2384
rect 6602 -2456 6704 -2418
rect 6602 -2490 6633 -2456
rect 6667 -2490 6704 -2456
rect 6602 -2528 6704 -2490
rect 6602 -2562 6633 -2528
rect 6667 -2562 6704 -2528
rect 6602 -2600 6704 -2562
rect 6602 -2634 6633 -2600
rect 6667 -2634 6704 -2600
rect 6602 -2672 6704 -2634
rect 6602 -2706 6633 -2672
rect 6667 -2706 6704 -2672
rect 6602 -2744 6704 -2706
rect 6602 -2778 6633 -2744
rect 6667 -2778 6704 -2744
rect 6602 -2816 6704 -2778
rect 6602 -2850 6633 -2816
rect 6667 -2850 6704 -2816
rect 6602 -2888 6704 -2850
rect 6602 -2922 6633 -2888
rect 6667 -2922 6704 -2888
rect 6602 -2960 6704 -2922
rect 5568 -3003 6538 -2986
rect 5568 -3037 5597 -3003
rect 5631 -3037 5682 -3003
rect 5716 -3037 5754 -3003
rect 5788 -3037 5826 -3003
rect 5860 -3037 5898 -3003
rect 5932 -3037 5970 -3003
rect 6004 -3037 6042 -3003
rect 6076 -3037 6114 -3003
rect 6148 -3037 6186 -3003
rect 6220 -3037 6258 -3003
rect 6292 -3037 6330 -3003
rect 6364 -3037 6402 -3003
rect 6436 -3004 6538 -3003
rect 6436 -3037 6487 -3004
rect 5568 -3038 6487 -3037
rect 6521 -3038 6538 -3004
rect 5568 -3054 6538 -3038
rect 6602 -2994 6633 -2960
rect 6667 -2994 6704 -2960
rect 6602 -3032 6704 -2994
rect 5568 -3056 5654 -3054
rect 6462 -3058 6536 -3054
rect 5408 -3114 5510 -3066
rect 6602 -3066 6633 -3032
rect 6667 -3066 6704 -3032
rect 6602 -3114 6704 -3066
rect 6822 -2094 6924 -2028
rect 6822 -2128 6861 -2094
rect 6895 -2128 6924 -2094
rect 6822 -2166 6924 -2128
rect 6988 -2109 7954 -2092
rect 6988 -2143 7021 -2109
rect 7055 -2143 7093 -2109
rect 7127 -2143 7165 -2109
rect 7199 -2143 7237 -2109
rect 7271 -2143 7309 -2109
rect 7343 -2143 7381 -2109
rect 7415 -2143 7453 -2109
rect 7487 -2143 7525 -2109
rect 7559 -2143 7597 -2109
rect 7631 -2143 7669 -2109
rect 7703 -2143 7741 -2109
rect 7775 -2143 7813 -2109
rect 7847 -2143 7954 -2109
rect 6988 -2152 7954 -2143
rect 6822 -2200 6861 -2166
rect 6895 -2200 6924 -2166
rect 6822 -2238 6924 -2200
rect 6986 -2160 7954 -2152
rect 8016 -2094 8118 -2028
rect 8016 -2128 8047 -2094
rect 8081 -2128 8118 -2094
rect 6986 -2195 7064 -2160
rect 6986 -2229 7011 -2195
rect 7045 -2229 7064 -2195
rect 7876 -2195 7950 -2160
rect 6986 -2232 7064 -2229
rect 6822 -2272 6861 -2238
rect 6895 -2272 6924 -2238
rect 6822 -2310 6924 -2272
rect 6822 -2344 6861 -2310
rect 6895 -2344 6924 -2310
rect 6822 -2382 6924 -2344
rect 6822 -2416 6861 -2382
rect 6895 -2416 6924 -2382
rect 6822 -2454 6924 -2416
rect 6822 -2488 6861 -2454
rect 6895 -2488 6924 -2454
rect 6822 -2526 6924 -2488
rect 6822 -2560 6861 -2526
rect 6895 -2560 6924 -2526
rect 6822 -2598 6924 -2560
rect 6822 -2632 6861 -2598
rect 6895 -2632 6924 -2598
rect 6822 -2670 6924 -2632
rect 6822 -2704 6861 -2670
rect 6895 -2704 6924 -2670
rect 6822 -2742 6924 -2704
rect 6822 -2776 6861 -2742
rect 6895 -2776 6924 -2742
rect 6822 -2814 6924 -2776
rect 6822 -2848 6861 -2814
rect 6895 -2848 6924 -2814
rect 6822 -2886 6924 -2848
rect 6822 -2920 6861 -2886
rect 6895 -2920 6924 -2886
rect 6822 -2958 6924 -2920
rect 6822 -2992 6861 -2958
rect 6895 -2992 6924 -2958
rect 6988 -2267 7062 -2232
rect 6988 -2301 7011 -2267
rect 7045 -2301 7062 -2267
rect 6988 -2339 7062 -2301
rect 6988 -2373 7011 -2339
rect 7045 -2373 7062 -2339
rect 6988 -2411 7062 -2373
rect 6988 -2445 7011 -2411
rect 7045 -2445 7062 -2411
rect 6988 -2483 7062 -2445
rect 6988 -2517 7011 -2483
rect 7045 -2517 7062 -2483
rect 6988 -2555 7062 -2517
rect 6988 -2589 7011 -2555
rect 7045 -2589 7062 -2555
rect 6988 -2627 7062 -2589
rect 6988 -2661 7011 -2627
rect 7045 -2661 7062 -2627
rect 6988 -2699 7062 -2661
rect 6988 -2733 7011 -2699
rect 7045 -2733 7062 -2699
rect 6988 -2771 7062 -2733
rect 6988 -2805 7011 -2771
rect 7045 -2805 7062 -2771
rect 6988 -2843 7062 -2805
rect 6988 -2877 7011 -2843
rect 7045 -2877 7062 -2843
rect 6988 -2915 7062 -2877
rect 7128 -2910 7810 -2220
rect 7876 -2229 7901 -2195
rect 7935 -2229 7950 -2195
rect 7876 -2267 7950 -2229
rect 7876 -2301 7901 -2267
rect 7935 -2301 7950 -2267
rect 7876 -2339 7950 -2301
rect 7876 -2373 7901 -2339
rect 7935 -2373 7950 -2339
rect 7876 -2411 7950 -2373
rect 7876 -2445 7901 -2411
rect 7935 -2445 7950 -2411
rect 7876 -2483 7950 -2445
rect 7876 -2517 7901 -2483
rect 7935 -2517 7950 -2483
rect 7876 -2555 7950 -2517
rect 7876 -2589 7901 -2555
rect 7935 -2589 7950 -2555
rect 7876 -2627 7950 -2589
rect 7876 -2661 7901 -2627
rect 7935 -2661 7950 -2627
rect 7876 -2699 7950 -2661
rect 7876 -2733 7901 -2699
rect 7935 -2733 7950 -2699
rect 7876 -2771 7950 -2733
rect 7876 -2805 7901 -2771
rect 7935 -2805 7950 -2771
rect 7876 -2843 7950 -2805
rect 7876 -2877 7901 -2843
rect 7935 -2877 7950 -2843
rect 6988 -2949 7011 -2915
rect 7045 -2949 7062 -2915
rect 6988 -2980 7062 -2949
rect 7876 -2915 7950 -2877
rect 7876 -2949 7901 -2915
rect 7935 -2949 7950 -2915
rect 6822 -3030 6924 -2992
rect 6822 -3064 6861 -3030
rect 6895 -3064 6924 -3030
rect 6982 -2984 7068 -2980
rect 7876 -2984 7950 -2949
rect 8016 -2166 8118 -2128
rect 8016 -2200 8047 -2166
rect 8081 -2200 8118 -2166
rect 8016 -2238 8118 -2200
rect 8016 -2272 8047 -2238
rect 8081 -2272 8118 -2238
rect 8016 -2310 8118 -2272
rect 8016 -2344 8047 -2310
rect 8081 -2344 8118 -2310
rect 8016 -2382 8118 -2344
rect 8016 -2416 8047 -2382
rect 8081 -2416 8118 -2382
rect 8016 -2454 8118 -2416
rect 8016 -2488 8047 -2454
rect 8081 -2488 8118 -2454
rect 8016 -2526 8118 -2488
rect 8016 -2560 8047 -2526
rect 8081 -2560 8118 -2526
rect 8016 -2598 8118 -2560
rect 8016 -2632 8047 -2598
rect 8081 -2632 8118 -2598
rect 8016 -2670 8118 -2632
rect 8016 -2704 8047 -2670
rect 8081 -2704 8118 -2670
rect 8016 -2742 8118 -2704
rect 8016 -2776 8047 -2742
rect 8081 -2776 8118 -2742
rect 8016 -2814 8118 -2776
rect 8016 -2848 8047 -2814
rect 8081 -2848 8118 -2814
rect 8016 -2886 8118 -2848
rect 8016 -2920 8047 -2886
rect 8081 -2920 8118 -2886
rect 8016 -2958 8118 -2920
rect 6982 -3001 7952 -2984
rect 6982 -3035 7011 -3001
rect 7045 -3035 7096 -3001
rect 7130 -3035 7168 -3001
rect 7202 -3035 7240 -3001
rect 7274 -3035 7312 -3001
rect 7346 -3035 7384 -3001
rect 7418 -3035 7456 -3001
rect 7490 -3035 7528 -3001
rect 7562 -3035 7600 -3001
rect 7634 -3035 7672 -3001
rect 7706 -3035 7744 -3001
rect 7778 -3035 7816 -3001
rect 7850 -3002 7952 -3001
rect 7850 -3035 7901 -3002
rect 6982 -3036 7901 -3035
rect 7935 -3036 7952 -3002
rect 6982 -3052 7952 -3036
rect 8016 -2992 8047 -2958
rect 8081 -2992 8118 -2958
rect 8016 -3030 8118 -2992
rect 6982 -3054 7068 -3052
rect 7876 -3056 7950 -3052
rect 6822 -3112 6924 -3064
rect 8016 -3064 8047 -3030
rect 8081 -3064 8118 -3030
rect 8016 -3112 8118 -3064
rect 5408 -3151 6706 -3114
rect 5408 -3185 5464 -3151
rect 5498 -3185 5536 -3151
rect 5570 -3185 5608 -3151
rect 5642 -3185 5680 -3151
rect 5714 -3185 5752 -3151
rect 5786 -3185 5824 -3151
rect 5858 -3185 5896 -3151
rect 5930 -3185 5968 -3151
rect 6002 -3185 6040 -3151
rect 6074 -3185 6112 -3151
rect 6146 -3185 6184 -3151
rect 6218 -3185 6256 -3151
rect 6290 -3185 6328 -3151
rect 6362 -3185 6400 -3151
rect 6434 -3185 6472 -3151
rect 6506 -3185 6544 -3151
rect 6578 -3185 6616 -3151
rect 6650 -3185 6706 -3151
rect 5408 -3194 6706 -3185
rect 6822 -3149 8120 -3112
rect 6822 -3183 6878 -3149
rect 6912 -3183 6950 -3149
rect 6984 -3183 7022 -3149
rect 7056 -3183 7094 -3149
rect 7128 -3183 7166 -3149
rect 7200 -3183 7238 -3149
rect 7272 -3183 7310 -3149
rect 7344 -3183 7382 -3149
rect 7416 -3183 7454 -3149
rect 7488 -3183 7526 -3149
rect 7560 -3183 7598 -3149
rect 7632 -3183 7670 -3149
rect 7704 -3183 7742 -3149
rect 7776 -3183 7814 -3149
rect 7848 -3183 7886 -3149
rect 7920 -3183 7958 -3149
rect 7992 -3183 8030 -3149
rect 8064 -3183 8120 -3149
rect 6822 -3192 8120 -3183
rect 9230 -3150 9270 -2108
rect 10136 -2260 10316 -2204
rect 10280 -2384 10316 -2260
rect 10280 -2420 10526 -2384
rect 9912 -2844 9960 -2662
rect 9912 -2896 10150 -2844
rect 10128 -3072 10180 -2954
rect 10128 -3074 10182 -3072
rect 9986 -3118 10182 -3074
rect 9230 -3188 9628 -3150
rect 9230 -3190 9380 -3188
rect 5406 -3220 6706 -3194
rect 6820 -3218 8120 -3192
rect 5406 -3228 5498 -3220
rect 6820 -3226 6910 -3218
rect 5408 -3262 5498 -3228
rect 5408 -3276 5504 -3262
rect 6822 -3268 6910 -3226
rect 6822 -3272 6920 -3268
rect 5408 -3329 6706 -3276
rect 5408 -3363 5464 -3329
rect 5498 -3363 5536 -3329
rect 5570 -3363 5608 -3329
rect 5642 -3363 5680 -3329
rect 5714 -3363 5752 -3329
rect 5786 -3363 5824 -3329
rect 5858 -3363 5896 -3329
rect 5930 -3363 5968 -3329
rect 6002 -3363 6040 -3329
rect 6074 -3363 6112 -3329
rect 6146 -3363 6184 -3329
rect 6218 -3363 6256 -3329
rect 6290 -3363 6328 -3329
rect 6362 -3363 6400 -3329
rect 6434 -3363 6472 -3329
rect 6506 -3363 6544 -3329
rect 6578 -3363 6616 -3329
rect 6650 -3363 6706 -3329
rect 5408 -3382 6706 -3363
rect 6824 -3282 6920 -3272
rect 6824 -3335 8122 -3282
rect 6824 -3369 6880 -3335
rect 6914 -3369 6952 -3335
rect 6986 -3369 7024 -3335
rect 7058 -3369 7096 -3335
rect 7130 -3369 7168 -3335
rect 7202 -3369 7240 -3335
rect 7274 -3369 7312 -3335
rect 7346 -3369 7384 -3335
rect 7418 -3369 7456 -3335
rect 7490 -3369 7528 -3335
rect 7562 -3369 7600 -3335
rect 7634 -3369 7672 -3335
rect 7706 -3369 7744 -3335
rect 7778 -3369 7816 -3335
rect 7850 -3369 7888 -3335
rect 7922 -3369 7960 -3335
rect 7994 -3369 8032 -3335
rect 8066 -3369 8122 -3335
rect 5408 -3448 5510 -3382
rect 5408 -3482 5447 -3448
rect 5481 -3482 5510 -3448
rect 5408 -3520 5510 -3482
rect 5574 -3463 6540 -3446
rect 5574 -3497 5607 -3463
rect 5641 -3497 5679 -3463
rect 5713 -3497 5751 -3463
rect 5785 -3497 5823 -3463
rect 5857 -3497 5895 -3463
rect 5929 -3497 5967 -3463
rect 6001 -3497 6039 -3463
rect 6073 -3497 6111 -3463
rect 6145 -3497 6183 -3463
rect 6217 -3497 6255 -3463
rect 6289 -3497 6327 -3463
rect 6361 -3497 6399 -3463
rect 6433 -3497 6540 -3463
rect 5574 -3506 6540 -3497
rect 5408 -3554 5447 -3520
rect 5481 -3554 5510 -3520
rect 5408 -3592 5510 -3554
rect 5572 -3514 6540 -3506
rect 6602 -3448 6704 -3382
rect 6602 -3482 6633 -3448
rect 6667 -3482 6704 -3448
rect 5572 -3549 5650 -3514
rect 5572 -3583 5597 -3549
rect 5631 -3583 5650 -3549
rect 6462 -3549 6536 -3514
rect 5572 -3586 5650 -3583
rect 5408 -3626 5447 -3592
rect 5481 -3626 5510 -3592
rect 5408 -3664 5510 -3626
rect 5408 -3698 5447 -3664
rect 5481 -3698 5510 -3664
rect 5408 -3736 5510 -3698
rect 5408 -3770 5447 -3736
rect 5481 -3770 5510 -3736
rect 5408 -3808 5510 -3770
rect 5408 -3842 5447 -3808
rect 5481 -3842 5510 -3808
rect 5408 -3880 5510 -3842
rect 5408 -3914 5447 -3880
rect 5481 -3914 5510 -3880
rect 5408 -3952 5510 -3914
rect 5408 -3986 5447 -3952
rect 5481 -3986 5510 -3952
rect 5408 -4024 5510 -3986
rect 5408 -4058 5447 -4024
rect 5481 -4058 5510 -4024
rect 5408 -4096 5510 -4058
rect 5408 -4130 5447 -4096
rect 5481 -4130 5510 -4096
rect 5408 -4168 5510 -4130
rect 5408 -4202 5447 -4168
rect 5481 -4202 5510 -4168
rect 5408 -4240 5510 -4202
rect 5408 -4274 5447 -4240
rect 5481 -4274 5510 -4240
rect 5408 -4312 5510 -4274
rect 5408 -4346 5447 -4312
rect 5481 -4346 5510 -4312
rect 5574 -3621 5648 -3586
rect 5574 -3655 5597 -3621
rect 5631 -3655 5648 -3621
rect 5574 -3693 5648 -3655
rect 5574 -3727 5597 -3693
rect 5631 -3727 5648 -3693
rect 5574 -3765 5648 -3727
rect 5574 -3799 5597 -3765
rect 5631 -3799 5648 -3765
rect 5574 -3837 5648 -3799
rect 5574 -3871 5597 -3837
rect 5631 -3871 5648 -3837
rect 5574 -3909 5648 -3871
rect 5574 -3943 5597 -3909
rect 5631 -3943 5648 -3909
rect 5574 -3981 5648 -3943
rect 5574 -4015 5597 -3981
rect 5631 -4015 5648 -3981
rect 5574 -4053 5648 -4015
rect 5574 -4087 5597 -4053
rect 5631 -4087 5648 -4053
rect 5574 -4125 5648 -4087
rect 5574 -4159 5597 -4125
rect 5631 -4159 5648 -4125
rect 5574 -4197 5648 -4159
rect 5574 -4231 5597 -4197
rect 5631 -4231 5648 -4197
rect 5574 -4269 5648 -4231
rect 5714 -4264 6396 -3574
rect 6462 -3583 6487 -3549
rect 6521 -3583 6536 -3549
rect 6462 -3621 6536 -3583
rect 6462 -3655 6487 -3621
rect 6521 -3655 6536 -3621
rect 6462 -3693 6536 -3655
rect 6462 -3727 6487 -3693
rect 6521 -3727 6536 -3693
rect 6462 -3765 6536 -3727
rect 6462 -3799 6487 -3765
rect 6521 -3799 6536 -3765
rect 6462 -3837 6536 -3799
rect 6462 -3871 6487 -3837
rect 6521 -3871 6536 -3837
rect 6462 -3909 6536 -3871
rect 6462 -3943 6487 -3909
rect 6521 -3943 6536 -3909
rect 6462 -3981 6536 -3943
rect 6462 -4015 6487 -3981
rect 6521 -4015 6536 -3981
rect 6462 -4053 6536 -4015
rect 6462 -4087 6487 -4053
rect 6521 -4087 6536 -4053
rect 6462 -4125 6536 -4087
rect 6462 -4159 6487 -4125
rect 6521 -4159 6536 -4125
rect 6462 -4197 6536 -4159
rect 6462 -4231 6487 -4197
rect 6521 -4231 6536 -4197
rect 5574 -4303 5597 -4269
rect 5631 -4303 5648 -4269
rect 5574 -4334 5648 -4303
rect 6462 -4269 6536 -4231
rect 6462 -4303 6487 -4269
rect 6521 -4303 6536 -4269
rect 5408 -4384 5510 -4346
rect 5408 -4418 5447 -4384
rect 5481 -4418 5510 -4384
rect 5568 -4338 5654 -4334
rect 6462 -4338 6536 -4303
rect 6602 -3520 6704 -3482
rect 6602 -3554 6633 -3520
rect 6667 -3554 6704 -3520
rect 6602 -3592 6704 -3554
rect 6602 -3626 6633 -3592
rect 6667 -3626 6704 -3592
rect 6602 -3664 6704 -3626
rect 6602 -3698 6633 -3664
rect 6667 -3698 6704 -3664
rect 6602 -3736 6704 -3698
rect 6602 -3770 6633 -3736
rect 6667 -3770 6704 -3736
rect 6602 -3808 6704 -3770
rect 6602 -3842 6633 -3808
rect 6667 -3842 6704 -3808
rect 6602 -3880 6704 -3842
rect 6602 -3914 6633 -3880
rect 6667 -3914 6704 -3880
rect 6602 -3952 6704 -3914
rect 6602 -3986 6633 -3952
rect 6667 -3986 6704 -3952
rect 6602 -4024 6704 -3986
rect 6602 -4058 6633 -4024
rect 6667 -4058 6704 -4024
rect 6602 -4096 6704 -4058
rect 6602 -4130 6633 -4096
rect 6667 -4130 6704 -4096
rect 6602 -4168 6704 -4130
rect 6602 -4202 6633 -4168
rect 6667 -4202 6704 -4168
rect 6602 -4240 6704 -4202
rect 6602 -4274 6633 -4240
rect 6667 -4274 6704 -4240
rect 6602 -4312 6704 -4274
rect 5568 -4355 6538 -4338
rect 5568 -4389 5597 -4355
rect 5631 -4389 5682 -4355
rect 5716 -4389 5754 -4355
rect 5788 -4389 5826 -4355
rect 5860 -4389 5898 -4355
rect 5932 -4389 5970 -4355
rect 6004 -4389 6042 -4355
rect 6076 -4389 6114 -4355
rect 6148 -4389 6186 -4355
rect 6220 -4389 6258 -4355
rect 6292 -4389 6330 -4355
rect 6364 -4389 6402 -4355
rect 6436 -4356 6538 -4355
rect 6436 -4389 6487 -4356
rect 5568 -4390 6487 -4389
rect 6521 -4390 6538 -4356
rect 5568 -4406 6538 -4390
rect 6602 -4346 6633 -4312
rect 6667 -4346 6704 -4312
rect 6602 -4384 6704 -4346
rect 5568 -4408 5654 -4406
rect 6462 -4410 6536 -4406
rect 5408 -4466 5510 -4418
rect 6602 -4418 6633 -4384
rect 6667 -4418 6704 -4384
rect 6602 -4466 6704 -4418
rect 6824 -3388 8122 -3369
rect 6824 -3454 6926 -3388
rect 6824 -3488 6863 -3454
rect 6897 -3488 6926 -3454
rect 6824 -3526 6926 -3488
rect 6990 -3469 7956 -3452
rect 6990 -3503 7023 -3469
rect 7057 -3503 7095 -3469
rect 7129 -3503 7167 -3469
rect 7201 -3503 7239 -3469
rect 7273 -3503 7311 -3469
rect 7345 -3503 7383 -3469
rect 7417 -3503 7455 -3469
rect 7489 -3503 7527 -3469
rect 7561 -3503 7599 -3469
rect 7633 -3503 7671 -3469
rect 7705 -3503 7743 -3469
rect 7777 -3503 7815 -3469
rect 7849 -3503 7956 -3469
rect 6990 -3512 7956 -3503
rect 6824 -3560 6863 -3526
rect 6897 -3560 6926 -3526
rect 6824 -3598 6926 -3560
rect 6988 -3520 7956 -3512
rect 8018 -3454 8120 -3388
rect 8018 -3488 8049 -3454
rect 8083 -3488 8120 -3454
rect 6988 -3555 7066 -3520
rect 6988 -3589 7013 -3555
rect 7047 -3589 7066 -3555
rect 7878 -3555 7952 -3520
rect 6988 -3592 7066 -3589
rect 6824 -3632 6863 -3598
rect 6897 -3632 6926 -3598
rect 6824 -3670 6926 -3632
rect 6824 -3704 6863 -3670
rect 6897 -3704 6926 -3670
rect 6824 -3742 6926 -3704
rect 6824 -3776 6863 -3742
rect 6897 -3776 6926 -3742
rect 6824 -3814 6926 -3776
rect 6824 -3848 6863 -3814
rect 6897 -3848 6926 -3814
rect 6824 -3886 6926 -3848
rect 6824 -3920 6863 -3886
rect 6897 -3920 6926 -3886
rect 6824 -3958 6926 -3920
rect 6824 -3992 6863 -3958
rect 6897 -3992 6926 -3958
rect 6824 -4030 6926 -3992
rect 6824 -4064 6863 -4030
rect 6897 -4064 6926 -4030
rect 6824 -4102 6926 -4064
rect 6824 -4136 6863 -4102
rect 6897 -4136 6926 -4102
rect 6824 -4174 6926 -4136
rect 6824 -4208 6863 -4174
rect 6897 -4208 6926 -4174
rect 6824 -4246 6926 -4208
rect 6824 -4280 6863 -4246
rect 6897 -4280 6926 -4246
rect 6824 -4318 6926 -4280
rect 6824 -4352 6863 -4318
rect 6897 -4352 6926 -4318
rect 6990 -3627 7064 -3592
rect 6990 -3661 7013 -3627
rect 7047 -3661 7064 -3627
rect 6990 -3699 7064 -3661
rect 6990 -3733 7013 -3699
rect 7047 -3733 7064 -3699
rect 6990 -3771 7064 -3733
rect 6990 -3805 7013 -3771
rect 7047 -3805 7064 -3771
rect 6990 -3843 7064 -3805
rect 6990 -3877 7013 -3843
rect 7047 -3877 7064 -3843
rect 6990 -3915 7064 -3877
rect 6990 -3949 7013 -3915
rect 7047 -3949 7064 -3915
rect 6990 -3987 7064 -3949
rect 6990 -4021 7013 -3987
rect 7047 -4021 7064 -3987
rect 6990 -4059 7064 -4021
rect 6990 -4093 7013 -4059
rect 7047 -4093 7064 -4059
rect 6990 -4131 7064 -4093
rect 6990 -4165 7013 -4131
rect 7047 -4165 7064 -4131
rect 6990 -4203 7064 -4165
rect 6990 -4237 7013 -4203
rect 7047 -4237 7064 -4203
rect 6990 -4275 7064 -4237
rect 7130 -4270 7812 -3580
rect 7878 -3589 7903 -3555
rect 7937 -3589 7952 -3555
rect 7878 -3627 7952 -3589
rect 7878 -3661 7903 -3627
rect 7937 -3661 7952 -3627
rect 7878 -3699 7952 -3661
rect 7878 -3733 7903 -3699
rect 7937 -3733 7952 -3699
rect 7878 -3771 7952 -3733
rect 7878 -3805 7903 -3771
rect 7937 -3805 7952 -3771
rect 7878 -3843 7952 -3805
rect 7878 -3877 7903 -3843
rect 7937 -3877 7952 -3843
rect 7878 -3915 7952 -3877
rect 7878 -3949 7903 -3915
rect 7937 -3949 7952 -3915
rect 7878 -3987 7952 -3949
rect 7878 -4021 7903 -3987
rect 7937 -4021 7952 -3987
rect 7878 -4059 7952 -4021
rect 7878 -4093 7903 -4059
rect 7937 -4093 7952 -4059
rect 7878 -4131 7952 -4093
rect 7878 -4165 7903 -4131
rect 7937 -4165 7952 -4131
rect 7878 -4203 7952 -4165
rect 7878 -4237 7903 -4203
rect 7937 -4237 7952 -4203
rect 6990 -4309 7013 -4275
rect 7047 -4309 7064 -4275
rect 6990 -4340 7064 -4309
rect 7878 -4275 7952 -4237
rect 7878 -4309 7903 -4275
rect 7937 -4309 7952 -4275
rect 6824 -4390 6926 -4352
rect 6824 -4424 6863 -4390
rect 6897 -4424 6926 -4390
rect 6984 -4344 7070 -4340
rect 7878 -4344 7952 -4309
rect 8018 -3526 8120 -3488
rect 8018 -3560 8049 -3526
rect 8083 -3560 8120 -3526
rect 8018 -3598 8120 -3560
rect 8018 -3632 8049 -3598
rect 8083 -3632 8120 -3598
rect 8018 -3670 8120 -3632
rect 8018 -3704 8049 -3670
rect 8083 -3704 8120 -3670
rect 8018 -3742 8120 -3704
rect 8018 -3776 8049 -3742
rect 8083 -3776 8120 -3742
rect 8018 -3814 8120 -3776
rect 8018 -3848 8049 -3814
rect 8083 -3848 8120 -3814
rect 8018 -3886 8120 -3848
rect 8018 -3920 8049 -3886
rect 8083 -3920 8120 -3886
rect 8018 -3958 8120 -3920
rect 8018 -3992 8049 -3958
rect 8083 -3992 8120 -3958
rect 8018 -4030 8120 -3992
rect 8018 -4064 8049 -4030
rect 8083 -4064 8120 -4030
rect 8018 -4102 8120 -4064
rect 8018 -4136 8049 -4102
rect 8083 -4136 8120 -4102
rect 8018 -4174 8120 -4136
rect 8018 -4208 8049 -4174
rect 8083 -4208 8120 -4174
rect 8018 -4246 8120 -4208
rect 8018 -4280 8049 -4246
rect 8083 -4280 8120 -4246
rect 8018 -4318 8120 -4280
rect 6984 -4361 7954 -4344
rect 6984 -4395 7013 -4361
rect 7047 -4395 7098 -4361
rect 7132 -4395 7170 -4361
rect 7204 -4395 7242 -4361
rect 7276 -4395 7314 -4361
rect 7348 -4395 7386 -4361
rect 7420 -4395 7458 -4361
rect 7492 -4395 7530 -4361
rect 7564 -4395 7602 -4361
rect 7636 -4395 7674 -4361
rect 7708 -4395 7746 -4361
rect 7780 -4395 7818 -4361
rect 7852 -4362 7954 -4361
rect 7852 -4395 7903 -4362
rect 6984 -4396 7903 -4395
rect 7937 -4396 7954 -4362
rect 6984 -4412 7954 -4396
rect 8018 -4352 8049 -4318
rect 8083 -4352 8120 -4318
rect 8018 -4390 8120 -4352
rect 6984 -4414 7070 -4412
rect 7878 -4416 7952 -4412
rect 5408 -4503 6706 -4466
rect 5408 -4537 5464 -4503
rect 5498 -4537 5536 -4503
rect 5570 -4537 5608 -4503
rect 5642 -4537 5680 -4503
rect 5714 -4537 5752 -4503
rect 5786 -4537 5824 -4503
rect 5858 -4537 5896 -4503
rect 5930 -4537 5968 -4503
rect 6002 -4537 6040 -4503
rect 6074 -4537 6112 -4503
rect 6146 -4537 6184 -4503
rect 6218 -4537 6256 -4503
rect 6290 -4537 6328 -4503
rect 6362 -4537 6400 -4503
rect 6434 -4537 6472 -4503
rect 6506 -4537 6544 -4503
rect 6578 -4537 6616 -4503
rect 6650 -4537 6706 -4503
rect 5408 -4546 6706 -4537
rect 5406 -4562 6706 -4546
rect 6824 -4472 6926 -4424
rect 8018 -4424 8049 -4390
rect 8083 -4424 8120 -4390
rect 8018 -4472 8120 -4424
rect 8702 -3962 8944 -3894
rect 6824 -4509 8122 -4472
rect 6824 -4543 6880 -4509
rect 6914 -4543 6952 -4509
rect 6986 -4543 7024 -4509
rect 7058 -4543 7096 -4509
rect 7130 -4543 7168 -4509
rect 7202 -4543 7240 -4509
rect 7274 -4543 7312 -4509
rect 7346 -4543 7384 -4509
rect 7418 -4543 7456 -4509
rect 7490 -4543 7528 -4509
rect 7562 -4543 7600 -4509
rect 7634 -4543 7672 -4509
rect 7706 -4543 7744 -4509
rect 7778 -4543 7816 -4509
rect 7850 -4543 7888 -4509
rect 7922 -4543 7960 -4509
rect 7994 -4543 8032 -4509
rect 8066 -4543 8122 -4509
rect 6824 -4552 8122 -4543
rect 5404 -4572 6706 -4562
rect 6822 -4572 8122 -4552
rect 5404 -4980 5496 -4572
rect 6818 -4578 8122 -4572
rect 6818 -4586 6912 -4578
rect 6818 -4980 6910 -4586
rect 8702 -4950 8756 -3962
rect 8702 -4980 8758 -4950
rect 9566 -4978 9628 -3188
rect 9986 -4950 10040 -3118
rect 10862 -3556 10916 34
rect 13390 -1124 13448 -1120
rect 12428 -2010 12486 -1162
rect 13382 -1956 13448 -1124
rect 14172 -1580 14238 -1174
rect 14048 -1660 14238 -1580
rect 14048 -1668 14110 -1660
rect 13382 -1984 13450 -1956
rect 11610 -2454 12216 -2390
rect 10860 -3620 11304 -3556
rect 9984 -4978 10042 -4950
rect 11246 -4978 11304 -3620
rect 11610 -3756 11676 -2454
rect 12430 -3552 12482 -2010
rect 13384 -2424 13450 -1984
rect 13158 -2494 13452 -2424
rect 11396 -3802 11676 -3756
rect 12214 -3594 12482 -3552
rect 13132 -3560 13186 -2606
rect 13922 -3560 13970 -2278
rect 12916 -3594 13186 -3560
rect 13706 -3594 13970 -3560
rect 14050 -3586 14110 -1668
rect 14048 -3594 14110 -3586
rect 11396 -4950 11460 -3802
rect 11394 -4978 11460 -4950
rect 12214 -4950 12262 -3594
rect 12916 -4950 12968 -3594
rect 12214 -4978 12266 -4950
rect 12916 -4978 12970 -4950
rect 13706 -4978 13754 -3594
rect 14048 -3730 14108 -3594
rect 13834 -3778 14108 -3730
rect 13834 -4978 13894 -3778
rect 9382 -4980 10288 -4978
rect 11246 -4980 11742 -4978
rect 12184 -4980 14022 -4978
rect -2110 -5005 14022 -4980
rect -2110 -5008 11122 -5005
rect -2110 -5009 9452 -5008
rect -2110 -5010 8385 -5009
rect -2110 -5180 -2079 -5010
rect -1841 -5011 1803 -5010
rect -1841 -5020 -1174 -5011
rect -1841 -5180 -1635 -5020
rect -2110 -5190 -1635 -5180
rect -1261 -5181 -1174 -5020
rect -868 -5180 1803 -5011
rect 2109 -5011 6663 -5010
rect 2109 -5015 5301 -5011
rect 2109 -5180 2193 -5015
rect 2499 -5038 5301 -5015
rect -868 -5181 2193 -5180
rect -1261 -5185 2193 -5181
rect 2499 -5140 4546 -5038
rect 5056 -5140 5301 -5038
rect 2499 -5181 5301 -5140
rect 5879 -5180 6663 -5011
rect 7241 -5179 8385 -5010
rect 9235 -5178 9452 -5009
rect 10166 -5175 11122 -5008
rect 11496 -5009 14022 -5005
rect 11496 -5175 12224 -5009
rect 10166 -5178 12224 -5175
rect 9235 -5179 12224 -5178
rect 12666 -5011 13632 -5009
rect 12666 -5179 12833 -5011
rect 7241 -5180 12833 -5179
rect 5879 -5181 12833 -5180
rect 13207 -5179 13632 -5011
rect 13938 -5179 14022 -5009
rect 13207 -5181 14022 -5179
rect 2499 -5185 14022 -5181
rect -1261 -5190 14022 -5185
rect -2110 -5206 14022 -5190
rect -2110 -5208 -1088 -5206
rect 6644 -5208 7260 -5206
<< viali >>
rect 6876 2069 6910 2103
rect 6948 2069 6982 2103
rect 7020 2069 7054 2103
rect 7092 2069 7126 2103
rect 7164 2069 7198 2103
rect 7236 2069 7270 2103
rect 7308 2069 7342 2103
rect 7380 2069 7414 2103
rect 7452 2069 7486 2103
rect 7524 2069 7558 2103
rect 7596 2069 7630 2103
rect 7668 2069 7702 2103
rect 7740 2069 7774 2103
rect 7812 2069 7846 2103
rect 7884 2069 7918 2103
rect 7956 2069 7990 2103
rect 8028 2069 8062 2103
rect 6859 1950 6893 1984
rect 7019 1935 7053 1969
rect 7091 1935 7125 1969
rect 7163 1935 7197 1969
rect 7235 1935 7269 1969
rect 7307 1935 7341 1969
rect 7379 1935 7413 1969
rect 7451 1935 7485 1969
rect 7523 1935 7557 1969
rect 7595 1935 7629 1969
rect 7667 1935 7701 1969
rect 7739 1935 7773 1969
rect 7811 1935 7845 1969
rect 6859 1878 6893 1912
rect 8045 1950 8079 1984
rect 7009 1849 7043 1883
rect 6859 1806 6893 1840
rect 6859 1734 6893 1768
rect 6859 1662 6893 1696
rect 6859 1590 6893 1624
rect 6859 1518 6893 1552
rect 6859 1446 6893 1480
rect 1911 448 1945 482
rect 1983 448 2017 482
rect 2055 448 2089 482
rect 2127 448 2161 482
rect 2199 448 2233 482
rect 2271 448 2305 482
rect 2343 448 2377 482
rect 2415 448 2449 482
rect 2487 448 2521 482
rect 2559 448 2593 482
rect 2631 448 2665 482
rect 2703 448 2737 482
rect 2775 448 2809 482
rect 2847 448 2881 482
rect 2919 448 2953 482
rect 2991 448 3025 482
rect 3063 448 3097 482
rect 1892 329 1926 363
rect 2053 315 2087 349
rect 2125 315 2159 349
rect 2197 315 2231 349
rect 2269 315 2303 349
rect 2341 315 2375 349
rect 2413 315 2447 349
rect 2485 315 2519 349
rect 2557 315 2591 349
rect 2629 315 2663 349
rect 2701 315 2735 349
rect 2773 315 2807 349
rect 2845 315 2879 349
rect 2917 315 2951 349
rect 1892 257 1926 291
rect 1892 185 1926 219
rect 1892 113 1926 147
rect 1892 41 1926 75
rect 1892 -31 1926 3
rect 1892 -103 1926 -69
rect 1892 -175 1926 -141
rect 1892 -247 1926 -213
rect 1892 -319 1926 -285
rect 1892 -391 1926 -357
rect 1892 -463 1926 -429
rect 1892 -535 1926 -501
rect 2042 229 2076 263
rect 2042 157 2076 191
rect 2042 85 2076 119
rect 2042 13 2076 47
rect 2042 -59 2076 -25
rect 2042 -131 2076 -97
rect 2042 -203 2076 -169
rect 2042 -275 2076 -241
rect 2042 -347 2076 -313
rect 2042 -419 2076 -385
rect 2042 -491 2076 -457
rect 2932 229 2966 263
rect 2932 157 2966 191
rect 2932 85 2966 119
rect 2932 13 2966 47
rect 2932 -59 2966 -25
rect 2932 -131 2966 -97
rect 2932 -203 2966 -169
rect 2932 -275 2966 -241
rect 2932 -347 2966 -313
rect 2932 -419 2966 -385
rect 2932 -491 2966 -457
rect 1892 -607 1926 -573
rect 2042 -577 2076 -543
rect 2127 -577 2161 -543
rect 2199 -577 2233 -543
rect 2271 -577 2305 -543
rect 2343 -577 2377 -543
rect 2415 -577 2449 -543
rect 2487 -577 2521 -543
rect 2559 -577 2593 -543
rect 2631 -577 2665 -543
rect 2703 -577 2737 -543
rect 2775 -577 2809 -543
rect 2847 -577 2881 -543
rect 2932 -577 2966 -543
rect 3082 329 3116 363
rect 3082 257 3116 291
rect 3082 185 3116 219
rect 3082 113 3116 147
rect 3082 41 3116 75
rect 3082 -31 3116 3
rect 3082 -103 3116 -69
rect 3082 -175 3116 -141
rect 3082 -247 3116 -213
rect 3082 -319 3116 -285
rect 3082 -391 3116 -357
rect 3082 -463 3116 -429
rect 3082 -535 3116 -501
rect 3082 -607 3116 -573
rect 1911 -726 1945 -692
rect 1983 -726 2017 -692
rect 2055 -726 2089 -692
rect 2127 -726 2161 -692
rect 2199 -726 2233 -692
rect 2271 -726 2305 -692
rect 2343 -726 2377 -692
rect 2415 -726 2449 -692
rect 2487 -726 2521 -692
rect 2559 -726 2593 -692
rect 2631 -726 2665 -692
rect 2703 -726 2737 -692
rect 2775 -726 2809 -692
rect 2847 -726 2881 -692
rect 2919 -726 2953 -692
rect 2991 -726 3025 -692
rect 3063 -726 3097 -692
rect 6859 1374 6893 1408
rect 6859 1302 6893 1336
rect 6859 1230 6893 1264
rect 6859 1158 6893 1192
rect 6859 1086 6893 1120
rect 7009 1777 7043 1811
rect 7009 1705 7043 1739
rect 7009 1633 7043 1667
rect 7009 1561 7043 1595
rect 7009 1489 7043 1523
rect 7009 1417 7043 1451
rect 7009 1345 7043 1379
rect 7009 1273 7043 1307
rect 7009 1201 7043 1235
rect 7899 1849 7933 1883
rect 7899 1777 7933 1811
rect 7899 1705 7933 1739
rect 7899 1633 7933 1667
rect 7899 1561 7933 1595
rect 7899 1489 7933 1523
rect 7899 1417 7933 1451
rect 7899 1345 7933 1379
rect 7899 1273 7933 1307
rect 7899 1201 7933 1235
rect 7009 1129 7043 1163
rect 7899 1129 7933 1163
rect 6859 1014 6893 1048
rect 8045 1878 8079 1912
rect 8045 1806 8079 1840
rect 8045 1734 8079 1768
rect 8045 1662 8079 1696
rect 8045 1590 8079 1624
rect 8045 1518 8079 1552
rect 8045 1446 8079 1480
rect 8045 1374 8079 1408
rect 8045 1302 8079 1336
rect 8045 1230 8079 1264
rect 8045 1158 8079 1192
rect 7009 1043 7043 1077
rect 7094 1043 7128 1077
rect 7166 1043 7200 1077
rect 7238 1043 7272 1077
rect 7310 1043 7344 1077
rect 7382 1043 7416 1077
rect 7454 1043 7488 1077
rect 7526 1043 7560 1077
rect 7598 1043 7632 1077
rect 7670 1043 7704 1077
rect 7742 1043 7776 1077
rect 7814 1043 7848 1077
rect 7899 1042 7933 1076
rect 8045 1086 8079 1120
rect 8045 1014 8079 1048
rect 6876 895 6910 929
rect 6948 895 6982 929
rect 7020 895 7054 929
rect 7092 895 7126 929
rect 7164 895 7198 929
rect 7236 895 7270 929
rect 7308 895 7342 929
rect 7380 895 7414 929
rect 7452 895 7486 929
rect 7524 895 7558 929
rect 7596 895 7630 929
rect 7668 895 7702 929
rect 7740 895 7774 929
rect 7812 895 7846 929
rect 7884 895 7918 929
rect 7956 895 7990 929
rect 8028 895 8062 929
rect 6880 713 6914 747
rect 6952 713 6986 747
rect 7024 713 7058 747
rect 7096 713 7130 747
rect 7168 713 7202 747
rect 7240 713 7274 747
rect 7312 713 7346 747
rect 7384 713 7418 747
rect 7456 713 7490 747
rect 7528 713 7562 747
rect 7600 713 7634 747
rect 7672 713 7706 747
rect 7744 713 7778 747
rect 7816 713 7850 747
rect 7888 713 7922 747
rect 7960 713 7994 747
rect 8032 713 8066 747
rect 6863 594 6897 628
rect 7023 579 7057 613
rect 7095 579 7129 613
rect 7167 579 7201 613
rect 7239 579 7273 613
rect 7311 579 7345 613
rect 7383 579 7417 613
rect 7455 579 7489 613
rect 7527 579 7561 613
rect 7599 579 7633 613
rect 7671 579 7705 613
rect 7743 579 7777 613
rect 7815 579 7849 613
rect 6863 522 6897 556
rect 8049 594 8083 628
rect 7013 493 7047 527
rect 6863 450 6897 484
rect 6863 378 6897 412
rect 6863 306 6897 340
rect 6863 234 6897 268
rect 6863 162 6897 196
rect 6863 90 6897 124
rect 6863 18 6897 52
rect 6863 -54 6897 -20
rect 6863 -126 6897 -92
rect 6863 -198 6897 -164
rect 6863 -270 6897 -236
rect 7013 421 7047 455
rect 7013 349 7047 383
rect 7013 277 7047 311
rect 7013 205 7047 239
rect 7013 133 7047 167
rect 7013 61 7047 95
rect 7013 -11 7047 23
rect 7013 -83 7047 -49
rect 7013 -155 7047 -121
rect 7903 493 7937 527
rect 7903 421 7937 455
rect 7903 349 7937 383
rect 7903 277 7937 311
rect 7903 205 7937 239
rect 7903 133 7937 167
rect 7903 61 7937 95
rect 7903 -11 7937 23
rect 7903 -83 7937 -49
rect 7903 -155 7937 -121
rect 7013 -227 7047 -193
rect 7903 -227 7937 -193
rect 6863 -342 6897 -308
rect 8049 522 8083 556
rect 8049 450 8083 484
rect 8049 378 8083 412
rect 8049 306 8083 340
rect 8049 234 8083 268
rect 8049 162 8083 196
rect 8049 90 8083 124
rect 8049 18 8083 52
rect 8049 -54 8083 -20
rect 8049 -126 8083 -92
rect 8049 -198 8083 -164
rect 7013 -313 7047 -279
rect 7098 -313 7132 -279
rect 7170 -313 7204 -279
rect 7242 -313 7276 -279
rect 7314 -313 7348 -279
rect 7386 -313 7420 -279
rect 7458 -313 7492 -279
rect 7530 -313 7564 -279
rect 7602 -313 7636 -279
rect 7674 -313 7708 -279
rect 7746 -313 7780 -279
rect 7818 -313 7852 -279
rect 7903 -314 7937 -280
rect 8049 -270 8083 -236
rect 8049 -342 8083 -308
rect 6880 -461 6914 -427
rect 6952 -461 6986 -427
rect 7024 -461 7058 -427
rect 7096 -461 7130 -427
rect 7168 -461 7202 -427
rect 7240 -461 7274 -427
rect 7312 -461 7346 -427
rect 7384 -461 7418 -427
rect 7456 -461 7490 -427
rect 7528 -461 7562 -427
rect 7600 -461 7634 -427
rect 7672 -461 7706 -427
rect 7744 -461 7778 -427
rect 7816 -461 7850 -427
rect 7888 -461 7922 -427
rect 7960 -461 7994 -427
rect 8032 -461 8066 -427
rect 5466 -655 5500 -621
rect 5538 -655 5572 -621
rect 5610 -655 5644 -621
rect 5682 -655 5716 -621
rect 5754 -655 5788 -621
rect 5826 -655 5860 -621
rect 5898 -655 5932 -621
rect 5970 -655 6004 -621
rect 6042 -655 6076 -621
rect 6114 -655 6148 -621
rect 6186 -655 6220 -621
rect 6258 -655 6292 -621
rect 6330 -655 6364 -621
rect 6402 -655 6436 -621
rect 6474 -655 6508 -621
rect 6546 -655 6580 -621
rect 6618 -655 6652 -621
rect 6876 -651 6910 -617
rect 6948 -651 6982 -617
rect 7020 -651 7054 -617
rect 7092 -651 7126 -617
rect 7164 -651 7198 -617
rect 7236 -651 7270 -617
rect 7308 -651 7342 -617
rect 7380 -651 7414 -617
rect 7452 -651 7486 -617
rect 7524 -651 7558 -617
rect 7596 -651 7630 -617
rect 7668 -651 7702 -617
rect 7740 -651 7774 -617
rect 7812 -651 7846 -617
rect 7884 -651 7918 -617
rect 7956 -651 7990 -617
rect 8028 -651 8062 -617
rect 5449 -774 5483 -740
rect 5609 -789 5643 -755
rect 5681 -789 5715 -755
rect 5753 -789 5787 -755
rect 5825 -789 5859 -755
rect 5897 -789 5931 -755
rect 5969 -789 6003 -755
rect 6041 -789 6075 -755
rect 6113 -789 6147 -755
rect 6185 -789 6219 -755
rect 6257 -789 6291 -755
rect 6329 -789 6363 -755
rect 6401 -789 6435 -755
rect 5449 -846 5483 -812
rect 6635 -774 6669 -740
rect 5599 -875 5633 -841
rect 5449 -918 5483 -884
rect 5449 -990 5483 -956
rect 5449 -1062 5483 -1028
rect 5449 -1134 5483 -1100
rect 5449 -1206 5483 -1172
rect 5449 -1278 5483 -1244
rect 5449 -1350 5483 -1316
rect 5449 -1422 5483 -1388
rect 5449 -1494 5483 -1460
rect 5449 -1566 5483 -1532
rect 5449 -1638 5483 -1604
rect 5599 -947 5633 -913
rect 5599 -1019 5633 -985
rect 5599 -1091 5633 -1057
rect 5599 -1163 5633 -1129
rect 5599 -1235 5633 -1201
rect 5599 -1307 5633 -1273
rect 5599 -1379 5633 -1345
rect 5599 -1451 5633 -1417
rect 5599 -1523 5633 -1489
rect 6489 -875 6523 -841
rect 6489 -947 6523 -913
rect 6489 -1019 6523 -985
rect 6489 -1091 6523 -1057
rect 6489 -1163 6523 -1129
rect 6489 -1235 6523 -1201
rect 6489 -1307 6523 -1273
rect 6489 -1379 6523 -1345
rect 6489 -1451 6523 -1417
rect 6489 -1523 6523 -1489
rect 5599 -1595 5633 -1561
rect 6489 -1595 6523 -1561
rect 5449 -1710 5483 -1676
rect 6635 -846 6669 -812
rect 6635 -918 6669 -884
rect 6635 -990 6669 -956
rect 6635 -1062 6669 -1028
rect 6635 -1134 6669 -1100
rect 6635 -1206 6669 -1172
rect 6635 -1278 6669 -1244
rect 6635 -1350 6669 -1316
rect 6635 -1422 6669 -1388
rect 6635 -1494 6669 -1460
rect 6635 -1566 6669 -1532
rect 5599 -1681 5633 -1647
rect 5684 -1681 5718 -1647
rect 5756 -1681 5790 -1647
rect 5828 -1681 5862 -1647
rect 5900 -1681 5934 -1647
rect 5972 -1681 6006 -1647
rect 6044 -1681 6078 -1647
rect 6116 -1681 6150 -1647
rect 6188 -1681 6222 -1647
rect 6260 -1681 6294 -1647
rect 6332 -1681 6366 -1647
rect 6404 -1681 6438 -1647
rect 6489 -1682 6523 -1648
rect 6635 -1638 6669 -1604
rect 6635 -1710 6669 -1676
rect 6859 -770 6893 -736
rect 7019 -785 7053 -751
rect 7091 -785 7125 -751
rect 7163 -785 7197 -751
rect 7235 -785 7269 -751
rect 7307 -785 7341 -751
rect 7379 -785 7413 -751
rect 7451 -785 7485 -751
rect 7523 -785 7557 -751
rect 7595 -785 7629 -751
rect 7667 -785 7701 -751
rect 7739 -785 7773 -751
rect 7811 -785 7845 -751
rect 6859 -842 6893 -808
rect 8045 -770 8079 -736
rect 7009 -871 7043 -837
rect 6859 -914 6893 -880
rect 6859 -986 6893 -952
rect 6859 -1058 6893 -1024
rect 6859 -1130 6893 -1096
rect 6859 -1202 6893 -1168
rect 6859 -1274 6893 -1240
rect 6859 -1346 6893 -1312
rect 6859 -1418 6893 -1384
rect 6859 -1490 6893 -1456
rect 6859 -1562 6893 -1528
rect 6859 -1634 6893 -1600
rect 7009 -943 7043 -909
rect 7009 -1015 7043 -981
rect 7009 -1087 7043 -1053
rect 7009 -1159 7043 -1125
rect 7009 -1231 7043 -1197
rect 7009 -1303 7043 -1269
rect 7009 -1375 7043 -1341
rect 7009 -1447 7043 -1413
rect 7009 -1519 7043 -1485
rect 7899 -871 7933 -837
rect 7899 -943 7933 -909
rect 7899 -1015 7933 -981
rect 7899 -1087 7933 -1053
rect 7899 -1159 7933 -1125
rect 7899 -1231 7933 -1197
rect 7899 -1303 7933 -1269
rect 7899 -1375 7933 -1341
rect 7899 -1447 7933 -1413
rect 7899 -1519 7933 -1485
rect 7009 -1591 7043 -1557
rect 7899 -1591 7933 -1557
rect 6859 -1706 6893 -1672
rect 8045 -842 8079 -808
rect 8045 -914 8079 -880
rect 8045 -986 8079 -952
rect 8045 -1058 8079 -1024
rect 8045 -1130 8079 -1096
rect 8045 -1202 8079 -1168
rect 8045 -1274 8079 -1240
rect 8045 -1346 8079 -1312
rect 8045 -1418 8079 -1384
rect 8045 -1490 8079 -1456
rect 8045 -1562 8079 -1528
rect 7009 -1677 7043 -1643
rect 7094 -1677 7128 -1643
rect 7166 -1677 7200 -1643
rect 7238 -1677 7272 -1643
rect 7310 -1677 7344 -1643
rect 7382 -1677 7416 -1643
rect 7454 -1677 7488 -1643
rect 7526 -1677 7560 -1643
rect 7598 -1677 7632 -1643
rect 7670 -1677 7704 -1643
rect 7742 -1677 7776 -1643
rect 7814 -1677 7848 -1643
rect 7899 -1678 7933 -1644
rect 8045 -1634 8079 -1600
rect 8045 -1706 8079 -1672
rect 5466 -1829 5500 -1795
rect 5538 -1829 5572 -1795
rect 5610 -1829 5644 -1795
rect 5682 -1829 5716 -1795
rect 5754 -1829 5788 -1795
rect 5826 -1829 5860 -1795
rect 5898 -1829 5932 -1795
rect 5970 -1829 6004 -1795
rect 6042 -1829 6076 -1795
rect 6114 -1829 6148 -1795
rect 6186 -1829 6220 -1795
rect 6258 -1829 6292 -1795
rect 6330 -1829 6364 -1795
rect 6402 -1829 6436 -1795
rect 6474 -1829 6508 -1795
rect 6546 -1829 6580 -1795
rect 6618 -1829 6652 -1795
rect 6876 -1825 6910 -1791
rect 6948 -1825 6982 -1791
rect 7020 -1825 7054 -1791
rect 7092 -1825 7126 -1791
rect 7164 -1825 7198 -1791
rect 7236 -1825 7270 -1791
rect 7308 -1825 7342 -1791
rect 7380 -1825 7414 -1791
rect 7452 -1825 7486 -1791
rect 7524 -1825 7558 -1791
rect 7596 -1825 7630 -1791
rect 7668 -1825 7702 -1791
rect 7740 -1825 7774 -1791
rect 7812 -1825 7846 -1791
rect 7884 -1825 7918 -1791
rect 7956 -1825 7990 -1791
rect 8028 -1825 8062 -1791
rect 5464 -2011 5498 -1977
rect 5536 -2011 5570 -1977
rect 5608 -2011 5642 -1977
rect 5680 -2011 5714 -1977
rect 5752 -2011 5786 -1977
rect 5824 -2011 5858 -1977
rect 5896 -2011 5930 -1977
rect 5968 -2011 6002 -1977
rect 6040 -2011 6074 -1977
rect 6112 -2011 6146 -1977
rect 6184 -2011 6218 -1977
rect 6256 -2011 6290 -1977
rect 6328 -2011 6362 -1977
rect 6400 -2011 6434 -1977
rect 6472 -2011 6506 -1977
rect 6544 -2011 6578 -1977
rect 6616 -2011 6650 -1977
rect 6878 -2009 6912 -1975
rect 6950 -2009 6984 -1975
rect 7022 -2009 7056 -1975
rect 7094 -2009 7128 -1975
rect 7166 -2009 7200 -1975
rect 7238 -2009 7272 -1975
rect 7310 -2009 7344 -1975
rect 7382 -2009 7416 -1975
rect 7454 -2009 7488 -1975
rect 7526 -2009 7560 -1975
rect 7598 -2009 7632 -1975
rect 7670 -2009 7704 -1975
rect 7742 -2009 7776 -1975
rect 7814 -2009 7848 -1975
rect 7886 -2009 7920 -1975
rect 7958 -2009 7992 -1975
rect 8030 -2009 8064 -1975
rect 5447 -2130 5481 -2096
rect 5607 -2145 5641 -2111
rect 5679 -2145 5713 -2111
rect 5751 -2145 5785 -2111
rect 5823 -2145 5857 -2111
rect 5895 -2145 5929 -2111
rect 5967 -2145 6001 -2111
rect 6039 -2145 6073 -2111
rect 6111 -2145 6145 -2111
rect 6183 -2145 6217 -2111
rect 6255 -2145 6289 -2111
rect 6327 -2145 6361 -2111
rect 6399 -2145 6433 -2111
rect 5447 -2202 5481 -2168
rect 6633 -2130 6667 -2096
rect 5597 -2231 5631 -2197
rect 5447 -2274 5481 -2240
rect 5447 -2346 5481 -2312
rect 5447 -2418 5481 -2384
rect 5447 -2490 5481 -2456
rect 5447 -2562 5481 -2528
rect 5447 -2634 5481 -2600
rect 5447 -2706 5481 -2672
rect 5447 -2778 5481 -2744
rect 5447 -2850 5481 -2816
rect 5447 -2922 5481 -2888
rect 5447 -2994 5481 -2960
rect 5597 -2303 5631 -2269
rect 5597 -2375 5631 -2341
rect 5597 -2447 5631 -2413
rect 5597 -2519 5631 -2485
rect 5597 -2591 5631 -2557
rect 5597 -2663 5631 -2629
rect 5597 -2735 5631 -2701
rect 5597 -2807 5631 -2773
rect 5597 -2879 5631 -2845
rect 6487 -2231 6521 -2197
rect 6487 -2303 6521 -2269
rect 6487 -2375 6521 -2341
rect 6487 -2447 6521 -2413
rect 6487 -2519 6521 -2485
rect 6487 -2591 6521 -2557
rect 6487 -2663 6521 -2629
rect 6487 -2735 6521 -2701
rect 6487 -2807 6521 -2773
rect 6487 -2879 6521 -2845
rect 5597 -2951 5631 -2917
rect 6487 -2951 6521 -2917
rect 5447 -3066 5481 -3032
rect 6633 -2202 6667 -2168
rect 6633 -2274 6667 -2240
rect 6633 -2346 6667 -2312
rect 6633 -2418 6667 -2384
rect 6633 -2490 6667 -2456
rect 6633 -2562 6667 -2528
rect 6633 -2634 6667 -2600
rect 6633 -2706 6667 -2672
rect 6633 -2778 6667 -2744
rect 6633 -2850 6667 -2816
rect 6633 -2922 6667 -2888
rect 5597 -3037 5631 -3003
rect 5682 -3037 5716 -3003
rect 5754 -3037 5788 -3003
rect 5826 -3037 5860 -3003
rect 5898 -3037 5932 -3003
rect 5970 -3037 6004 -3003
rect 6042 -3037 6076 -3003
rect 6114 -3037 6148 -3003
rect 6186 -3037 6220 -3003
rect 6258 -3037 6292 -3003
rect 6330 -3037 6364 -3003
rect 6402 -3037 6436 -3003
rect 6487 -3038 6521 -3004
rect 6633 -2994 6667 -2960
rect 6633 -3066 6667 -3032
rect 6861 -2128 6895 -2094
rect 7021 -2143 7055 -2109
rect 7093 -2143 7127 -2109
rect 7165 -2143 7199 -2109
rect 7237 -2143 7271 -2109
rect 7309 -2143 7343 -2109
rect 7381 -2143 7415 -2109
rect 7453 -2143 7487 -2109
rect 7525 -2143 7559 -2109
rect 7597 -2143 7631 -2109
rect 7669 -2143 7703 -2109
rect 7741 -2143 7775 -2109
rect 7813 -2143 7847 -2109
rect 6861 -2200 6895 -2166
rect 8047 -2128 8081 -2094
rect 7011 -2229 7045 -2195
rect 6861 -2272 6895 -2238
rect 6861 -2344 6895 -2310
rect 6861 -2416 6895 -2382
rect 6861 -2488 6895 -2454
rect 6861 -2560 6895 -2526
rect 6861 -2632 6895 -2598
rect 6861 -2704 6895 -2670
rect 6861 -2776 6895 -2742
rect 6861 -2848 6895 -2814
rect 6861 -2920 6895 -2886
rect 6861 -2992 6895 -2958
rect 7011 -2301 7045 -2267
rect 7011 -2373 7045 -2339
rect 7011 -2445 7045 -2411
rect 7011 -2517 7045 -2483
rect 7011 -2589 7045 -2555
rect 7011 -2661 7045 -2627
rect 7011 -2733 7045 -2699
rect 7011 -2805 7045 -2771
rect 7011 -2877 7045 -2843
rect 7901 -2229 7935 -2195
rect 7901 -2301 7935 -2267
rect 7901 -2373 7935 -2339
rect 7901 -2445 7935 -2411
rect 7901 -2517 7935 -2483
rect 7901 -2589 7935 -2555
rect 7901 -2661 7935 -2627
rect 7901 -2733 7935 -2699
rect 7901 -2805 7935 -2771
rect 7901 -2877 7935 -2843
rect 7011 -2949 7045 -2915
rect 7901 -2949 7935 -2915
rect 6861 -3064 6895 -3030
rect 8047 -2200 8081 -2166
rect 8047 -2272 8081 -2238
rect 8047 -2344 8081 -2310
rect 8047 -2416 8081 -2382
rect 8047 -2488 8081 -2454
rect 8047 -2560 8081 -2526
rect 8047 -2632 8081 -2598
rect 8047 -2704 8081 -2670
rect 8047 -2776 8081 -2742
rect 8047 -2848 8081 -2814
rect 8047 -2920 8081 -2886
rect 7011 -3035 7045 -3001
rect 7096 -3035 7130 -3001
rect 7168 -3035 7202 -3001
rect 7240 -3035 7274 -3001
rect 7312 -3035 7346 -3001
rect 7384 -3035 7418 -3001
rect 7456 -3035 7490 -3001
rect 7528 -3035 7562 -3001
rect 7600 -3035 7634 -3001
rect 7672 -3035 7706 -3001
rect 7744 -3035 7778 -3001
rect 7816 -3035 7850 -3001
rect 7901 -3036 7935 -3002
rect 8047 -2992 8081 -2958
rect 8047 -3064 8081 -3030
rect 5464 -3185 5498 -3151
rect 5536 -3185 5570 -3151
rect 5608 -3185 5642 -3151
rect 5680 -3185 5714 -3151
rect 5752 -3185 5786 -3151
rect 5824 -3185 5858 -3151
rect 5896 -3185 5930 -3151
rect 5968 -3185 6002 -3151
rect 6040 -3185 6074 -3151
rect 6112 -3185 6146 -3151
rect 6184 -3185 6218 -3151
rect 6256 -3185 6290 -3151
rect 6328 -3185 6362 -3151
rect 6400 -3185 6434 -3151
rect 6472 -3185 6506 -3151
rect 6544 -3185 6578 -3151
rect 6616 -3185 6650 -3151
rect 6878 -3183 6912 -3149
rect 6950 -3183 6984 -3149
rect 7022 -3183 7056 -3149
rect 7094 -3183 7128 -3149
rect 7166 -3183 7200 -3149
rect 7238 -3183 7272 -3149
rect 7310 -3183 7344 -3149
rect 7382 -3183 7416 -3149
rect 7454 -3183 7488 -3149
rect 7526 -3183 7560 -3149
rect 7598 -3183 7632 -3149
rect 7670 -3183 7704 -3149
rect 7742 -3183 7776 -3149
rect 7814 -3183 7848 -3149
rect 7886 -3183 7920 -3149
rect 7958 -3183 7992 -3149
rect 8030 -3183 8064 -3149
rect 5464 -3363 5498 -3329
rect 5536 -3363 5570 -3329
rect 5608 -3363 5642 -3329
rect 5680 -3363 5714 -3329
rect 5752 -3363 5786 -3329
rect 5824 -3363 5858 -3329
rect 5896 -3363 5930 -3329
rect 5968 -3363 6002 -3329
rect 6040 -3363 6074 -3329
rect 6112 -3363 6146 -3329
rect 6184 -3363 6218 -3329
rect 6256 -3363 6290 -3329
rect 6328 -3363 6362 -3329
rect 6400 -3363 6434 -3329
rect 6472 -3363 6506 -3329
rect 6544 -3363 6578 -3329
rect 6616 -3363 6650 -3329
rect 6880 -3369 6914 -3335
rect 6952 -3369 6986 -3335
rect 7024 -3369 7058 -3335
rect 7096 -3369 7130 -3335
rect 7168 -3369 7202 -3335
rect 7240 -3369 7274 -3335
rect 7312 -3369 7346 -3335
rect 7384 -3369 7418 -3335
rect 7456 -3369 7490 -3335
rect 7528 -3369 7562 -3335
rect 7600 -3369 7634 -3335
rect 7672 -3369 7706 -3335
rect 7744 -3369 7778 -3335
rect 7816 -3369 7850 -3335
rect 7888 -3369 7922 -3335
rect 7960 -3369 7994 -3335
rect 8032 -3369 8066 -3335
rect 5447 -3482 5481 -3448
rect 5607 -3497 5641 -3463
rect 5679 -3497 5713 -3463
rect 5751 -3497 5785 -3463
rect 5823 -3497 5857 -3463
rect 5895 -3497 5929 -3463
rect 5967 -3497 6001 -3463
rect 6039 -3497 6073 -3463
rect 6111 -3497 6145 -3463
rect 6183 -3497 6217 -3463
rect 6255 -3497 6289 -3463
rect 6327 -3497 6361 -3463
rect 6399 -3497 6433 -3463
rect 5447 -3554 5481 -3520
rect 6633 -3482 6667 -3448
rect 5597 -3583 5631 -3549
rect 5447 -3626 5481 -3592
rect 5447 -3698 5481 -3664
rect 5447 -3770 5481 -3736
rect 5447 -3842 5481 -3808
rect 5447 -3914 5481 -3880
rect 5447 -3986 5481 -3952
rect 5447 -4058 5481 -4024
rect 5447 -4130 5481 -4096
rect 5447 -4202 5481 -4168
rect 5447 -4274 5481 -4240
rect 5447 -4346 5481 -4312
rect 5597 -3655 5631 -3621
rect 5597 -3727 5631 -3693
rect 5597 -3799 5631 -3765
rect 5597 -3871 5631 -3837
rect 5597 -3943 5631 -3909
rect 5597 -4015 5631 -3981
rect 5597 -4087 5631 -4053
rect 5597 -4159 5631 -4125
rect 5597 -4231 5631 -4197
rect 6487 -3583 6521 -3549
rect 6487 -3655 6521 -3621
rect 6487 -3727 6521 -3693
rect 6487 -3799 6521 -3765
rect 6487 -3871 6521 -3837
rect 6487 -3943 6521 -3909
rect 6487 -4015 6521 -3981
rect 6487 -4087 6521 -4053
rect 6487 -4159 6521 -4125
rect 6487 -4231 6521 -4197
rect 5597 -4303 5631 -4269
rect 6487 -4303 6521 -4269
rect 5447 -4418 5481 -4384
rect 6633 -3554 6667 -3520
rect 6633 -3626 6667 -3592
rect 6633 -3698 6667 -3664
rect 6633 -3770 6667 -3736
rect 6633 -3842 6667 -3808
rect 6633 -3914 6667 -3880
rect 6633 -3986 6667 -3952
rect 6633 -4058 6667 -4024
rect 6633 -4130 6667 -4096
rect 6633 -4202 6667 -4168
rect 6633 -4274 6667 -4240
rect 5597 -4389 5631 -4355
rect 5682 -4389 5716 -4355
rect 5754 -4389 5788 -4355
rect 5826 -4389 5860 -4355
rect 5898 -4389 5932 -4355
rect 5970 -4389 6004 -4355
rect 6042 -4389 6076 -4355
rect 6114 -4389 6148 -4355
rect 6186 -4389 6220 -4355
rect 6258 -4389 6292 -4355
rect 6330 -4389 6364 -4355
rect 6402 -4389 6436 -4355
rect 6487 -4390 6521 -4356
rect 6633 -4346 6667 -4312
rect 6633 -4418 6667 -4384
rect 6863 -3488 6897 -3454
rect 7023 -3503 7057 -3469
rect 7095 -3503 7129 -3469
rect 7167 -3503 7201 -3469
rect 7239 -3503 7273 -3469
rect 7311 -3503 7345 -3469
rect 7383 -3503 7417 -3469
rect 7455 -3503 7489 -3469
rect 7527 -3503 7561 -3469
rect 7599 -3503 7633 -3469
rect 7671 -3503 7705 -3469
rect 7743 -3503 7777 -3469
rect 7815 -3503 7849 -3469
rect 6863 -3560 6897 -3526
rect 8049 -3488 8083 -3454
rect 7013 -3589 7047 -3555
rect 6863 -3632 6897 -3598
rect 6863 -3704 6897 -3670
rect 6863 -3776 6897 -3742
rect 6863 -3848 6897 -3814
rect 6863 -3920 6897 -3886
rect 6863 -3992 6897 -3958
rect 6863 -4064 6897 -4030
rect 6863 -4136 6897 -4102
rect 6863 -4208 6897 -4174
rect 6863 -4280 6897 -4246
rect 6863 -4352 6897 -4318
rect 7013 -3661 7047 -3627
rect 7013 -3733 7047 -3699
rect 7013 -3805 7047 -3771
rect 7013 -3877 7047 -3843
rect 7013 -3949 7047 -3915
rect 7013 -4021 7047 -3987
rect 7013 -4093 7047 -4059
rect 7013 -4165 7047 -4131
rect 7013 -4237 7047 -4203
rect 7903 -3589 7937 -3555
rect 7903 -3661 7937 -3627
rect 7903 -3733 7937 -3699
rect 7903 -3805 7937 -3771
rect 7903 -3877 7937 -3843
rect 7903 -3949 7937 -3915
rect 7903 -4021 7937 -3987
rect 7903 -4093 7937 -4059
rect 7903 -4165 7937 -4131
rect 7903 -4237 7937 -4203
rect 7013 -4309 7047 -4275
rect 7903 -4309 7937 -4275
rect 6863 -4424 6897 -4390
rect 8049 -3560 8083 -3526
rect 8049 -3632 8083 -3598
rect 8049 -3704 8083 -3670
rect 8049 -3776 8083 -3742
rect 8049 -3848 8083 -3814
rect 8049 -3920 8083 -3886
rect 8049 -3992 8083 -3958
rect 8049 -4064 8083 -4030
rect 8049 -4136 8083 -4102
rect 8049 -4208 8083 -4174
rect 8049 -4280 8083 -4246
rect 7013 -4395 7047 -4361
rect 7098 -4395 7132 -4361
rect 7170 -4395 7204 -4361
rect 7242 -4395 7276 -4361
rect 7314 -4395 7348 -4361
rect 7386 -4395 7420 -4361
rect 7458 -4395 7492 -4361
rect 7530 -4395 7564 -4361
rect 7602 -4395 7636 -4361
rect 7674 -4395 7708 -4361
rect 7746 -4395 7780 -4361
rect 7818 -4395 7852 -4361
rect 7903 -4396 7937 -4362
rect 8049 -4352 8083 -4318
rect 5464 -4537 5498 -4503
rect 5536 -4537 5570 -4503
rect 5608 -4537 5642 -4503
rect 5680 -4537 5714 -4503
rect 5752 -4537 5786 -4503
rect 5824 -4537 5858 -4503
rect 5896 -4537 5930 -4503
rect 5968 -4537 6002 -4503
rect 6040 -4537 6074 -4503
rect 6112 -4537 6146 -4503
rect 6184 -4537 6218 -4503
rect 6256 -4537 6290 -4503
rect 6328 -4537 6362 -4503
rect 6400 -4537 6434 -4503
rect 6472 -4537 6506 -4503
rect 6544 -4537 6578 -4503
rect 6616 -4537 6650 -4503
rect 8049 -4424 8083 -4390
rect 6880 -4543 6914 -4509
rect 6952 -4543 6986 -4509
rect 7024 -4543 7058 -4509
rect 7096 -4543 7130 -4509
rect 7168 -4543 7202 -4509
rect 7240 -4543 7274 -4509
rect 7312 -4543 7346 -4509
rect 7384 -4543 7418 -4509
rect 7456 -4543 7490 -4509
rect 7528 -4543 7562 -4509
rect 7600 -4543 7634 -4509
rect 7672 -4543 7706 -4509
rect 7744 -4543 7778 -4509
rect 7816 -4543 7850 -4509
rect 7888 -4543 7922 -4509
rect 7960 -4543 7994 -4509
rect 8032 -4543 8066 -4509
rect 2316 -5126 2350 -5092
rect 5585 -5127 5619 -5093
rect 7002 -5091 7036 -5057
<< metal1 >>
rect 526 8276 566 8546
rect 2478 8332 2512 8532
rect 524 8206 566 8276
rect 2476 8260 2514 8332
rect 3826 8260 3860 8530
rect 5462 8340 5496 8562
rect 2472 8214 2512 8260
rect 3822 8214 3860 8260
rect 5458 8260 5496 8340
rect 5458 8214 5492 8260
rect 5916 8214 5950 8488
rect 6948 8342 6986 8560
rect 522 7158 566 8206
rect 2470 7158 2512 8214
rect 3820 7158 3862 8214
rect 522 5444 564 7158
rect 2470 5444 2510 7158
rect 522 5308 560 5444
rect 332 5270 562 5308
rect 332 5064 376 5270
rect 2470 5220 2508 5444
rect 2472 5086 2506 5220
rect 3820 5214 3858 7158
rect 5456 7154 5492 8214
rect 5914 7154 5950 8214
rect 6946 8278 6986 8342
rect 8004 8306 8036 8440
rect 8868 8306 8900 8454
rect 6946 8266 6984 8278
rect 6946 8198 6982 8266
rect 8004 8202 8038 8306
rect 8868 8208 8902 8306
rect 6946 7954 6980 8198
rect 8004 8050 8040 8202
rect 8866 8056 8902 8208
rect 9716 8202 9754 8452
rect 9716 8198 9752 8202
rect 9718 8060 9752 8198
rect 5456 7048 5490 7154
rect 5914 7064 5948 7154
rect 5946 7056 5948 7064
rect 3818 5090 3858 5214
rect -1166 4712 -1086 4796
rect 10290 4280 10506 4322
rect 10290 4278 10342 4280
rect 798 4138 1362 4194
rect 4280 3252 5096 3328
rect 4280 3250 4362 3252
rect 4468 3100 4790 3144
rect 3390 1190 3392 1200
rect 800 1132 944 1188
rect 1626 1146 2048 1184
rect 3220 1180 3362 1190
rect 2922 1169 2982 1178
rect 686 1050 774 1054
rect 686 998 704 1050
rect 756 998 774 1050
rect 686 994 774 998
rect 686 992 720 994
rect -1848 -1660 -1784 682
rect 896 -84 942 1132
rect 1142 1048 1222 1056
rect 1142 996 1162 1048
rect 1214 996 1222 1048
rect 1142 992 1222 996
rect 1136 915 1220 950
rect 1136 863 1152 915
rect 1204 863 1220 915
rect 1136 844 1220 863
rect 1920 730 1960 1146
rect 2922 1117 2926 1169
rect 2978 1117 2982 1169
rect 2922 1106 2982 1117
rect 3220 1128 3239 1180
rect 3291 1128 3362 1180
rect 3220 1116 3362 1128
rect 3364 1120 3392 1190
rect 3562 1071 3676 1082
rect 2240 1054 2320 1056
rect 2240 950 2310 1054
rect 2706 1024 3468 1058
rect 3562 1019 3594 1071
rect 3646 1019 3676 1071
rect 4150 1064 4240 1070
rect 3562 1008 3676 1019
rect 3980 950 4040 1036
rect 4150 1012 4169 1064
rect 4221 1012 4240 1064
rect 4150 1004 4240 1012
rect 2240 942 4040 950
rect 2240 890 2254 942
rect 2306 890 4040 942
rect 2240 880 4040 890
rect 4468 844 4544 3100
rect 4736 3044 4790 3100
rect 5026 2750 5096 3252
rect 7402 3172 7462 3178
rect 7400 3155 7462 3172
rect 10164 3168 10230 3170
rect 7400 3103 7407 3155
rect 7459 3103 7462 3155
rect 9308 3154 9368 3162
rect 7400 3094 7462 3103
rect 8446 3142 8506 3148
rect 8446 3090 8454 3142
rect 9308 3102 9316 3154
rect 10164 3116 10172 3168
rect 10224 3116 10230 3168
rect 10164 3106 10230 3116
rect 9308 3092 9368 3102
rect 8446 3080 8506 3090
rect 5610 3052 5680 3060
rect 5610 3000 5620 3052
rect 5672 3000 5680 3052
rect 9340 3044 9798 3046
rect 8636 3040 8960 3044
rect 5610 2990 5680 3000
rect 5876 3034 7472 3036
rect 8420 3034 8960 3040
rect 5876 2998 8120 3034
rect 5876 2996 7472 2998
rect 7994 2996 8120 2998
rect 8330 2996 8960 3034
rect 9272 3032 9798 3044
rect 9030 3000 9798 3032
rect 9030 2998 9498 3000
rect 8400 2994 8960 2996
rect 8420 2988 8960 2994
rect 5026 2692 8190 2750
rect 5026 2690 5286 2692
rect 5026 2594 5096 2690
rect 4926 2590 5228 2594
rect 4926 2534 5890 2590
rect 5834 1545 5890 2534
rect 8140 2586 8190 2692
rect 8698 2588 9676 2590
rect 8698 2586 9736 2588
rect 10290 2586 10340 4278
rect 8140 2518 10340 2586
rect 8140 2516 9736 2518
rect 8140 2514 9676 2516
rect 6820 2156 6916 2170
rect 6820 2103 8118 2156
rect 6820 2069 6876 2103
rect 6910 2069 6948 2103
rect 6982 2069 7020 2103
rect 7054 2069 7092 2103
rect 7126 2069 7164 2103
rect 7198 2069 7236 2103
rect 7270 2069 7308 2103
rect 7342 2069 7380 2103
rect 7414 2069 7452 2103
rect 7486 2069 7524 2103
rect 7558 2069 7596 2103
rect 7630 2069 7668 2103
rect 7702 2069 7740 2103
rect 7774 2069 7812 2103
rect 7846 2069 7884 2103
rect 7918 2069 7956 2103
rect 7990 2069 8028 2103
rect 8062 2069 8118 2103
rect 6820 2050 8118 2069
rect 6820 1984 6922 2050
rect 6820 1950 6859 1984
rect 6893 1950 6922 1984
rect 6820 1912 6922 1950
rect 6986 1969 7952 1986
rect 6986 1935 7019 1969
rect 7053 1935 7091 1969
rect 7125 1935 7163 1969
rect 7197 1935 7235 1969
rect 7269 1935 7307 1969
rect 7341 1935 7379 1969
rect 7413 1935 7451 1969
rect 7485 1935 7523 1969
rect 7557 1935 7595 1969
rect 7629 1935 7667 1969
rect 7701 1935 7739 1969
rect 7773 1935 7811 1969
rect 7845 1935 7952 1969
rect 6986 1926 7952 1935
rect 6820 1878 6859 1912
rect 6893 1878 6922 1912
rect 6522 1736 6558 1864
rect 6820 1840 6922 1878
rect 6984 1918 7952 1926
rect 8014 1984 8116 2050
rect 8014 1950 8045 1984
rect 8079 1950 8116 1984
rect 6984 1883 7062 1918
rect 6984 1849 7009 1883
rect 7043 1849 7062 1883
rect 7874 1883 7948 1918
rect 6984 1846 7062 1849
rect 6820 1806 6859 1840
rect 6893 1806 6922 1840
rect 6820 1768 6922 1806
rect 5834 1124 6370 1545
rect 6520 1432 6562 1736
rect 6820 1734 6859 1768
rect 6893 1734 6922 1768
rect 6820 1696 6922 1734
rect 6820 1662 6859 1696
rect 6893 1662 6922 1696
rect 6820 1624 6922 1662
rect 6820 1590 6859 1624
rect 6893 1590 6922 1624
rect 6820 1552 6922 1590
rect 6820 1518 6859 1552
rect 6893 1518 6922 1552
rect 6820 1480 6922 1518
rect 6820 1446 6859 1480
rect 6893 1446 6922 1480
rect 3220 831 4544 844
rect 3220 779 3244 831
rect 3296 828 4544 831
rect 3296 779 3595 828
rect 3220 776 3595 779
rect 3647 776 4544 828
rect 3220 766 4544 776
rect 4700 972 4744 1006
rect 1618 712 1684 720
rect 1618 660 1626 712
rect 1678 660 1684 712
rect 1920 690 3510 730
rect 1618 652 1684 660
rect 1660 650 1684 652
rect 3300 542 3368 552
rect 1890 522 3150 528
rect 1862 482 3150 522
rect 1862 448 1911 482
rect 1945 448 1983 482
rect 2017 448 2055 482
rect 2089 448 2127 482
rect 2161 448 2199 482
rect 2233 448 2271 482
rect 2305 448 2343 482
rect 2377 448 2415 482
rect 2449 448 2487 482
rect 2521 448 2559 482
rect 2593 448 2631 482
rect 2665 448 2703 482
rect 2737 448 2775 482
rect 2809 448 2847 482
rect 2881 448 2919 482
rect 2953 448 2991 482
rect 3025 448 3063 482
rect 3097 448 3150 482
rect 3300 490 3310 542
rect 3362 490 3368 542
rect 3300 480 3368 490
rect 1862 428 3150 448
rect 1862 363 1954 428
rect 1862 329 1892 363
rect 1926 329 1954 363
rect 1862 291 1954 329
rect 2022 349 2986 368
rect 2022 315 2053 349
rect 2087 315 2125 349
rect 2159 315 2197 349
rect 2231 315 2269 349
rect 2303 315 2341 349
rect 2375 315 2413 349
rect 2447 315 2485 349
rect 2519 315 2557 349
rect 2591 315 2629 349
rect 2663 315 2701 349
rect 2735 315 2773 349
rect 2807 315 2845 349
rect 2879 315 2917 349
rect 2951 315 2986 349
rect 2022 312 2986 315
rect 1862 257 1892 291
rect 1926 257 1954 291
rect 1862 219 1954 257
rect 1616 171 1690 192
rect 1616 119 1624 171
rect 1676 119 1690 171
rect 1616 88 1690 119
rect 1862 185 1892 219
rect 1926 185 1954 219
rect 1862 147 1954 185
rect 1862 113 1892 147
rect 1926 113 1954 147
rect 892 -196 942 -84
rect 1862 75 1954 113
rect 1862 41 1892 75
rect 1926 41 1954 75
rect 1862 3 1954 41
rect 1862 -31 1892 3
rect 1926 -31 1954 3
rect 1862 -69 1954 -31
rect 1862 -103 1892 -69
rect 1926 -103 1954 -69
rect 1862 -141 1954 -103
rect 1862 -175 1892 -141
rect 1926 -175 1954 -141
rect 892 -244 1266 -196
rect 1862 -213 1954 -175
rect 892 -446 940 -244
rect -910 -498 -860 -488
rect -910 -666 -836 -498
rect 1216 -582 1264 -244
rect 1862 -247 1892 -213
rect 1926 -247 1954 -213
rect 1862 -285 1954 -247
rect 1862 -319 1892 -285
rect 1926 -319 1954 -285
rect 1862 -357 1954 -319
rect 1862 -391 1892 -357
rect 1926 -391 1954 -357
rect 1862 -429 1954 -391
rect 1862 -463 1892 -429
rect 1926 -463 1954 -429
rect 1862 -501 1954 -463
rect 1862 -535 1892 -501
rect 1926 -535 1954 -501
rect 2020 298 2986 312
rect 2020 263 2090 298
rect 2020 229 2042 263
rect 2076 229 2090 263
rect 2916 263 2986 298
rect 2020 191 2090 229
rect 2020 157 2042 191
rect 2076 157 2090 191
rect 2020 119 2090 157
rect 2020 85 2042 119
rect 2076 85 2090 119
rect 2020 47 2090 85
rect 2020 13 2042 47
rect 2076 13 2090 47
rect 2020 -25 2090 13
rect 2020 -59 2042 -25
rect 2076 -59 2090 -25
rect 2020 -97 2090 -59
rect 2020 -131 2042 -97
rect 2076 -131 2090 -97
rect 2020 -169 2090 -131
rect 2020 -203 2042 -169
rect 2076 -203 2090 -169
rect 2020 -241 2090 -203
rect 2020 -275 2042 -241
rect 2076 -275 2090 -241
rect 2020 -313 2090 -275
rect 2020 -347 2042 -313
rect 2076 -347 2090 -313
rect 2020 -385 2090 -347
rect 2020 -419 2042 -385
rect 2076 -419 2090 -385
rect 2020 -457 2090 -419
rect 2020 -491 2042 -457
rect 2076 -491 2090 -457
rect 2154 173 2844 230
rect 2154 -391 2224 173
rect 2788 -391 2844 173
rect 2154 -462 2844 -391
rect 2916 229 2932 263
rect 2966 229 2986 263
rect 2916 191 2986 229
rect 2916 157 2932 191
rect 2966 157 2986 191
rect 2916 119 2986 157
rect 2916 85 2932 119
rect 2966 85 2986 119
rect 2916 47 2986 85
rect 2916 13 2932 47
rect 2966 13 2986 47
rect 2916 -25 2986 13
rect 2916 -59 2932 -25
rect 2966 -59 2986 -25
rect 2916 -97 2986 -59
rect 2916 -131 2932 -97
rect 2966 -131 2986 -97
rect 2916 -169 2986 -131
rect 2916 -203 2932 -169
rect 2966 -203 2986 -169
rect 2916 -241 2986 -203
rect 2916 -275 2932 -241
rect 2966 -275 2986 -241
rect 2916 -313 2986 -275
rect 2916 -347 2932 -313
rect 2966 -347 2986 -313
rect 2916 -385 2986 -347
rect 2916 -419 2932 -385
rect 2966 -419 2986 -385
rect 2916 -457 2986 -419
rect 2020 -526 2090 -491
rect 2916 -491 2932 -457
rect 2966 -491 2986 -457
rect 2916 -526 2986 -491
rect 1862 -573 1954 -535
rect 1862 -607 1892 -573
rect 1926 -607 1954 -573
rect 2018 -538 2986 -526
rect 2018 -590 2031 -538
rect 2083 -543 2986 -538
rect 2083 -577 2127 -543
rect 2161 -577 2199 -543
rect 2233 -577 2271 -543
rect 2305 -577 2343 -543
rect 2377 -577 2415 -543
rect 2449 -577 2487 -543
rect 2521 -577 2559 -543
rect 2593 -577 2631 -543
rect 2665 -577 2703 -543
rect 2737 -577 2775 -543
rect 2809 -577 2847 -543
rect 2881 -577 2932 -543
rect 2966 -577 2986 -543
rect 2083 -590 2986 -577
rect 2018 -596 2986 -590
rect 3052 363 3144 428
rect 3052 329 3082 363
rect 3116 329 3144 363
rect 3052 291 3144 329
rect 3052 257 3082 291
rect 3116 257 3144 291
rect 3052 219 3144 257
rect 3052 185 3082 219
rect 3116 185 3144 219
rect 3052 147 3144 185
rect 3052 113 3082 147
rect 3116 113 3144 147
rect 3052 75 3144 113
rect 3052 41 3082 75
rect 3116 41 3144 75
rect 3052 3 3144 41
rect 3052 -31 3082 3
rect 3116 -31 3144 3
rect 3052 -69 3144 -31
rect 3052 -103 3082 -69
rect 3116 -103 3144 -69
rect 3052 -141 3144 -103
rect 3052 -175 3082 -141
rect 3116 -175 3144 -141
rect 3052 -213 3144 -175
rect 3052 -247 3082 -213
rect 3116 -247 3144 -213
rect 3052 -285 3144 -247
rect 3052 -319 3082 -285
rect 3116 -319 3144 -285
rect 3052 -357 3144 -319
rect 3052 -391 3082 -357
rect 3116 -391 3144 -357
rect 3052 -429 3144 -391
rect 3052 -463 3082 -429
rect 3116 -463 3144 -429
rect 3052 -501 3144 -463
rect 3052 -535 3082 -501
rect 3116 -535 3144 -501
rect 3052 -573 3144 -535
rect 2018 -598 2100 -596
rect 1862 -660 1954 -607
rect 3052 -607 3082 -573
rect 3116 -607 3144 -573
rect 3052 -660 3144 -607
rect -2022 -1736 -1782 -1660
rect -2020 -3420 -1950 -1736
rect -1166 -2236 -1090 -1820
rect -1378 -3136 -1328 -2946
rect -2018 -4950 -1950 -3420
rect -1588 -3186 -1328 -3136
rect -1588 -4950 -1532 -3186
rect -1158 -3540 -1090 -3286
rect -1374 -3594 -1090 -3540
rect -910 -3566 -860 -666
rect 1860 -692 3144 -660
rect 1860 -726 1911 -692
rect 1945 -726 1983 -692
rect 2017 -726 2055 -692
rect 2089 -726 2127 -692
rect 2161 -726 2199 -692
rect 2233 -726 2271 -692
rect 2305 -726 2343 -692
rect 2377 -726 2415 -692
rect 2449 -726 2487 -692
rect 2521 -726 2559 -692
rect 2593 -726 2631 -692
rect 2665 -726 2703 -692
rect 2737 -726 2775 -692
rect 2809 -726 2847 -692
rect 2881 -726 2919 -692
rect 2953 -726 2991 -692
rect 3025 -726 3063 -692
rect 3097 -726 3144 -692
rect 1860 -754 3144 -726
rect 1860 -760 3120 -754
rect 1888 -1358 1952 -760
rect 3304 -826 3368 480
rect 2392 -884 3368 -826
rect 2392 -1096 2430 -884
rect 3460 -988 3510 690
rect 4700 660 4742 972
rect 3930 630 4742 660
rect 3930 608 4740 630
rect 3930 400 3980 608
rect 4150 512 4252 514
rect 4150 460 4178 512
rect 4230 460 4252 512
rect 4150 450 4252 460
rect 3928 352 4094 400
rect 3928 350 4066 352
rect 3932 -818 3976 350
rect 4580 156 5092 158
rect 6120 156 6154 274
rect 4580 122 6154 156
rect 4580 120 5096 122
rect 6120 120 6154 122
rect 3932 -864 4536 -818
rect 3932 -866 3976 -864
rect 3460 -1012 3508 -988
rect 4502 -1074 4536 -864
rect 2392 -1144 2452 -1096
rect 4482 -1110 4536 -1074
rect -912 -3570 -860 -3566
rect -1374 -4922 -1298 -3594
rect -912 -3748 -858 -3570
rect -1126 -3792 -858 -3748
rect -2018 -5148 -1948 -4950
rect -1590 -5104 -1530 -4950
rect -1374 -5112 -1296 -4922
rect -1126 -4950 -1078 -3792
rect 1890 -4950 1950 -1358
rect -1374 -5114 -1306 -5112
rect -1126 -5184 -1076 -4950
rect 1890 -5178 1954 -4950
rect 2296 -5081 2374 -5060
rect 2296 -5133 2309 -5081
rect 2361 -5133 2374 -5081
rect 4582 -5102 4644 120
rect 6520 0 6560 1432
rect 6820 1408 6922 1446
rect 6820 1374 6859 1408
rect 6893 1374 6922 1408
rect 6820 1336 6922 1374
rect 6820 1302 6859 1336
rect 6893 1302 6922 1336
rect 6820 1264 6922 1302
rect 6820 1230 6859 1264
rect 6893 1230 6922 1264
rect 6820 1192 6922 1230
rect 6820 1158 6859 1192
rect 6893 1158 6922 1192
rect 6820 1120 6922 1158
rect 6820 1086 6859 1120
rect 6893 1086 6922 1120
rect 6986 1811 7060 1846
rect 6986 1777 7009 1811
rect 7043 1777 7060 1811
rect 6986 1739 7060 1777
rect 6986 1705 7009 1739
rect 7043 1705 7060 1739
rect 6986 1667 7060 1705
rect 6986 1633 7009 1667
rect 7043 1633 7060 1667
rect 6986 1595 7060 1633
rect 6986 1561 7009 1595
rect 7043 1561 7060 1595
rect 6986 1523 7060 1561
rect 6986 1489 7009 1523
rect 7043 1489 7060 1523
rect 6986 1451 7060 1489
rect 6986 1417 7009 1451
rect 7043 1417 7060 1451
rect 6986 1379 7060 1417
rect 6986 1345 7009 1379
rect 7043 1345 7060 1379
rect 6986 1307 7060 1345
rect 6986 1273 7009 1307
rect 7043 1273 7060 1307
rect 6986 1235 7060 1273
rect 6986 1201 7009 1235
rect 7043 1201 7060 1235
rect 6986 1163 7060 1201
rect 7126 1786 7808 1858
rect 7126 1222 7188 1786
rect 7752 1222 7808 1786
rect 7126 1168 7808 1222
rect 7874 1849 7899 1883
rect 7933 1849 7948 1883
rect 7874 1811 7948 1849
rect 7874 1777 7899 1811
rect 7933 1777 7948 1811
rect 7874 1739 7948 1777
rect 7874 1705 7899 1739
rect 7933 1705 7948 1739
rect 7874 1667 7948 1705
rect 7874 1633 7899 1667
rect 7933 1633 7948 1667
rect 7874 1595 7948 1633
rect 7874 1561 7899 1595
rect 7933 1561 7948 1595
rect 7874 1523 7948 1561
rect 7874 1489 7899 1523
rect 7933 1489 7948 1523
rect 7874 1451 7948 1489
rect 7874 1417 7899 1451
rect 7933 1417 7948 1451
rect 7874 1379 7948 1417
rect 7874 1345 7899 1379
rect 7933 1345 7948 1379
rect 7874 1307 7948 1345
rect 7874 1273 7899 1307
rect 7933 1273 7948 1307
rect 7874 1235 7948 1273
rect 7874 1201 7899 1235
rect 7933 1201 7948 1235
rect 6986 1129 7009 1163
rect 7043 1129 7060 1163
rect 6986 1098 7060 1129
rect 7874 1163 7948 1201
rect 7874 1129 7899 1163
rect 7933 1129 7948 1163
rect 6820 1048 6922 1086
rect 6820 1014 6859 1048
rect 6893 1014 6922 1048
rect 6980 1094 7066 1098
rect 7874 1094 7948 1129
rect 8014 1912 8116 1950
rect 8014 1878 8045 1912
rect 8079 1878 8116 1912
rect 8014 1840 8116 1878
rect 8014 1806 8045 1840
rect 8079 1806 8116 1840
rect 8014 1768 8116 1806
rect 8014 1734 8045 1768
rect 8079 1734 8116 1768
rect 8014 1696 8116 1734
rect 8014 1662 8045 1696
rect 8079 1662 8116 1696
rect 8014 1624 8116 1662
rect 8014 1590 8045 1624
rect 8079 1590 8116 1624
rect 8014 1552 8116 1590
rect 8014 1518 8045 1552
rect 8079 1518 8116 1552
rect 8900 1622 8992 1660
rect 8900 1570 8920 1622
rect 8972 1570 8992 1622
rect 8900 1542 8992 1570
rect 8014 1480 8116 1518
rect 8014 1446 8045 1480
rect 8079 1446 8116 1480
rect 8014 1408 8116 1446
rect 8014 1374 8045 1408
rect 8079 1374 8116 1408
rect 8014 1336 8116 1374
rect 8014 1302 8045 1336
rect 8079 1302 8116 1336
rect 8014 1264 8116 1302
rect 8014 1230 8045 1264
rect 8079 1230 8116 1264
rect 8014 1192 8116 1230
rect 12158 1302 12278 1334
rect 12158 1250 12184 1302
rect 12236 1250 12278 1302
rect 12158 1216 12278 1250
rect 8014 1158 8045 1192
rect 8079 1158 8116 1192
rect 8014 1120 8116 1158
rect 6980 1084 7950 1094
rect 6980 1032 6997 1084
rect 7049 1077 7950 1084
rect 7049 1043 7094 1077
rect 7128 1043 7166 1077
rect 7200 1043 7238 1077
rect 7272 1043 7310 1077
rect 7344 1043 7382 1077
rect 7416 1043 7454 1077
rect 7488 1043 7526 1077
rect 7560 1043 7598 1077
rect 7632 1043 7670 1077
rect 7704 1043 7742 1077
rect 7776 1043 7814 1077
rect 7848 1076 7950 1077
rect 7848 1043 7899 1076
rect 7049 1042 7899 1043
rect 7933 1042 7950 1076
rect 7049 1032 7950 1042
rect 6980 1026 7950 1032
rect 8014 1086 8045 1120
rect 8079 1086 8116 1120
rect 8014 1048 8116 1086
rect 6980 1024 7066 1026
rect 7874 1022 7948 1026
rect 6820 966 6922 1014
rect 8014 1014 8045 1048
rect 8079 1014 8116 1048
rect 8014 966 8116 1014
rect 6820 929 8118 966
rect 6820 895 6876 929
rect 6910 895 6948 929
rect 6982 895 7020 929
rect 7054 895 7092 929
rect 7126 895 7164 929
rect 7198 895 7236 929
rect 7270 895 7308 929
rect 7342 895 7380 929
rect 7414 895 7452 929
rect 7486 895 7524 929
rect 7558 895 7596 929
rect 7630 895 7668 929
rect 7702 895 7740 929
rect 7774 895 7812 929
rect 7846 895 7884 929
rect 7918 895 7956 929
rect 7990 895 8028 929
rect 8062 895 8118 929
rect 6820 886 8118 895
rect 13110 894 13216 898
rect 6818 860 8118 886
rect 13104 878 13216 894
rect 6818 852 6920 860
rect 6820 812 6920 852
rect 13104 826 13136 878
rect 13188 826 13216 878
rect 13104 820 13216 826
rect 4928 -42 6560 0
rect 4930 -66 6560 -42
rect 4930 -5100 5002 -66
rect 6520 -72 6560 -66
rect 6824 800 6920 812
rect 13110 804 13216 820
rect 6824 747 8122 800
rect 6824 713 6880 747
rect 6914 713 6952 747
rect 6986 713 7024 747
rect 7058 713 7096 747
rect 7130 713 7168 747
rect 7202 713 7240 747
rect 7274 713 7312 747
rect 7346 713 7384 747
rect 7418 713 7456 747
rect 7490 713 7528 747
rect 7562 713 7600 747
rect 7634 713 7672 747
rect 7706 713 7744 747
rect 7778 713 7816 747
rect 7850 713 7888 747
rect 7922 713 7960 747
rect 7994 713 8032 747
rect 8066 713 8122 747
rect 6824 694 8122 713
rect 13900 723 13988 726
rect 6824 628 6926 694
rect 6824 594 6863 628
rect 6897 594 6926 628
rect 6824 556 6926 594
rect 6990 613 7956 630
rect 6990 579 7023 613
rect 7057 579 7095 613
rect 7129 579 7167 613
rect 7201 579 7239 613
rect 7273 579 7311 613
rect 7345 579 7383 613
rect 7417 579 7455 613
rect 7489 579 7527 613
rect 7561 579 7599 613
rect 7633 579 7671 613
rect 7705 579 7743 613
rect 7777 579 7815 613
rect 7849 579 7956 613
rect 6990 578 7956 579
rect 6990 570 7004 578
rect 6824 522 6863 556
rect 6897 522 6926 556
rect 6824 484 6926 522
rect 6988 526 7004 570
rect 7056 562 7956 578
rect 8018 628 8120 694
rect 13900 671 13919 723
rect 13971 671 13988 723
rect 13900 664 13988 671
rect 8018 594 8049 628
rect 8083 594 8120 628
rect 7056 526 7066 562
rect 6988 493 7013 526
rect 7047 493 7066 526
rect 7878 527 7952 562
rect 6988 490 7066 493
rect 6824 450 6863 484
rect 6897 450 6926 484
rect 6824 412 6926 450
rect 6824 378 6863 412
rect 6897 378 6926 412
rect 6824 340 6926 378
rect 6824 306 6863 340
rect 6897 306 6926 340
rect 6824 268 6926 306
rect 6824 234 6863 268
rect 6897 234 6926 268
rect 6824 196 6926 234
rect 6824 162 6863 196
rect 6897 162 6926 196
rect 6824 124 6926 162
rect 6824 90 6863 124
rect 6897 90 6926 124
rect 6824 52 6926 90
rect 6824 18 6863 52
rect 6897 18 6926 52
rect 6824 -20 6926 18
rect 6824 -54 6863 -20
rect 6897 -54 6926 -20
rect 6824 -92 6926 -54
rect 6824 -126 6863 -92
rect 6897 -126 6926 -92
rect 6824 -164 6926 -126
rect 6824 -198 6863 -164
rect 6897 -198 6926 -164
rect 6824 -236 6926 -198
rect 6824 -270 6863 -236
rect 6897 -270 6926 -236
rect 6990 455 7064 490
rect 6990 421 7013 455
rect 7047 421 7064 455
rect 6990 383 7064 421
rect 6990 349 7013 383
rect 7047 349 7064 383
rect 6990 311 7064 349
rect 6990 277 7013 311
rect 7047 277 7064 311
rect 6990 239 7064 277
rect 6990 205 7013 239
rect 7047 205 7064 239
rect 6990 167 7064 205
rect 6990 133 7013 167
rect 7047 133 7064 167
rect 6990 95 7064 133
rect 6990 61 7013 95
rect 7047 61 7064 95
rect 6990 23 7064 61
rect 6990 -11 7013 23
rect 7047 -11 7064 23
rect 6990 -49 7064 -11
rect 6990 -83 7013 -49
rect 7047 -83 7064 -49
rect 6990 -121 7064 -83
rect 6990 -155 7013 -121
rect 7047 -155 7064 -121
rect 6990 -193 7064 -155
rect 7130 430 7812 502
rect 7130 -134 7192 430
rect 7756 -134 7812 430
rect 7130 -188 7812 -134
rect 7878 493 7903 527
rect 7937 493 7952 527
rect 7878 455 7952 493
rect 7878 421 7903 455
rect 7937 421 7952 455
rect 7878 383 7952 421
rect 7878 349 7903 383
rect 7937 349 7952 383
rect 7878 311 7952 349
rect 7878 277 7903 311
rect 7937 277 7952 311
rect 7878 239 7952 277
rect 7878 205 7903 239
rect 7937 205 7952 239
rect 7878 167 7952 205
rect 7878 133 7903 167
rect 7937 133 7952 167
rect 7878 95 7952 133
rect 7878 61 7903 95
rect 7937 61 7952 95
rect 7878 23 7952 61
rect 7878 -11 7903 23
rect 7937 -11 7952 23
rect 7878 -49 7952 -11
rect 7878 -83 7903 -49
rect 7937 -83 7952 -49
rect 7878 -121 7952 -83
rect 7878 -155 7903 -121
rect 7937 -155 7952 -121
rect 6990 -227 7013 -193
rect 7047 -227 7064 -193
rect 6990 -258 7064 -227
rect 7878 -193 7952 -155
rect 7878 -227 7903 -193
rect 7937 -227 7952 -193
rect 6824 -308 6926 -270
rect 6824 -342 6863 -308
rect 6897 -342 6926 -308
rect 6984 -262 7070 -258
rect 7878 -262 7952 -227
rect 8018 556 8120 594
rect 8018 522 8049 556
rect 8083 522 8120 556
rect 8018 484 8120 522
rect 8018 450 8049 484
rect 8083 450 8120 484
rect 8018 412 8120 450
rect 8018 378 8049 412
rect 8083 378 8120 412
rect 8018 340 8120 378
rect 8018 306 8049 340
rect 8083 306 8120 340
rect 8018 268 8120 306
rect 8018 234 8049 268
rect 8083 234 8120 268
rect 8018 196 8120 234
rect 8018 162 8049 196
rect 8083 162 8120 196
rect 8018 124 8120 162
rect 8018 90 8049 124
rect 8083 90 8120 124
rect 8018 52 8120 90
rect 8018 18 8049 52
rect 8083 18 8120 52
rect 8018 -20 8120 18
rect 8018 -54 8049 -20
rect 8083 -54 8120 -20
rect 8018 -92 8120 -54
rect 8018 -126 8049 -92
rect 8083 -126 8120 -92
rect 8018 -164 8120 -126
rect 8018 -198 8049 -164
rect 8083 -198 8120 -164
rect 8018 -236 8120 -198
rect 6984 -272 7954 -262
rect 6984 -324 7001 -272
rect 7053 -279 7954 -272
rect 7053 -313 7098 -279
rect 7132 -313 7170 -279
rect 7204 -313 7242 -279
rect 7276 -313 7314 -279
rect 7348 -313 7386 -279
rect 7420 -313 7458 -279
rect 7492 -313 7530 -279
rect 7564 -313 7602 -279
rect 7636 -313 7674 -279
rect 7708 -313 7746 -279
rect 7780 -313 7818 -279
rect 7852 -280 7954 -279
rect 7852 -313 7903 -280
rect 7053 -314 7903 -313
rect 7937 -314 7954 -280
rect 7053 -324 7954 -314
rect 6984 -330 7954 -324
rect 8018 -270 8049 -236
rect 8083 -270 8120 -236
rect 8018 -308 8120 -270
rect 6984 -332 7070 -330
rect 7878 -334 7952 -330
rect 6824 -390 6926 -342
rect 8018 -342 8049 -308
rect 8083 -342 8120 -308
rect 8018 -390 8120 -342
rect 6824 -427 8122 -390
rect 6824 -461 6880 -427
rect 6914 -461 6952 -427
rect 6986 -461 7024 -427
rect 7058 -461 7096 -427
rect 7130 -461 7168 -427
rect 7202 -461 7240 -427
rect 7274 -461 7312 -427
rect 7346 -461 7384 -427
rect 7418 -461 7456 -427
rect 7490 -461 7528 -427
rect 7562 -461 7600 -427
rect 7634 -461 7672 -427
rect 7706 -461 7744 -427
rect 7778 -461 7816 -427
rect 7850 -461 7888 -427
rect 7922 -461 7960 -427
rect 7994 -461 8032 -427
rect 8066 -461 8122 -427
rect 6824 -470 8122 -461
rect 6822 -494 8122 -470
rect 6820 -496 8122 -494
rect 6820 -550 6914 -496
rect 5410 -568 5506 -554
rect 6820 -564 6916 -550
rect 5410 -621 6708 -568
rect 5410 -655 5466 -621
rect 5500 -655 5538 -621
rect 5572 -655 5610 -621
rect 5644 -655 5682 -621
rect 5716 -655 5754 -621
rect 5788 -655 5826 -621
rect 5860 -655 5898 -621
rect 5932 -655 5970 -621
rect 6004 -655 6042 -621
rect 6076 -655 6114 -621
rect 6148 -655 6186 -621
rect 6220 -655 6258 -621
rect 6292 -655 6330 -621
rect 6364 -655 6402 -621
rect 6436 -655 6474 -621
rect 6508 -655 6546 -621
rect 6580 -655 6618 -621
rect 6652 -655 6708 -621
rect 5410 -674 6708 -655
rect 6820 -617 8118 -564
rect 6820 -651 6876 -617
rect 6910 -651 6948 -617
rect 6982 -651 7020 -617
rect 7054 -651 7092 -617
rect 7126 -651 7164 -617
rect 7198 -651 7236 -617
rect 7270 -651 7308 -617
rect 7342 -651 7380 -617
rect 7414 -651 7452 -617
rect 7486 -651 7524 -617
rect 7558 -651 7596 -617
rect 7630 -651 7668 -617
rect 7702 -651 7740 -617
rect 7774 -651 7812 -617
rect 7846 -651 7884 -617
rect 7918 -651 7956 -617
rect 7990 -651 8028 -617
rect 8062 -651 8118 -617
rect 6820 -670 8118 -651
rect 5410 -740 5512 -674
rect 5410 -774 5449 -740
rect 5483 -774 5512 -740
rect 5410 -812 5512 -774
rect 5576 -755 6542 -738
rect 5576 -789 5609 -755
rect 5643 -789 5681 -755
rect 5715 -789 5753 -755
rect 5787 -789 5825 -755
rect 5859 -789 5897 -755
rect 5931 -789 5969 -755
rect 6003 -789 6041 -755
rect 6075 -789 6113 -755
rect 6147 -789 6185 -755
rect 6219 -789 6257 -755
rect 6291 -789 6329 -755
rect 6363 -789 6401 -755
rect 6435 -789 6542 -755
rect 5576 -798 6542 -789
rect 5410 -846 5449 -812
rect 5483 -846 5512 -812
rect 5410 -884 5512 -846
rect 5574 -806 6542 -798
rect 6604 -740 6706 -674
rect 6604 -774 6635 -740
rect 6669 -774 6706 -740
rect 5574 -841 5652 -806
rect 5574 -875 5599 -841
rect 5633 -875 5652 -841
rect 6464 -841 6538 -806
rect 5574 -878 5652 -875
rect 5410 -918 5449 -884
rect 5483 -918 5512 -884
rect 5410 -956 5512 -918
rect 5410 -990 5449 -956
rect 5483 -990 5512 -956
rect 5410 -1028 5512 -990
rect 5410 -1062 5449 -1028
rect 5483 -1062 5512 -1028
rect 5410 -1100 5512 -1062
rect 5410 -1134 5449 -1100
rect 5483 -1134 5512 -1100
rect 5410 -1172 5512 -1134
rect 5410 -1206 5449 -1172
rect 5483 -1206 5512 -1172
rect 5410 -1244 5512 -1206
rect 5410 -1278 5449 -1244
rect 5483 -1278 5512 -1244
rect 5410 -1316 5512 -1278
rect 5410 -1350 5449 -1316
rect 5483 -1350 5512 -1316
rect 5410 -1388 5512 -1350
rect 5410 -1422 5449 -1388
rect 5483 -1422 5512 -1388
rect 5410 -1460 5512 -1422
rect 5410 -1494 5449 -1460
rect 5483 -1494 5512 -1460
rect 5410 -1532 5512 -1494
rect 5410 -1566 5449 -1532
rect 5483 -1566 5512 -1532
rect 5410 -1604 5512 -1566
rect 5410 -1638 5449 -1604
rect 5483 -1638 5512 -1604
rect 5576 -913 5650 -878
rect 5576 -947 5599 -913
rect 5633 -947 5650 -913
rect 5576 -985 5650 -947
rect 5576 -1019 5599 -985
rect 5633 -1019 5650 -985
rect 5576 -1057 5650 -1019
rect 5576 -1091 5599 -1057
rect 5633 -1091 5650 -1057
rect 5576 -1129 5650 -1091
rect 5576 -1163 5599 -1129
rect 5633 -1163 5650 -1129
rect 5576 -1201 5650 -1163
rect 5576 -1235 5599 -1201
rect 5633 -1235 5650 -1201
rect 5576 -1273 5650 -1235
rect 5576 -1307 5599 -1273
rect 5633 -1307 5650 -1273
rect 5576 -1345 5650 -1307
rect 5576 -1379 5599 -1345
rect 5633 -1379 5650 -1345
rect 5576 -1417 5650 -1379
rect 5576 -1451 5599 -1417
rect 5633 -1451 5650 -1417
rect 5576 -1489 5650 -1451
rect 5576 -1523 5599 -1489
rect 5633 -1523 5650 -1489
rect 5576 -1561 5650 -1523
rect 5716 -938 6398 -866
rect 5716 -1502 5778 -938
rect 6342 -1502 6398 -938
rect 5716 -1556 6398 -1502
rect 6464 -875 6489 -841
rect 6523 -875 6538 -841
rect 6464 -913 6538 -875
rect 6464 -947 6489 -913
rect 6523 -947 6538 -913
rect 6464 -985 6538 -947
rect 6464 -1019 6489 -985
rect 6523 -1019 6538 -985
rect 6464 -1057 6538 -1019
rect 6464 -1091 6489 -1057
rect 6523 -1091 6538 -1057
rect 6464 -1129 6538 -1091
rect 6464 -1163 6489 -1129
rect 6523 -1163 6538 -1129
rect 6464 -1201 6538 -1163
rect 6464 -1235 6489 -1201
rect 6523 -1235 6538 -1201
rect 6464 -1273 6538 -1235
rect 6464 -1307 6489 -1273
rect 6523 -1307 6538 -1273
rect 6464 -1345 6538 -1307
rect 6464 -1379 6489 -1345
rect 6523 -1379 6538 -1345
rect 6464 -1417 6538 -1379
rect 6464 -1451 6489 -1417
rect 6523 -1451 6538 -1417
rect 6464 -1489 6538 -1451
rect 6464 -1523 6489 -1489
rect 6523 -1523 6538 -1489
rect 5576 -1595 5599 -1561
rect 5633 -1595 5650 -1561
rect 5576 -1626 5650 -1595
rect 6464 -1561 6538 -1523
rect 6464 -1595 6489 -1561
rect 6523 -1595 6538 -1561
rect 5410 -1676 5512 -1638
rect 5410 -1710 5449 -1676
rect 5483 -1710 5512 -1676
rect 5570 -1630 5656 -1626
rect 6464 -1630 6538 -1595
rect 6604 -812 6706 -774
rect 6604 -846 6635 -812
rect 6669 -846 6706 -812
rect 6604 -884 6706 -846
rect 6604 -918 6635 -884
rect 6669 -918 6706 -884
rect 6604 -956 6706 -918
rect 6604 -990 6635 -956
rect 6669 -990 6706 -956
rect 6604 -1028 6706 -990
rect 6604 -1062 6635 -1028
rect 6669 -1062 6706 -1028
rect 6604 -1100 6706 -1062
rect 6604 -1134 6635 -1100
rect 6669 -1134 6706 -1100
rect 6604 -1172 6706 -1134
rect 6604 -1206 6635 -1172
rect 6669 -1206 6706 -1172
rect 6604 -1244 6706 -1206
rect 6604 -1278 6635 -1244
rect 6669 -1278 6706 -1244
rect 6604 -1316 6706 -1278
rect 6604 -1350 6635 -1316
rect 6669 -1350 6706 -1316
rect 6604 -1388 6706 -1350
rect 6604 -1422 6635 -1388
rect 6669 -1422 6706 -1388
rect 6604 -1460 6706 -1422
rect 6604 -1494 6635 -1460
rect 6669 -1494 6706 -1460
rect 6604 -1532 6706 -1494
rect 6604 -1566 6635 -1532
rect 6669 -1566 6706 -1532
rect 6604 -1604 6706 -1566
rect 5570 -1640 6540 -1630
rect 5570 -1692 5587 -1640
rect 5639 -1647 6540 -1640
rect 5639 -1681 5684 -1647
rect 5718 -1681 5756 -1647
rect 5790 -1681 5828 -1647
rect 5862 -1681 5900 -1647
rect 5934 -1681 5972 -1647
rect 6006 -1681 6044 -1647
rect 6078 -1681 6116 -1647
rect 6150 -1681 6188 -1647
rect 6222 -1681 6260 -1647
rect 6294 -1681 6332 -1647
rect 6366 -1681 6404 -1647
rect 6438 -1648 6540 -1647
rect 6438 -1681 6489 -1648
rect 5639 -1682 6489 -1681
rect 6523 -1682 6540 -1648
rect 5639 -1692 6540 -1682
rect 5570 -1698 6540 -1692
rect 6604 -1638 6635 -1604
rect 6669 -1638 6706 -1604
rect 6604 -1676 6706 -1638
rect 5570 -1700 5656 -1698
rect 6464 -1702 6538 -1698
rect 5410 -1758 5512 -1710
rect 6604 -1710 6635 -1676
rect 6669 -1710 6706 -1676
rect 6604 -1758 6706 -1710
rect 6820 -736 6922 -670
rect 6820 -770 6859 -736
rect 6893 -770 6922 -736
rect 6820 -808 6922 -770
rect 6986 -751 7952 -734
rect 6986 -785 7019 -751
rect 7053 -785 7091 -751
rect 7125 -785 7163 -751
rect 7197 -785 7235 -751
rect 7269 -785 7307 -751
rect 7341 -785 7379 -751
rect 7413 -785 7451 -751
rect 7485 -785 7523 -751
rect 7557 -785 7595 -751
rect 7629 -785 7667 -751
rect 7701 -785 7739 -751
rect 7773 -785 7811 -751
rect 7845 -785 7952 -751
rect 6986 -786 7952 -785
rect 6986 -794 7002 -786
rect 6820 -842 6859 -808
rect 6893 -842 6922 -808
rect 6820 -880 6922 -842
rect 6984 -838 7002 -794
rect 7054 -802 7952 -786
rect 8014 -736 8116 -670
rect 8014 -770 8045 -736
rect 8079 -770 8116 -736
rect 7054 -838 7062 -802
rect 6984 -871 7009 -838
rect 7043 -871 7062 -838
rect 7874 -837 7948 -802
rect 6984 -874 7062 -871
rect 6820 -914 6859 -880
rect 6893 -914 6922 -880
rect 6820 -952 6922 -914
rect 6820 -986 6859 -952
rect 6893 -986 6922 -952
rect 6820 -1024 6922 -986
rect 6820 -1058 6859 -1024
rect 6893 -1058 6922 -1024
rect 6820 -1096 6922 -1058
rect 6820 -1130 6859 -1096
rect 6893 -1130 6922 -1096
rect 6820 -1168 6922 -1130
rect 6820 -1202 6859 -1168
rect 6893 -1202 6922 -1168
rect 6820 -1240 6922 -1202
rect 6820 -1274 6859 -1240
rect 6893 -1274 6922 -1240
rect 6820 -1312 6922 -1274
rect 6820 -1346 6859 -1312
rect 6893 -1346 6922 -1312
rect 6820 -1384 6922 -1346
rect 6820 -1418 6859 -1384
rect 6893 -1418 6922 -1384
rect 6820 -1456 6922 -1418
rect 6820 -1490 6859 -1456
rect 6893 -1490 6922 -1456
rect 6820 -1528 6922 -1490
rect 6820 -1562 6859 -1528
rect 6893 -1562 6922 -1528
rect 6820 -1600 6922 -1562
rect 6820 -1634 6859 -1600
rect 6893 -1634 6922 -1600
rect 6986 -909 7060 -874
rect 6986 -943 7009 -909
rect 7043 -943 7060 -909
rect 6986 -981 7060 -943
rect 6986 -1015 7009 -981
rect 7043 -1015 7060 -981
rect 6986 -1053 7060 -1015
rect 6986 -1087 7009 -1053
rect 7043 -1087 7060 -1053
rect 6986 -1125 7060 -1087
rect 6986 -1159 7009 -1125
rect 7043 -1159 7060 -1125
rect 6986 -1197 7060 -1159
rect 6986 -1231 7009 -1197
rect 7043 -1231 7060 -1197
rect 6986 -1269 7060 -1231
rect 6986 -1303 7009 -1269
rect 7043 -1303 7060 -1269
rect 6986 -1341 7060 -1303
rect 6986 -1375 7009 -1341
rect 7043 -1375 7060 -1341
rect 6986 -1413 7060 -1375
rect 6986 -1447 7009 -1413
rect 7043 -1447 7060 -1413
rect 6986 -1485 7060 -1447
rect 6986 -1519 7009 -1485
rect 7043 -1519 7060 -1485
rect 6986 -1557 7060 -1519
rect 7126 -934 7808 -862
rect 7126 -1498 7188 -934
rect 7752 -1498 7808 -934
rect 7126 -1552 7808 -1498
rect 7874 -871 7899 -837
rect 7933 -871 7948 -837
rect 7874 -909 7948 -871
rect 7874 -943 7899 -909
rect 7933 -943 7948 -909
rect 7874 -981 7948 -943
rect 7874 -1015 7899 -981
rect 7933 -1015 7948 -981
rect 7874 -1053 7948 -1015
rect 7874 -1087 7899 -1053
rect 7933 -1087 7948 -1053
rect 7874 -1125 7948 -1087
rect 7874 -1159 7899 -1125
rect 7933 -1159 7948 -1125
rect 7874 -1197 7948 -1159
rect 7874 -1231 7899 -1197
rect 7933 -1231 7948 -1197
rect 7874 -1269 7948 -1231
rect 7874 -1303 7899 -1269
rect 7933 -1303 7948 -1269
rect 7874 -1341 7948 -1303
rect 7874 -1375 7899 -1341
rect 7933 -1375 7948 -1341
rect 7874 -1413 7948 -1375
rect 7874 -1447 7899 -1413
rect 7933 -1447 7948 -1413
rect 7874 -1485 7948 -1447
rect 7874 -1519 7899 -1485
rect 7933 -1519 7948 -1485
rect 6986 -1591 7009 -1557
rect 7043 -1591 7060 -1557
rect 6986 -1622 7060 -1591
rect 7874 -1557 7948 -1519
rect 7874 -1591 7899 -1557
rect 7933 -1591 7948 -1557
rect 6820 -1672 6922 -1634
rect 6820 -1706 6859 -1672
rect 6893 -1706 6922 -1672
rect 6980 -1626 7066 -1622
rect 7874 -1626 7948 -1591
rect 8014 -808 8116 -770
rect 8014 -842 8045 -808
rect 8079 -842 8116 -808
rect 8014 -880 8116 -842
rect 8014 -914 8045 -880
rect 8079 -914 8116 -880
rect 8014 -952 8116 -914
rect 8014 -986 8045 -952
rect 8079 -986 8116 -952
rect 8014 -1024 8116 -986
rect 8014 -1058 8045 -1024
rect 8079 -1058 8116 -1024
rect 8014 -1096 8116 -1058
rect 8014 -1130 8045 -1096
rect 8079 -1130 8116 -1096
rect 8014 -1168 8116 -1130
rect 8014 -1202 8045 -1168
rect 8079 -1202 8116 -1168
rect 8014 -1240 8116 -1202
rect 8014 -1274 8045 -1240
rect 8079 -1274 8116 -1240
rect 8014 -1312 8116 -1274
rect 8014 -1346 8045 -1312
rect 8079 -1346 8116 -1312
rect 8014 -1384 8116 -1346
rect 8014 -1418 8045 -1384
rect 8079 -1418 8116 -1384
rect 8014 -1456 8116 -1418
rect 8014 -1490 8045 -1456
rect 8079 -1490 8116 -1456
rect 8014 -1528 8116 -1490
rect 8014 -1562 8045 -1528
rect 8079 -1562 8116 -1528
rect 8014 -1600 8116 -1562
rect 6980 -1636 7950 -1626
rect 6980 -1688 6997 -1636
rect 7049 -1643 7950 -1636
rect 7049 -1677 7094 -1643
rect 7128 -1677 7166 -1643
rect 7200 -1677 7238 -1643
rect 7272 -1677 7310 -1643
rect 7344 -1677 7382 -1643
rect 7416 -1677 7454 -1643
rect 7488 -1677 7526 -1643
rect 7560 -1677 7598 -1643
rect 7632 -1677 7670 -1643
rect 7704 -1677 7742 -1643
rect 7776 -1677 7814 -1643
rect 7848 -1644 7950 -1643
rect 7848 -1677 7899 -1644
rect 7049 -1678 7899 -1677
rect 7933 -1678 7950 -1644
rect 7049 -1688 7950 -1678
rect 6980 -1694 7950 -1688
rect 8014 -1634 8045 -1600
rect 8079 -1634 8116 -1600
rect 8014 -1672 8116 -1634
rect 6980 -1696 7066 -1694
rect 7874 -1698 7948 -1694
rect 6820 -1754 6922 -1706
rect 8014 -1706 8045 -1672
rect 8079 -1706 8116 -1672
rect 8014 -1754 8116 -1706
rect 5410 -1795 6708 -1758
rect 5410 -1829 5466 -1795
rect 5500 -1829 5538 -1795
rect 5572 -1829 5610 -1795
rect 5644 -1829 5682 -1795
rect 5716 -1829 5754 -1795
rect 5788 -1829 5826 -1795
rect 5860 -1829 5898 -1795
rect 5932 -1829 5970 -1795
rect 6004 -1829 6042 -1795
rect 6076 -1829 6114 -1795
rect 6148 -1829 6186 -1795
rect 6220 -1829 6258 -1795
rect 6292 -1829 6330 -1795
rect 6364 -1829 6402 -1795
rect 6436 -1829 6474 -1795
rect 6508 -1829 6546 -1795
rect 6580 -1829 6618 -1795
rect 6652 -1829 6708 -1795
rect 5410 -1838 6708 -1829
rect 6820 -1791 8118 -1754
rect 6820 -1825 6876 -1791
rect 6910 -1825 6948 -1791
rect 6982 -1825 7020 -1791
rect 7054 -1825 7092 -1791
rect 7126 -1825 7164 -1791
rect 7198 -1825 7236 -1791
rect 7270 -1825 7308 -1791
rect 7342 -1825 7380 -1791
rect 7414 -1825 7452 -1791
rect 7486 -1825 7524 -1791
rect 7558 -1825 7596 -1791
rect 7630 -1825 7668 -1791
rect 7702 -1825 7740 -1791
rect 7774 -1825 7812 -1791
rect 7846 -1825 7884 -1791
rect 7918 -1825 7956 -1791
rect 7990 -1825 8028 -1791
rect 8062 -1825 8118 -1791
rect 6820 -1834 8118 -1825
rect 5408 -1864 6708 -1838
rect 6818 -1860 8118 -1834
rect 5408 -1872 5500 -1864
rect 6818 -1868 6916 -1860
rect 5410 -1910 5500 -1872
rect 6820 -1908 6916 -1868
rect 6820 -1910 6918 -1908
rect 5408 -1924 5504 -1910
rect 6822 -1922 6918 -1910
rect 5408 -1977 6706 -1924
rect 5408 -2011 5464 -1977
rect 5498 -2011 5536 -1977
rect 5570 -2011 5608 -1977
rect 5642 -2011 5680 -1977
rect 5714 -2011 5752 -1977
rect 5786 -2011 5824 -1977
rect 5858 -2011 5896 -1977
rect 5930 -2011 5968 -1977
rect 6002 -2011 6040 -1977
rect 6074 -2011 6112 -1977
rect 6146 -2011 6184 -1977
rect 6218 -2011 6256 -1977
rect 6290 -2011 6328 -1977
rect 6362 -2011 6400 -1977
rect 6434 -2011 6472 -1977
rect 6506 -2011 6544 -1977
rect 6578 -2011 6616 -1977
rect 6650 -2011 6706 -1977
rect 5408 -2030 6706 -2011
rect 6822 -1975 8120 -1922
rect 6822 -2009 6878 -1975
rect 6912 -2009 6950 -1975
rect 6984 -2009 7022 -1975
rect 7056 -2009 7094 -1975
rect 7128 -2009 7166 -1975
rect 7200 -2009 7238 -1975
rect 7272 -2009 7310 -1975
rect 7344 -2009 7382 -1975
rect 7416 -2009 7454 -1975
rect 7488 -2009 7526 -1975
rect 7560 -2009 7598 -1975
rect 7632 -2009 7670 -1975
rect 7704 -2009 7742 -1975
rect 7776 -2009 7814 -1975
rect 7848 -2009 7886 -1975
rect 7920 -2009 7958 -1975
rect 7992 -2009 8030 -1975
rect 8064 -2009 8120 -1975
rect 6822 -2028 8120 -2009
rect 5408 -2096 5510 -2030
rect 5408 -2130 5447 -2096
rect 5481 -2130 5510 -2096
rect 5408 -2168 5510 -2130
rect 5574 -2111 6540 -2094
rect 5574 -2145 5607 -2111
rect 5641 -2145 5679 -2111
rect 5713 -2145 5751 -2111
rect 5785 -2145 5823 -2111
rect 5857 -2145 5895 -2111
rect 5929 -2145 5967 -2111
rect 6001 -2145 6039 -2111
rect 6073 -2145 6111 -2111
rect 6145 -2145 6183 -2111
rect 6217 -2145 6255 -2111
rect 6289 -2145 6327 -2111
rect 6361 -2145 6399 -2111
rect 6433 -2145 6540 -2111
rect 5574 -2150 6540 -2145
rect 5574 -2154 5590 -2150
rect 5408 -2202 5447 -2168
rect 5481 -2202 5510 -2168
rect 5408 -2240 5510 -2202
rect 5572 -2202 5590 -2154
rect 5642 -2162 6540 -2150
rect 6602 -2096 6704 -2030
rect 6602 -2130 6633 -2096
rect 6667 -2130 6704 -2096
rect 5642 -2202 5650 -2162
rect 5572 -2231 5597 -2202
rect 5631 -2231 5650 -2202
rect 6462 -2197 6536 -2162
rect 5572 -2234 5650 -2231
rect 5408 -2274 5447 -2240
rect 5481 -2274 5510 -2240
rect 5408 -2312 5510 -2274
rect 5408 -2346 5447 -2312
rect 5481 -2346 5510 -2312
rect 5408 -2384 5510 -2346
rect 5408 -2418 5447 -2384
rect 5481 -2418 5510 -2384
rect 5408 -2456 5510 -2418
rect 5408 -2490 5447 -2456
rect 5481 -2490 5510 -2456
rect 5408 -2528 5510 -2490
rect 5408 -2562 5447 -2528
rect 5481 -2562 5510 -2528
rect 5408 -2600 5510 -2562
rect 5408 -2634 5447 -2600
rect 5481 -2634 5510 -2600
rect 5408 -2672 5510 -2634
rect 5408 -2706 5447 -2672
rect 5481 -2706 5510 -2672
rect 5408 -2744 5510 -2706
rect 5408 -2778 5447 -2744
rect 5481 -2778 5510 -2744
rect 5408 -2816 5510 -2778
rect 5408 -2850 5447 -2816
rect 5481 -2850 5510 -2816
rect 5408 -2888 5510 -2850
rect 5408 -2922 5447 -2888
rect 5481 -2922 5510 -2888
rect 5408 -2960 5510 -2922
rect 5408 -2994 5447 -2960
rect 5481 -2994 5510 -2960
rect 5574 -2269 5648 -2234
rect 5574 -2303 5597 -2269
rect 5631 -2303 5648 -2269
rect 5574 -2341 5648 -2303
rect 5574 -2375 5597 -2341
rect 5631 -2375 5648 -2341
rect 5574 -2413 5648 -2375
rect 5574 -2447 5597 -2413
rect 5631 -2447 5648 -2413
rect 5574 -2485 5648 -2447
rect 5574 -2519 5597 -2485
rect 5631 -2519 5648 -2485
rect 5574 -2557 5648 -2519
rect 5574 -2591 5597 -2557
rect 5631 -2591 5648 -2557
rect 5574 -2629 5648 -2591
rect 5574 -2663 5597 -2629
rect 5631 -2663 5648 -2629
rect 5574 -2701 5648 -2663
rect 5574 -2735 5597 -2701
rect 5631 -2735 5648 -2701
rect 5574 -2773 5648 -2735
rect 5574 -2807 5597 -2773
rect 5631 -2807 5648 -2773
rect 5574 -2845 5648 -2807
rect 5574 -2879 5597 -2845
rect 5631 -2879 5648 -2845
rect 5574 -2917 5648 -2879
rect 5714 -2294 6396 -2222
rect 5714 -2858 5776 -2294
rect 6340 -2858 6396 -2294
rect 5714 -2912 6396 -2858
rect 6462 -2231 6487 -2197
rect 6521 -2231 6536 -2197
rect 6462 -2269 6536 -2231
rect 6462 -2303 6487 -2269
rect 6521 -2303 6536 -2269
rect 6462 -2341 6536 -2303
rect 6462 -2375 6487 -2341
rect 6521 -2375 6536 -2341
rect 6462 -2413 6536 -2375
rect 6462 -2447 6487 -2413
rect 6521 -2447 6536 -2413
rect 6462 -2485 6536 -2447
rect 6462 -2519 6487 -2485
rect 6521 -2519 6536 -2485
rect 6462 -2557 6536 -2519
rect 6462 -2591 6487 -2557
rect 6521 -2591 6536 -2557
rect 6462 -2629 6536 -2591
rect 6462 -2663 6487 -2629
rect 6521 -2663 6536 -2629
rect 6462 -2701 6536 -2663
rect 6462 -2735 6487 -2701
rect 6521 -2735 6536 -2701
rect 6462 -2773 6536 -2735
rect 6462 -2807 6487 -2773
rect 6521 -2807 6536 -2773
rect 6462 -2845 6536 -2807
rect 6462 -2879 6487 -2845
rect 6521 -2879 6536 -2845
rect 5574 -2951 5597 -2917
rect 5631 -2951 5648 -2917
rect 5574 -2982 5648 -2951
rect 6462 -2917 6536 -2879
rect 6462 -2951 6487 -2917
rect 6521 -2951 6536 -2917
rect 5408 -3032 5510 -2994
rect 5408 -3066 5447 -3032
rect 5481 -3066 5510 -3032
rect 5570 -2986 5652 -2982
rect 6462 -2986 6536 -2951
rect 6602 -2168 6704 -2130
rect 6602 -2202 6633 -2168
rect 6667 -2202 6704 -2168
rect 6602 -2240 6704 -2202
rect 6602 -2274 6633 -2240
rect 6667 -2274 6704 -2240
rect 6602 -2312 6704 -2274
rect 6602 -2346 6633 -2312
rect 6667 -2346 6704 -2312
rect 6602 -2384 6704 -2346
rect 6602 -2418 6633 -2384
rect 6667 -2418 6704 -2384
rect 6602 -2456 6704 -2418
rect 6602 -2490 6633 -2456
rect 6667 -2490 6704 -2456
rect 6602 -2528 6704 -2490
rect 6602 -2562 6633 -2528
rect 6667 -2562 6704 -2528
rect 6602 -2600 6704 -2562
rect 6602 -2634 6633 -2600
rect 6667 -2634 6704 -2600
rect 6602 -2672 6704 -2634
rect 6602 -2706 6633 -2672
rect 6667 -2706 6704 -2672
rect 6602 -2744 6704 -2706
rect 6602 -2778 6633 -2744
rect 6667 -2778 6704 -2744
rect 6602 -2816 6704 -2778
rect 6602 -2850 6633 -2816
rect 6667 -2850 6704 -2816
rect 6602 -2888 6704 -2850
rect 6602 -2922 6633 -2888
rect 6667 -2922 6704 -2888
rect 6602 -2960 6704 -2922
rect 5570 -2996 6538 -2986
rect 5570 -3048 5585 -2996
rect 5637 -3003 6538 -2996
rect 5637 -3037 5682 -3003
rect 5716 -3037 5754 -3003
rect 5788 -3037 5826 -3003
rect 5860 -3037 5898 -3003
rect 5932 -3037 5970 -3003
rect 6004 -3037 6042 -3003
rect 6076 -3037 6114 -3003
rect 6148 -3037 6186 -3003
rect 6220 -3037 6258 -3003
rect 6292 -3037 6330 -3003
rect 6364 -3037 6402 -3003
rect 6436 -3004 6538 -3003
rect 6436 -3037 6487 -3004
rect 5637 -3038 6487 -3037
rect 6521 -3038 6538 -3004
rect 5637 -3048 6538 -3038
rect 5570 -3054 6538 -3048
rect 6602 -2994 6633 -2960
rect 6667 -2994 6704 -2960
rect 6602 -3032 6704 -2994
rect 6462 -3058 6536 -3054
rect 5408 -3114 5510 -3066
rect 6602 -3066 6633 -3032
rect 6667 -3066 6704 -3032
rect 6602 -3114 6704 -3066
rect 6822 -2094 6924 -2028
rect 6822 -2128 6861 -2094
rect 6895 -2128 6924 -2094
rect 6822 -2166 6924 -2128
rect 6988 -2109 7954 -2092
rect 6988 -2143 7021 -2109
rect 7055 -2143 7093 -2109
rect 7127 -2143 7165 -2109
rect 7199 -2143 7237 -2109
rect 7271 -2143 7309 -2109
rect 7343 -2143 7381 -2109
rect 7415 -2143 7453 -2109
rect 7487 -2143 7525 -2109
rect 7559 -2143 7597 -2109
rect 7631 -2143 7669 -2109
rect 7703 -2143 7741 -2109
rect 7775 -2143 7813 -2109
rect 7847 -2143 7954 -2109
rect 6988 -2152 7954 -2143
rect 6822 -2200 6861 -2166
rect 6895 -2200 6924 -2166
rect 6822 -2238 6924 -2200
rect 6986 -2154 7954 -2152
rect 6986 -2206 7000 -2154
rect 7052 -2160 7954 -2154
rect 8016 -2094 8118 -2028
rect 8016 -2128 8047 -2094
rect 8081 -2128 8118 -2094
rect 7052 -2206 7064 -2160
rect 6986 -2229 7011 -2206
rect 7045 -2229 7064 -2206
rect 7876 -2195 7950 -2160
rect 6986 -2232 7064 -2229
rect 6822 -2272 6861 -2238
rect 6895 -2272 6924 -2238
rect 6822 -2310 6924 -2272
rect 6822 -2344 6861 -2310
rect 6895 -2344 6924 -2310
rect 6822 -2382 6924 -2344
rect 6822 -2416 6861 -2382
rect 6895 -2416 6924 -2382
rect 6822 -2454 6924 -2416
rect 6822 -2488 6861 -2454
rect 6895 -2488 6924 -2454
rect 6822 -2526 6924 -2488
rect 6822 -2560 6861 -2526
rect 6895 -2560 6924 -2526
rect 6822 -2598 6924 -2560
rect 6822 -2632 6861 -2598
rect 6895 -2632 6924 -2598
rect 6822 -2670 6924 -2632
rect 6822 -2704 6861 -2670
rect 6895 -2704 6924 -2670
rect 6822 -2742 6924 -2704
rect 6822 -2776 6861 -2742
rect 6895 -2776 6924 -2742
rect 6822 -2814 6924 -2776
rect 6822 -2848 6861 -2814
rect 6895 -2848 6924 -2814
rect 6822 -2886 6924 -2848
rect 6822 -2920 6861 -2886
rect 6895 -2920 6924 -2886
rect 6822 -2958 6924 -2920
rect 6822 -2992 6861 -2958
rect 6895 -2992 6924 -2958
rect 6988 -2267 7062 -2232
rect 6988 -2301 7011 -2267
rect 7045 -2301 7062 -2267
rect 6988 -2339 7062 -2301
rect 6988 -2373 7011 -2339
rect 7045 -2373 7062 -2339
rect 6988 -2411 7062 -2373
rect 6988 -2445 7011 -2411
rect 7045 -2445 7062 -2411
rect 6988 -2483 7062 -2445
rect 6988 -2517 7011 -2483
rect 7045 -2517 7062 -2483
rect 6988 -2555 7062 -2517
rect 6988 -2589 7011 -2555
rect 7045 -2589 7062 -2555
rect 6988 -2627 7062 -2589
rect 6988 -2661 7011 -2627
rect 7045 -2661 7062 -2627
rect 6988 -2699 7062 -2661
rect 6988 -2733 7011 -2699
rect 7045 -2733 7062 -2699
rect 6988 -2771 7062 -2733
rect 6988 -2805 7011 -2771
rect 7045 -2805 7062 -2771
rect 6988 -2843 7062 -2805
rect 6988 -2877 7011 -2843
rect 7045 -2877 7062 -2843
rect 6988 -2915 7062 -2877
rect 7128 -2292 7810 -2220
rect 7128 -2856 7190 -2292
rect 7754 -2856 7810 -2292
rect 7128 -2910 7810 -2856
rect 7876 -2229 7901 -2195
rect 7935 -2229 7950 -2195
rect 7876 -2267 7950 -2229
rect 7876 -2301 7901 -2267
rect 7935 -2301 7950 -2267
rect 7876 -2339 7950 -2301
rect 7876 -2373 7901 -2339
rect 7935 -2373 7950 -2339
rect 7876 -2411 7950 -2373
rect 7876 -2445 7901 -2411
rect 7935 -2445 7950 -2411
rect 7876 -2483 7950 -2445
rect 7876 -2517 7901 -2483
rect 7935 -2517 7950 -2483
rect 7876 -2555 7950 -2517
rect 7876 -2589 7901 -2555
rect 7935 -2589 7950 -2555
rect 7876 -2627 7950 -2589
rect 7876 -2661 7901 -2627
rect 7935 -2661 7950 -2627
rect 7876 -2699 7950 -2661
rect 7876 -2733 7901 -2699
rect 7935 -2733 7950 -2699
rect 7876 -2771 7950 -2733
rect 7876 -2805 7901 -2771
rect 7935 -2805 7950 -2771
rect 7876 -2843 7950 -2805
rect 7876 -2877 7901 -2843
rect 7935 -2877 7950 -2843
rect 6988 -2949 7011 -2915
rect 7045 -2949 7062 -2915
rect 6988 -2980 7062 -2949
rect 7876 -2915 7950 -2877
rect 7876 -2949 7901 -2915
rect 7935 -2949 7950 -2915
rect 6822 -3030 6924 -2992
rect 6822 -3064 6861 -3030
rect 6895 -3064 6924 -3030
rect 6982 -2984 7068 -2980
rect 7876 -2984 7950 -2949
rect 8016 -2166 8118 -2128
rect 8016 -2200 8047 -2166
rect 8081 -2200 8118 -2166
rect 8016 -2238 8118 -2200
rect 8016 -2272 8047 -2238
rect 8081 -2272 8118 -2238
rect 8016 -2310 8118 -2272
rect 8016 -2344 8047 -2310
rect 8081 -2344 8118 -2310
rect 8016 -2382 8118 -2344
rect 8016 -2416 8047 -2382
rect 8081 -2416 8118 -2382
rect 8016 -2454 8118 -2416
rect 8016 -2488 8047 -2454
rect 8081 -2488 8118 -2454
rect 8016 -2526 8118 -2488
rect 8016 -2560 8047 -2526
rect 8081 -2560 8118 -2526
rect 8016 -2598 8118 -2560
rect 8016 -2632 8047 -2598
rect 8081 -2632 8118 -2598
rect 8016 -2670 8118 -2632
rect 8016 -2704 8047 -2670
rect 8081 -2704 8118 -2670
rect 8016 -2742 8118 -2704
rect 8016 -2776 8047 -2742
rect 8081 -2776 8118 -2742
rect 8016 -2814 8118 -2776
rect 8016 -2848 8047 -2814
rect 8081 -2848 8118 -2814
rect 8016 -2886 8118 -2848
rect 8016 -2920 8047 -2886
rect 8081 -2920 8118 -2886
rect 8016 -2958 8118 -2920
rect 6982 -2994 7952 -2984
rect 6982 -3046 6999 -2994
rect 7051 -3001 7952 -2994
rect 7051 -3035 7096 -3001
rect 7130 -3035 7168 -3001
rect 7202 -3035 7240 -3001
rect 7274 -3035 7312 -3001
rect 7346 -3035 7384 -3001
rect 7418 -3035 7456 -3001
rect 7490 -3035 7528 -3001
rect 7562 -3035 7600 -3001
rect 7634 -3035 7672 -3001
rect 7706 -3035 7744 -3001
rect 7778 -3035 7816 -3001
rect 7850 -3002 7952 -3001
rect 7850 -3035 7901 -3002
rect 7051 -3036 7901 -3035
rect 7935 -3036 7952 -3002
rect 7051 -3046 7952 -3036
rect 6982 -3052 7952 -3046
rect 8016 -2992 8047 -2958
rect 8081 -2992 8118 -2958
rect 8016 -3030 8118 -2992
rect 6982 -3054 7068 -3052
rect 7876 -3056 7950 -3052
rect 6822 -3112 6924 -3064
rect 8016 -3064 8047 -3030
rect 8081 -3064 8118 -3030
rect 8016 -3112 8118 -3064
rect 5408 -3151 6706 -3114
rect 5408 -3185 5464 -3151
rect 5498 -3185 5536 -3151
rect 5570 -3185 5608 -3151
rect 5642 -3185 5680 -3151
rect 5714 -3185 5752 -3151
rect 5786 -3185 5824 -3151
rect 5858 -3185 5896 -3151
rect 5930 -3185 5968 -3151
rect 6002 -3185 6040 -3151
rect 6074 -3185 6112 -3151
rect 6146 -3185 6184 -3151
rect 6218 -3185 6256 -3151
rect 6290 -3185 6328 -3151
rect 6362 -3185 6400 -3151
rect 6434 -3185 6472 -3151
rect 6506 -3185 6544 -3151
rect 6578 -3185 6616 -3151
rect 6650 -3185 6706 -3151
rect 5408 -3194 6706 -3185
rect 6822 -3149 8120 -3112
rect 6822 -3183 6878 -3149
rect 6912 -3183 6950 -3149
rect 6984 -3183 7022 -3149
rect 7056 -3183 7094 -3149
rect 7128 -3183 7166 -3149
rect 7200 -3183 7238 -3149
rect 7272 -3183 7310 -3149
rect 7344 -3183 7382 -3149
rect 7416 -3183 7454 -3149
rect 7488 -3183 7526 -3149
rect 7560 -3183 7598 -3149
rect 7632 -3183 7670 -3149
rect 7704 -3183 7742 -3149
rect 7776 -3183 7814 -3149
rect 7848 -3183 7886 -3149
rect 7920 -3183 7958 -3149
rect 7992 -3183 8030 -3149
rect 8064 -3183 8120 -3149
rect 6822 -3192 8120 -3183
rect 9230 -3150 9270 -2108
rect 10136 -2260 10316 -2204
rect 10280 -2384 10316 -2260
rect 10280 -2420 10526 -2384
rect 9912 -2844 9960 -2662
rect 9912 -2896 10150 -2844
rect 10128 -3072 10180 -2954
rect 10128 -3074 10182 -3072
rect 9986 -3118 10182 -3074
rect 9230 -3188 9628 -3150
rect 9230 -3190 9380 -3188
rect 5406 -3220 6706 -3194
rect 6820 -3218 8120 -3192
rect 5406 -3228 5498 -3220
rect 6820 -3226 6910 -3218
rect 5408 -3262 5498 -3228
rect 5408 -3276 5504 -3262
rect 6822 -3268 6910 -3226
rect 6822 -3272 6920 -3268
rect 5408 -3329 6706 -3276
rect 5408 -3363 5464 -3329
rect 5498 -3363 5536 -3329
rect 5570 -3363 5608 -3329
rect 5642 -3363 5680 -3329
rect 5714 -3363 5752 -3329
rect 5786 -3363 5824 -3329
rect 5858 -3363 5896 -3329
rect 5930 -3363 5968 -3329
rect 6002 -3363 6040 -3329
rect 6074 -3363 6112 -3329
rect 6146 -3363 6184 -3329
rect 6218 -3363 6256 -3329
rect 6290 -3363 6328 -3329
rect 6362 -3363 6400 -3329
rect 6434 -3363 6472 -3329
rect 6506 -3363 6544 -3329
rect 6578 -3363 6616 -3329
rect 6650 -3363 6706 -3329
rect 5408 -3382 6706 -3363
rect 6824 -3282 6920 -3272
rect 6824 -3335 8122 -3282
rect 6824 -3369 6880 -3335
rect 6914 -3369 6952 -3335
rect 6986 -3369 7024 -3335
rect 7058 -3369 7096 -3335
rect 7130 -3369 7168 -3335
rect 7202 -3369 7240 -3335
rect 7274 -3369 7312 -3335
rect 7346 -3369 7384 -3335
rect 7418 -3369 7456 -3335
rect 7490 -3369 7528 -3335
rect 7562 -3369 7600 -3335
rect 7634 -3369 7672 -3335
rect 7706 -3369 7744 -3335
rect 7778 -3369 7816 -3335
rect 7850 -3369 7888 -3335
rect 7922 -3369 7960 -3335
rect 7994 -3369 8032 -3335
rect 8066 -3369 8122 -3335
rect 5408 -3448 5510 -3382
rect 5408 -3482 5447 -3448
rect 5481 -3482 5510 -3448
rect 5408 -3520 5510 -3482
rect 5574 -3463 6540 -3446
rect 5574 -3497 5607 -3463
rect 5641 -3497 5679 -3463
rect 5713 -3497 5751 -3463
rect 5785 -3497 5823 -3463
rect 5857 -3497 5895 -3463
rect 5929 -3497 5967 -3463
rect 6001 -3497 6039 -3463
rect 6073 -3497 6111 -3463
rect 6145 -3497 6183 -3463
rect 6217 -3497 6255 -3463
rect 6289 -3497 6327 -3463
rect 6361 -3497 6399 -3463
rect 6433 -3497 6540 -3463
rect 5574 -3506 6540 -3497
rect 5408 -3554 5447 -3520
rect 5481 -3554 5510 -3520
rect 5408 -3592 5510 -3554
rect 5572 -3558 5586 -3506
rect 5638 -3514 6540 -3506
rect 6602 -3448 6704 -3382
rect 6602 -3482 6633 -3448
rect 6667 -3482 6704 -3448
rect 5638 -3558 5650 -3514
rect 5572 -3583 5597 -3558
rect 5631 -3583 5650 -3558
rect 6462 -3549 6536 -3514
rect 5572 -3586 5650 -3583
rect 5408 -3626 5447 -3592
rect 5481 -3626 5510 -3592
rect 5408 -3664 5510 -3626
rect 5408 -3698 5447 -3664
rect 5481 -3698 5510 -3664
rect 5408 -3736 5510 -3698
rect 5408 -3770 5447 -3736
rect 5481 -3770 5510 -3736
rect 5408 -3808 5510 -3770
rect 5408 -3842 5447 -3808
rect 5481 -3842 5510 -3808
rect 5408 -3880 5510 -3842
rect 5408 -3914 5447 -3880
rect 5481 -3914 5510 -3880
rect 5408 -3952 5510 -3914
rect 5408 -3986 5447 -3952
rect 5481 -3986 5510 -3952
rect 5408 -4024 5510 -3986
rect 5408 -4058 5447 -4024
rect 5481 -4058 5510 -4024
rect 5408 -4096 5510 -4058
rect 5408 -4130 5447 -4096
rect 5481 -4130 5510 -4096
rect 5408 -4168 5510 -4130
rect 5408 -4202 5447 -4168
rect 5481 -4202 5510 -4168
rect 5408 -4240 5510 -4202
rect 5408 -4274 5447 -4240
rect 5481 -4274 5510 -4240
rect 5408 -4312 5510 -4274
rect 5408 -4346 5447 -4312
rect 5481 -4346 5510 -4312
rect 5574 -3621 5648 -3586
rect 5574 -3655 5597 -3621
rect 5631 -3655 5648 -3621
rect 5574 -3693 5648 -3655
rect 5574 -3727 5597 -3693
rect 5631 -3727 5648 -3693
rect 5574 -3765 5648 -3727
rect 5574 -3799 5597 -3765
rect 5631 -3799 5648 -3765
rect 5574 -3837 5648 -3799
rect 5574 -3871 5597 -3837
rect 5631 -3871 5648 -3837
rect 5574 -3909 5648 -3871
rect 5574 -3943 5597 -3909
rect 5631 -3943 5648 -3909
rect 5574 -3981 5648 -3943
rect 5574 -4015 5597 -3981
rect 5631 -4015 5648 -3981
rect 5574 -4053 5648 -4015
rect 5574 -4087 5597 -4053
rect 5631 -4087 5648 -4053
rect 5574 -4125 5648 -4087
rect 5574 -4159 5597 -4125
rect 5631 -4159 5648 -4125
rect 5574 -4197 5648 -4159
rect 5574 -4231 5597 -4197
rect 5631 -4231 5648 -4197
rect 5574 -4269 5648 -4231
rect 5714 -3646 6396 -3574
rect 5714 -4210 5776 -3646
rect 6340 -4210 6396 -3646
rect 5714 -4264 6396 -4210
rect 6462 -3583 6487 -3549
rect 6521 -3583 6536 -3549
rect 6462 -3621 6536 -3583
rect 6462 -3655 6487 -3621
rect 6521 -3655 6536 -3621
rect 6462 -3693 6536 -3655
rect 6462 -3727 6487 -3693
rect 6521 -3727 6536 -3693
rect 6462 -3765 6536 -3727
rect 6462 -3799 6487 -3765
rect 6521 -3799 6536 -3765
rect 6462 -3837 6536 -3799
rect 6462 -3871 6487 -3837
rect 6521 -3871 6536 -3837
rect 6462 -3909 6536 -3871
rect 6462 -3943 6487 -3909
rect 6521 -3943 6536 -3909
rect 6462 -3981 6536 -3943
rect 6462 -4015 6487 -3981
rect 6521 -4015 6536 -3981
rect 6462 -4053 6536 -4015
rect 6462 -4087 6487 -4053
rect 6521 -4087 6536 -4053
rect 6462 -4125 6536 -4087
rect 6462 -4159 6487 -4125
rect 6521 -4159 6536 -4125
rect 6462 -4197 6536 -4159
rect 6462 -4231 6487 -4197
rect 6521 -4231 6536 -4197
rect 5574 -4303 5597 -4269
rect 5631 -4303 5648 -4269
rect 5574 -4334 5648 -4303
rect 6462 -4269 6536 -4231
rect 6462 -4303 6487 -4269
rect 6521 -4303 6536 -4269
rect 5408 -4384 5510 -4346
rect 5408 -4418 5447 -4384
rect 5481 -4418 5510 -4384
rect 5568 -4338 5654 -4334
rect 6462 -4338 6536 -4303
rect 6602 -3520 6704 -3482
rect 6602 -3554 6633 -3520
rect 6667 -3554 6704 -3520
rect 6602 -3592 6704 -3554
rect 6602 -3626 6633 -3592
rect 6667 -3626 6704 -3592
rect 6602 -3664 6704 -3626
rect 6602 -3698 6633 -3664
rect 6667 -3698 6704 -3664
rect 6602 -3736 6704 -3698
rect 6602 -3770 6633 -3736
rect 6667 -3770 6704 -3736
rect 6602 -3808 6704 -3770
rect 6602 -3842 6633 -3808
rect 6667 -3842 6704 -3808
rect 6602 -3880 6704 -3842
rect 6602 -3914 6633 -3880
rect 6667 -3914 6704 -3880
rect 6602 -3952 6704 -3914
rect 6602 -3986 6633 -3952
rect 6667 -3986 6704 -3952
rect 6602 -4024 6704 -3986
rect 6602 -4058 6633 -4024
rect 6667 -4058 6704 -4024
rect 6602 -4096 6704 -4058
rect 6602 -4130 6633 -4096
rect 6667 -4130 6704 -4096
rect 6602 -4168 6704 -4130
rect 6602 -4202 6633 -4168
rect 6667 -4202 6704 -4168
rect 6602 -4240 6704 -4202
rect 6602 -4274 6633 -4240
rect 6667 -4274 6704 -4240
rect 6602 -4312 6704 -4274
rect 5568 -4348 6538 -4338
rect 5568 -4400 5585 -4348
rect 5637 -4355 6538 -4348
rect 5637 -4389 5682 -4355
rect 5716 -4389 5754 -4355
rect 5788 -4389 5826 -4355
rect 5860 -4389 5898 -4355
rect 5932 -4389 5970 -4355
rect 6004 -4389 6042 -4355
rect 6076 -4389 6114 -4355
rect 6148 -4389 6186 -4355
rect 6220 -4389 6258 -4355
rect 6292 -4389 6330 -4355
rect 6364 -4389 6402 -4355
rect 6436 -4356 6538 -4355
rect 6436 -4389 6487 -4356
rect 5637 -4390 6487 -4389
rect 6521 -4390 6538 -4356
rect 5637 -4400 6538 -4390
rect 5568 -4406 6538 -4400
rect 6602 -4346 6633 -4312
rect 6667 -4346 6704 -4312
rect 6602 -4384 6704 -4346
rect 5568 -4408 5654 -4406
rect 6462 -4410 6536 -4406
rect 5408 -4466 5510 -4418
rect 6602 -4418 6633 -4384
rect 6667 -4418 6704 -4384
rect 6602 -4466 6704 -4418
rect 6824 -3388 8122 -3369
rect 6824 -3454 6926 -3388
rect 6824 -3488 6863 -3454
rect 6897 -3488 6926 -3454
rect 6824 -3526 6926 -3488
rect 6990 -3469 7956 -3452
rect 6990 -3503 7023 -3469
rect 7057 -3503 7095 -3469
rect 7129 -3503 7167 -3469
rect 7201 -3503 7239 -3469
rect 7273 -3503 7311 -3469
rect 7345 -3503 7383 -3469
rect 7417 -3503 7455 -3469
rect 7489 -3503 7527 -3469
rect 7561 -3503 7599 -3469
rect 7633 -3503 7671 -3469
rect 7705 -3503 7743 -3469
rect 7777 -3503 7815 -3469
rect 7849 -3503 7956 -3469
rect 6990 -3508 7956 -3503
rect 6990 -3512 7011 -3508
rect 6824 -3560 6863 -3526
rect 6897 -3560 6926 -3526
rect 6824 -3598 6926 -3560
rect 6988 -3560 7011 -3512
rect 7063 -3520 7956 -3508
rect 8018 -3454 8120 -3388
rect 8018 -3488 8049 -3454
rect 8083 -3488 8120 -3454
rect 7063 -3560 7066 -3520
rect 6988 -3589 7013 -3560
rect 7047 -3589 7066 -3560
rect 7878 -3555 7952 -3520
rect 6988 -3592 7066 -3589
rect 6824 -3632 6863 -3598
rect 6897 -3632 6926 -3598
rect 6824 -3670 6926 -3632
rect 6824 -3704 6863 -3670
rect 6897 -3704 6926 -3670
rect 6824 -3742 6926 -3704
rect 6824 -3776 6863 -3742
rect 6897 -3776 6926 -3742
rect 6824 -3814 6926 -3776
rect 6824 -3848 6863 -3814
rect 6897 -3848 6926 -3814
rect 6824 -3886 6926 -3848
rect 6824 -3920 6863 -3886
rect 6897 -3920 6926 -3886
rect 6824 -3958 6926 -3920
rect 6824 -3992 6863 -3958
rect 6897 -3992 6926 -3958
rect 6824 -4030 6926 -3992
rect 6824 -4064 6863 -4030
rect 6897 -4064 6926 -4030
rect 6824 -4102 6926 -4064
rect 6824 -4136 6863 -4102
rect 6897 -4136 6926 -4102
rect 6824 -4174 6926 -4136
rect 6824 -4208 6863 -4174
rect 6897 -4208 6926 -4174
rect 6824 -4246 6926 -4208
rect 6824 -4280 6863 -4246
rect 6897 -4280 6926 -4246
rect 6824 -4318 6926 -4280
rect 6824 -4352 6863 -4318
rect 6897 -4352 6926 -4318
rect 6990 -3627 7064 -3592
rect 6990 -3661 7013 -3627
rect 7047 -3661 7064 -3627
rect 6990 -3699 7064 -3661
rect 6990 -3733 7013 -3699
rect 7047 -3733 7064 -3699
rect 6990 -3771 7064 -3733
rect 6990 -3805 7013 -3771
rect 7047 -3805 7064 -3771
rect 6990 -3843 7064 -3805
rect 6990 -3877 7013 -3843
rect 7047 -3877 7064 -3843
rect 6990 -3915 7064 -3877
rect 6990 -3949 7013 -3915
rect 7047 -3949 7064 -3915
rect 6990 -3987 7064 -3949
rect 6990 -4021 7013 -3987
rect 7047 -4021 7064 -3987
rect 6990 -4059 7064 -4021
rect 6990 -4093 7013 -4059
rect 7047 -4093 7064 -4059
rect 6990 -4131 7064 -4093
rect 6990 -4165 7013 -4131
rect 7047 -4165 7064 -4131
rect 6990 -4203 7064 -4165
rect 6990 -4237 7013 -4203
rect 7047 -4237 7064 -4203
rect 6990 -4275 7064 -4237
rect 7130 -3652 7812 -3580
rect 7130 -4216 7192 -3652
rect 7756 -4216 7812 -3652
rect 7130 -4270 7812 -4216
rect 7878 -3589 7903 -3555
rect 7937 -3589 7952 -3555
rect 7878 -3627 7952 -3589
rect 7878 -3661 7903 -3627
rect 7937 -3661 7952 -3627
rect 7878 -3699 7952 -3661
rect 7878 -3733 7903 -3699
rect 7937 -3733 7952 -3699
rect 7878 -3771 7952 -3733
rect 7878 -3805 7903 -3771
rect 7937 -3805 7952 -3771
rect 7878 -3843 7952 -3805
rect 7878 -3877 7903 -3843
rect 7937 -3877 7952 -3843
rect 7878 -3915 7952 -3877
rect 7878 -3949 7903 -3915
rect 7937 -3949 7952 -3915
rect 7878 -3987 7952 -3949
rect 7878 -4021 7903 -3987
rect 7937 -4021 7952 -3987
rect 7878 -4059 7952 -4021
rect 7878 -4093 7903 -4059
rect 7937 -4093 7952 -4059
rect 7878 -4131 7952 -4093
rect 7878 -4165 7903 -4131
rect 7937 -4165 7952 -4131
rect 7878 -4203 7952 -4165
rect 7878 -4237 7903 -4203
rect 7937 -4237 7952 -4203
rect 6990 -4309 7013 -4275
rect 7047 -4309 7064 -4275
rect 6990 -4340 7064 -4309
rect 7878 -4275 7952 -4237
rect 7878 -4309 7903 -4275
rect 7937 -4309 7952 -4275
rect 6824 -4390 6926 -4352
rect 6824 -4424 6863 -4390
rect 6897 -4424 6926 -4390
rect 6984 -4344 7070 -4340
rect 7878 -4344 7952 -4309
rect 8018 -3526 8120 -3488
rect 8018 -3560 8049 -3526
rect 8083 -3560 8120 -3526
rect 8018 -3598 8120 -3560
rect 8018 -3632 8049 -3598
rect 8083 -3632 8120 -3598
rect 8018 -3670 8120 -3632
rect 8018 -3704 8049 -3670
rect 8083 -3704 8120 -3670
rect 8018 -3742 8120 -3704
rect 8018 -3776 8049 -3742
rect 8083 -3776 8120 -3742
rect 8018 -3814 8120 -3776
rect 8018 -3848 8049 -3814
rect 8083 -3848 8120 -3814
rect 8018 -3886 8120 -3848
rect 8018 -3920 8049 -3886
rect 8083 -3920 8120 -3886
rect 8018 -3958 8120 -3920
rect 8018 -3992 8049 -3958
rect 8083 -3992 8120 -3958
rect 8018 -4030 8120 -3992
rect 8018 -4064 8049 -4030
rect 8083 -4064 8120 -4030
rect 8018 -4102 8120 -4064
rect 8018 -4136 8049 -4102
rect 8083 -4136 8120 -4102
rect 8018 -4174 8120 -4136
rect 8018 -4208 8049 -4174
rect 8083 -4208 8120 -4174
rect 8018 -4246 8120 -4208
rect 8018 -4280 8049 -4246
rect 8083 -4280 8120 -4246
rect 8018 -4318 8120 -4280
rect 6984 -4354 7954 -4344
rect 6984 -4406 7001 -4354
rect 7053 -4361 7954 -4354
rect 7053 -4395 7098 -4361
rect 7132 -4395 7170 -4361
rect 7204 -4395 7242 -4361
rect 7276 -4395 7314 -4361
rect 7348 -4395 7386 -4361
rect 7420 -4395 7458 -4361
rect 7492 -4395 7530 -4361
rect 7564 -4395 7602 -4361
rect 7636 -4395 7674 -4361
rect 7708 -4395 7746 -4361
rect 7780 -4395 7818 -4361
rect 7852 -4362 7954 -4361
rect 7852 -4395 7903 -4362
rect 7053 -4396 7903 -4395
rect 7937 -4396 7954 -4362
rect 7053 -4406 7954 -4396
rect 6984 -4412 7954 -4406
rect 8018 -4352 8049 -4318
rect 8083 -4352 8120 -4318
rect 8018 -4390 8120 -4352
rect 6984 -4414 7070 -4412
rect 7878 -4416 7952 -4412
rect 5408 -4503 6706 -4466
rect 5408 -4537 5464 -4503
rect 5498 -4537 5536 -4503
rect 5570 -4537 5608 -4503
rect 5642 -4537 5680 -4503
rect 5714 -4537 5752 -4503
rect 5786 -4537 5824 -4503
rect 5858 -4537 5896 -4503
rect 5930 -4537 5968 -4503
rect 6002 -4537 6040 -4503
rect 6074 -4537 6112 -4503
rect 6146 -4537 6184 -4503
rect 6218 -4537 6256 -4503
rect 6290 -4537 6328 -4503
rect 6362 -4537 6400 -4503
rect 6434 -4537 6472 -4503
rect 6506 -4537 6544 -4503
rect 6578 -4537 6616 -4503
rect 6650 -4537 6706 -4503
rect 5408 -4546 6706 -4537
rect 5406 -4562 6706 -4546
rect 6824 -4472 6926 -4424
rect 8018 -4424 8049 -4390
rect 8083 -4424 8120 -4390
rect 8018 -4472 8120 -4424
rect 8702 -3962 8944 -3894
rect 6824 -4509 8122 -4472
rect 6824 -4543 6880 -4509
rect 6914 -4543 6952 -4509
rect 6986 -4543 7024 -4509
rect 7058 -4543 7096 -4509
rect 7130 -4543 7168 -4509
rect 7202 -4543 7240 -4509
rect 7274 -4543 7312 -4509
rect 7346 -4543 7384 -4509
rect 7418 -4543 7456 -4509
rect 7490 -4543 7528 -4509
rect 7562 -4543 7600 -4509
rect 7634 -4543 7672 -4509
rect 7706 -4543 7744 -4509
rect 7778 -4543 7816 -4509
rect 7850 -4543 7888 -4509
rect 7922 -4543 7960 -4509
rect 7994 -4543 8032 -4509
rect 8066 -4543 8122 -4509
rect 6824 -4552 8122 -4543
rect 5404 -4572 6706 -4562
rect 6822 -4572 8122 -4552
rect 2296 -5148 2374 -5133
rect 5404 -5160 5496 -4572
rect 6818 -4578 8122 -4572
rect 6818 -4586 6912 -4578
rect 6818 -5068 6910 -4586
rect 8702 -4950 8756 -3962
rect 6980 -5046 7064 -5026
rect 5560 -5082 5648 -5080
rect 5560 -5134 5579 -5082
rect 5631 -5134 5648 -5082
rect 6980 -5098 6994 -5046
rect 7046 -5098 7064 -5046
rect 6980 -5108 7064 -5098
rect 8702 -5134 8758 -4950
rect 9566 -4996 9628 -3188
rect 9986 -4950 10040 -3118
rect 10862 -3556 10916 34
rect 13390 -1124 13448 -1120
rect 12428 -2010 12486 -1162
rect 13382 -1956 13448 -1124
rect 14172 -1580 14238 -1174
rect 14048 -1660 14238 -1580
rect 14048 -1668 14110 -1660
rect 13382 -1984 13450 -1956
rect 11610 -2454 12216 -2390
rect 10860 -3620 11304 -3556
rect 9984 -4996 10042 -4950
rect 5560 -5146 5648 -5134
rect 9570 -5182 9626 -4996
rect 9986 -5180 10042 -4996
rect 11246 -5122 11304 -3620
rect 11610 -3756 11676 -2454
rect 12430 -3552 12482 -2010
rect 13384 -2424 13450 -1984
rect 13158 -2494 13452 -2424
rect 11396 -3802 11676 -3756
rect 12214 -3594 12482 -3552
rect 13132 -3560 13186 -2606
rect 13922 -3560 13970 -2278
rect 12916 -3594 13186 -3560
rect 13706 -3594 13970 -3560
rect 14050 -3586 14110 -1668
rect 14048 -3594 14110 -3586
rect 11396 -4950 11460 -3802
rect 11394 -5132 11460 -4950
rect 12214 -4950 12262 -3594
rect 12916 -4950 12968 -3594
rect 12214 -5126 12266 -4950
rect 12916 -5170 12970 -4950
rect 13706 -5170 13754 -3594
rect 14048 -3730 14108 -3594
rect 13834 -3778 14108 -3730
rect 13834 -5108 13894 -3778
<< via1 >>
rect 704 998 756 1050
rect 1162 996 1214 1048
rect 1152 863 1204 915
rect 2926 1117 2978 1169
rect 3239 1128 3291 1180
rect 3594 1019 3646 1071
rect 4169 1012 4221 1064
rect 2254 890 2306 942
rect 7407 3103 7459 3155
rect 8454 3090 8506 3142
rect 9316 3102 9368 3154
rect 10172 3116 10224 3168
rect 5620 3000 5672 3052
rect 3244 779 3296 831
rect 3595 776 3647 828
rect 1626 660 1678 712
rect 3310 490 3362 542
rect 1624 119 1676 171
rect 2224 -391 2788 173
rect 2031 -543 2083 -538
rect 2031 -577 2042 -543
rect 2042 -577 2076 -543
rect 2076 -577 2083 -543
rect 2031 -590 2083 -577
rect 4178 460 4230 512
rect 2309 -5092 2361 -5081
rect 2309 -5126 2316 -5092
rect 2316 -5126 2350 -5092
rect 2350 -5126 2361 -5092
rect 2309 -5133 2361 -5126
rect 7188 1222 7752 1786
rect 8920 1570 8972 1622
rect 12184 1250 12236 1302
rect 6997 1077 7049 1084
rect 6997 1043 7009 1077
rect 7009 1043 7043 1077
rect 7043 1043 7049 1077
rect 6997 1032 7049 1043
rect 13136 826 13188 878
rect 7004 527 7056 578
rect 13919 671 13971 723
rect 7004 526 7013 527
rect 7013 526 7047 527
rect 7047 526 7056 527
rect 7192 -134 7756 430
rect 7001 -279 7053 -272
rect 7001 -313 7013 -279
rect 7013 -313 7047 -279
rect 7047 -313 7053 -279
rect 7001 -324 7053 -313
rect 5778 -1502 6342 -938
rect 5587 -1647 5639 -1640
rect 5587 -1681 5599 -1647
rect 5599 -1681 5633 -1647
rect 5633 -1681 5639 -1647
rect 5587 -1692 5639 -1681
rect 7002 -837 7054 -786
rect 7002 -838 7009 -837
rect 7009 -838 7043 -837
rect 7043 -838 7054 -837
rect 7188 -1498 7752 -934
rect 6997 -1643 7049 -1636
rect 6997 -1677 7009 -1643
rect 7009 -1677 7043 -1643
rect 7043 -1677 7049 -1643
rect 6997 -1688 7049 -1677
rect 5590 -2197 5642 -2150
rect 5590 -2202 5597 -2197
rect 5597 -2202 5631 -2197
rect 5631 -2202 5642 -2197
rect 5776 -2858 6340 -2294
rect 5585 -3003 5637 -2996
rect 5585 -3037 5597 -3003
rect 5597 -3037 5631 -3003
rect 5631 -3037 5637 -3003
rect 5585 -3048 5637 -3037
rect 7000 -2195 7052 -2154
rect 7000 -2206 7011 -2195
rect 7011 -2206 7045 -2195
rect 7045 -2206 7052 -2195
rect 7190 -2856 7754 -2292
rect 6999 -3001 7051 -2994
rect 6999 -3035 7011 -3001
rect 7011 -3035 7045 -3001
rect 7045 -3035 7051 -3001
rect 6999 -3046 7051 -3035
rect 5586 -3549 5638 -3506
rect 5586 -3558 5597 -3549
rect 5597 -3558 5631 -3549
rect 5631 -3558 5638 -3549
rect 5776 -4210 6340 -3646
rect 5585 -4355 5637 -4348
rect 5585 -4389 5597 -4355
rect 5597 -4389 5631 -4355
rect 5631 -4389 5637 -4355
rect 5585 -4400 5637 -4389
rect 7011 -3555 7063 -3508
rect 7011 -3560 7013 -3555
rect 7013 -3560 7047 -3555
rect 7047 -3560 7063 -3555
rect 7192 -4216 7756 -3652
rect 7001 -4361 7053 -4354
rect 7001 -4395 7013 -4361
rect 7013 -4395 7047 -4361
rect 7047 -4395 7053 -4361
rect 7001 -4406 7053 -4395
rect 5579 -5093 5631 -5082
rect 5579 -5127 5585 -5093
rect 5585 -5127 5619 -5093
rect 5619 -5127 5631 -5093
rect 5579 -5134 5631 -5127
rect 6994 -5057 7046 -5046
rect 6994 -5091 7002 -5057
rect 7002 -5091 7036 -5057
rect 7036 -5091 7046 -5057
rect 6994 -5098 7046 -5091
<< metal2 >>
rect -1168 4712 -522 4798
rect -580 2966 -522 4712
rect 10164 3174 10388 3176
rect 10164 3168 10390 3174
rect 7400 3162 7462 3168
rect 7398 3160 7462 3162
rect 7398 3155 7932 3160
rect 7398 3103 7407 3155
rect 7459 3103 7932 3155
rect 9308 3154 9496 3162
rect 7398 3096 7932 3103
rect 7398 3094 7462 3096
rect 5610 3052 5680 3060
rect 5610 3000 5620 3052
rect 5672 3000 5680 3052
rect -580 722 -510 2966
rect 5610 2920 5680 3000
rect 4382 2880 5680 2920
rect 2924 1180 2966 1182
rect 3220 1180 3310 1190
rect 2924 1169 3120 1180
rect 2924 1117 2926 1169
rect 2978 1117 3120 1169
rect 2924 1102 3120 1117
rect 2924 1100 2966 1102
rect 1142 1054 1222 1056
rect 686 1050 1222 1054
rect 686 998 704 1050
rect 756 1048 1222 1050
rect 756 998 1162 1048
rect 686 996 1162 998
rect 1214 996 1222 1048
rect 686 992 1222 996
rect 3050 950 3120 1102
rect 1136 948 3120 950
rect 3220 1128 3239 1180
rect 3291 1128 3310 1180
rect 1136 942 3122 948
rect 1136 915 2254 942
rect 1136 863 1152 915
rect 1204 890 2254 915
rect 2306 890 3122 942
rect 1204 863 3122 890
rect 1136 846 3122 863
rect 3220 926 3310 1128
rect 3560 1071 3680 1082
rect 3560 1019 3594 1071
rect 3646 1019 3680 1071
rect 1136 844 3120 846
rect 1714 842 3120 844
rect -580 712 1684 722
rect -580 660 1626 712
rect 1678 660 1684 712
rect -580 650 1684 660
rect 3050 570 3120 842
rect 3220 831 3312 926
rect 3220 779 3244 831
rect 3296 779 3312 831
rect 3220 766 3312 779
rect 3560 828 3680 1019
rect 4150 1064 4240 1070
rect 4150 1012 4169 1064
rect 4221 1012 4240 1064
rect 4150 970 4240 1012
rect 4382 970 4420 2880
rect 7892 2422 7932 3096
rect 8446 3142 8636 3150
rect 8446 3090 8454 3142
rect 8506 3090 8636 3142
rect 9308 3102 9316 3154
rect 9368 3102 9496 3154
rect 10164 3116 10172 3168
rect 10224 3116 10390 3168
rect 10164 3106 10390 3116
rect 9308 3092 9496 3102
rect 8446 3080 8636 3090
rect 8596 2770 8636 3080
rect 9456 2902 9496 3092
rect 9456 2900 9642 2902
rect 9456 2860 10160 2900
rect 8596 2730 10020 2770
rect 8290 2424 8330 2426
rect 8290 2422 8650 2424
rect 7892 2382 8650 2422
rect 7120 1786 7806 2286
rect 8574 2156 8650 2382
rect 9980 2288 10020 2730
rect 8574 2054 9012 2156
rect 8570 2052 9012 2054
rect 8570 2025 8690 2052
rect 8570 1969 8598 2025
rect 8654 1969 8690 2025
rect 8570 1934 8690 1969
rect 7120 1222 7188 1786
rect 7752 1222 7806 1786
rect 8890 1622 9012 2052
rect 8890 1570 8920 1622
rect 8972 1570 9012 1622
rect 8890 1542 9012 1570
rect 4150 930 4420 970
rect 3560 776 3595 828
rect 3647 800 3680 828
rect 3647 776 4260 800
rect 3560 740 4260 776
rect 3926 738 4260 740
rect 3052 554 3120 570
rect 3052 550 3192 554
rect 3052 542 3368 550
rect 3052 490 3310 542
rect 3362 490 3368 542
rect 3052 480 3368 490
rect 4150 512 4260 738
rect 3052 476 3192 480
rect 4150 460 4178 512
rect 4230 460 4260 512
rect 4150 450 4260 460
rect 7120 430 7806 1222
rect 9980 1262 10018 2288
rect 10120 1452 10160 2860
rect 10346 1570 10390 3106
rect 10346 1530 13610 1570
rect 10346 1528 10390 1530
rect 12328 1452 12872 1454
rect 10120 1408 12872 1452
rect 10120 1406 10160 1408
rect 12158 1307 12278 1334
rect 12158 1302 12186 1307
rect 12158 1262 12184 1302
rect 9980 1250 12184 1262
rect 12242 1251 12278 1307
rect 12236 1250 12278 1251
rect 9980 1220 12278 1250
rect 12158 1216 12278 1220
rect 12778 1210 12872 1408
rect 12778 922 12870 1210
rect 12778 900 13198 922
rect 12778 879 13220 900
rect 12778 832 13134 879
rect 13102 823 13134 832
rect 13190 823 13220 879
rect 13102 810 13220 823
rect 13106 788 13220 810
rect 13500 752 13610 1530
rect 13890 752 14000 754
rect 13500 731 14002 752
rect 13500 675 13916 731
rect 13972 675 14002 731
rect 13500 671 13919 675
rect 13971 671 14002 675
rect 13500 644 14002 671
rect 13888 642 14002 644
rect 1616 173 2844 231
rect 1616 171 2224 173
rect 1616 119 1624 171
rect 1676 119 2224 171
rect 1616 -391 2224 119
rect 2788 -391 2844 173
rect 7120 -134 7192 430
rect 7756 -134 7806 430
rect 1616 -409 2844 -391
rect 2154 -462 2844 -409
rect 2016 -538 2104 -526
rect 2016 -590 2031 -538
rect 2083 -590 2104 -538
rect 2016 -884 2104 -590
rect 2014 -886 2104 -884
rect 2014 -1004 2098 -886
rect 5710 -938 6396 -862
rect 2014 -1114 2096 -1004
rect 2014 -1174 2362 -1114
rect 2298 -4950 2362 -1174
rect 5710 -1502 5778 -938
rect 6342 -1502 6396 -938
rect 5710 -1556 6396 -1502
rect 7120 -934 7806 -134
rect 7120 -1498 7188 -934
rect 7752 -1498 7806 -934
rect 5570 -1640 5654 -1628
rect 5570 -1692 5587 -1640
rect 5639 -1692 5654 -1640
rect 5570 -1844 5654 -1692
rect 5568 -1872 5654 -1844
rect 5572 -2150 5652 -1872
rect 5572 -2202 5590 -2150
rect 5642 -2202 5652 -2150
rect 5572 -2212 5652 -2202
rect 5710 -2219 6395 -1556
rect 5710 -2294 6394 -2219
rect 5710 -2858 5776 -2294
rect 6340 -2858 6394 -2294
rect 5570 -2996 5652 -2984
rect 5570 -3048 5585 -2996
rect 5637 -3048 5652 -2996
rect 5570 -3506 5652 -3048
rect 5570 -3558 5586 -3506
rect 5638 -3558 5652 -3506
rect 5570 -3582 5652 -3558
rect 5710 -3568 6394 -2858
rect 7120 -2292 7806 -1498
rect 7120 -2856 7190 -2292
rect 7754 -2856 7806 -2292
rect 5708 -3646 6394 -3568
rect 5708 -4210 5776 -3646
rect 6340 -3648 6394 -3646
rect 7120 -3648 7806 -2856
rect 6340 -3652 7810 -3648
rect 6340 -4210 7192 -3652
rect 5708 -4216 7192 -4210
rect 7756 -4216 7810 -3652
rect 5708 -4230 7810 -4216
rect 5712 -4270 7810 -4230
rect 5568 -4348 5652 -4336
rect 5568 -4400 5585 -4348
rect 5637 -4400 5652 -4348
rect 5568 -4552 5652 -4400
rect 6984 -4354 7068 -4342
rect 6984 -4406 7001 -4354
rect 7053 -4406 7068 -4354
rect 6984 -4552 7068 -4406
rect 5566 -4562 5652 -4552
rect 5564 -4580 5652 -4562
rect 2296 -5081 2376 -4950
rect 2296 -5133 2309 -5081
rect 2361 -5133 2376 -5081
rect 2296 -5150 2376 -5133
rect 5564 -5082 5648 -4580
rect 5564 -5134 5579 -5082
rect 5631 -5134 5648 -5082
rect 6978 -4586 7068 -4552
rect 6978 -5046 7066 -4586
rect 6978 -5098 6994 -5046
rect 7046 -5098 7066 -5046
rect 6978 -5108 7066 -5098
rect 5564 -5146 5648 -5134
<< via2 >>
rect 8598 1969 8654 2025
rect 12186 1302 12242 1307
rect 12186 1251 12236 1302
rect 12236 1251 12242 1302
rect 13134 878 13190 879
rect 13134 826 13136 878
rect 13136 826 13188 878
rect 13188 826 13190 878
rect 13134 823 13190 826
rect 13916 723 13972 731
rect 13916 675 13919 723
rect 13919 675 13971 723
rect 13971 675 13972 723
<< metal3 >>
rect 8572 2030 8684 2046
rect 8572 1966 8594 2030
rect 8658 1966 8684 2030
rect 8572 1944 8684 1966
rect 12160 1312 12272 1328
rect 12160 1248 12182 1312
rect 12246 1248 12272 1312
rect 12160 1226 12272 1248
rect 13108 884 13220 900
rect 13108 820 13130 884
rect 13194 820 13220 884
rect 13108 798 13220 820
rect 13890 736 14002 752
rect 13890 672 13912 736
rect 13976 672 14002 736
rect 13890 650 14002 672
<< via3 >>
rect 8594 2025 8658 2030
rect 8594 1969 8598 2025
rect 8598 1969 8654 2025
rect 8654 1969 8658 2025
rect 8594 1966 8658 1969
rect 12182 1307 12246 1312
rect 12182 1251 12186 1307
rect 12186 1251 12242 1307
rect 12242 1251 12246 1307
rect 12182 1248 12246 1251
rect 13130 879 13194 884
rect 13130 823 13134 879
rect 13134 823 13190 879
rect 13190 823 13194 879
rect 13130 820 13194 823
rect 13912 731 13976 736
rect 13912 675 13916 731
rect 13916 675 13972 731
rect 13972 675 13976 731
rect 13912 672 13976 675
<< metal4 >>
rect 8572 2030 8684 2046
rect 8572 1966 8594 2030
rect 8658 1966 8684 2030
rect 8572 1948 8684 1966
rect 8570 1858 8684 1948
rect 13978 1858 14200 2120
rect 8570 1798 14200 1858
rect 14280 1328 14530 1612
rect 12158 1312 14530 1328
rect 12158 1248 12182 1312
rect 12246 1248 14530 1312
rect 12158 1216 14530 1248
rect 14970 920 15220 1244
rect 13106 884 15220 920
rect 13106 820 13130 884
rect 13194 860 15220 884
rect 13194 858 13810 860
rect 13194 820 13220 858
rect 13106 788 13220 820
rect 13888 736 14002 752
rect 13888 672 13912 736
rect 13976 702 14002 736
rect 15462 702 15700 956
rect 13976 672 15700 702
rect 13888 642 15700 672
use 298k  R1
timestamp 1669522153
transform 1 0 6899 0 1 335
box 0 0 1 1
use 52k  R2
timestamp 1669522153
transform 1 0 6895 0 1 335
box 0 0 1 1
use 485k  R3
timestamp 1669522153
transform 1 0 6896 0 1 335
box 0 0 1 1
use 520k  R4
timestamp 1669522153
transform 1 0 6897 0 1 335
box 0 0 1 1
use 520k  R5
timestamp 1669522153
transform 1 0 6898 0 1 335
box 0 0 1 1
use 295k  R6
timestamp 1669522153
transform 1 0 8517 0 1 176
box 0 0 1 1
use 298k  R7
timestamp 1669522153
transform 1 0 8518 0 1 176
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_E8XWE6  XM7
timestamp 1669522153
transform 1 0 4066 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__nfet_01v8_B2EJVN  XM8
timestamp 1669522153
transform 1 0 3468 0 1 -1129
box -1084 -157 1084 157
use sky130_fd_pr__nfet_01v8_2HQT3D  XM10
timestamp 1669522153
transform 1 0 5106 0 1 361
box -1084 -157 1084 157
use sky130_fd_pr__pfet_01v8_KVG9ZD  XM11
timestamp 1669522153
transform 1 0 7194 0 1 5504
box -294 -2514 294 2548
use sky130_fd_pr__pfet_01v8_E8XWA6  XM12
timestamp 1669522153
transform 1 0 2260 0 1 3068
box -294 -2064 294 2098
use res2_529K  res2_529K_0
timestamp 1669522153
transform 1 0 10116 0 1 -3116
box -284 0 72 1254
use res2_529K  res2_529K_1
timestamp 1669522153
transform 1 0 -1162 0 1 -3420
box -284 0 72 1254
use res52_504  res52_504_0
timestamp 1669522153
transform -1 0 6382 0 -1 3244
box -228 662 50 2126
use res69_646K  res69_646K_0
timestamp 1669522153
transform -1 0 13978 0 -1 774
box -340 0 72 3264
use res81_075K  res81_075K_0
timestamp 1669522153
transform -1 0 13192 0 -1 922
box -322 0 72 3664
use res92_504K  res92_504K_0
timestamp 1669522153
transform -1 0 12256 0 -1 1346
box -374 0 72 4064
use res141_475K  res141_475K_0
timestamp 1669522153
transform -1 0 8980 0 -1 1626
box -424 0 72 5778
use res172_504K  res172_504K_0
timestamp 1669522153
transform 1 0 -1162 0 1 -1918
box -754 0 72 6864
use res172_504K  res172_504K_1
timestamp 1669522153
transform -1 0 10550 0 -1 4342
box -754 0 72 6864
use sky130_fd_pr__nfet_01v8_7ZFCMD  sky130_fd_pr__nfet_01v8_7ZFCMD_0
timestamp 1669522153
transform 1 0 176 0 1 -588
box -1084 -188 1084 188
use sky130_fd_pr__nfet_01v8_7ZFCMD  sky130_fd_pr__nfet_01v8_7ZFCMD_1
timestamp 1669522153
transform 0 -1 4786 1 0 2020
box -1084 -188 1084 188
use sky130_fd_pr__pfet_01v8_A42UEE  sky130_fd_pr__pfet_01v8_A42UEE_0
timestamp 1669522153
transform 1 0 580 0 1 3056
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8AXA6  sky130_fd_pr__pfet_01v8_E8AXA6_0
timestamp 1669522153
transform 1 0 8248 0 1 5542
box -294 -2564 294 2598
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_0
timestamp 1669522153
transform 1 0 5702 0 1 5044
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_1
timestamp 1669522153
transform 1 0 3608 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_2
timestamp 1669522153
transform 1 0 2718 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_EZH9H8  sky130_fd_pr__pfet_01v8_EZH9H8_0
timestamp 1669522153
transform 1 0 1416 0 1 2068
box -294 -2100 294 2100
use sky130_fd_pr__pfet_01v8_WN8SF2  sky130_fd_pr__pfet_01v8_WN8SF2_0
timestamp 1669522153
transform 1 0 9960 0 1 5554
box -294 -2564 294 2598
use sky130_fd_pr__pfet_01v8_WN8SF2  sky130_fd_pr__pfet_01v8_WN8SF2_1
timestamp 1669522153
transform 1 0 9112 0 1 5550
box -294 -2564 294 2598
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0
timestamp 1669522153
transform 1 0 6808 0 1 848
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1669522153
transform 1 0 6806 0 1 -518
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1669522153
transform 1 0 1834 0 1 -786
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1669522153
transform 1 0 6804 0 1 -1882
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1669522153
transform 1 0 5394 0 1 -1886
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1669522153
transform 1 0 6804 0 1 -3240
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1669522153
transform 1 0 5394 0 1 -3240
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1669522153
transform 1 0 5394 0 1 -4590
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1669522153
transform 1 0 6808 0 1 -4596
box 0 0 1340 1340
<< labels >>
rlabel locali s 3256 -5140 3574 -5020 4 GND
port 1 nsew
rlabel locali s 4384 8406 4706 8560 4 Vdd
port 2 nsew
rlabel metal4 s 15036 912 15128 1078 4 Vref2
port 3 nsew
rlabel metal4 s 14326 1352 14490 1562 4 Vref1
port 4 nsew
rlabel metal4 s 15500 672 15620 828 4 Vref3
port 5 nsew
rlabel metal4 s 14018 1848 14140 2008 4 Vout
port 6 nsew
rlabel metal1 s 2388 702 2476 726 4 G9
port 7 nsew
rlabel metal1 s 3792 894 3914 942 4 G11
port 8 nsew
rlabel metal1 s 898 -244 932 -204 4 G1
port 9 nsew
rlabel metal1 s 10206 -2250 10280 -2218 4 R2
port 10 nsew
rlabel metal1 s 4334 616 4406 648 4 SM9
port 11 nsew
rlabel metal1 s -1158 -2110 -1098 -2006 4 R7
port 12 nsew
rlabel metal1 s 4570 3258 4762 3312 4 SM7
port 13 nsew
rlabel metal2 s 7164 2310 7164 2310 4 Q2
port 14 nsew
rlabel metal2 s 4174 678 4244 750 4 G10
port 15 nsew
<< end >>
