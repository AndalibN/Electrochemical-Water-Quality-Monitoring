magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect 19 122 77 128
rect 19 88 31 122
rect 19 82 77 88
<< pwell >>
rect -151 -76 151 76
<< nmos >>
rect -63 -50 -33 50
rect 33 -50 63 50
<< ndiff >>
rect -125 17 -63 50
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -50 -63 -17
rect -33 17 33 50
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -50 33 -17
rect 63 17 125 50
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -50 125 -17
<< ndiffc >>
rect -113 -17 -79 17
rect -17 -17 17 17
rect 79 -17 113 17
<< poly >>
rect -63 122 81 138
rect -63 88 31 122
rect 65 88 81 122
rect -63 72 81 88
rect -63 50 -33 72
rect 33 50 63 72
rect -63 -76 -33 -50
rect 33 -76 63 -50
<< polycont >>
rect 31 88 65 122
<< locali >>
rect 15 88 31 122
rect 65 88 81 122
rect -113 17 -79 54
rect -113 -54 -79 -17
rect -17 17 17 54
rect -17 -54 17 -17
rect 79 17 113 54
rect 79 -54 113 -17
<< viali >>
rect 31 88 65 122
rect -113 -17 -79 17
rect -17 -17 17 17
rect 79 -17 113 17
<< metal1 >>
rect 19 122 77 128
rect 19 88 31 122
rect 65 88 77 122
rect 19 82 77 88
rect -119 17 -73 50
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -50 -73 -17
rect -23 17 23 50
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -50 23 -17
rect 73 17 119 50
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -50 119 -17
<< end >>
