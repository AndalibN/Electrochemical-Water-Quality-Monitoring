magic
tech sky130A
magscale 1 2
timestamp 1662683859
<< error_p >>
rect 19 122 77 128
rect 19 88 31 122
rect 19 82 77 88
<< nmos >>
rect -63 -50 -33 50
rect 33 -50 63 50
<< ndiff >>
rect -125 38 -63 50
rect -125 -38 -113 38
rect -79 -38 -63 38
rect -125 -50 -63 -38
rect -33 38 33 50
rect -33 -38 -17 38
rect 17 -38 33 38
rect -33 -50 33 -38
rect 63 38 125 50
rect 63 -38 79 38
rect 113 -38 125 38
rect 63 -50 125 -38
<< ndiffc >>
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
<< poly >>
rect 15 122 81 138
rect -63 88 31 122
rect 65 88 81 122
rect -63 50 -33 88
rect 15 72 81 88
rect 33 50 63 72
rect -63 -76 -33 -50
rect 33 -76 63 -50
<< polycont >>
rect 31 88 65 122
<< locali >>
rect 15 88 31 122
rect 65 88 81 122
rect -113 38 -79 54
rect -113 -54 -79 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 79 38 113 54
rect 79 -54 113 -38
<< viali >>
rect 31 88 65 122
rect -113 -38 -79 38
rect -17 -38 17 38
rect 79 -38 113 38
<< metal1 >>
rect 19 122 77 128
rect 19 88 31 122
rect 65 88 77 122
rect 19 82 77 88
rect -119 38 -73 50
rect -119 -38 -113 38
rect -79 -38 -73 38
rect -119 -50 -73 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 73 38 119 50
rect 73 -38 79 38
rect 113 -38 119 38
rect 73 -50 119 -38
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
