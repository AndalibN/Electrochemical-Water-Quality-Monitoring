magic
tech sky130A
magscale 1 2
timestamp 1668796479
<< metal1 >>
rect -28540 -38846 28540 -34879
rect -28540 -39300 -7600 -38846
rect -28540 -51342 -28488 -39300
rect -28494 -51384 -28488 -51342
rect -12628 -40616 -7600 -39300
rect 7600 -39238 28540 -38846
rect 7600 -40616 12628 -39238
rect -12628 -40706 12628 -40616
rect -12628 -41236 -7600 -40706
rect 7600 -41236 12628 -40706
rect -12628 -41326 12628 -41236
rect -12628 -41856 -7600 -41326
rect 7600 -41856 12628 -41326
rect -12628 -41946 12628 -41856
rect -12628 -42476 -7600 -41946
rect 7600 -42476 12628 -41946
rect -12628 -42566 12628 -42476
rect -12628 -43096 -7600 -42566
rect 7600 -43096 12628 -42566
rect -12628 -43186 12628 -43096
rect -12628 -43716 -7600 -43186
rect 7600 -43716 12628 -43186
rect -12628 -43806 12628 -43716
rect -12628 -44336 -7600 -43806
rect 7600 -44336 12628 -43806
rect -12628 -44426 12628 -44336
rect -12628 -44956 -7600 -44426
rect 7600 -44956 12628 -44426
rect -12628 -45046 12628 -44956
rect -12628 -45576 -7600 -45046
rect 7600 -45576 12628 -45046
rect -12628 -45666 12628 -45576
rect -12628 -46196 -7600 -45666
rect 7600 -46196 12628 -45666
rect -12628 -46286 12628 -46196
rect -12628 -46816 -7600 -46286
rect 7600 -46816 12628 -46286
rect -12628 -46906 12628 -46816
rect -12628 -47436 -7600 -46906
rect 7600 -47436 12628 -46906
rect -12628 -47526 12628 -47436
rect -12628 -48056 -7600 -47526
rect 7600 -48056 12628 -47526
rect -12628 -48146 12628 -48056
rect -12628 -48676 -7600 -48146
rect 7600 -48676 12628 -48146
rect -12628 -48766 12628 -48676
rect -12628 -49296 -7600 -48766
rect 7600 -49296 12628 -48766
rect -12628 -49386 12628 -49296
rect -12628 -49916 -7600 -49386
rect 7600 -49916 12628 -49386
rect -12628 -50006 12628 -49916
rect -12628 -50536 -7600 -50006
rect 7600 -50536 12628 -50006
rect -12628 -50626 12628 -50536
rect -12628 -51156 -7600 -50626
rect 7600 -51156 12628 -50626
rect -12628 -51246 12628 -51156
rect -12628 -51342 -7600 -51246
rect 7600 -51322 12628 -51246
rect 28488 -51322 28540 -39238
rect 7600 -51342 28540 -51322
rect -12628 -51384 -12622 -51342
rect -28494 -51390 -12622 -51384
<< via1 >>
rect -28488 -51384 -12628 -39300
rect 12628 -51322 28488 -39238
<< metal2 >>
rect 12622 -39238 28494 -39232
rect 12622 -39243 12628 -39238
rect 12601 -39252 12628 -39243
rect 28488 -39243 28494 -39238
rect 28488 -39252 28515 -39243
rect -28494 -39300 -12622 -39294
rect -28494 -39305 -28488 -39300
rect -28515 -39314 -28488 -39305
rect -12628 -39305 -12622 -39300
rect -12628 -39314 -12601 -39305
rect -28515 -51370 -28506 -39314
rect -12610 -51370 -12601 -39314
rect 12601 -51308 12610 -39252
rect 28506 -51308 28515 -39252
rect 12601 -51317 12628 -51308
rect 12622 -51322 12628 -51317
rect 28488 -51317 28515 -51308
rect 28488 -51322 28494 -51317
rect 12622 -51328 28494 -51322
rect -28515 -51379 -28488 -51370
rect -28494 -51384 -28488 -51379
rect -12628 -51379 -12601 -51370
rect -12628 -51384 -12622 -51379
rect -28494 -51390 -12622 -51384
<< via2 >>
rect -28506 -51370 -28488 -39314
rect -28488 -51370 -12628 -39314
rect -12628 -51370 -12610 -39314
rect 12610 -51308 12628 -39252
rect 12628 -51308 28488 -39252
rect 28488 -51308 28506 -39252
<< metal3 >>
rect 12600 -39248 28516 -39242
rect -28516 -39310 -12600 -39304
rect -28516 -51374 -28510 -39310
rect -12606 -51374 -12600 -39310
rect 12600 -51312 12606 -39248
rect 28510 -51312 28516 -39248
rect 12600 -51318 28516 -51312
rect -28516 -51380 -12600 -51374
<< via3 >>
rect -28510 -39314 -12606 -39310
rect -28510 -51370 -28506 -39314
rect -28506 -51370 -12610 -39314
rect -12610 -51370 -12606 -39314
rect -28510 -51374 -12606 -51370
rect 12606 -39252 28510 -39248
rect 12606 -51308 12610 -39252
rect 12610 -51308 28506 -39252
rect 28506 -51308 28510 -39252
rect 12606 -51312 28510 -51308
<< via4 >>
rect 12600 -39248 28516 -39242
rect -28516 -39310 -12600 -39304
rect -28516 -51374 -28510 -39310
rect -28510 -51374 -12606 -39310
rect -12606 -51374 -12600 -39310
rect 12600 -51312 12606 -39248
rect 12606 -51312 28510 -39248
rect 28510 -51312 28516 -39248
rect 12600 -51318 28516 -51312
rect -28516 -51380 -12600 -51374
<< metal5 >>
rect -28540 -39304 -12576 -39280
rect -28540 -51380 -28516 -39304
rect -12600 -51380 -12576 -39304
rect -650 -39342 650 -34514
rect 12576 -39242 28540 -39218
tri -4600 -41342 -2600 -39342 se
rect -2600 -41342 2600 -39342
tri 2600 -41342 4600 -39342 sw
rect -4600 -49342 4600 -41342
tri -4600 -51342 -2600 -49342 ne
rect -2600 -51342 2600 -49342
tri 2600 -51342 4600 -49342 nw
rect 12576 -51318 12600 -39242
rect 28516 -51318 28540 -39242
rect 12576 -51342 28540 -51318
rect -28540 -51404 -12576 -51380
<< fillblock >>
rect -28540 -51404 28540 -34514
<< end >>
