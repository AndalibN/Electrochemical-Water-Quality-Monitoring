magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -852 -1100 858 1100
rect -852 -1112 802 -1100
<< pmos >>
rect -758 -1000 -658 1000
rect -600 -1000 -500 1000
rect -442 -1000 -342 1000
rect -284 -1000 -184 1000
rect -126 -1000 -26 1000
rect 32 -1000 132 1000
rect 190 -1000 290 1000
rect 348 -1000 448 1000
rect 506 -1000 606 1000
rect 664 -1000 764 1000
<< pdiff >>
rect -816 969 -758 1000
rect -816 935 -804 969
rect -770 935 -758 969
rect -816 901 -758 935
rect -816 867 -804 901
rect -770 867 -758 901
rect -816 833 -758 867
rect -816 799 -804 833
rect -770 799 -758 833
rect -816 765 -758 799
rect -816 731 -804 765
rect -770 731 -758 765
rect -816 697 -758 731
rect -816 663 -804 697
rect -770 663 -758 697
rect -816 629 -758 663
rect -816 595 -804 629
rect -770 595 -758 629
rect -816 561 -758 595
rect -816 527 -804 561
rect -770 527 -758 561
rect -816 493 -758 527
rect -816 459 -804 493
rect -770 459 -758 493
rect -816 425 -758 459
rect -816 391 -804 425
rect -770 391 -758 425
rect -816 357 -758 391
rect -816 323 -804 357
rect -770 323 -758 357
rect -816 289 -758 323
rect -816 255 -804 289
rect -770 255 -758 289
rect -816 221 -758 255
rect -816 187 -804 221
rect -770 187 -758 221
rect -816 153 -758 187
rect -816 119 -804 153
rect -770 119 -758 153
rect -816 85 -758 119
rect -816 51 -804 85
rect -770 51 -758 85
rect -816 17 -758 51
rect -816 -17 -804 17
rect -770 -17 -758 17
rect -816 -51 -758 -17
rect -816 -85 -804 -51
rect -770 -85 -758 -51
rect -816 -119 -758 -85
rect -816 -153 -804 -119
rect -770 -153 -758 -119
rect -816 -187 -758 -153
rect -816 -221 -804 -187
rect -770 -221 -758 -187
rect -816 -255 -758 -221
rect -816 -289 -804 -255
rect -770 -289 -758 -255
rect -816 -323 -758 -289
rect -816 -357 -804 -323
rect -770 -357 -758 -323
rect -816 -391 -758 -357
rect -816 -425 -804 -391
rect -770 -425 -758 -391
rect -816 -459 -758 -425
rect -816 -493 -804 -459
rect -770 -493 -758 -459
rect -816 -527 -758 -493
rect -816 -561 -804 -527
rect -770 -561 -758 -527
rect -816 -595 -758 -561
rect -816 -629 -804 -595
rect -770 -629 -758 -595
rect -816 -663 -758 -629
rect -816 -697 -804 -663
rect -770 -697 -758 -663
rect -816 -731 -758 -697
rect -816 -765 -804 -731
rect -770 -765 -758 -731
rect -816 -799 -758 -765
rect -816 -833 -804 -799
rect -770 -833 -758 -799
rect -816 -867 -758 -833
rect -816 -901 -804 -867
rect -770 -901 -758 -867
rect -816 -935 -758 -901
rect -816 -969 -804 -935
rect -770 -969 -758 -935
rect -816 -1000 -758 -969
rect -658 969 -600 1000
rect -658 935 -646 969
rect -612 935 -600 969
rect -658 901 -600 935
rect -658 867 -646 901
rect -612 867 -600 901
rect -658 833 -600 867
rect -658 799 -646 833
rect -612 799 -600 833
rect -658 765 -600 799
rect -658 731 -646 765
rect -612 731 -600 765
rect -658 697 -600 731
rect -658 663 -646 697
rect -612 663 -600 697
rect -658 629 -600 663
rect -658 595 -646 629
rect -612 595 -600 629
rect -658 561 -600 595
rect -658 527 -646 561
rect -612 527 -600 561
rect -658 493 -600 527
rect -658 459 -646 493
rect -612 459 -600 493
rect -658 425 -600 459
rect -658 391 -646 425
rect -612 391 -600 425
rect -658 357 -600 391
rect -658 323 -646 357
rect -612 323 -600 357
rect -658 289 -600 323
rect -658 255 -646 289
rect -612 255 -600 289
rect -658 221 -600 255
rect -658 187 -646 221
rect -612 187 -600 221
rect -658 153 -600 187
rect -658 119 -646 153
rect -612 119 -600 153
rect -658 85 -600 119
rect -658 51 -646 85
rect -612 51 -600 85
rect -658 17 -600 51
rect -658 -17 -646 17
rect -612 -17 -600 17
rect -658 -51 -600 -17
rect -658 -85 -646 -51
rect -612 -85 -600 -51
rect -658 -119 -600 -85
rect -658 -153 -646 -119
rect -612 -153 -600 -119
rect -658 -187 -600 -153
rect -658 -221 -646 -187
rect -612 -221 -600 -187
rect -658 -255 -600 -221
rect -658 -289 -646 -255
rect -612 -289 -600 -255
rect -658 -323 -600 -289
rect -658 -357 -646 -323
rect -612 -357 -600 -323
rect -658 -391 -600 -357
rect -658 -425 -646 -391
rect -612 -425 -600 -391
rect -658 -459 -600 -425
rect -658 -493 -646 -459
rect -612 -493 -600 -459
rect -658 -527 -600 -493
rect -658 -561 -646 -527
rect -612 -561 -600 -527
rect -658 -595 -600 -561
rect -658 -629 -646 -595
rect -612 -629 -600 -595
rect -658 -663 -600 -629
rect -658 -697 -646 -663
rect -612 -697 -600 -663
rect -658 -731 -600 -697
rect -658 -765 -646 -731
rect -612 -765 -600 -731
rect -658 -799 -600 -765
rect -658 -833 -646 -799
rect -612 -833 -600 -799
rect -658 -867 -600 -833
rect -658 -901 -646 -867
rect -612 -901 -600 -867
rect -658 -935 -600 -901
rect -658 -969 -646 -935
rect -612 -969 -600 -935
rect -658 -1000 -600 -969
rect -500 969 -442 1000
rect -500 935 -488 969
rect -454 935 -442 969
rect -500 901 -442 935
rect -500 867 -488 901
rect -454 867 -442 901
rect -500 833 -442 867
rect -500 799 -488 833
rect -454 799 -442 833
rect -500 765 -442 799
rect -500 731 -488 765
rect -454 731 -442 765
rect -500 697 -442 731
rect -500 663 -488 697
rect -454 663 -442 697
rect -500 629 -442 663
rect -500 595 -488 629
rect -454 595 -442 629
rect -500 561 -442 595
rect -500 527 -488 561
rect -454 527 -442 561
rect -500 493 -442 527
rect -500 459 -488 493
rect -454 459 -442 493
rect -500 425 -442 459
rect -500 391 -488 425
rect -454 391 -442 425
rect -500 357 -442 391
rect -500 323 -488 357
rect -454 323 -442 357
rect -500 289 -442 323
rect -500 255 -488 289
rect -454 255 -442 289
rect -500 221 -442 255
rect -500 187 -488 221
rect -454 187 -442 221
rect -500 153 -442 187
rect -500 119 -488 153
rect -454 119 -442 153
rect -500 85 -442 119
rect -500 51 -488 85
rect -454 51 -442 85
rect -500 17 -442 51
rect -500 -17 -488 17
rect -454 -17 -442 17
rect -500 -51 -442 -17
rect -500 -85 -488 -51
rect -454 -85 -442 -51
rect -500 -119 -442 -85
rect -500 -153 -488 -119
rect -454 -153 -442 -119
rect -500 -187 -442 -153
rect -500 -221 -488 -187
rect -454 -221 -442 -187
rect -500 -255 -442 -221
rect -500 -289 -488 -255
rect -454 -289 -442 -255
rect -500 -323 -442 -289
rect -500 -357 -488 -323
rect -454 -357 -442 -323
rect -500 -391 -442 -357
rect -500 -425 -488 -391
rect -454 -425 -442 -391
rect -500 -459 -442 -425
rect -500 -493 -488 -459
rect -454 -493 -442 -459
rect -500 -527 -442 -493
rect -500 -561 -488 -527
rect -454 -561 -442 -527
rect -500 -595 -442 -561
rect -500 -629 -488 -595
rect -454 -629 -442 -595
rect -500 -663 -442 -629
rect -500 -697 -488 -663
rect -454 -697 -442 -663
rect -500 -731 -442 -697
rect -500 -765 -488 -731
rect -454 -765 -442 -731
rect -500 -799 -442 -765
rect -500 -833 -488 -799
rect -454 -833 -442 -799
rect -500 -867 -442 -833
rect -500 -901 -488 -867
rect -454 -901 -442 -867
rect -500 -935 -442 -901
rect -500 -969 -488 -935
rect -454 -969 -442 -935
rect -500 -1000 -442 -969
rect -342 969 -284 1000
rect -342 935 -330 969
rect -296 935 -284 969
rect -342 901 -284 935
rect -342 867 -330 901
rect -296 867 -284 901
rect -342 833 -284 867
rect -342 799 -330 833
rect -296 799 -284 833
rect -342 765 -284 799
rect -342 731 -330 765
rect -296 731 -284 765
rect -342 697 -284 731
rect -342 663 -330 697
rect -296 663 -284 697
rect -342 629 -284 663
rect -342 595 -330 629
rect -296 595 -284 629
rect -342 561 -284 595
rect -342 527 -330 561
rect -296 527 -284 561
rect -342 493 -284 527
rect -342 459 -330 493
rect -296 459 -284 493
rect -342 425 -284 459
rect -342 391 -330 425
rect -296 391 -284 425
rect -342 357 -284 391
rect -342 323 -330 357
rect -296 323 -284 357
rect -342 289 -284 323
rect -342 255 -330 289
rect -296 255 -284 289
rect -342 221 -284 255
rect -342 187 -330 221
rect -296 187 -284 221
rect -342 153 -284 187
rect -342 119 -330 153
rect -296 119 -284 153
rect -342 85 -284 119
rect -342 51 -330 85
rect -296 51 -284 85
rect -342 17 -284 51
rect -342 -17 -330 17
rect -296 -17 -284 17
rect -342 -51 -284 -17
rect -342 -85 -330 -51
rect -296 -85 -284 -51
rect -342 -119 -284 -85
rect -342 -153 -330 -119
rect -296 -153 -284 -119
rect -342 -187 -284 -153
rect -342 -221 -330 -187
rect -296 -221 -284 -187
rect -342 -255 -284 -221
rect -342 -289 -330 -255
rect -296 -289 -284 -255
rect -342 -323 -284 -289
rect -342 -357 -330 -323
rect -296 -357 -284 -323
rect -342 -391 -284 -357
rect -342 -425 -330 -391
rect -296 -425 -284 -391
rect -342 -459 -284 -425
rect -342 -493 -330 -459
rect -296 -493 -284 -459
rect -342 -527 -284 -493
rect -342 -561 -330 -527
rect -296 -561 -284 -527
rect -342 -595 -284 -561
rect -342 -629 -330 -595
rect -296 -629 -284 -595
rect -342 -663 -284 -629
rect -342 -697 -330 -663
rect -296 -697 -284 -663
rect -342 -731 -284 -697
rect -342 -765 -330 -731
rect -296 -765 -284 -731
rect -342 -799 -284 -765
rect -342 -833 -330 -799
rect -296 -833 -284 -799
rect -342 -867 -284 -833
rect -342 -901 -330 -867
rect -296 -901 -284 -867
rect -342 -935 -284 -901
rect -342 -969 -330 -935
rect -296 -969 -284 -935
rect -342 -1000 -284 -969
rect -184 969 -126 1000
rect -184 935 -172 969
rect -138 935 -126 969
rect -184 901 -126 935
rect -184 867 -172 901
rect -138 867 -126 901
rect -184 833 -126 867
rect -184 799 -172 833
rect -138 799 -126 833
rect -184 765 -126 799
rect -184 731 -172 765
rect -138 731 -126 765
rect -184 697 -126 731
rect -184 663 -172 697
rect -138 663 -126 697
rect -184 629 -126 663
rect -184 595 -172 629
rect -138 595 -126 629
rect -184 561 -126 595
rect -184 527 -172 561
rect -138 527 -126 561
rect -184 493 -126 527
rect -184 459 -172 493
rect -138 459 -126 493
rect -184 425 -126 459
rect -184 391 -172 425
rect -138 391 -126 425
rect -184 357 -126 391
rect -184 323 -172 357
rect -138 323 -126 357
rect -184 289 -126 323
rect -184 255 -172 289
rect -138 255 -126 289
rect -184 221 -126 255
rect -184 187 -172 221
rect -138 187 -126 221
rect -184 153 -126 187
rect -184 119 -172 153
rect -138 119 -126 153
rect -184 85 -126 119
rect -184 51 -172 85
rect -138 51 -126 85
rect -184 17 -126 51
rect -184 -17 -172 17
rect -138 -17 -126 17
rect -184 -51 -126 -17
rect -184 -85 -172 -51
rect -138 -85 -126 -51
rect -184 -119 -126 -85
rect -184 -153 -172 -119
rect -138 -153 -126 -119
rect -184 -187 -126 -153
rect -184 -221 -172 -187
rect -138 -221 -126 -187
rect -184 -255 -126 -221
rect -184 -289 -172 -255
rect -138 -289 -126 -255
rect -184 -323 -126 -289
rect -184 -357 -172 -323
rect -138 -357 -126 -323
rect -184 -391 -126 -357
rect -184 -425 -172 -391
rect -138 -425 -126 -391
rect -184 -459 -126 -425
rect -184 -493 -172 -459
rect -138 -493 -126 -459
rect -184 -527 -126 -493
rect -184 -561 -172 -527
rect -138 -561 -126 -527
rect -184 -595 -126 -561
rect -184 -629 -172 -595
rect -138 -629 -126 -595
rect -184 -663 -126 -629
rect -184 -697 -172 -663
rect -138 -697 -126 -663
rect -184 -731 -126 -697
rect -184 -765 -172 -731
rect -138 -765 -126 -731
rect -184 -799 -126 -765
rect -184 -833 -172 -799
rect -138 -833 -126 -799
rect -184 -867 -126 -833
rect -184 -901 -172 -867
rect -138 -901 -126 -867
rect -184 -935 -126 -901
rect -184 -969 -172 -935
rect -138 -969 -126 -935
rect -184 -1000 -126 -969
rect -26 969 32 1000
rect -26 935 -14 969
rect 20 935 32 969
rect -26 901 32 935
rect -26 867 -14 901
rect 20 867 32 901
rect -26 833 32 867
rect -26 799 -14 833
rect 20 799 32 833
rect -26 765 32 799
rect -26 731 -14 765
rect 20 731 32 765
rect -26 697 32 731
rect -26 663 -14 697
rect 20 663 32 697
rect -26 629 32 663
rect -26 595 -14 629
rect 20 595 32 629
rect -26 561 32 595
rect -26 527 -14 561
rect 20 527 32 561
rect -26 493 32 527
rect -26 459 -14 493
rect 20 459 32 493
rect -26 425 32 459
rect -26 391 -14 425
rect 20 391 32 425
rect -26 357 32 391
rect -26 323 -14 357
rect 20 323 32 357
rect -26 289 32 323
rect -26 255 -14 289
rect 20 255 32 289
rect -26 221 32 255
rect -26 187 -14 221
rect 20 187 32 221
rect -26 153 32 187
rect -26 119 -14 153
rect 20 119 32 153
rect -26 85 32 119
rect -26 51 -14 85
rect 20 51 32 85
rect -26 17 32 51
rect -26 -17 -14 17
rect 20 -17 32 17
rect -26 -51 32 -17
rect -26 -85 -14 -51
rect 20 -85 32 -51
rect -26 -119 32 -85
rect -26 -153 -14 -119
rect 20 -153 32 -119
rect -26 -187 32 -153
rect -26 -221 -14 -187
rect 20 -221 32 -187
rect -26 -255 32 -221
rect -26 -289 -14 -255
rect 20 -289 32 -255
rect -26 -323 32 -289
rect -26 -357 -14 -323
rect 20 -357 32 -323
rect -26 -391 32 -357
rect -26 -425 -14 -391
rect 20 -425 32 -391
rect -26 -459 32 -425
rect -26 -493 -14 -459
rect 20 -493 32 -459
rect -26 -527 32 -493
rect -26 -561 -14 -527
rect 20 -561 32 -527
rect -26 -595 32 -561
rect -26 -629 -14 -595
rect 20 -629 32 -595
rect -26 -663 32 -629
rect -26 -697 -14 -663
rect 20 -697 32 -663
rect -26 -731 32 -697
rect -26 -765 -14 -731
rect 20 -765 32 -731
rect -26 -799 32 -765
rect -26 -833 -14 -799
rect 20 -833 32 -799
rect -26 -867 32 -833
rect -26 -901 -14 -867
rect 20 -901 32 -867
rect -26 -935 32 -901
rect -26 -969 -14 -935
rect 20 -969 32 -935
rect -26 -1000 32 -969
rect 132 969 190 1000
rect 132 935 144 969
rect 178 935 190 969
rect 132 901 190 935
rect 132 867 144 901
rect 178 867 190 901
rect 132 833 190 867
rect 132 799 144 833
rect 178 799 190 833
rect 132 765 190 799
rect 132 731 144 765
rect 178 731 190 765
rect 132 697 190 731
rect 132 663 144 697
rect 178 663 190 697
rect 132 629 190 663
rect 132 595 144 629
rect 178 595 190 629
rect 132 561 190 595
rect 132 527 144 561
rect 178 527 190 561
rect 132 493 190 527
rect 132 459 144 493
rect 178 459 190 493
rect 132 425 190 459
rect 132 391 144 425
rect 178 391 190 425
rect 132 357 190 391
rect 132 323 144 357
rect 178 323 190 357
rect 132 289 190 323
rect 132 255 144 289
rect 178 255 190 289
rect 132 221 190 255
rect 132 187 144 221
rect 178 187 190 221
rect 132 153 190 187
rect 132 119 144 153
rect 178 119 190 153
rect 132 85 190 119
rect 132 51 144 85
rect 178 51 190 85
rect 132 17 190 51
rect 132 -17 144 17
rect 178 -17 190 17
rect 132 -51 190 -17
rect 132 -85 144 -51
rect 178 -85 190 -51
rect 132 -119 190 -85
rect 132 -153 144 -119
rect 178 -153 190 -119
rect 132 -187 190 -153
rect 132 -221 144 -187
rect 178 -221 190 -187
rect 132 -255 190 -221
rect 132 -289 144 -255
rect 178 -289 190 -255
rect 132 -323 190 -289
rect 132 -357 144 -323
rect 178 -357 190 -323
rect 132 -391 190 -357
rect 132 -425 144 -391
rect 178 -425 190 -391
rect 132 -459 190 -425
rect 132 -493 144 -459
rect 178 -493 190 -459
rect 132 -527 190 -493
rect 132 -561 144 -527
rect 178 -561 190 -527
rect 132 -595 190 -561
rect 132 -629 144 -595
rect 178 -629 190 -595
rect 132 -663 190 -629
rect 132 -697 144 -663
rect 178 -697 190 -663
rect 132 -731 190 -697
rect 132 -765 144 -731
rect 178 -765 190 -731
rect 132 -799 190 -765
rect 132 -833 144 -799
rect 178 -833 190 -799
rect 132 -867 190 -833
rect 132 -901 144 -867
rect 178 -901 190 -867
rect 132 -935 190 -901
rect 132 -969 144 -935
rect 178 -969 190 -935
rect 132 -1000 190 -969
rect 290 969 348 1000
rect 290 935 302 969
rect 336 935 348 969
rect 290 901 348 935
rect 290 867 302 901
rect 336 867 348 901
rect 290 833 348 867
rect 290 799 302 833
rect 336 799 348 833
rect 290 765 348 799
rect 290 731 302 765
rect 336 731 348 765
rect 290 697 348 731
rect 290 663 302 697
rect 336 663 348 697
rect 290 629 348 663
rect 290 595 302 629
rect 336 595 348 629
rect 290 561 348 595
rect 290 527 302 561
rect 336 527 348 561
rect 290 493 348 527
rect 290 459 302 493
rect 336 459 348 493
rect 290 425 348 459
rect 290 391 302 425
rect 336 391 348 425
rect 290 357 348 391
rect 290 323 302 357
rect 336 323 348 357
rect 290 289 348 323
rect 290 255 302 289
rect 336 255 348 289
rect 290 221 348 255
rect 290 187 302 221
rect 336 187 348 221
rect 290 153 348 187
rect 290 119 302 153
rect 336 119 348 153
rect 290 85 348 119
rect 290 51 302 85
rect 336 51 348 85
rect 290 17 348 51
rect 290 -17 302 17
rect 336 -17 348 17
rect 290 -51 348 -17
rect 290 -85 302 -51
rect 336 -85 348 -51
rect 290 -119 348 -85
rect 290 -153 302 -119
rect 336 -153 348 -119
rect 290 -187 348 -153
rect 290 -221 302 -187
rect 336 -221 348 -187
rect 290 -255 348 -221
rect 290 -289 302 -255
rect 336 -289 348 -255
rect 290 -323 348 -289
rect 290 -357 302 -323
rect 336 -357 348 -323
rect 290 -391 348 -357
rect 290 -425 302 -391
rect 336 -425 348 -391
rect 290 -459 348 -425
rect 290 -493 302 -459
rect 336 -493 348 -459
rect 290 -527 348 -493
rect 290 -561 302 -527
rect 336 -561 348 -527
rect 290 -595 348 -561
rect 290 -629 302 -595
rect 336 -629 348 -595
rect 290 -663 348 -629
rect 290 -697 302 -663
rect 336 -697 348 -663
rect 290 -731 348 -697
rect 290 -765 302 -731
rect 336 -765 348 -731
rect 290 -799 348 -765
rect 290 -833 302 -799
rect 336 -833 348 -799
rect 290 -867 348 -833
rect 290 -901 302 -867
rect 336 -901 348 -867
rect 290 -935 348 -901
rect 290 -969 302 -935
rect 336 -969 348 -935
rect 290 -1000 348 -969
rect 448 969 506 1000
rect 448 935 460 969
rect 494 935 506 969
rect 448 901 506 935
rect 448 867 460 901
rect 494 867 506 901
rect 448 833 506 867
rect 448 799 460 833
rect 494 799 506 833
rect 448 765 506 799
rect 448 731 460 765
rect 494 731 506 765
rect 448 697 506 731
rect 448 663 460 697
rect 494 663 506 697
rect 448 629 506 663
rect 448 595 460 629
rect 494 595 506 629
rect 448 561 506 595
rect 448 527 460 561
rect 494 527 506 561
rect 448 493 506 527
rect 448 459 460 493
rect 494 459 506 493
rect 448 425 506 459
rect 448 391 460 425
rect 494 391 506 425
rect 448 357 506 391
rect 448 323 460 357
rect 494 323 506 357
rect 448 289 506 323
rect 448 255 460 289
rect 494 255 506 289
rect 448 221 506 255
rect 448 187 460 221
rect 494 187 506 221
rect 448 153 506 187
rect 448 119 460 153
rect 494 119 506 153
rect 448 85 506 119
rect 448 51 460 85
rect 494 51 506 85
rect 448 17 506 51
rect 448 -17 460 17
rect 494 -17 506 17
rect 448 -51 506 -17
rect 448 -85 460 -51
rect 494 -85 506 -51
rect 448 -119 506 -85
rect 448 -153 460 -119
rect 494 -153 506 -119
rect 448 -187 506 -153
rect 448 -221 460 -187
rect 494 -221 506 -187
rect 448 -255 506 -221
rect 448 -289 460 -255
rect 494 -289 506 -255
rect 448 -323 506 -289
rect 448 -357 460 -323
rect 494 -357 506 -323
rect 448 -391 506 -357
rect 448 -425 460 -391
rect 494 -425 506 -391
rect 448 -459 506 -425
rect 448 -493 460 -459
rect 494 -493 506 -459
rect 448 -527 506 -493
rect 448 -561 460 -527
rect 494 -561 506 -527
rect 448 -595 506 -561
rect 448 -629 460 -595
rect 494 -629 506 -595
rect 448 -663 506 -629
rect 448 -697 460 -663
rect 494 -697 506 -663
rect 448 -731 506 -697
rect 448 -765 460 -731
rect 494 -765 506 -731
rect 448 -799 506 -765
rect 448 -833 460 -799
rect 494 -833 506 -799
rect 448 -867 506 -833
rect 448 -901 460 -867
rect 494 -901 506 -867
rect 448 -935 506 -901
rect 448 -969 460 -935
rect 494 -969 506 -935
rect 448 -1000 506 -969
rect 606 969 664 1000
rect 606 935 618 969
rect 652 935 664 969
rect 606 901 664 935
rect 606 867 618 901
rect 652 867 664 901
rect 606 833 664 867
rect 606 799 618 833
rect 652 799 664 833
rect 606 765 664 799
rect 606 731 618 765
rect 652 731 664 765
rect 606 697 664 731
rect 606 663 618 697
rect 652 663 664 697
rect 606 629 664 663
rect 606 595 618 629
rect 652 595 664 629
rect 606 561 664 595
rect 606 527 618 561
rect 652 527 664 561
rect 606 493 664 527
rect 606 459 618 493
rect 652 459 664 493
rect 606 425 664 459
rect 606 391 618 425
rect 652 391 664 425
rect 606 357 664 391
rect 606 323 618 357
rect 652 323 664 357
rect 606 289 664 323
rect 606 255 618 289
rect 652 255 664 289
rect 606 221 664 255
rect 606 187 618 221
rect 652 187 664 221
rect 606 153 664 187
rect 606 119 618 153
rect 652 119 664 153
rect 606 85 664 119
rect 606 51 618 85
rect 652 51 664 85
rect 606 17 664 51
rect 606 -17 618 17
rect 652 -17 664 17
rect 606 -51 664 -17
rect 606 -85 618 -51
rect 652 -85 664 -51
rect 606 -119 664 -85
rect 606 -153 618 -119
rect 652 -153 664 -119
rect 606 -187 664 -153
rect 606 -221 618 -187
rect 652 -221 664 -187
rect 606 -255 664 -221
rect 606 -289 618 -255
rect 652 -289 664 -255
rect 606 -323 664 -289
rect 606 -357 618 -323
rect 652 -357 664 -323
rect 606 -391 664 -357
rect 606 -425 618 -391
rect 652 -425 664 -391
rect 606 -459 664 -425
rect 606 -493 618 -459
rect 652 -493 664 -459
rect 606 -527 664 -493
rect 606 -561 618 -527
rect 652 -561 664 -527
rect 606 -595 664 -561
rect 606 -629 618 -595
rect 652 -629 664 -595
rect 606 -663 664 -629
rect 606 -697 618 -663
rect 652 -697 664 -663
rect 606 -731 664 -697
rect 606 -765 618 -731
rect 652 -765 664 -731
rect 606 -799 664 -765
rect 606 -833 618 -799
rect 652 -833 664 -799
rect 606 -867 664 -833
rect 606 -901 618 -867
rect 652 -901 664 -867
rect 606 -935 664 -901
rect 606 -969 618 -935
rect 652 -969 664 -935
rect 606 -1000 664 -969
rect 764 969 822 1000
rect 764 935 776 969
rect 810 935 822 969
rect 764 901 822 935
rect 764 867 776 901
rect 810 867 822 901
rect 764 833 822 867
rect 764 799 776 833
rect 810 799 822 833
rect 764 765 822 799
rect 764 731 776 765
rect 810 731 822 765
rect 764 697 822 731
rect 764 663 776 697
rect 810 663 822 697
rect 764 629 822 663
rect 764 595 776 629
rect 810 595 822 629
rect 764 561 822 595
rect 764 527 776 561
rect 810 527 822 561
rect 764 493 822 527
rect 764 459 776 493
rect 810 459 822 493
rect 764 425 822 459
rect 764 391 776 425
rect 810 391 822 425
rect 764 357 822 391
rect 764 323 776 357
rect 810 323 822 357
rect 764 289 822 323
rect 764 255 776 289
rect 810 255 822 289
rect 764 221 822 255
rect 764 187 776 221
rect 810 187 822 221
rect 764 153 822 187
rect 764 119 776 153
rect 810 119 822 153
rect 764 85 822 119
rect 764 51 776 85
rect 810 51 822 85
rect 764 17 822 51
rect 764 -17 776 17
rect 810 -17 822 17
rect 764 -51 822 -17
rect 764 -85 776 -51
rect 810 -85 822 -51
rect 764 -119 822 -85
rect 764 -153 776 -119
rect 810 -153 822 -119
rect 764 -187 822 -153
rect 764 -221 776 -187
rect 810 -221 822 -187
rect 764 -255 822 -221
rect 764 -289 776 -255
rect 810 -289 822 -255
rect 764 -323 822 -289
rect 764 -357 776 -323
rect 810 -357 822 -323
rect 764 -391 822 -357
rect 764 -425 776 -391
rect 810 -425 822 -391
rect 764 -459 822 -425
rect 764 -493 776 -459
rect 810 -493 822 -459
rect 764 -527 822 -493
rect 764 -561 776 -527
rect 810 -561 822 -527
rect 764 -595 822 -561
rect 764 -629 776 -595
rect 810 -629 822 -595
rect 764 -663 822 -629
rect 764 -697 776 -663
rect 810 -697 822 -663
rect 764 -731 822 -697
rect 764 -765 776 -731
rect 810 -765 822 -731
rect 764 -799 822 -765
rect 764 -833 776 -799
rect 810 -833 822 -799
rect 764 -867 822 -833
rect 764 -901 776 -867
rect 810 -901 822 -867
rect 764 -935 822 -901
rect 764 -969 776 -935
rect 810 -969 822 -935
rect 764 -1000 822 -969
<< pdiffc >>
rect -804 935 -770 969
rect -804 867 -770 901
rect -804 799 -770 833
rect -804 731 -770 765
rect -804 663 -770 697
rect -804 595 -770 629
rect -804 527 -770 561
rect -804 459 -770 493
rect -804 391 -770 425
rect -804 323 -770 357
rect -804 255 -770 289
rect -804 187 -770 221
rect -804 119 -770 153
rect -804 51 -770 85
rect -804 -17 -770 17
rect -804 -85 -770 -51
rect -804 -153 -770 -119
rect -804 -221 -770 -187
rect -804 -289 -770 -255
rect -804 -357 -770 -323
rect -804 -425 -770 -391
rect -804 -493 -770 -459
rect -804 -561 -770 -527
rect -804 -629 -770 -595
rect -804 -697 -770 -663
rect -804 -765 -770 -731
rect -804 -833 -770 -799
rect -804 -901 -770 -867
rect -804 -969 -770 -935
rect -646 935 -612 969
rect -646 867 -612 901
rect -646 799 -612 833
rect -646 731 -612 765
rect -646 663 -612 697
rect -646 595 -612 629
rect -646 527 -612 561
rect -646 459 -612 493
rect -646 391 -612 425
rect -646 323 -612 357
rect -646 255 -612 289
rect -646 187 -612 221
rect -646 119 -612 153
rect -646 51 -612 85
rect -646 -17 -612 17
rect -646 -85 -612 -51
rect -646 -153 -612 -119
rect -646 -221 -612 -187
rect -646 -289 -612 -255
rect -646 -357 -612 -323
rect -646 -425 -612 -391
rect -646 -493 -612 -459
rect -646 -561 -612 -527
rect -646 -629 -612 -595
rect -646 -697 -612 -663
rect -646 -765 -612 -731
rect -646 -833 -612 -799
rect -646 -901 -612 -867
rect -646 -969 -612 -935
rect -488 935 -454 969
rect -488 867 -454 901
rect -488 799 -454 833
rect -488 731 -454 765
rect -488 663 -454 697
rect -488 595 -454 629
rect -488 527 -454 561
rect -488 459 -454 493
rect -488 391 -454 425
rect -488 323 -454 357
rect -488 255 -454 289
rect -488 187 -454 221
rect -488 119 -454 153
rect -488 51 -454 85
rect -488 -17 -454 17
rect -488 -85 -454 -51
rect -488 -153 -454 -119
rect -488 -221 -454 -187
rect -488 -289 -454 -255
rect -488 -357 -454 -323
rect -488 -425 -454 -391
rect -488 -493 -454 -459
rect -488 -561 -454 -527
rect -488 -629 -454 -595
rect -488 -697 -454 -663
rect -488 -765 -454 -731
rect -488 -833 -454 -799
rect -488 -901 -454 -867
rect -488 -969 -454 -935
rect -330 935 -296 969
rect -330 867 -296 901
rect -330 799 -296 833
rect -330 731 -296 765
rect -330 663 -296 697
rect -330 595 -296 629
rect -330 527 -296 561
rect -330 459 -296 493
rect -330 391 -296 425
rect -330 323 -296 357
rect -330 255 -296 289
rect -330 187 -296 221
rect -330 119 -296 153
rect -330 51 -296 85
rect -330 -17 -296 17
rect -330 -85 -296 -51
rect -330 -153 -296 -119
rect -330 -221 -296 -187
rect -330 -289 -296 -255
rect -330 -357 -296 -323
rect -330 -425 -296 -391
rect -330 -493 -296 -459
rect -330 -561 -296 -527
rect -330 -629 -296 -595
rect -330 -697 -296 -663
rect -330 -765 -296 -731
rect -330 -833 -296 -799
rect -330 -901 -296 -867
rect -330 -969 -296 -935
rect -172 935 -138 969
rect -172 867 -138 901
rect -172 799 -138 833
rect -172 731 -138 765
rect -172 663 -138 697
rect -172 595 -138 629
rect -172 527 -138 561
rect -172 459 -138 493
rect -172 391 -138 425
rect -172 323 -138 357
rect -172 255 -138 289
rect -172 187 -138 221
rect -172 119 -138 153
rect -172 51 -138 85
rect -172 -17 -138 17
rect -172 -85 -138 -51
rect -172 -153 -138 -119
rect -172 -221 -138 -187
rect -172 -289 -138 -255
rect -172 -357 -138 -323
rect -172 -425 -138 -391
rect -172 -493 -138 -459
rect -172 -561 -138 -527
rect -172 -629 -138 -595
rect -172 -697 -138 -663
rect -172 -765 -138 -731
rect -172 -833 -138 -799
rect -172 -901 -138 -867
rect -172 -969 -138 -935
rect -14 935 20 969
rect -14 867 20 901
rect -14 799 20 833
rect -14 731 20 765
rect -14 663 20 697
rect -14 595 20 629
rect -14 527 20 561
rect -14 459 20 493
rect -14 391 20 425
rect -14 323 20 357
rect -14 255 20 289
rect -14 187 20 221
rect -14 119 20 153
rect -14 51 20 85
rect -14 -17 20 17
rect -14 -85 20 -51
rect -14 -153 20 -119
rect -14 -221 20 -187
rect -14 -289 20 -255
rect -14 -357 20 -323
rect -14 -425 20 -391
rect -14 -493 20 -459
rect -14 -561 20 -527
rect -14 -629 20 -595
rect -14 -697 20 -663
rect -14 -765 20 -731
rect -14 -833 20 -799
rect -14 -901 20 -867
rect -14 -969 20 -935
rect 144 935 178 969
rect 144 867 178 901
rect 144 799 178 833
rect 144 731 178 765
rect 144 663 178 697
rect 144 595 178 629
rect 144 527 178 561
rect 144 459 178 493
rect 144 391 178 425
rect 144 323 178 357
rect 144 255 178 289
rect 144 187 178 221
rect 144 119 178 153
rect 144 51 178 85
rect 144 -17 178 17
rect 144 -85 178 -51
rect 144 -153 178 -119
rect 144 -221 178 -187
rect 144 -289 178 -255
rect 144 -357 178 -323
rect 144 -425 178 -391
rect 144 -493 178 -459
rect 144 -561 178 -527
rect 144 -629 178 -595
rect 144 -697 178 -663
rect 144 -765 178 -731
rect 144 -833 178 -799
rect 144 -901 178 -867
rect 144 -969 178 -935
rect 302 935 336 969
rect 302 867 336 901
rect 302 799 336 833
rect 302 731 336 765
rect 302 663 336 697
rect 302 595 336 629
rect 302 527 336 561
rect 302 459 336 493
rect 302 391 336 425
rect 302 323 336 357
rect 302 255 336 289
rect 302 187 336 221
rect 302 119 336 153
rect 302 51 336 85
rect 302 -17 336 17
rect 302 -85 336 -51
rect 302 -153 336 -119
rect 302 -221 336 -187
rect 302 -289 336 -255
rect 302 -357 336 -323
rect 302 -425 336 -391
rect 302 -493 336 -459
rect 302 -561 336 -527
rect 302 -629 336 -595
rect 302 -697 336 -663
rect 302 -765 336 -731
rect 302 -833 336 -799
rect 302 -901 336 -867
rect 302 -969 336 -935
rect 460 935 494 969
rect 460 867 494 901
rect 460 799 494 833
rect 460 731 494 765
rect 460 663 494 697
rect 460 595 494 629
rect 460 527 494 561
rect 460 459 494 493
rect 460 391 494 425
rect 460 323 494 357
rect 460 255 494 289
rect 460 187 494 221
rect 460 119 494 153
rect 460 51 494 85
rect 460 -17 494 17
rect 460 -85 494 -51
rect 460 -153 494 -119
rect 460 -221 494 -187
rect 460 -289 494 -255
rect 460 -357 494 -323
rect 460 -425 494 -391
rect 460 -493 494 -459
rect 460 -561 494 -527
rect 460 -629 494 -595
rect 460 -697 494 -663
rect 460 -765 494 -731
rect 460 -833 494 -799
rect 460 -901 494 -867
rect 460 -969 494 -935
rect 618 935 652 969
rect 618 867 652 901
rect 618 799 652 833
rect 618 731 652 765
rect 618 663 652 697
rect 618 595 652 629
rect 618 527 652 561
rect 618 459 652 493
rect 618 391 652 425
rect 618 323 652 357
rect 618 255 652 289
rect 618 187 652 221
rect 618 119 652 153
rect 618 51 652 85
rect 618 -17 652 17
rect 618 -85 652 -51
rect 618 -153 652 -119
rect 618 -221 652 -187
rect 618 -289 652 -255
rect 618 -357 652 -323
rect 618 -425 652 -391
rect 618 -493 652 -459
rect 618 -561 652 -527
rect 618 -629 652 -595
rect 618 -697 652 -663
rect 618 -765 652 -731
rect 618 -833 652 -799
rect 618 -901 652 -867
rect 618 -969 652 -935
rect 776 935 810 969
rect 776 867 810 901
rect 776 799 810 833
rect 776 731 810 765
rect 776 663 810 697
rect 776 595 810 629
rect 776 527 810 561
rect 776 459 810 493
rect 776 391 810 425
rect 776 323 810 357
rect 776 255 810 289
rect 776 187 810 221
rect 776 119 810 153
rect 776 51 810 85
rect 776 -17 810 17
rect 776 -85 810 -51
rect 776 -153 810 -119
rect 776 -221 810 -187
rect 776 -289 810 -255
rect 776 -357 810 -323
rect 776 -425 810 -391
rect 776 -493 810 -459
rect 776 -561 810 -527
rect 776 -629 810 -595
rect 776 -697 810 -663
rect 776 -765 810 -731
rect 776 -833 810 -799
rect 776 -901 810 -867
rect 776 -969 810 -935
<< poly >>
rect -758 1046 764 1098
rect -758 1000 -658 1046
rect -600 1000 -500 1046
rect -442 1000 -342 1046
rect -284 1000 -184 1046
rect -126 1000 -26 1046
rect 32 1000 132 1046
rect 190 1000 290 1046
rect 348 1000 448 1046
rect 506 1000 606 1046
rect 664 1000 764 1046
rect -758 -1056 -658 -1000
rect -600 -1056 -500 -1000
rect -442 -1056 -342 -1000
rect -284 -1056 -184 -1000
rect -126 -1056 -26 -1000
rect 32 -1056 132 -1000
rect 190 -1056 290 -1000
rect 348 -1056 448 -1000
rect 506 -1056 606 -1000
rect 664 -1056 764 -1000
rect -758 -1108 764 -1056
<< locali >>
rect -804 969 -770 1004
rect -804 901 -770 919
rect -804 833 -770 847
rect -804 765 -770 775
rect -804 697 -770 703
rect -804 629 -770 631
rect -804 593 -770 595
rect -804 521 -770 527
rect -804 449 -770 459
rect -804 377 -770 391
rect -804 305 -770 323
rect -804 233 -770 255
rect -804 161 -770 187
rect -804 89 -770 119
rect -804 17 -770 51
rect -804 -51 -770 -17
rect -804 -119 -770 -89
rect -804 -187 -770 -161
rect -804 -255 -770 -233
rect -804 -323 -770 -305
rect -804 -391 -770 -377
rect -804 -459 -770 -449
rect -804 -527 -770 -521
rect -804 -595 -770 -593
rect -804 -631 -770 -629
rect -804 -703 -770 -697
rect -804 -775 -770 -765
rect -804 -847 -770 -833
rect -804 -919 -770 -901
rect -804 -1004 -770 -969
rect -646 969 -612 1004
rect -646 901 -612 919
rect -646 833 -612 847
rect -646 765 -612 775
rect -646 697 -612 703
rect -646 629 -612 631
rect -646 593 -612 595
rect -646 521 -612 527
rect -646 449 -612 459
rect -646 377 -612 391
rect -646 305 -612 323
rect -646 233 -612 255
rect -646 161 -612 187
rect -646 89 -612 119
rect -646 17 -612 51
rect -646 -51 -612 -17
rect -646 -119 -612 -89
rect -646 -187 -612 -161
rect -646 -255 -612 -233
rect -646 -323 -612 -305
rect -646 -391 -612 -377
rect -646 -459 -612 -449
rect -646 -527 -612 -521
rect -646 -595 -612 -593
rect -646 -631 -612 -629
rect -646 -703 -612 -697
rect -646 -775 -612 -765
rect -646 -847 -612 -833
rect -646 -919 -612 -901
rect -646 -1004 -612 -969
rect -488 969 -454 1004
rect -488 901 -454 919
rect -488 833 -454 847
rect -488 765 -454 775
rect -488 697 -454 703
rect -488 629 -454 631
rect -488 593 -454 595
rect -488 521 -454 527
rect -488 449 -454 459
rect -488 377 -454 391
rect -488 305 -454 323
rect -488 233 -454 255
rect -488 161 -454 187
rect -488 89 -454 119
rect -488 17 -454 51
rect -488 -51 -454 -17
rect -488 -119 -454 -89
rect -488 -187 -454 -161
rect -488 -255 -454 -233
rect -488 -323 -454 -305
rect -488 -391 -454 -377
rect -488 -459 -454 -449
rect -488 -527 -454 -521
rect -488 -595 -454 -593
rect -488 -631 -454 -629
rect -488 -703 -454 -697
rect -488 -775 -454 -765
rect -488 -847 -454 -833
rect -488 -919 -454 -901
rect -488 -1004 -454 -969
rect -330 969 -296 1004
rect -330 901 -296 919
rect -330 833 -296 847
rect -330 765 -296 775
rect -330 697 -296 703
rect -330 629 -296 631
rect -330 593 -296 595
rect -330 521 -296 527
rect -330 449 -296 459
rect -330 377 -296 391
rect -330 305 -296 323
rect -330 233 -296 255
rect -330 161 -296 187
rect -330 89 -296 119
rect -330 17 -296 51
rect -330 -51 -296 -17
rect -330 -119 -296 -89
rect -330 -187 -296 -161
rect -330 -255 -296 -233
rect -330 -323 -296 -305
rect -330 -391 -296 -377
rect -330 -459 -296 -449
rect -330 -527 -296 -521
rect -330 -595 -296 -593
rect -330 -631 -296 -629
rect -330 -703 -296 -697
rect -330 -775 -296 -765
rect -330 -847 -296 -833
rect -330 -919 -296 -901
rect -330 -1004 -296 -969
rect -172 969 -138 1004
rect -172 901 -138 919
rect -172 833 -138 847
rect -172 765 -138 775
rect -172 697 -138 703
rect -172 629 -138 631
rect -172 593 -138 595
rect -172 521 -138 527
rect -172 449 -138 459
rect -172 377 -138 391
rect -172 305 -138 323
rect -172 233 -138 255
rect -172 161 -138 187
rect -172 89 -138 119
rect -172 17 -138 51
rect -172 -51 -138 -17
rect -172 -119 -138 -89
rect -172 -187 -138 -161
rect -172 -255 -138 -233
rect -172 -323 -138 -305
rect -172 -391 -138 -377
rect -172 -459 -138 -449
rect -172 -527 -138 -521
rect -172 -595 -138 -593
rect -172 -631 -138 -629
rect -172 -703 -138 -697
rect -172 -775 -138 -765
rect -172 -847 -138 -833
rect -172 -919 -138 -901
rect -172 -1004 -138 -969
rect -14 969 20 1004
rect -14 901 20 919
rect -14 833 20 847
rect -14 765 20 775
rect -14 697 20 703
rect -14 629 20 631
rect -14 593 20 595
rect -14 521 20 527
rect -14 449 20 459
rect -14 377 20 391
rect -14 305 20 323
rect -14 233 20 255
rect -14 161 20 187
rect -14 89 20 119
rect -14 17 20 51
rect -14 -51 20 -17
rect -14 -119 20 -89
rect -14 -187 20 -161
rect -14 -255 20 -233
rect -14 -323 20 -305
rect -14 -391 20 -377
rect -14 -459 20 -449
rect -14 -527 20 -521
rect -14 -595 20 -593
rect -14 -631 20 -629
rect -14 -703 20 -697
rect -14 -775 20 -765
rect -14 -847 20 -833
rect -14 -919 20 -901
rect -14 -1004 20 -969
rect 144 969 178 1004
rect 144 901 178 919
rect 144 833 178 847
rect 144 765 178 775
rect 144 697 178 703
rect 144 629 178 631
rect 144 593 178 595
rect 144 521 178 527
rect 144 449 178 459
rect 144 377 178 391
rect 144 305 178 323
rect 144 233 178 255
rect 144 161 178 187
rect 144 89 178 119
rect 144 17 178 51
rect 144 -51 178 -17
rect 144 -119 178 -89
rect 144 -187 178 -161
rect 144 -255 178 -233
rect 144 -323 178 -305
rect 144 -391 178 -377
rect 144 -459 178 -449
rect 144 -527 178 -521
rect 144 -595 178 -593
rect 144 -631 178 -629
rect 144 -703 178 -697
rect 144 -775 178 -765
rect 144 -847 178 -833
rect 144 -919 178 -901
rect 144 -1004 178 -969
rect 302 969 336 1004
rect 302 901 336 919
rect 302 833 336 847
rect 302 765 336 775
rect 302 697 336 703
rect 302 629 336 631
rect 302 593 336 595
rect 302 521 336 527
rect 302 449 336 459
rect 302 377 336 391
rect 302 305 336 323
rect 302 233 336 255
rect 302 161 336 187
rect 302 89 336 119
rect 302 17 336 51
rect 302 -51 336 -17
rect 302 -119 336 -89
rect 302 -187 336 -161
rect 302 -255 336 -233
rect 302 -323 336 -305
rect 302 -391 336 -377
rect 302 -459 336 -449
rect 302 -527 336 -521
rect 302 -595 336 -593
rect 302 -631 336 -629
rect 302 -703 336 -697
rect 302 -775 336 -765
rect 302 -847 336 -833
rect 302 -919 336 -901
rect 302 -1004 336 -969
rect 460 969 494 1004
rect 460 901 494 919
rect 460 833 494 847
rect 460 765 494 775
rect 460 697 494 703
rect 460 629 494 631
rect 460 593 494 595
rect 460 521 494 527
rect 460 449 494 459
rect 460 377 494 391
rect 460 305 494 323
rect 460 233 494 255
rect 460 161 494 187
rect 460 89 494 119
rect 460 17 494 51
rect 460 -51 494 -17
rect 460 -119 494 -89
rect 460 -187 494 -161
rect 460 -255 494 -233
rect 460 -323 494 -305
rect 460 -391 494 -377
rect 460 -459 494 -449
rect 460 -527 494 -521
rect 460 -595 494 -593
rect 460 -631 494 -629
rect 460 -703 494 -697
rect 460 -775 494 -765
rect 460 -847 494 -833
rect 460 -919 494 -901
rect 460 -1004 494 -969
rect 618 969 652 1004
rect 618 901 652 919
rect 618 833 652 847
rect 618 765 652 775
rect 618 697 652 703
rect 618 629 652 631
rect 618 593 652 595
rect 618 521 652 527
rect 618 449 652 459
rect 618 377 652 391
rect 618 305 652 323
rect 618 233 652 255
rect 618 161 652 187
rect 618 89 652 119
rect 618 17 652 51
rect 618 -51 652 -17
rect 618 -119 652 -89
rect 618 -187 652 -161
rect 618 -255 652 -233
rect 618 -323 652 -305
rect 618 -391 652 -377
rect 618 -459 652 -449
rect 618 -527 652 -521
rect 618 -595 652 -593
rect 618 -631 652 -629
rect 618 -703 652 -697
rect 618 -775 652 -765
rect 618 -847 652 -833
rect 618 -919 652 -901
rect 618 -1004 652 -969
rect 776 969 810 1004
rect 776 901 810 919
rect 776 833 810 847
rect 776 765 810 775
rect 776 697 810 703
rect 776 629 810 631
rect 776 593 810 595
rect 776 521 810 527
rect 776 449 810 459
rect 776 377 810 391
rect 776 305 810 323
rect 776 233 810 255
rect 776 161 810 187
rect 776 89 810 119
rect 776 17 810 51
rect 776 -51 810 -17
rect 776 -119 810 -89
rect 776 -187 810 -161
rect 776 -255 810 -233
rect 776 -323 810 -305
rect 776 -391 810 -377
rect 776 -459 810 -449
rect 776 -527 810 -521
rect 776 -595 810 -593
rect 776 -631 810 -629
rect 776 -703 810 -697
rect 776 -775 810 -765
rect 776 -847 810 -833
rect 776 -919 810 -901
rect 776 -1004 810 -969
<< viali >>
rect -804 935 -770 953
rect -804 919 -770 935
rect -804 867 -770 881
rect -804 847 -770 867
rect -804 799 -770 809
rect -804 775 -770 799
rect -804 731 -770 737
rect -804 703 -770 731
rect -804 663 -770 665
rect -804 631 -770 663
rect -804 561 -770 593
rect -804 559 -770 561
rect -804 493 -770 521
rect -804 487 -770 493
rect -804 425 -770 449
rect -804 415 -770 425
rect -804 357 -770 377
rect -804 343 -770 357
rect -804 289 -770 305
rect -804 271 -770 289
rect -804 221 -770 233
rect -804 199 -770 221
rect -804 153 -770 161
rect -804 127 -770 153
rect -804 85 -770 89
rect -804 55 -770 85
rect -804 -17 -770 17
rect -804 -85 -770 -55
rect -804 -89 -770 -85
rect -804 -153 -770 -127
rect -804 -161 -770 -153
rect -804 -221 -770 -199
rect -804 -233 -770 -221
rect -804 -289 -770 -271
rect -804 -305 -770 -289
rect -804 -357 -770 -343
rect -804 -377 -770 -357
rect -804 -425 -770 -415
rect -804 -449 -770 -425
rect -804 -493 -770 -487
rect -804 -521 -770 -493
rect -804 -561 -770 -559
rect -804 -593 -770 -561
rect -804 -663 -770 -631
rect -804 -665 -770 -663
rect -804 -731 -770 -703
rect -804 -737 -770 -731
rect -804 -799 -770 -775
rect -804 -809 -770 -799
rect -804 -867 -770 -847
rect -804 -881 -770 -867
rect -804 -935 -770 -919
rect -804 -953 -770 -935
rect -646 935 -612 953
rect -646 919 -612 935
rect -646 867 -612 881
rect -646 847 -612 867
rect -646 799 -612 809
rect -646 775 -612 799
rect -646 731 -612 737
rect -646 703 -612 731
rect -646 663 -612 665
rect -646 631 -612 663
rect -646 561 -612 593
rect -646 559 -612 561
rect -646 493 -612 521
rect -646 487 -612 493
rect -646 425 -612 449
rect -646 415 -612 425
rect -646 357 -612 377
rect -646 343 -612 357
rect -646 289 -612 305
rect -646 271 -612 289
rect -646 221 -612 233
rect -646 199 -612 221
rect -646 153 -612 161
rect -646 127 -612 153
rect -646 85 -612 89
rect -646 55 -612 85
rect -646 -17 -612 17
rect -646 -85 -612 -55
rect -646 -89 -612 -85
rect -646 -153 -612 -127
rect -646 -161 -612 -153
rect -646 -221 -612 -199
rect -646 -233 -612 -221
rect -646 -289 -612 -271
rect -646 -305 -612 -289
rect -646 -357 -612 -343
rect -646 -377 -612 -357
rect -646 -425 -612 -415
rect -646 -449 -612 -425
rect -646 -493 -612 -487
rect -646 -521 -612 -493
rect -646 -561 -612 -559
rect -646 -593 -612 -561
rect -646 -663 -612 -631
rect -646 -665 -612 -663
rect -646 -731 -612 -703
rect -646 -737 -612 -731
rect -646 -799 -612 -775
rect -646 -809 -612 -799
rect -646 -867 -612 -847
rect -646 -881 -612 -867
rect -646 -935 -612 -919
rect -646 -953 -612 -935
rect -488 935 -454 953
rect -488 919 -454 935
rect -488 867 -454 881
rect -488 847 -454 867
rect -488 799 -454 809
rect -488 775 -454 799
rect -488 731 -454 737
rect -488 703 -454 731
rect -488 663 -454 665
rect -488 631 -454 663
rect -488 561 -454 593
rect -488 559 -454 561
rect -488 493 -454 521
rect -488 487 -454 493
rect -488 425 -454 449
rect -488 415 -454 425
rect -488 357 -454 377
rect -488 343 -454 357
rect -488 289 -454 305
rect -488 271 -454 289
rect -488 221 -454 233
rect -488 199 -454 221
rect -488 153 -454 161
rect -488 127 -454 153
rect -488 85 -454 89
rect -488 55 -454 85
rect -488 -17 -454 17
rect -488 -85 -454 -55
rect -488 -89 -454 -85
rect -488 -153 -454 -127
rect -488 -161 -454 -153
rect -488 -221 -454 -199
rect -488 -233 -454 -221
rect -488 -289 -454 -271
rect -488 -305 -454 -289
rect -488 -357 -454 -343
rect -488 -377 -454 -357
rect -488 -425 -454 -415
rect -488 -449 -454 -425
rect -488 -493 -454 -487
rect -488 -521 -454 -493
rect -488 -561 -454 -559
rect -488 -593 -454 -561
rect -488 -663 -454 -631
rect -488 -665 -454 -663
rect -488 -731 -454 -703
rect -488 -737 -454 -731
rect -488 -799 -454 -775
rect -488 -809 -454 -799
rect -488 -867 -454 -847
rect -488 -881 -454 -867
rect -488 -935 -454 -919
rect -488 -953 -454 -935
rect -330 935 -296 953
rect -330 919 -296 935
rect -330 867 -296 881
rect -330 847 -296 867
rect -330 799 -296 809
rect -330 775 -296 799
rect -330 731 -296 737
rect -330 703 -296 731
rect -330 663 -296 665
rect -330 631 -296 663
rect -330 561 -296 593
rect -330 559 -296 561
rect -330 493 -296 521
rect -330 487 -296 493
rect -330 425 -296 449
rect -330 415 -296 425
rect -330 357 -296 377
rect -330 343 -296 357
rect -330 289 -296 305
rect -330 271 -296 289
rect -330 221 -296 233
rect -330 199 -296 221
rect -330 153 -296 161
rect -330 127 -296 153
rect -330 85 -296 89
rect -330 55 -296 85
rect -330 -17 -296 17
rect -330 -85 -296 -55
rect -330 -89 -296 -85
rect -330 -153 -296 -127
rect -330 -161 -296 -153
rect -330 -221 -296 -199
rect -330 -233 -296 -221
rect -330 -289 -296 -271
rect -330 -305 -296 -289
rect -330 -357 -296 -343
rect -330 -377 -296 -357
rect -330 -425 -296 -415
rect -330 -449 -296 -425
rect -330 -493 -296 -487
rect -330 -521 -296 -493
rect -330 -561 -296 -559
rect -330 -593 -296 -561
rect -330 -663 -296 -631
rect -330 -665 -296 -663
rect -330 -731 -296 -703
rect -330 -737 -296 -731
rect -330 -799 -296 -775
rect -330 -809 -296 -799
rect -330 -867 -296 -847
rect -330 -881 -296 -867
rect -330 -935 -296 -919
rect -330 -953 -296 -935
rect -172 935 -138 953
rect -172 919 -138 935
rect -172 867 -138 881
rect -172 847 -138 867
rect -172 799 -138 809
rect -172 775 -138 799
rect -172 731 -138 737
rect -172 703 -138 731
rect -172 663 -138 665
rect -172 631 -138 663
rect -172 561 -138 593
rect -172 559 -138 561
rect -172 493 -138 521
rect -172 487 -138 493
rect -172 425 -138 449
rect -172 415 -138 425
rect -172 357 -138 377
rect -172 343 -138 357
rect -172 289 -138 305
rect -172 271 -138 289
rect -172 221 -138 233
rect -172 199 -138 221
rect -172 153 -138 161
rect -172 127 -138 153
rect -172 85 -138 89
rect -172 55 -138 85
rect -172 -17 -138 17
rect -172 -85 -138 -55
rect -172 -89 -138 -85
rect -172 -153 -138 -127
rect -172 -161 -138 -153
rect -172 -221 -138 -199
rect -172 -233 -138 -221
rect -172 -289 -138 -271
rect -172 -305 -138 -289
rect -172 -357 -138 -343
rect -172 -377 -138 -357
rect -172 -425 -138 -415
rect -172 -449 -138 -425
rect -172 -493 -138 -487
rect -172 -521 -138 -493
rect -172 -561 -138 -559
rect -172 -593 -138 -561
rect -172 -663 -138 -631
rect -172 -665 -138 -663
rect -172 -731 -138 -703
rect -172 -737 -138 -731
rect -172 -799 -138 -775
rect -172 -809 -138 -799
rect -172 -867 -138 -847
rect -172 -881 -138 -867
rect -172 -935 -138 -919
rect -172 -953 -138 -935
rect -14 935 20 953
rect -14 919 20 935
rect -14 867 20 881
rect -14 847 20 867
rect -14 799 20 809
rect -14 775 20 799
rect -14 731 20 737
rect -14 703 20 731
rect -14 663 20 665
rect -14 631 20 663
rect -14 561 20 593
rect -14 559 20 561
rect -14 493 20 521
rect -14 487 20 493
rect -14 425 20 449
rect -14 415 20 425
rect -14 357 20 377
rect -14 343 20 357
rect -14 289 20 305
rect -14 271 20 289
rect -14 221 20 233
rect -14 199 20 221
rect -14 153 20 161
rect -14 127 20 153
rect -14 85 20 89
rect -14 55 20 85
rect -14 -17 20 17
rect -14 -85 20 -55
rect -14 -89 20 -85
rect -14 -153 20 -127
rect -14 -161 20 -153
rect -14 -221 20 -199
rect -14 -233 20 -221
rect -14 -289 20 -271
rect -14 -305 20 -289
rect -14 -357 20 -343
rect -14 -377 20 -357
rect -14 -425 20 -415
rect -14 -449 20 -425
rect -14 -493 20 -487
rect -14 -521 20 -493
rect -14 -561 20 -559
rect -14 -593 20 -561
rect -14 -663 20 -631
rect -14 -665 20 -663
rect -14 -731 20 -703
rect -14 -737 20 -731
rect -14 -799 20 -775
rect -14 -809 20 -799
rect -14 -867 20 -847
rect -14 -881 20 -867
rect -14 -935 20 -919
rect -14 -953 20 -935
rect 144 935 178 953
rect 144 919 178 935
rect 144 867 178 881
rect 144 847 178 867
rect 144 799 178 809
rect 144 775 178 799
rect 144 731 178 737
rect 144 703 178 731
rect 144 663 178 665
rect 144 631 178 663
rect 144 561 178 593
rect 144 559 178 561
rect 144 493 178 521
rect 144 487 178 493
rect 144 425 178 449
rect 144 415 178 425
rect 144 357 178 377
rect 144 343 178 357
rect 144 289 178 305
rect 144 271 178 289
rect 144 221 178 233
rect 144 199 178 221
rect 144 153 178 161
rect 144 127 178 153
rect 144 85 178 89
rect 144 55 178 85
rect 144 -17 178 17
rect 144 -85 178 -55
rect 144 -89 178 -85
rect 144 -153 178 -127
rect 144 -161 178 -153
rect 144 -221 178 -199
rect 144 -233 178 -221
rect 144 -289 178 -271
rect 144 -305 178 -289
rect 144 -357 178 -343
rect 144 -377 178 -357
rect 144 -425 178 -415
rect 144 -449 178 -425
rect 144 -493 178 -487
rect 144 -521 178 -493
rect 144 -561 178 -559
rect 144 -593 178 -561
rect 144 -663 178 -631
rect 144 -665 178 -663
rect 144 -731 178 -703
rect 144 -737 178 -731
rect 144 -799 178 -775
rect 144 -809 178 -799
rect 144 -867 178 -847
rect 144 -881 178 -867
rect 144 -935 178 -919
rect 144 -953 178 -935
rect 302 935 336 953
rect 302 919 336 935
rect 302 867 336 881
rect 302 847 336 867
rect 302 799 336 809
rect 302 775 336 799
rect 302 731 336 737
rect 302 703 336 731
rect 302 663 336 665
rect 302 631 336 663
rect 302 561 336 593
rect 302 559 336 561
rect 302 493 336 521
rect 302 487 336 493
rect 302 425 336 449
rect 302 415 336 425
rect 302 357 336 377
rect 302 343 336 357
rect 302 289 336 305
rect 302 271 336 289
rect 302 221 336 233
rect 302 199 336 221
rect 302 153 336 161
rect 302 127 336 153
rect 302 85 336 89
rect 302 55 336 85
rect 302 -17 336 17
rect 302 -85 336 -55
rect 302 -89 336 -85
rect 302 -153 336 -127
rect 302 -161 336 -153
rect 302 -221 336 -199
rect 302 -233 336 -221
rect 302 -289 336 -271
rect 302 -305 336 -289
rect 302 -357 336 -343
rect 302 -377 336 -357
rect 302 -425 336 -415
rect 302 -449 336 -425
rect 302 -493 336 -487
rect 302 -521 336 -493
rect 302 -561 336 -559
rect 302 -593 336 -561
rect 302 -663 336 -631
rect 302 -665 336 -663
rect 302 -731 336 -703
rect 302 -737 336 -731
rect 302 -799 336 -775
rect 302 -809 336 -799
rect 302 -867 336 -847
rect 302 -881 336 -867
rect 302 -935 336 -919
rect 302 -953 336 -935
rect 460 935 494 953
rect 460 919 494 935
rect 460 867 494 881
rect 460 847 494 867
rect 460 799 494 809
rect 460 775 494 799
rect 460 731 494 737
rect 460 703 494 731
rect 460 663 494 665
rect 460 631 494 663
rect 460 561 494 593
rect 460 559 494 561
rect 460 493 494 521
rect 460 487 494 493
rect 460 425 494 449
rect 460 415 494 425
rect 460 357 494 377
rect 460 343 494 357
rect 460 289 494 305
rect 460 271 494 289
rect 460 221 494 233
rect 460 199 494 221
rect 460 153 494 161
rect 460 127 494 153
rect 460 85 494 89
rect 460 55 494 85
rect 460 -17 494 17
rect 460 -85 494 -55
rect 460 -89 494 -85
rect 460 -153 494 -127
rect 460 -161 494 -153
rect 460 -221 494 -199
rect 460 -233 494 -221
rect 460 -289 494 -271
rect 460 -305 494 -289
rect 460 -357 494 -343
rect 460 -377 494 -357
rect 460 -425 494 -415
rect 460 -449 494 -425
rect 460 -493 494 -487
rect 460 -521 494 -493
rect 460 -561 494 -559
rect 460 -593 494 -561
rect 460 -663 494 -631
rect 460 -665 494 -663
rect 460 -731 494 -703
rect 460 -737 494 -731
rect 460 -799 494 -775
rect 460 -809 494 -799
rect 460 -867 494 -847
rect 460 -881 494 -867
rect 460 -935 494 -919
rect 460 -953 494 -935
rect 618 935 652 953
rect 618 919 652 935
rect 618 867 652 881
rect 618 847 652 867
rect 618 799 652 809
rect 618 775 652 799
rect 618 731 652 737
rect 618 703 652 731
rect 618 663 652 665
rect 618 631 652 663
rect 618 561 652 593
rect 618 559 652 561
rect 618 493 652 521
rect 618 487 652 493
rect 618 425 652 449
rect 618 415 652 425
rect 618 357 652 377
rect 618 343 652 357
rect 618 289 652 305
rect 618 271 652 289
rect 618 221 652 233
rect 618 199 652 221
rect 618 153 652 161
rect 618 127 652 153
rect 618 85 652 89
rect 618 55 652 85
rect 618 -17 652 17
rect 618 -85 652 -55
rect 618 -89 652 -85
rect 618 -153 652 -127
rect 618 -161 652 -153
rect 618 -221 652 -199
rect 618 -233 652 -221
rect 618 -289 652 -271
rect 618 -305 652 -289
rect 618 -357 652 -343
rect 618 -377 652 -357
rect 618 -425 652 -415
rect 618 -449 652 -425
rect 618 -493 652 -487
rect 618 -521 652 -493
rect 618 -561 652 -559
rect 618 -593 652 -561
rect 618 -663 652 -631
rect 618 -665 652 -663
rect 618 -731 652 -703
rect 618 -737 652 -731
rect 618 -799 652 -775
rect 618 -809 652 -799
rect 618 -867 652 -847
rect 618 -881 652 -867
rect 618 -935 652 -919
rect 618 -953 652 -935
rect 776 935 810 953
rect 776 919 810 935
rect 776 867 810 881
rect 776 847 810 867
rect 776 799 810 809
rect 776 775 810 799
rect 776 731 810 737
rect 776 703 810 731
rect 776 663 810 665
rect 776 631 810 663
rect 776 561 810 593
rect 776 559 810 561
rect 776 493 810 521
rect 776 487 810 493
rect 776 425 810 449
rect 776 415 810 425
rect 776 357 810 377
rect 776 343 810 357
rect 776 289 810 305
rect 776 271 810 289
rect 776 221 810 233
rect 776 199 810 221
rect 776 153 810 161
rect 776 127 810 153
rect 776 85 810 89
rect 776 55 810 85
rect 776 -17 810 17
rect 776 -85 810 -55
rect 776 -89 810 -85
rect 776 -153 810 -127
rect 776 -161 810 -153
rect 776 -221 810 -199
rect 776 -233 810 -221
rect 776 -289 810 -271
rect 776 -305 810 -289
rect 776 -357 810 -343
rect 776 -377 810 -357
rect 776 -425 810 -415
rect 776 -449 810 -425
rect 776 -493 810 -487
rect 776 -521 810 -493
rect 776 -561 810 -559
rect 776 -593 810 -561
rect 776 -663 810 -631
rect 776 -665 810 -663
rect 776 -731 810 -703
rect 776 -737 810 -731
rect 776 -799 810 -775
rect 776 -809 810 -799
rect 776 -867 810 -847
rect 776 -881 810 -867
rect 776 -935 810 -919
rect 776 -953 810 -935
<< metal1 >>
rect -26 1152 32 1174
rect -810 1106 816 1152
rect -810 953 -764 1106
rect -810 919 -804 953
rect -770 919 -764 953
rect -810 881 -764 919
rect -810 847 -804 881
rect -770 847 -764 881
rect -810 809 -764 847
rect -810 775 -804 809
rect -770 775 -764 809
rect -810 737 -764 775
rect -810 703 -804 737
rect -770 703 -764 737
rect -810 665 -764 703
rect -810 631 -804 665
rect -770 631 -764 665
rect -810 593 -764 631
rect -810 559 -804 593
rect -770 559 -764 593
rect -810 521 -764 559
rect -810 487 -804 521
rect -770 487 -764 521
rect -810 449 -764 487
rect -810 415 -804 449
rect -770 415 -764 449
rect -810 377 -764 415
rect -810 343 -804 377
rect -770 343 -764 377
rect -810 305 -764 343
rect -810 271 -804 305
rect -770 271 -764 305
rect -810 233 -764 271
rect -810 199 -804 233
rect -770 199 -764 233
rect -810 161 -764 199
rect -810 127 -804 161
rect -770 127 -764 161
rect -810 89 -764 127
rect -810 55 -804 89
rect -770 55 -764 89
rect -810 17 -764 55
rect -810 -17 -804 17
rect -770 -17 -764 17
rect -810 -55 -764 -17
rect -810 -89 -804 -55
rect -770 -89 -764 -55
rect -810 -127 -764 -89
rect -810 -161 -804 -127
rect -770 -161 -764 -127
rect -810 -199 -764 -161
rect -810 -233 -804 -199
rect -770 -233 -764 -199
rect -810 -271 -764 -233
rect -810 -305 -804 -271
rect -770 -305 -764 -271
rect -810 -343 -764 -305
rect -810 -377 -804 -343
rect -770 -377 -764 -343
rect -810 -415 -764 -377
rect -810 -449 -804 -415
rect -770 -449 -764 -415
rect -810 -487 -764 -449
rect -810 -521 -804 -487
rect -770 -521 -764 -487
rect -810 -559 -764 -521
rect -810 -593 -804 -559
rect -770 -593 -764 -559
rect -810 -631 -764 -593
rect -810 -665 -804 -631
rect -770 -665 -764 -631
rect -810 -703 -764 -665
rect -810 -737 -804 -703
rect -770 -737 -764 -703
rect -810 -775 -764 -737
rect -810 -809 -804 -775
rect -770 -809 -764 -775
rect -810 -847 -764 -809
rect -810 -881 -804 -847
rect -770 -881 -764 -847
rect -810 -919 -764 -881
rect -810 -953 -804 -919
rect -770 -953 -764 -919
rect -810 -1000 -764 -953
rect -652 953 -606 1000
rect -652 919 -646 953
rect -612 919 -606 953
rect -652 881 -606 919
rect -652 847 -646 881
rect -612 847 -606 881
rect -652 809 -606 847
rect -652 775 -646 809
rect -612 775 -606 809
rect -652 737 -606 775
rect -652 703 -646 737
rect -612 703 -606 737
rect -652 665 -606 703
rect -652 631 -646 665
rect -612 631 -606 665
rect -652 593 -606 631
rect -652 559 -646 593
rect -612 559 -606 593
rect -652 521 -606 559
rect -652 487 -646 521
rect -612 487 -606 521
rect -652 449 -606 487
rect -652 415 -646 449
rect -612 415 -606 449
rect -652 377 -606 415
rect -652 343 -646 377
rect -612 343 -606 377
rect -652 305 -606 343
rect -652 271 -646 305
rect -612 271 -606 305
rect -652 233 -606 271
rect -652 199 -646 233
rect -612 199 -606 233
rect -652 161 -606 199
rect -652 127 -646 161
rect -612 127 -606 161
rect -652 89 -606 127
rect -652 55 -646 89
rect -612 55 -606 89
rect -652 17 -606 55
rect -652 -17 -646 17
rect -612 -17 -606 17
rect -652 -55 -606 -17
rect -652 -89 -646 -55
rect -612 -89 -606 -55
rect -652 -127 -606 -89
rect -652 -161 -646 -127
rect -612 -161 -606 -127
rect -652 -199 -606 -161
rect -652 -233 -646 -199
rect -612 -233 -606 -199
rect -652 -271 -606 -233
rect -652 -305 -646 -271
rect -612 -305 -606 -271
rect -652 -343 -606 -305
rect -652 -377 -646 -343
rect -612 -377 -606 -343
rect -652 -415 -606 -377
rect -652 -449 -646 -415
rect -612 -449 -606 -415
rect -652 -487 -606 -449
rect -652 -521 -646 -487
rect -612 -521 -606 -487
rect -652 -559 -606 -521
rect -652 -593 -646 -559
rect -612 -593 -606 -559
rect -652 -631 -606 -593
rect -652 -665 -646 -631
rect -612 -665 -606 -631
rect -652 -703 -606 -665
rect -652 -737 -646 -703
rect -612 -737 -606 -703
rect -652 -775 -606 -737
rect -652 -809 -646 -775
rect -612 -809 -606 -775
rect -652 -847 -606 -809
rect -652 -881 -646 -847
rect -612 -881 -606 -847
rect -652 -919 -606 -881
rect -652 -953 -646 -919
rect -612 -953 -606 -919
rect -652 -1118 -606 -953
rect -494 953 -448 1106
rect -494 919 -488 953
rect -454 919 -448 953
rect -494 881 -448 919
rect -494 847 -488 881
rect -454 847 -448 881
rect -494 809 -448 847
rect -494 775 -488 809
rect -454 775 -448 809
rect -494 737 -448 775
rect -494 703 -488 737
rect -454 703 -448 737
rect -494 665 -448 703
rect -494 631 -488 665
rect -454 631 -448 665
rect -494 593 -448 631
rect -494 559 -488 593
rect -454 559 -448 593
rect -494 521 -448 559
rect -494 487 -488 521
rect -454 487 -448 521
rect -494 449 -448 487
rect -494 415 -488 449
rect -454 415 -448 449
rect -494 377 -448 415
rect -494 343 -488 377
rect -454 343 -448 377
rect -494 305 -448 343
rect -494 271 -488 305
rect -454 271 -448 305
rect -494 233 -448 271
rect -494 199 -488 233
rect -454 199 -448 233
rect -494 161 -448 199
rect -494 127 -488 161
rect -454 127 -448 161
rect -494 89 -448 127
rect -494 55 -488 89
rect -454 55 -448 89
rect -494 17 -448 55
rect -494 -17 -488 17
rect -454 -17 -448 17
rect -494 -55 -448 -17
rect -494 -89 -488 -55
rect -454 -89 -448 -55
rect -494 -127 -448 -89
rect -494 -161 -488 -127
rect -454 -161 -448 -127
rect -494 -199 -448 -161
rect -494 -233 -488 -199
rect -454 -233 -448 -199
rect -494 -271 -448 -233
rect -494 -305 -488 -271
rect -454 -305 -448 -271
rect -494 -343 -448 -305
rect -494 -377 -488 -343
rect -454 -377 -448 -343
rect -494 -415 -448 -377
rect -494 -449 -488 -415
rect -454 -449 -448 -415
rect -494 -487 -448 -449
rect -494 -521 -488 -487
rect -454 -521 -448 -487
rect -494 -559 -448 -521
rect -494 -593 -488 -559
rect -454 -593 -448 -559
rect -494 -631 -448 -593
rect -494 -665 -488 -631
rect -454 -665 -448 -631
rect -494 -703 -448 -665
rect -494 -737 -488 -703
rect -454 -737 -448 -703
rect -494 -775 -448 -737
rect -494 -809 -488 -775
rect -454 -809 -448 -775
rect -494 -847 -448 -809
rect -494 -881 -488 -847
rect -454 -881 -448 -847
rect -494 -919 -448 -881
rect -494 -953 -488 -919
rect -454 -953 -448 -919
rect -494 -1000 -448 -953
rect -336 953 -290 1000
rect -336 919 -330 953
rect -296 919 -290 953
rect -336 881 -290 919
rect -336 847 -330 881
rect -296 847 -290 881
rect -336 809 -290 847
rect -336 775 -330 809
rect -296 775 -290 809
rect -336 737 -290 775
rect -336 703 -330 737
rect -296 703 -290 737
rect -336 665 -290 703
rect -336 631 -330 665
rect -296 631 -290 665
rect -336 593 -290 631
rect -336 559 -330 593
rect -296 559 -290 593
rect -336 521 -290 559
rect -336 487 -330 521
rect -296 487 -290 521
rect -336 449 -290 487
rect -336 415 -330 449
rect -296 415 -290 449
rect -336 377 -290 415
rect -336 343 -330 377
rect -296 343 -290 377
rect -336 305 -290 343
rect -336 271 -330 305
rect -296 271 -290 305
rect -336 233 -290 271
rect -336 199 -330 233
rect -296 199 -290 233
rect -336 161 -290 199
rect -336 127 -330 161
rect -296 127 -290 161
rect -336 89 -290 127
rect -336 55 -330 89
rect -296 55 -290 89
rect -336 17 -290 55
rect -336 -17 -330 17
rect -296 -17 -290 17
rect -336 -55 -290 -17
rect -336 -89 -330 -55
rect -296 -89 -290 -55
rect -336 -127 -290 -89
rect -336 -161 -330 -127
rect -296 -161 -290 -127
rect -336 -199 -290 -161
rect -336 -233 -330 -199
rect -296 -233 -290 -199
rect -336 -271 -290 -233
rect -336 -305 -330 -271
rect -296 -305 -290 -271
rect -336 -343 -290 -305
rect -336 -377 -330 -343
rect -296 -377 -290 -343
rect -336 -415 -290 -377
rect -336 -449 -330 -415
rect -296 -449 -290 -415
rect -336 -487 -290 -449
rect -336 -521 -330 -487
rect -296 -521 -290 -487
rect -336 -559 -290 -521
rect -336 -593 -330 -559
rect -296 -593 -290 -559
rect -336 -631 -290 -593
rect -336 -665 -330 -631
rect -296 -665 -290 -631
rect -336 -703 -290 -665
rect -336 -737 -330 -703
rect -296 -737 -290 -703
rect -336 -775 -290 -737
rect -336 -809 -330 -775
rect -296 -809 -290 -775
rect -336 -847 -290 -809
rect -336 -881 -330 -847
rect -296 -881 -290 -847
rect -336 -919 -290 -881
rect -336 -953 -330 -919
rect -296 -953 -290 -919
rect -336 -1118 -290 -953
rect -178 953 -132 1106
rect -178 919 -172 953
rect -138 919 -132 953
rect -178 881 -132 919
rect -178 847 -172 881
rect -138 847 -132 881
rect -178 809 -132 847
rect -178 775 -172 809
rect -138 775 -132 809
rect -178 737 -132 775
rect -178 703 -172 737
rect -138 703 -132 737
rect -178 665 -132 703
rect -178 631 -172 665
rect -138 631 -132 665
rect -178 593 -132 631
rect -178 559 -172 593
rect -138 559 -132 593
rect -178 521 -132 559
rect -178 487 -172 521
rect -138 487 -132 521
rect -178 449 -132 487
rect -178 415 -172 449
rect -138 415 -132 449
rect -178 377 -132 415
rect -178 343 -172 377
rect -138 343 -132 377
rect -178 305 -132 343
rect -178 271 -172 305
rect -138 271 -132 305
rect -178 233 -132 271
rect -178 199 -172 233
rect -138 199 -132 233
rect -178 161 -132 199
rect -178 127 -172 161
rect -138 127 -132 161
rect -178 89 -132 127
rect -178 55 -172 89
rect -138 55 -132 89
rect -178 17 -132 55
rect -178 -17 -172 17
rect -138 -17 -132 17
rect -178 -55 -132 -17
rect -178 -89 -172 -55
rect -138 -89 -132 -55
rect -178 -127 -132 -89
rect -178 -161 -172 -127
rect -138 -161 -132 -127
rect -178 -199 -132 -161
rect -178 -233 -172 -199
rect -138 -233 -132 -199
rect -178 -271 -132 -233
rect -178 -305 -172 -271
rect -138 -305 -132 -271
rect -178 -343 -132 -305
rect -178 -377 -172 -343
rect -138 -377 -132 -343
rect -178 -415 -132 -377
rect -178 -449 -172 -415
rect -138 -449 -132 -415
rect -178 -487 -132 -449
rect -178 -521 -172 -487
rect -138 -521 -132 -487
rect -178 -559 -132 -521
rect -178 -593 -172 -559
rect -138 -593 -132 -559
rect -178 -631 -132 -593
rect -178 -665 -172 -631
rect -138 -665 -132 -631
rect -178 -703 -132 -665
rect -178 -737 -172 -703
rect -138 -737 -132 -703
rect -178 -775 -132 -737
rect -178 -809 -172 -775
rect -138 -809 -132 -775
rect -178 -847 -132 -809
rect -178 -881 -172 -847
rect -138 -881 -132 -847
rect -178 -919 -132 -881
rect -178 -953 -172 -919
rect -138 -953 -132 -919
rect -178 -1000 -132 -953
rect -20 953 26 1000
rect -20 919 -14 953
rect 20 919 26 953
rect -20 881 26 919
rect -20 847 -14 881
rect 20 847 26 881
rect -20 809 26 847
rect -20 775 -14 809
rect 20 775 26 809
rect -20 737 26 775
rect -20 703 -14 737
rect 20 703 26 737
rect -20 665 26 703
rect -20 631 -14 665
rect 20 631 26 665
rect -20 593 26 631
rect -20 559 -14 593
rect 20 559 26 593
rect -20 521 26 559
rect -20 487 -14 521
rect 20 487 26 521
rect -20 449 26 487
rect -20 415 -14 449
rect 20 415 26 449
rect -20 377 26 415
rect -20 343 -14 377
rect 20 343 26 377
rect -20 305 26 343
rect -20 271 -14 305
rect 20 271 26 305
rect -20 233 26 271
rect -20 199 -14 233
rect 20 199 26 233
rect -20 161 26 199
rect -20 127 -14 161
rect 20 127 26 161
rect -20 89 26 127
rect -20 55 -14 89
rect 20 55 26 89
rect -20 17 26 55
rect -20 -17 -14 17
rect 20 -17 26 17
rect -20 -55 26 -17
rect -20 -89 -14 -55
rect 20 -89 26 -55
rect -20 -127 26 -89
rect -20 -161 -14 -127
rect 20 -161 26 -127
rect -20 -199 26 -161
rect -20 -233 -14 -199
rect 20 -233 26 -199
rect -20 -271 26 -233
rect -20 -305 -14 -271
rect 20 -305 26 -271
rect -20 -343 26 -305
rect -20 -377 -14 -343
rect 20 -377 26 -343
rect -20 -415 26 -377
rect -20 -449 -14 -415
rect 20 -449 26 -415
rect -20 -487 26 -449
rect -20 -521 -14 -487
rect 20 -521 26 -487
rect -20 -559 26 -521
rect -20 -593 -14 -559
rect 20 -593 26 -559
rect -20 -631 26 -593
rect -20 -665 -14 -631
rect 20 -665 26 -631
rect -20 -703 26 -665
rect -20 -737 -14 -703
rect 20 -737 26 -703
rect -20 -775 26 -737
rect -20 -809 -14 -775
rect 20 -809 26 -775
rect -20 -847 26 -809
rect -20 -881 -14 -847
rect 20 -881 26 -847
rect -20 -919 26 -881
rect -20 -953 -14 -919
rect 20 -953 26 -919
rect -20 -1118 26 -953
rect 138 953 184 1106
rect 138 919 144 953
rect 178 919 184 953
rect 138 881 184 919
rect 138 847 144 881
rect 178 847 184 881
rect 138 809 184 847
rect 138 775 144 809
rect 178 775 184 809
rect 138 737 184 775
rect 138 703 144 737
rect 178 703 184 737
rect 138 665 184 703
rect 138 631 144 665
rect 178 631 184 665
rect 138 593 184 631
rect 138 559 144 593
rect 178 559 184 593
rect 138 521 184 559
rect 138 487 144 521
rect 178 487 184 521
rect 138 449 184 487
rect 138 415 144 449
rect 178 415 184 449
rect 138 377 184 415
rect 138 343 144 377
rect 178 343 184 377
rect 138 305 184 343
rect 138 271 144 305
rect 178 271 184 305
rect 138 233 184 271
rect 138 199 144 233
rect 178 199 184 233
rect 138 161 184 199
rect 138 127 144 161
rect 178 127 184 161
rect 138 89 184 127
rect 138 55 144 89
rect 178 55 184 89
rect 138 17 184 55
rect 138 -17 144 17
rect 178 -17 184 17
rect 138 -55 184 -17
rect 138 -89 144 -55
rect 178 -89 184 -55
rect 138 -127 184 -89
rect 138 -161 144 -127
rect 178 -161 184 -127
rect 138 -199 184 -161
rect 138 -233 144 -199
rect 178 -233 184 -199
rect 138 -271 184 -233
rect 138 -305 144 -271
rect 178 -305 184 -271
rect 138 -343 184 -305
rect 138 -377 144 -343
rect 178 -377 184 -343
rect 138 -415 184 -377
rect 138 -449 144 -415
rect 178 -449 184 -415
rect 138 -487 184 -449
rect 138 -521 144 -487
rect 178 -521 184 -487
rect 138 -559 184 -521
rect 138 -593 144 -559
rect 178 -593 184 -559
rect 138 -631 184 -593
rect 138 -665 144 -631
rect 178 -665 184 -631
rect 138 -703 184 -665
rect 138 -737 144 -703
rect 178 -737 184 -703
rect 138 -775 184 -737
rect 138 -809 144 -775
rect 178 -809 184 -775
rect 138 -847 184 -809
rect 138 -881 144 -847
rect 178 -881 184 -847
rect 138 -919 184 -881
rect 138 -953 144 -919
rect 178 -953 184 -919
rect 138 -1000 184 -953
rect 296 953 342 1000
rect 296 919 302 953
rect 336 919 342 953
rect 296 881 342 919
rect 296 847 302 881
rect 336 847 342 881
rect 296 809 342 847
rect 296 775 302 809
rect 336 775 342 809
rect 296 737 342 775
rect 296 703 302 737
rect 336 703 342 737
rect 296 665 342 703
rect 296 631 302 665
rect 336 631 342 665
rect 296 593 342 631
rect 296 559 302 593
rect 336 559 342 593
rect 296 521 342 559
rect 296 487 302 521
rect 336 487 342 521
rect 296 449 342 487
rect 296 415 302 449
rect 336 415 342 449
rect 296 377 342 415
rect 296 343 302 377
rect 336 343 342 377
rect 296 305 342 343
rect 296 271 302 305
rect 336 271 342 305
rect 296 233 342 271
rect 296 199 302 233
rect 336 199 342 233
rect 296 161 342 199
rect 296 127 302 161
rect 336 127 342 161
rect 296 89 342 127
rect 296 55 302 89
rect 336 55 342 89
rect 296 17 342 55
rect 296 -17 302 17
rect 336 -17 342 17
rect 296 -55 342 -17
rect 296 -89 302 -55
rect 336 -89 342 -55
rect 296 -127 342 -89
rect 296 -161 302 -127
rect 336 -161 342 -127
rect 296 -199 342 -161
rect 296 -233 302 -199
rect 336 -233 342 -199
rect 296 -271 342 -233
rect 296 -305 302 -271
rect 336 -305 342 -271
rect 296 -343 342 -305
rect 296 -377 302 -343
rect 336 -377 342 -343
rect 296 -415 342 -377
rect 296 -449 302 -415
rect 336 -449 342 -415
rect 296 -487 342 -449
rect 296 -521 302 -487
rect 336 -521 342 -487
rect 296 -559 342 -521
rect 296 -593 302 -559
rect 336 -593 342 -559
rect 296 -631 342 -593
rect 296 -665 302 -631
rect 336 -665 342 -631
rect 296 -703 342 -665
rect 296 -737 302 -703
rect 336 -737 342 -703
rect 296 -775 342 -737
rect 296 -809 302 -775
rect 336 -809 342 -775
rect 296 -847 342 -809
rect 296 -881 302 -847
rect 336 -881 342 -847
rect 296 -919 342 -881
rect 296 -953 302 -919
rect 336 -953 342 -919
rect 296 -1118 342 -953
rect 454 953 500 1106
rect 454 919 460 953
rect 494 919 500 953
rect 454 881 500 919
rect 454 847 460 881
rect 494 847 500 881
rect 454 809 500 847
rect 454 775 460 809
rect 494 775 500 809
rect 454 737 500 775
rect 454 703 460 737
rect 494 703 500 737
rect 454 665 500 703
rect 454 631 460 665
rect 494 631 500 665
rect 454 593 500 631
rect 454 559 460 593
rect 494 559 500 593
rect 454 521 500 559
rect 454 487 460 521
rect 494 487 500 521
rect 454 449 500 487
rect 454 415 460 449
rect 494 415 500 449
rect 454 377 500 415
rect 454 343 460 377
rect 494 343 500 377
rect 454 305 500 343
rect 454 271 460 305
rect 494 271 500 305
rect 454 233 500 271
rect 454 199 460 233
rect 494 199 500 233
rect 454 161 500 199
rect 454 127 460 161
rect 494 127 500 161
rect 454 89 500 127
rect 454 55 460 89
rect 494 55 500 89
rect 454 17 500 55
rect 454 -17 460 17
rect 494 -17 500 17
rect 454 -55 500 -17
rect 454 -89 460 -55
rect 494 -89 500 -55
rect 454 -127 500 -89
rect 454 -161 460 -127
rect 494 -161 500 -127
rect 454 -199 500 -161
rect 454 -233 460 -199
rect 494 -233 500 -199
rect 454 -271 500 -233
rect 454 -305 460 -271
rect 494 -305 500 -271
rect 454 -343 500 -305
rect 454 -377 460 -343
rect 494 -377 500 -343
rect 454 -415 500 -377
rect 454 -449 460 -415
rect 494 -449 500 -415
rect 454 -487 500 -449
rect 454 -521 460 -487
rect 494 -521 500 -487
rect 454 -559 500 -521
rect 454 -593 460 -559
rect 494 -593 500 -559
rect 454 -631 500 -593
rect 454 -665 460 -631
rect 494 -665 500 -631
rect 454 -703 500 -665
rect 454 -737 460 -703
rect 494 -737 500 -703
rect 454 -775 500 -737
rect 454 -809 460 -775
rect 494 -809 500 -775
rect 454 -847 500 -809
rect 454 -881 460 -847
rect 494 -881 500 -847
rect 454 -919 500 -881
rect 454 -953 460 -919
rect 494 -953 500 -919
rect 454 -1000 500 -953
rect 612 953 658 1000
rect 612 919 618 953
rect 652 919 658 953
rect 612 881 658 919
rect 612 847 618 881
rect 652 847 658 881
rect 612 809 658 847
rect 612 775 618 809
rect 652 775 658 809
rect 612 737 658 775
rect 612 703 618 737
rect 652 703 658 737
rect 612 665 658 703
rect 612 631 618 665
rect 652 631 658 665
rect 612 593 658 631
rect 612 559 618 593
rect 652 559 658 593
rect 612 521 658 559
rect 612 487 618 521
rect 652 487 658 521
rect 612 449 658 487
rect 612 415 618 449
rect 652 415 658 449
rect 612 377 658 415
rect 612 343 618 377
rect 652 343 658 377
rect 612 305 658 343
rect 612 271 618 305
rect 652 271 658 305
rect 612 233 658 271
rect 612 199 618 233
rect 652 199 658 233
rect 612 161 658 199
rect 612 127 618 161
rect 652 127 658 161
rect 612 89 658 127
rect 612 55 618 89
rect 652 55 658 89
rect 612 17 658 55
rect 612 -17 618 17
rect 652 -17 658 17
rect 612 -55 658 -17
rect 612 -89 618 -55
rect 652 -89 658 -55
rect 612 -127 658 -89
rect 612 -161 618 -127
rect 652 -161 658 -127
rect 612 -199 658 -161
rect 612 -233 618 -199
rect 652 -233 658 -199
rect 612 -271 658 -233
rect 612 -305 618 -271
rect 652 -305 658 -271
rect 612 -343 658 -305
rect 612 -377 618 -343
rect 652 -377 658 -343
rect 612 -415 658 -377
rect 612 -449 618 -415
rect 652 -449 658 -415
rect 612 -487 658 -449
rect 612 -521 618 -487
rect 652 -521 658 -487
rect 612 -559 658 -521
rect 612 -593 618 -559
rect 652 -593 658 -559
rect 612 -631 658 -593
rect 612 -665 618 -631
rect 652 -665 658 -631
rect 612 -703 658 -665
rect 612 -737 618 -703
rect 652 -737 658 -703
rect 612 -775 658 -737
rect 612 -809 618 -775
rect 652 -809 658 -775
rect 612 -847 658 -809
rect 612 -881 618 -847
rect 652 -881 658 -847
rect 612 -919 658 -881
rect 612 -953 618 -919
rect 652 -953 658 -919
rect 612 -1118 658 -953
rect 770 953 816 1106
rect 770 919 776 953
rect 810 919 816 953
rect 770 881 816 919
rect 770 847 776 881
rect 810 847 816 881
rect 770 809 816 847
rect 770 775 776 809
rect 810 775 816 809
rect 770 737 816 775
rect 770 703 776 737
rect 810 703 816 737
rect 770 665 816 703
rect 770 631 776 665
rect 810 631 816 665
rect 770 593 816 631
rect 770 559 776 593
rect 810 559 816 593
rect 770 521 816 559
rect 770 487 776 521
rect 810 487 816 521
rect 770 449 816 487
rect 770 415 776 449
rect 810 415 816 449
rect 770 377 816 415
rect 770 343 776 377
rect 810 343 816 377
rect 770 305 816 343
rect 770 271 776 305
rect 810 271 816 305
rect 770 233 816 271
rect 770 199 776 233
rect 810 199 816 233
rect 770 161 816 199
rect 770 127 776 161
rect 810 127 816 161
rect 770 89 816 127
rect 770 55 776 89
rect 810 55 816 89
rect 770 17 816 55
rect 770 -17 776 17
rect 810 -17 816 17
rect 770 -55 816 -17
rect 770 -89 776 -55
rect 810 -89 816 -55
rect 770 -127 816 -89
rect 770 -161 776 -127
rect 810 -161 816 -127
rect 770 -199 816 -161
rect 770 -233 776 -199
rect 810 -233 816 -199
rect 770 -271 816 -233
rect 770 -305 776 -271
rect 810 -305 816 -271
rect 770 -343 816 -305
rect 770 -377 776 -343
rect 810 -377 816 -343
rect 770 -415 816 -377
rect 770 -449 776 -415
rect 810 -449 816 -415
rect 770 -487 816 -449
rect 770 -521 776 -487
rect 810 -521 816 -487
rect 770 -559 816 -521
rect 770 -593 776 -559
rect 810 -593 816 -559
rect 770 -631 816 -593
rect 770 -665 776 -631
rect 810 -665 816 -631
rect 770 -703 816 -665
rect 770 -737 776 -703
rect 810 -737 816 -703
rect 770 -775 816 -737
rect 770 -809 776 -775
rect 810 -809 816 -775
rect 770 -847 816 -809
rect 770 -881 776 -847
rect 810 -881 816 -847
rect 770 -919 816 -881
rect 770 -953 776 -919
rect 810 -953 816 -919
rect 770 -1000 816 -953
rect -652 -1164 658 -1118
rect -20 -1174 26 -1164
<< end >>
