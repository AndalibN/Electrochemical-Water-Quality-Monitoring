magic
tech sky130A
magscale 1 2
timestamp 1666815582
<< checkpaint >>
rect 7329 -1773 21875 1347
<< error_s >>
rect 3419 2739 3481 2745
rect 3419 2705 3431 2739
rect 3419 2699 3481 2705
rect 7918 2156 7980 2162
rect 7918 2122 7930 2156
rect 7918 2116 7980 2122
rect 338 2063 373 2097
rect 339 2044 373 2063
rect 147 1995 209 2001
rect 147 1961 159 1995
rect 147 1955 209 1961
rect 147 719 209 725
rect 147 685 159 719
rect 147 679 209 685
rect 358 583 373 2044
rect 392 2010 427 2044
rect 392 583 426 2010
rect 556 1942 618 1948
rect 556 1908 568 1942
rect 556 1902 618 1908
rect 1974 1869 2009 1903
rect 1975 1850 2009 1869
rect 1783 1801 1845 1807
rect 1783 1767 1795 1801
rect 1783 1761 1845 1767
rect 748 1213 782 1267
rect 556 666 618 672
rect 556 632 568 666
rect 556 626 618 632
rect 392 549 407 583
rect 767 530 782 1213
rect 801 1179 836 1213
rect 801 530 835 1179
rect 965 1111 1027 1117
rect 965 1077 977 1111
rect 965 1071 1027 1077
rect 1157 858 1191 912
rect 1619 894 1653 912
rect 965 613 1027 619
rect 965 579 977 613
rect 965 573 1027 579
rect 801 496 816 530
rect 1176 477 1191 858
rect 1210 824 1245 858
rect 1210 477 1244 824
rect 1374 756 1436 762
rect 1374 722 1386 756
rect 1374 716 1436 722
rect 1374 560 1436 566
rect 1374 526 1386 560
rect 1374 520 1436 526
rect 1210 443 1225 477
rect 1583 424 1653 894
rect 1783 507 1845 513
rect 1783 473 1795 507
rect 1783 467 1845 473
rect 1583 388 1636 424
rect 1994 371 2009 1850
rect 2028 1816 2063 1850
rect 2028 371 2062 1816
rect 2192 1748 2254 1754
rect 2192 1714 2204 1748
rect 2192 1708 2254 1714
rect 2384 1019 2418 1073
rect 2846 1055 2880 1073
rect 2192 454 2254 460
rect 2192 420 2204 454
rect 2192 414 2254 420
rect 2028 337 2043 371
rect 2403 318 2418 1019
rect 2437 985 2472 1019
rect 2437 318 2471 985
rect 2601 917 2663 923
rect 2601 883 2613 917
rect 2601 877 2663 883
rect 2601 401 2663 407
rect 2601 367 2613 401
rect 2601 361 2663 367
rect 2437 284 2452 318
rect 2810 265 2880 1055
rect 3010 1040 3072 1046
rect 3010 1006 3022 1040
rect 3010 1000 3072 1006
rect 3010 348 3072 354
rect 3010 314 3022 348
rect 3010 308 3072 314
rect 2810 229 2863 265
rect 3221 212 3236 1142
rect 3255 212 3289 1196
rect 4428 1163 4463 1197
rect 4429 1144 4463 1163
rect 4237 1095 4299 1101
rect 3611 1036 3645 1090
rect 4073 1072 4107 1090
rect 3419 295 3481 301
rect 3419 261 3431 295
rect 3419 255 3481 261
rect 3255 178 3270 212
rect 3630 159 3645 1036
rect 3664 1002 3699 1036
rect 3664 159 3698 1002
rect 3828 934 3890 940
rect 3828 900 3840 934
rect 3828 894 3890 900
rect 3828 242 3890 248
rect 3828 208 3840 242
rect 3828 202 3890 208
rect 3664 125 3679 159
rect 4037 106 4107 1072
rect 4237 1061 4249 1095
rect 4237 1055 4299 1061
rect 4237 189 4299 195
rect 4237 155 4249 189
rect 4237 149 4299 155
rect 4037 70 4090 106
rect 4448 53 4463 1144
rect 4482 1110 4517 1144
rect 4837 1110 4872 1144
rect 4482 53 4516 1110
rect 4838 1091 4872 1110
rect 4646 1042 4708 1048
rect 4646 1008 4658 1042
rect 4646 1002 4708 1008
rect 4646 136 4708 142
rect 4646 102 4658 136
rect 4646 96 4708 102
rect 4482 19 4497 53
rect 4857 0 4872 1091
rect 4891 1057 4926 1091
rect 5246 1057 5281 1091
rect 4891 0 4925 1057
rect 5247 1038 5281 1057
rect 5055 989 5117 995
rect 5055 955 5067 989
rect 5055 949 5117 955
rect 5055 83 5117 89
rect 5055 49 5067 83
rect 5055 43 5117 49
rect 4891 -34 4906 0
rect 5266 -53 5281 1038
rect 5300 1004 5335 1038
rect 5655 1004 5690 1038
rect 5300 -53 5334 1004
rect 5656 985 5690 1004
rect 5464 936 5526 942
rect 5464 902 5476 936
rect 5464 896 5526 902
rect 5464 30 5526 36
rect 5464 -4 5476 30
rect 5464 -10 5526 -4
rect 5300 -87 5315 -53
rect 5675 -106 5690 985
rect 5709 951 5744 985
rect 6064 951 6099 985
rect 5709 -106 5743 951
rect 6065 932 6099 951
rect 5873 883 5935 889
rect 5873 849 5885 883
rect 5873 843 5935 849
rect 5873 -23 5935 -17
rect 5873 -57 5885 -23
rect 5873 -63 5935 -57
rect 5709 -140 5724 -106
rect 6084 -159 6099 932
rect 6118 898 6153 932
rect 6473 898 6508 932
rect 6118 -159 6152 898
rect 6474 879 6508 898
rect 6282 830 6344 836
rect 6282 796 6294 830
rect 6282 790 6344 796
rect 6282 -76 6344 -70
rect 6282 -110 6294 -76
rect 6282 -116 6344 -110
rect 6118 -193 6133 -159
rect 6493 -212 6508 879
rect 6527 845 6562 879
rect 6882 845 6917 879
rect 6527 -212 6561 845
rect 6883 826 6917 845
rect 6691 777 6753 783
rect 6691 743 6703 777
rect 6691 737 6753 743
rect 6691 -129 6753 -123
rect 6691 -163 6703 -129
rect 6691 -169 6753 -163
rect 6527 -246 6542 -212
rect 6902 -265 6917 826
rect 6936 792 6971 826
rect 6936 -265 6970 792
rect 7100 724 7162 730
rect 7100 690 7112 724
rect 7100 684 7162 690
rect 7292 595 7326 613
rect 7292 559 7362 595
rect 7309 525 7380 559
rect 7100 -182 7162 -176
rect 7100 -216 7112 -182
rect 7100 -222 7162 -216
rect 6936 -299 6951 -265
rect 7309 -318 7379 525
rect 7509 457 7571 463
rect 7509 423 7521 457
rect 7509 417 7571 423
rect 7509 -235 7571 -229
rect 7509 -269 7521 -235
rect 7509 -275 7571 -269
rect 7309 -354 7362 -318
rect 7720 -371 7735 559
rect 7754 -371 7788 613
rect 8110 453 8144 507
rect 7918 -288 7980 -282
rect 7918 -322 7930 -288
rect 7918 -328 7980 -322
rect 7754 -405 7769 -371
rect 8129 -424 8144 453
rect 8163 419 8198 453
rect 8163 -424 8197 419
rect 8327 351 8389 357
rect 8327 317 8339 351
rect 8327 311 8389 317
rect 8327 -341 8389 -335
rect 8327 -375 8339 -341
rect 8327 -381 8389 -375
rect 8163 -458 8178 -424
use sky130_fd_pr__cap_mim_m3_1_MTBYP6  XC1
timestamp 0
transform 1 0 11596 0 1 -213
box -3007 -300 3006 300
use sky130_fd_pr__cap_mim_m3_1_MTBYP6  XC2
timestamp 0
transform 1 0 17609 0 1 -213
box -3007 -300 3006 300
use sky130_fd_pr__pfet_01v8_lvt_E7VWN7  XM1
timestamp 0
transform 1 0 1814 0 1 1137
box -231 -802 231 802
use sky130_fd_pr__pfet_01v8_lvt_E7VWN7  XM2
timestamp 0
transform 1 0 2223 0 1 1084
box -231 -802 231 802
use sky130_fd_pr__nfet_01v8_lvt_U66HNY  XM3
timestamp 0
transform 1 0 996 0 1 845
box -231 -404 231 404
use sky130_fd_pr__nfet_01v8_lvt_Y7U3JD  XM4
timestamp 0
transform 1 0 587 0 1 1287
box -231 -793 231 793
use sky130_fd_pr__pfet_01v8_lvt_4YYSM3  XM5
timestamp 0
transform 1 0 2632 0 1 642
box -231 -413 231 413
use sky130_fd_pr__nfet_01v8_lvt_Y7U3JD  XM6
timestamp 0
transform 1 0 178 0 1 1340
box -231 -793 231 793
use sky130_fd_pr__nfet_01v8_lvt_CN6LX3  XM7
timestamp 0
transform 1 0 1405 0 1 641
box -231 -253 231 253
use sky130_fd_pr__nfet_01v8_lvt_86CZ93  XM8
timestamp 0
transform 1 0 3041 0 1 677
box -231 -501 231 501
use sky130_fd_pr__nfet_01v8_lvt_KRU4ZZ  XM9
timestamp 0
transform 1 0 3450 0 1 1500
box -231 -1377 231 1377
use sky130_fd_pr__nfet_01v8_lvt_86CZ93  XM10
timestamp 0
transform 1 0 3859 0 1 571
box -231 -501 231 501
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM11
timestamp 0
transform 1 0 4268 0 1 625
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM12
timestamp 0
transform 1 0 4677 0 1 572
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM13
timestamp 0
transform 1 0 5495 0 1 466
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM14
timestamp 0
transform 1 0 5904 0 1 413
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM15
timestamp 0
transform 1 0 5086 0 1 519
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM16
timestamp 0
transform 1 0 6313 0 1 360
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM17
timestamp 0
transform 1 0 6722 0 1 307
box -231 -608 231 608
use sky130_fd_pr__pfet_01v8_lvt_4JSEF6  XM18
timestamp 0
transform 1 0 7131 0 1 254
box -231 -608 231 608
use sky130_fd_pr__nfet_01v8_lvt_86CZ93  XM19
timestamp 0
transform 1 0 7540 0 1 94
box -231 -501 231 501
use sky130_fd_pr__nfet_01v8_lvt_KRU4ZZ  XM20
timestamp 0
transform 1 0 7949 0 1 917
box -231 -1377 231 1377
use sky130_fd_pr__nfet_01v8_lvt_86CZ93  XM21
timestamp 0
transform 1 0 8358 0 1 -12
box -231 -501 231 501
<< end >>
