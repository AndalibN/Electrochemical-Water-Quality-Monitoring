magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -1084 -126 1084 126
<< nmos >>
rect -1000 -100 1000 100
<< ndiff >>
rect -1058 85 -1000 100
rect -1058 51 -1046 85
rect -1012 51 -1000 85
rect -1058 17 -1000 51
rect -1058 -17 -1046 17
rect -1012 -17 -1000 17
rect -1058 -51 -1000 -17
rect -1058 -85 -1046 -51
rect -1012 -85 -1000 -51
rect -1058 -100 -1000 -85
rect 1000 85 1058 100
rect 1000 51 1012 85
rect 1046 51 1058 85
rect 1000 17 1058 51
rect 1000 -17 1012 17
rect 1046 -17 1058 17
rect 1000 -51 1058 -17
rect 1000 -85 1012 -51
rect 1046 -85 1058 -51
rect 1000 -100 1058 -85
<< ndiffc >>
rect -1046 51 -1012 85
rect -1046 -17 -1012 17
rect -1046 -85 -1012 -51
rect 1012 51 1046 85
rect 1012 -17 1046 17
rect 1012 -85 1046 -51
<< poly >>
rect -1000 172 1000 188
rect -1000 138 -969 172
rect -935 138 -901 172
rect -867 138 -833 172
rect -799 138 -765 172
rect -731 138 -697 172
rect -663 138 -629 172
rect -595 138 -561 172
rect -527 138 -493 172
rect -459 138 -425 172
rect -391 138 -357 172
rect -323 138 -289 172
rect -255 138 -221 172
rect -187 138 -153 172
rect -119 138 -85 172
rect -51 138 -17 172
rect 17 138 51 172
rect 85 138 119 172
rect 153 138 187 172
rect 221 138 255 172
rect 289 138 323 172
rect 357 138 391 172
rect 425 138 459 172
rect 493 138 527 172
rect 561 138 595 172
rect 629 138 663 172
rect 697 138 731 172
rect 765 138 799 172
rect 833 138 867 172
rect 901 138 935 172
rect 969 138 1000 172
rect -1000 100 1000 138
rect -1000 -138 1000 -100
rect -1000 -172 -969 -138
rect -935 -172 -901 -138
rect -867 -172 -833 -138
rect -799 -172 -765 -138
rect -731 -172 -697 -138
rect -663 -172 -629 -138
rect -595 -172 -561 -138
rect -527 -172 -493 -138
rect -459 -172 -425 -138
rect -391 -172 -357 -138
rect -323 -172 -289 -138
rect -255 -172 -221 -138
rect -187 -172 -153 -138
rect -119 -172 -85 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 85 -172 119 -138
rect 153 -172 187 -138
rect 221 -172 255 -138
rect 289 -172 323 -138
rect 357 -172 391 -138
rect 425 -172 459 -138
rect 493 -172 527 -138
rect 561 -172 595 -138
rect 629 -172 663 -138
rect 697 -172 731 -138
rect 765 -172 799 -138
rect 833 -172 867 -138
rect 901 -172 935 -138
rect 969 -172 1000 -138
rect -1000 -188 1000 -172
<< polycont >>
rect -969 138 -935 172
rect -901 138 -867 172
rect -833 138 -799 172
rect -765 138 -731 172
rect -697 138 -663 172
rect -629 138 -595 172
rect -561 138 -527 172
rect -493 138 -459 172
rect -425 138 -391 172
rect -357 138 -323 172
rect -289 138 -255 172
rect -221 138 -187 172
rect -153 138 -119 172
rect -85 138 -51 172
rect -17 138 17 172
rect 51 138 85 172
rect 119 138 153 172
rect 187 138 221 172
rect 255 138 289 172
rect 323 138 357 172
rect 391 138 425 172
rect 459 138 493 172
rect 527 138 561 172
rect 595 138 629 172
rect 663 138 697 172
rect 731 138 765 172
rect 799 138 833 172
rect 867 138 901 172
rect 935 138 969 172
rect -969 -172 -935 -138
rect -901 -172 -867 -138
rect -833 -172 -799 -138
rect -765 -172 -731 -138
rect -697 -172 -663 -138
rect -629 -172 -595 -138
rect -561 -172 -527 -138
rect -493 -172 -459 -138
rect -425 -172 -391 -138
rect -357 -172 -323 -138
rect -289 -172 -255 -138
rect -221 -172 -187 -138
rect -153 -172 -119 -138
rect -85 -172 -51 -138
rect -17 -172 17 -138
rect 51 -172 85 -138
rect 119 -172 153 -138
rect 187 -172 221 -138
rect 255 -172 289 -138
rect 323 -172 357 -138
rect 391 -172 425 -138
rect 459 -172 493 -138
rect 527 -172 561 -138
rect 595 -172 629 -138
rect 663 -172 697 -138
rect 731 -172 765 -138
rect 799 -172 833 -138
rect 867 -172 901 -138
rect 935 -172 969 -138
<< locali >>
rect -1000 138 -969 172
rect -919 138 -901 172
rect -847 138 -833 172
rect -775 138 -765 172
rect -703 138 -697 172
rect -631 138 -629 172
rect -595 138 -593 172
rect -527 138 -521 172
rect -459 138 -449 172
rect -391 138 -377 172
rect -323 138 -305 172
rect -255 138 -233 172
rect -187 138 -161 172
rect -119 138 -89 172
rect -51 138 -17 172
rect 17 138 51 172
rect 89 138 119 172
rect 161 138 187 172
rect 233 138 255 172
rect 305 138 323 172
rect 377 138 391 172
rect 449 138 459 172
rect 521 138 527 172
rect 593 138 595 172
rect 629 138 631 172
rect 697 138 703 172
rect 765 138 775 172
rect 833 138 847 172
rect 901 138 919 172
rect 969 138 1000 172
rect -1046 85 -1012 104
rect -1046 17 -1012 19
rect -1046 -19 -1012 -17
rect -1046 -104 -1012 -85
rect 1012 85 1046 104
rect 1012 17 1046 19
rect 1012 -19 1046 -17
rect 1012 -104 1046 -85
rect -1000 -172 -969 -138
rect -919 -172 -901 -138
rect -847 -172 -833 -138
rect -775 -172 -765 -138
rect -703 -172 -697 -138
rect -631 -172 -629 -138
rect -595 -172 -593 -138
rect -527 -172 -521 -138
rect -459 -172 -449 -138
rect -391 -172 -377 -138
rect -323 -172 -305 -138
rect -255 -172 -233 -138
rect -187 -172 -161 -138
rect -119 -172 -89 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 89 -172 119 -138
rect 161 -172 187 -138
rect 233 -172 255 -138
rect 305 -172 323 -138
rect 377 -172 391 -138
rect 449 -172 459 -138
rect 521 -172 527 -138
rect 593 -172 595 -138
rect 629 -172 631 -138
rect 697 -172 703 -138
rect 765 -172 775 -138
rect 833 -172 847 -138
rect 901 -172 919 -138
rect 969 -172 1000 -138
<< viali >>
rect -953 138 -935 172
rect -935 138 -919 172
rect -881 138 -867 172
rect -867 138 -847 172
rect -809 138 -799 172
rect -799 138 -775 172
rect -737 138 -731 172
rect -731 138 -703 172
rect -665 138 -663 172
rect -663 138 -631 172
rect -593 138 -561 172
rect -561 138 -559 172
rect -521 138 -493 172
rect -493 138 -487 172
rect -449 138 -425 172
rect -425 138 -415 172
rect -377 138 -357 172
rect -357 138 -343 172
rect -305 138 -289 172
rect -289 138 -271 172
rect -233 138 -221 172
rect -221 138 -199 172
rect -161 138 -153 172
rect -153 138 -127 172
rect -89 138 -85 172
rect -85 138 -55 172
rect -17 138 17 172
rect 55 138 85 172
rect 85 138 89 172
rect 127 138 153 172
rect 153 138 161 172
rect 199 138 221 172
rect 221 138 233 172
rect 271 138 289 172
rect 289 138 305 172
rect 343 138 357 172
rect 357 138 377 172
rect 415 138 425 172
rect 425 138 449 172
rect 487 138 493 172
rect 493 138 521 172
rect 559 138 561 172
rect 561 138 593 172
rect 631 138 663 172
rect 663 138 665 172
rect 703 138 731 172
rect 731 138 737 172
rect 775 138 799 172
rect 799 138 809 172
rect 847 138 867 172
rect 867 138 881 172
rect 919 138 935 172
rect 935 138 953 172
rect -1046 51 -1012 53
rect -1046 19 -1012 51
rect -1046 -51 -1012 -19
rect -1046 -53 -1012 -51
rect 1012 51 1046 53
rect 1012 19 1046 51
rect 1012 -51 1046 -19
rect 1012 -53 1046 -51
rect -953 -172 -935 -138
rect -935 -172 -919 -138
rect -881 -172 -867 -138
rect -867 -172 -847 -138
rect -809 -172 -799 -138
rect -799 -172 -775 -138
rect -737 -172 -731 -138
rect -731 -172 -703 -138
rect -665 -172 -663 -138
rect -663 -172 -631 -138
rect -593 -172 -561 -138
rect -561 -172 -559 -138
rect -521 -172 -493 -138
rect -493 -172 -487 -138
rect -449 -172 -425 -138
rect -425 -172 -415 -138
rect -377 -172 -357 -138
rect -357 -172 -343 -138
rect -305 -172 -289 -138
rect -289 -172 -271 -138
rect -233 -172 -221 -138
rect -221 -172 -199 -138
rect -161 -172 -153 -138
rect -153 -172 -127 -138
rect -89 -172 -85 -138
rect -85 -172 -55 -138
rect -17 -172 17 -138
rect 55 -172 85 -138
rect 85 -172 89 -138
rect 127 -172 153 -138
rect 153 -172 161 -138
rect 199 -172 221 -138
rect 221 -172 233 -138
rect 271 -172 289 -138
rect 289 -172 305 -138
rect 343 -172 357 -138
rect 357 -172 377 -138
rect 415 -172 425 -138
rect 425 -172 449 -138
rect 487 -172 493 -138
rect 493 -172 521 -138
rect 559 -172 561 -138
rect 561 -172 593 -138
rect 631 -172 663 -138
rect 663 -172 665 -138
rect 703 -172 731 -138
rect 731 -172 737 -138
rect 775 -172 799 -138
rect 799 -172 809 -138
rect 847 -172 867 -138
rect 867 -172 881 -138
rect 919 -172 935 -138
rect 935 -172 953 -138
<< metal1 >>
rect -996 172 996 178
rect -996 138 -953 172
rect -919 138 -881 172
rect -847 138 -809 172
rect -775 138 -737 172
rect -703 138 -665 172
rect -631 138 -593 172
rect -559 138 -521 172
rect -487 138 -449 172
rect -415 138 -377 172
rect -343 138 -305 172
rect -271 138 -233 172
rect -199 138 -161 172
rect -127 138 -89 172
rect -55 138 -17 172
rect 17 138 55 172
rect 89 138 127 172
rect 161 138 199 172
rect 233 138 271 172
rect 305 138 343 172
rect 377 138 415 172
rect 449 138 487 172
rect 521 138 559 172
rect 593 138 631 172
rect 665 138 703 172
rect 737 138 775 172
rect 809 138 847 172
rect 881 138 919 172
rect 953 138 996 172
rect -996 132 996 138
rect -1052 53 -1006 100
rect -1052 19 -1046 53
rect -1012 19 -1006 53
rect -1052 -19 -1006 19
rect -1052 -53 -1046 -19
rect -1012 -53 -1006 -19
rect -1052 -100 -1006 -53
rect 1006 53 1052 100
rect 1006 19 1012 53
rect 1046 19 1052 53
rect 1006 -19 1052 19
rect 1006 -53 1012 -19
rect 1046 -53 1052 -19
rect 1006 -100 1052 -53
rect -996 -138 996 -132
rect -996 -172 -953 -138
rect -919 -172 -881 -138
rect -847 -172 -809 -138
rect -775 -172 -737 -138
rect -703 -172 -665 -138
rect -631 -172 -593 -138
rect -559 -172 -521 -138
rect -487 -172 -449 -138
rect -415 -172 -377 -138
rect -343 -172 -305 -138
rect -271 -172 -233 -138
rect -199 -172 -161 -138
rect -127 -172 -89 -138
rect -55 -172 -17 -138
rect 17 -172 55 -138
rect 89 -172 127 -138
rect 161 -172 199 -138
rect 233 -172 271 -138
rect 305 -172 343 -138
rect 377 -172 415 -138
rect 449 -172 487 -138
rect 521 -172 559 -138
rect 593 -172 631 -138
rect 665 -172 703 -138
rect 737 -172 775 -138
rect 809 -172 847 -138
rect 881 -172 919 -138
rect 953 -172 996 -138
rect -996 -178 996 -172
<< end >>
