magic
tech sky130B
timestamp 1668220879
<< metal4 >>
rect 2700 -3550 3200 7000
rect 2700 -3700 2750 -3550
rect 2900 -3700 2950 -3550
rect 3100 -3700 3200 -3550
rect 2700 -3750 3200 -3700
rect 2700 -3900 2800 -3750
rect 2950 -3900 3000 -3750
rect 3150 -3900 3200 -3750
rect 2700 -4000 3200 -3900
<< via4 >>
rect 2750 -3700 2900 -3550
rect 2950 -3700 3100 -3550
rect 2800 -3900 2950 -3750
rect 3000 -3900 3150 -3750
<< metal5 >>
rect -4650 6400 17900 6900
rect -6900 5600 17100 6100
rect -6900 -17400 -6400 5600
rect -6100 4800 16300 5300
rect -6100 -16600 -5600 4800
rect -5300 4000 15500 4500
rect -5300 -15800 -4800 4000
rect -4500 3200 14700 3700
rect -4500 -15000 -4000 3200
rect -3700 2400 13900 2900
rect -3700 -14200 -3200 2400
rect -2900 1600 13100 2100
rect -2900 -13400 -2400 1600
rect -2100 800 12300 1300
rect -2100 -12600 -1600 800
rect -1300 0 11500 500
rect -1300 -11800 -800 0
rect -500 -800 10700 -300
rect -500 -11000 0 -800
rect 300 -1600 9900 -1100
rect 300 -10200 800 -1600
rect 1100 -2400 9100 -1900
rect 1100 -9400 1600 -2400
rect 1900 -3200 8300 -2700
rect 1900 -8600 2400 -3200
rect 2700 -3550 3200 -3500
rect 2700 -3700 2750 -3550
rect 2900 -3700 2950 -3550
rect 3100 -3700 3200 -3550
rect 2700 -3750 3200 -3700
rect 2700 -3900 2800 -3750
rect 2950 -3900 3000 -3750
rect 3150 -3900 3200 -3750
rect 2700 -7800 3200 -3900
rect 7800 -7800 8300 -3200
rect 2700 -8300 8300 -7800
rect 8600 -8600 9100 -2400
rect 1900 -9100 9100 -8600
rect 9400 -9400 9900 -1600
rect 1100 -9900 9900 -9400
rect 10200 -10200 10700 -800
rect 300 -10700 10700 -10200
rect 11000 -11000 11500 0
rect -500 -11500 11500 -11000
rect 11800 -11800 12300 800
rect -1300 -12300 12300 -11800
rect 12600 -12600 13100 1600
rect -2100 -13100 13100 -12600
rect 13400 -13400 13900 2400
rect -2900 -13900 13900 -13400
rect 14200 -14200 14700 3200
rect -3700 -14700 14700 -14200
rect 15000 -15000 15500 4000
rect -4500 -15500 15500 -15000
rect 15800 -15800 16300 4800
rect -5300 -16300 16300 -15800
rect 16600 -16600 17100 5600
rect -6100 -17100 17100 -16600
rect 17400 -17400 17900 6400
rect -6900 -17900 17900 -17400
<< end >>
