magic
tech sky130A
magscale 1 2
timestamp 1667444884
<< nwell >>
rect -323 -1500 323 1500
<< pmos >>
rect -229 -1400 -29 1400
rect 29 -1400 229 1400
<< pdiff >>
rect -287 1388 -229 1400
rect -287 -1388 -275 1388
rect -241 -1388 -229 1388
rect -287 -1400 -229 -1388
rect -29 1388 29 1400
rect -29 -1388 -17 1388
rect 17 -1388 29 1388
rect -29 -1400 29 -1388
rect 229 1388 287 1400
rect 229 -1388 241 1388
rect 275 -1388 287 1388
rect 229 -1400 287 -1388
<< pdiffc >>
rect -275 -1388 -241 1388
rect -17 -1388 17 1388
rect 241 -1388 275 1388
<< poly >>
rect -229 1481 -29 1497
rect -229 1447 -213 1481
rect -45 1447 -29 1481
rect -229 1400 -29 1447
rect 29 1481 229 1497
rect 29 1447 45 1481
rect 213 1447 229 1481
rect 29 1400 229 1447
rect -229 -1447 -29 -1400
rect -229 -1481 -213 -1447
rect -45 -1481 -29 -1447
rect -229 -1497 -29 -1481
rect 29 -1447 229 -1400
rect 29 -1481 45 -1447
rect 213 -1481 229 -1447
rect 29 -1497 229 -1481
<< polycont >>
rect -213 1447 -45 1481
rect 45 1447 213 1481
rect -213 -1481 -45 -1447
rect 45 -1481 213 -1447
<< locali >>
rect -229 1447 -213 1481
rect -45 1447 -29 1481
rect 29 1447 45 1481
rect 213 1447 229 1481
rect -275 1388 -241 1404
rect -275 -1404 -241 -1388
rect -17 1388 17 1404
rect -17 -1404 17 -1388
rect 241 1388 275 1404
rect 241 -1404 275 -1388
rect -229 -1481 -213 -1447
rect -45 -1481 -29 -1447
rect 29 -1481 45 -1447
rect 213 -1481 229 -1447
<< viali >>
rect -213 1447 -45 1481
rect 45 1447 213 1481
rect -275 -1388 -241 1388
rect -17 -1388 17 1388
rect 241 -1388 275 1388
rect -213 -1481 -45 -1447
rect 45 -1481 213 -1447
<< metal1 >>
rect -225 1481 -33 1487
rect -225 1447 -213 1481
rect -45 1447 -33 1481
rect -225 1441 -33 1447
rect 33 1481 225 1487
rect 33 1447 45 1481
rect 213 1447 225 1481
rect 33 1441 225 1447
rect -281 1388 -235 1400
rect -281 -1388 -275 1388
rect -241 -1388 -235 1388
rect -281 -1400 -235 -1388
rect -23 1388 23 1400
rect -23 -1388 -17 1388
rect 17 -1388 23 1388
rect -23 -1400 23 -1388
rect 235 1388 281 1400
rect 235 -1388 241 1388
rect 275 -1388 281 1388
rect 235 -1400 281 -1388
rect -225 -1447 -33 -1441
rect -225 -1481 -213 -1447
rect -45 -1481 -33 -1447
rect -225 -1487 -33 -1481
rect 33 -1447 225 -1441
rect 33 -1481 45 -1447
rect 213 -1481 225 -1447
rect 33 -1487 225 -1481
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 14.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
