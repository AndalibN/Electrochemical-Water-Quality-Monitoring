magic
tech sky130A
magscale 1 2
timestamp 1667263279
<< xpolycontact >>
rect -35 175 35 607
rect -35 -607 35 -175
<< ppolyres >>
rect -35 -175 35 175
<< viali >>
rect -19 192 19 589
rect -19 -589 19 -192
<< metal1 >>
rect -25 589 25 601
rect -25 192 -19 589
rect 19 192 25 589
rect -25 180 25 192
rect -25 -192 25 -180
rect -25 -589 -19 -192
rect 19 -589 25 -192
rect -25 -601 25 -589
<< res0p35 >>
rect -37 -177 37 177
<< properties >>
string gencell sky130_fd_pr__res_high_po_0p35
string library sky130
string parameters w 0.350 l 1.75 m 1 nx 1 wmin 0.350 lmin 0.50 rho 319.8 val 2.712k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 0.350 vias 1 n_guard 0 hv_guard 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
