magic
tech sky130A
magscale 1 2
timestamp 1666894475
<< error_p >>
rect -200 2912 -142 2918
rect -86 2912 -28 2918
rect 28 2912 86 2918
rect 142 2912 200 2918
rect -200 2878 -188 2912
rect -86 2878 -74 2912
rect 28 2878 40 2912
rect 142 2878 154 2912
rect -200 2872 -142 2878
rect -86 2872 -28 2878
rect 28 2872 86 2878
rect 142 2872 200 2878
rect -200 -2878 -142 -2872
rect -86 -2878 -28 -2872
rect 28 -2878 86 -2872
rect 142 -2878 200 -2872
rect -200 -2912 -188 -2878
rect -86 -2912 -74 -2878
rect 28 -2912 40 -2878
rect 142 -2912 154 -2878
rect -200 -2918 -142 -2912
rect -86 -2918 -28 -2912
rect 28 -2918 86 -2912
rect 142 -2918 200 -2912
<< pwell >>
rect -395 -3050 395 3050
<< nmos >>
rect -199 -2840 -143 2840
rect -85 -2840 -29 2840
rect 29 -2840 85 2840
rect 143 -2840 199 2840
<< ndiff >>
rect -257 2828 -199 2840
rect -257 -2828 -245 2828
rect -211 -2828 -199 2828
rect -257 -2840 -199 -2828
rect -143 2828 -85 2840
rect -143 -2828 -131 2828
rect -97 -2828 -85 2828
rect -143 -2840 -85 -2828
rect -29 2828 29 2840
rect -29 -2828 -17 2828
rect 17 -2828 29 2828
rect -29 -2840 29 -2828
rect 85 2828 143 2840
rect 85 -2828 97 2828
rect 131 -2828 143 2828
rect 85 -2840 143 -2828
rect 199 2828 257 2840
rect 199 -2828 211 2828
rect 245 -2828 257 2828
rect 199 -2840 257 -2828
<< ndiffc >>
rect -245 -2828 -211 2828
rect -131 -2828 -97 2828
rect -17 -2828 17 2828
rect 97 -2828 131 2828
rect 211 -2828 245 2828
<< psubdiff >>
rect -359 2980 -263 3014
rect 263 2980 359 3014
rect -359 2918 -325 2980
rect 325 2918 359 2980
rect -359 -2980 -325 -2918
rect 325 -2980 359 -2918
rect -359 -3014 -263 -2980
rect 263 -3014 359 -2980
<< psubdiffcont >>
rect -263 2980 263 3014
rect -359 -2918 -325 2918
rect 325 -2918 359 2918
rect -263 -3014 263 -2980
<< poly >>
rect -204 2912 -138 2928
rect -204 2878 -188 2912
rect -154 2878 -138 2912
rect -204 2862 -138 2878
rect -90 2912 -24 2928
rect -90 2878 -74 2912
rect -40 2878 -24 2912
rect -90 2862 -24 2878
rect 24 2912 90 2928
rect 24 2878 40 2912
rect 74 2878 90 2912
rect 24 2862 90 2878
rect 138 2912 204 2928
rect 138 2878 154 2912
rect 188 2878 204 2912
rect 138 2862 204 2878
rect -199 2840 -143 2862
rect -85 2840 -29 2862
rect 29 2840 85 2862
rect 143 2840 199 2862
rect -199 -2862 -143 -2840
rect -85 -2862 -29 -2840
rect 29 -2862 85 -2840
rect 143 -2862 199 -2840
rect -204 -2878 -138 -2862
rect -204 -2912 -188 -2878
rect -154 -2912 -138 -2878
rect -204 -2928 -138 -2912
rect -90 -2878 -24 -2862
rect -90 -2912 -74 -2878
rect -40 -2912 -24 -2878
rect -90 -2928 -24 -2912
rect 24 -2878 90 -2862
rect 24 -2912 40 -2878
rect 74 -2912 90 -2878
rect 24 -2928 90 -2912
rect 138 -2878 204 -2862
rect 138 -2912 154 -2878
rect 188 -2912 204 -2878
rect 138 -2928 204 -2912
<< polycont >>
rect -188 2878 -154 2912
rect -74 2878 -40 2912
rect 40 2878 74 2912
rect 154 2878 188 2912
rect -188 -2912 -154 -2878
rect -74 -2912 -40 -2878
rect 40 -2912 74 -2878
rect 154 -2912 188 -2878
<< locali >>
rect -359 2980 -263 3014
rect 263 2980 359 3014
rect -359 2918 -325 2980
rect 325 2918 359 2980
rect -204 2878 -188 2912
rect -154 2878 -138 2912
rect -90 2878 -74 2912
rect -40 2878 -24 2912
rect 24 2878 40 2912
rect 74 2878 90 2912
rect 138 2878 154 2912
rect 188 2878 204 2912
rect -245 2828 -211 2844
rect -245 -2844 -211 -2828
rect -131 2828 -97 2844
rect -131 -2844 -97 -2828
rect -17 2828 17 2844
rect -17 -2844 17 -2828
rect 97 2828 131 2844
rect 97 -2844 131 -2828
rect 211 2828 245 2844
rect 211 -2844 245 -2828
rect -204 -2912 -188 -2878
rect -154 -2912 -138 -2878
rect -90 -2912 -74 -2878
rect -40 -2912 -24 -2878
rect 24 -2912 40 -2878
rect 74 -2912 90 -2878
rect 138 -2912 154 -2878
rect 188 -2912 204 -2878
rect -359 -2980 -325 -2918
rect 325 -2980 359 -2918
rect -359 -3014 -263 -2980
rect 263 -3014 359 -2980
<< viali >>
rect -188 2878 -154 2912
rect -74 2878 -40 2912
rect 40 2878 74 2912
rect 154 2878 188 2912
rect -245 -2828 -211 2828
rect -131 -2828 -97 2828
rect -17 -2828 17 2828
rect 97 -2828 131 2828
rect 211 -2828 245 2828
rect -188 -2912 -154 -2878
rect -74 -2912 -40 -2878
rect 40 -2912 74 -2878
rect 154 -2912 188 -2878
<< metal1 >>
rect -200 2912 -142 2918
rect -200 2878 -188 2912
rect -154 2878 -142 2912
rect -200 2872 -142 2878
rect -86 2912 -28 2918
rect -86 2878 -74 2912
rect -40 2878 -28 2912
rect -86 2872 -28 2878
rect 28 2912 86 2918
rect 28 2878 40 2912
rect 74 2878 86 2912
rect 28 2872 86 2878
rect 142 2912 200 2918
rect 142 2878 154 2912
rect 188 2878 200 2912
rect 142 2872 200 2878
rect -251 2828 -205 2840
rect -251 -2828 -245 2828
rect -211 -2828 -205 2828
rect -251 -2840 -205 -2828
rect -137 2828 -91 2840
rect -137 -2828 -131 2828
rect -97 -2828 -91 2828
rect -137 -2840 -91 -2828
rect -23 2828 23 2840
rect -23 -2828 -17 2828
rect 17 -2828 23 2828
rect -23 -2840 23 -2828
rect 91 2828 137 2840
rect 91 -2828 97 2828
rect 131 -2828 137 2828
rect 91 -2840 137 -2828
rect 205 2828 251 2840
rect 205 -2828 211 2828
rect 245 -2828 251 2828
rect 205 -2840 251 -2828
rect -200 -2878 -142 -2872
rect -200 -2912 -188 -2878
rect -154 -2912 -142 -2878
rect -200 -2918 -142 -2912
rect -86 -2878 -28 -2872
rect -86 -2912 -74 -2878
rect -40 -2912 -28 -2878
rect -86 -2918 -28 -2912
rect 28 -2878 86 -2872
rect 28 -2912 40 -2878
rect 74 -2912 86 -2878
rect 28 -2918 86 -2912
rect 142 -2878 200 -2872
rect 142 -2912 154 -2878
rect 188 -2912 200 -2878
rect 142 -2918 200 -2912
<< properties >>
string FIXED_BBOX -342 -2997 342 2997
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 28.4 l 0.28 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
