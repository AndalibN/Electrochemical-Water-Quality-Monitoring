magic
tech sky130A
magscale 1 2
timestamp 1667488624
<< error_p >>
rect -941 1993 -883 1999
rect -749 1993 -691 1999
rect -557 1993 -499 1999
rect -365 1993 -307 1999
rect -173 1993 -115 1999
rect 19 1993 77 1999
rect 211 1993 269 1999
rect 403 1993 461 1999
rect 595 1993 653 1999
rect 787 1993 845 1999
rect -941 1959 -929 1993
rect -749 1959 -737 1993
rect -557 1959 -545 1993
rect -365 1959 -353 1993
rect -173 1959 -161 1993
rect 19 1959 31 1993
rect 211 1959 223 1993
rect 403 1959 415 1993
rect 595 1959 607 1993
rect 787 1959 799 1993
rect -941 1953 -883 1959
rect -749 1953 -691 1959
rect -557 1953 -499 1959
rect -365 1953 -307 1959
rect -173 1953 -115 1959
rect 19 1953 77 1959
rect 211 1953 269 1959
rect 403 1953 461 1959
rect 595 1953 653 1959
rect 787 1953 845 1959
rect -845 1695 -787 1701
rect -653 1695 -595 1701
rect -461 1695 -403 1701
rect -269 1695 -211 1701
rect -77 1695 -19 1701
rect 115 1695 173 1701
rect 307 1695 365 1701
rect 499 1695 557 1701
rect 691 1695 749 1701
rect 883 1695 941 1701
rect -845 1661 -833 1695
rect -653 1661 -641 1695
rect -461 1661 -449 1695
rect -269 1661 -257 1695
rect -77 1661 -65 1695
rect 115 1661 127 1695
rect 307 1661 319 1695
rect 499 1661 511 1695
rect 691 1661 703 1695
rect 883 1661 895 1695
rect -845 1655 -787 1661
rect -653 1655 -595 1661
rect -461 1655 -403 1661
rect -269 1655 -211 1661
rect -77 1655 -19 1661
rect 115 1655 173 1661
rect 307 1655 365 1661
rect 499 1655 557 1661
rect 691 1655 749 1661
rect 883 1655 941 1661
rect -845 1587 -787 1593
rect -653 1587 -595 1593
rect -461 1587 -403 1593
rect -269 1587 -211 1593
rect -77 1587 -19 1593
rect 115 1587 173 1593
rect 307 1587 365 1593
rect 499 1587 557 1593
rect 691 1587 749 1593
rect 883 1587 941 1593
rect -845 1553 -833 1587
rect -653 1553 -641 1587
rect -461 1553 -449 1587
rect -269 1553 -257 1587
rect -77 1553 -65 1587
rect 115 1553 127 1587
rect 307 1553 319 1587
rect 499 1553 511 1587
rect 691 1553 703 1587
rect 883 1553 895 1587
rect -845 1547 -787 1553
rect -653 1547 -595 1553
rect -461 1547 -403 1553
rect -269 1547 -211 1553
rect -77 1547 -19 1553
rect 115 1547 173 1553
rect 307 1547 365 1553
rect 499 1547 557 1553
rect 691 1547 749 1553
rect 883 1547 941 1553
rect -941 1289 -883 1295
rect -749 1289 -691 1295
rect -557 1289 -499 1295
rect -365 1289 -307 1295
rect -173 1289 -115 1295
rect 19 1289 77 1295
rect 211 1289 269 1295
rect 403 1289 461 1295
rect 595 1289 653 1295
rect 787 1289 845 1295
rect -941 1255 -929 1289
rect -749 1255 -737 1289
rect -557 1255 -545 1289
rect -365 1255 -353 1289
rect -173 1255 -161 1289
rect 19 1255 31 1289
rect 211 1255 223 1289
rect 403 1255 415 1289
rect 595 1255 607 1289
rect 787 1255 799 1289
rect -941 1249 -883 1255
rect -749 1249 -691 1255
rect -557 1249 -499 1255
rect -365 1249 -307 1255
rect -173 1249 -115 1255
rect 19 1249 77 1255
rect 211 1249 269 1255
rect 403 1249 461 1255
rect 595 1249 653 1255
rect 787 1249 845 1255
rect -941 1181 -883 1187
rect -749 1181 -691 1187
rect -557 1181 -499 1187
rect -365 1181 -307 1187
rect -173 1181 -115 1187
rect 19 1181 77 1187
rect 211 1181 269 1187
rect 403 1181 461 1187
rect 595 1181 653 1187
rect 787 1181 845 1187
rect -941 1147 -929 1181
rect -749 1147 -737 1181
rect -557 1147 -545 1181
rect -365 1147 -353 1181
rect -173 1147 -161 1181
rect 19 1147 31 1181
rect 211 1147 223 1181
rect 403 1147 415 1181
rect 595 1147 607 1181
rect 787 1147 799 1181
rect -941 1141 -883 1147
rect -749 1141 -691 1147
rect -557 1141 -499 1147
rect -365 1141 -307 1147
rect -173 1141 -115 1147
rect 19 1141 77 1147
rect 211 1141 269 1147
rect 403 1141 461 1147
rect 595 1141 653 1147
rect 787 1141 845 1147
rect -845 883 -787 889
rect -653 883 -595 889
rect -461 883 -403 889
rect -269 883 -211 889
rect -77 883 -19 889
rect 115 883 173 889
rect 307 883 365 889
rect 499 883 557 889
rect 691 883 749 889
rect 883 883 941 889
rect -845 849 -833 883
rect -653 849 -641 883
rect -461 849 -449 883
rect -269 849 -257 883
rect -77 849 -65 883
rect 115 849 127 883
rect 307 849 319 883
rect 499 849 511 883
rect 691 849 703 883
rect 883 849 895 883
rect -845 843 -787 849
rect -653 843 -595 849
rect -461 843 -403 849
rect -269 843 -211 849
rect -77 843 -19 849
rect 115 843 173 849
rect 307 843 365 849
rect 499 843 557 849
rect 691 843 749 849
rect 883 843 941 849
rect -845 775 -787 781
rect -653 775 -595 781
rect -461 775 -403 781
rect -269 775 -211 781
rect -77 775 -19 781
rect 115 775 173 781
rect 307 775 365 781
rect 499 775 557 781
rect 691 775 749 781
rect 883 775 941 781
rect -845 741 -833 775
rect -653 741 -641 775
rect -461 741 -449 775
rect -269 741 -257 775
rect -77 741 -65 775
rect 115 741 127 775
rect 307 741 319 775
rect 499 741 511 775
rect 691 741 703 775
rect 883 741 895 775
rect -845 735 -787 741
rect -653 735 -595 741
rect -461 735 -403 741
rect -269 735 -211 741
rect -77 735 -19 741
rect 115 735 173 741
rect 307 735 365 741
rect 499 735 557 741
rect 691 735 749 741
rect 883 735 941 741
rect -941 477 -883 483
rect -749 477 -691 483
rect -557 477 -499 483
rect -365 477 -307 483
rect -173 477 -115 483
rect 19 477 77 483
rect 211 477 269 483
rect 403 477 461 483
rect 595 477 653 483
rect 787 477 845 483
rect -941 443 -929 477
rect -749 443 -737 477
rect -557 443 -545 477
rect -365 443 -353 477
rect -173 443 -161 477
rect 19 443 31 477
rect 211 443 223 477
rect 403 443 415 477
rect 595 443 607 477
rect 787 443 799 477
rect -941 437 -883 443
rect -749 437 -691 443
rect -557 437 -499 443
rect -365 437 -307 443
rect -173 437 -115 443
rect 19 437 77 443
rect 211 437 269 443
rect 403 437 461 443
rect 595 437 653 443
rect 787 437 845 443
rect -941 369 -883 375
rect -749 369 -691 375
rect -557 369 -499 375
rect -365 369 -307 375
rect -173 369 -115 375
rect 19 369 77 375
rect 211 369 269 375
rect 403 369 461 375
rect 595 369 653 375
rect 787 369 845 375
rect -941 335 -929 369
rect -749 335 -737 369
rect -557 335 -545 369
rect -365 335 -353 369
rect -173 335 -161 369
rect 19 335 31 369
rect 211 335 223 369
rect 403 335 415 369
rect 595 335 607 369
rect 787 335 799 369
rect -941 329 -883 335
rect -749 329 -691 335
rect -557 329 -499 335
rect -365 329 -307 335
rect -173 329 -115 335
rect 19 329 77 335
rect 211 329 269 335
rect 403 329 461 335
rect 595 329 653 335
rect 787 329 845 335
rect -845 71 -787 77
rect -653 71 -595 77
rect -461 71 -403 77
rect -269 71 -211 77
rect -77 71 -19 77
rect 115 71 173 77
rect 307 71 365 77
rect 499 71 557 77
rect 691 71 749 77
rect 883 71 941 77
rect -845 37 -833 71
rect -653 37 -641 71
rect -461 37 -449 71
rect -269 37 -257 71
rect -77 37 -65 71
rect 115 37 127 71
rect 307 37 319 71
rect 499 37 511 71
rect 691 37 703 71
rect 883 37 895 71
rect -845 31 -787 37
rect -653 31 -595 37
rect -461 31 -403 37
rect -269 31 -211 37
rect -77 31 -19 37
rect 115 31 173 37
rect 307 31 365 37
rect 499 31 557 37
rect 691 31 749 37
rect 883 31 941 37
rect -845 -37 -787 -31
rect -653 -37 -595 -31
rect -461 -37 -403 -31
rect -269 -37 -211 -31
rect -77 -37 -19 -31
rect 115 -37 173 -31
rect 307 -37 365 -31
rect 499 -37 557 -31
rect 691 -37 749 -31
rect 883 -37 941 -31
rect -845 -71 -833 -37
rect -653 -71 -641 -37
rect -461 -71 -449 -37
rect -269 -71 -257 -37
rect -77 -71 -65 -37
rect 115 -71 127 -37
rect 307 -71 319 -37
rect 499 -71 511 -37
rect 691 -71 703 -37
rect 883 -71 895 -37
rect -845 -77 -787 -71
rect -653 -77 -595 -71
rect -461 -77 -403 -71
rect -269 -77 -211 -71
rect -77 -77 -19 -71
rect 115 -77 173 -71
rect 307 -77 365 -71
rect 499 -77 557 -71
rect 691 -77 749 -71
rect 883 -77 941 -71
rect -941 -335 -883 -329
rect -749 -335 -691 -329
rect -557 -335 -499 -329
rect -365 -335 -307 -329
rect -173 -335 -115 -329
rect 19 -335 77 -329
rect 211 -335 269 -329
rect 403 -335 461 -329
rect 595 -335 653 -329
rect 787 -335 845 -329
rect -941 -369 -929 -335
rect -749 -369 -737 -335
rect -557 -369 -545 -335
rect -365 -369 -353 -335
rect -173 -369 -161 -335
rect 19 -369 31 -335
rect 211 -369 223 -335
rect 403 -369 415 -335
rect 595 -369 607 -335
rect 787 -369 799 -335
rect -941 -375 -883 -369
rect -749 -375 -691 -369
rect -557 -375 -499 -369
rect -365 -375 -307 -369
rect -173 -375 -115 -369
rect 19 -375 77 -369
rect 211 -375 269 -369
rect 403 -375 461 -369
rect 595 -375 653 -369
rect 787 -375 845 -369
rect -941 -443 -883 -437
rect -749 -443 -691 -437
rect -557 -443 -499 -437
rect -365 -443 -307 -437
rect -173 -443 -115 -437
rect 19 -443 77 -437
rect 211 -443 269 -437
rect 403 -443 461 -437
rect 595 -443 653 -437
rect 787 -443 845 -437
rect -941 -477 -929 -443
rect -749 -477 -737 -443
rect -557 -477 -545 -443
rect -365 -477 -353 -443
rect -173 -477 -161 -443
rect 19 -477 31 -443
rect 211 -477 223 -443
rect 403 -477 415 -443
rect 595 -477 607 -443
rect 787 -477 799 -443
rect -941 -483 -883 -477
rect -749 -483 -691 -477
rect -557 -483 -499 -477
rect -365 -483 -307 -477
rect -173 -483 -115 -477
rect 19 -483 77 -477
rect 211 -483 269 -477
rect 403 -483 461 -477
rect 595 -483 653 -477
rect 787 -483 845 -477
rect -845 -741 -787 -735
rect -653 -741 -595 -735
rect -461 -741 -403 -735
rect -269 -741 -211 -735
rect -77 -741 -19 -735
rect 115 -741 173 -735
rect 307 -741 365 -735
rect 499 -741 557 -735
rect 691 -741 749 -735
rect 883 -741 941 -735
rect -845 -775 -833 -741
rect -653 -775 -641 -741
rect -461 -775 -449 -741
rect -269 -775 -257 -741
rect -77 -775 -65 -741
rect 115 -775 127 -741
rect 307 -775 319 -741
rect 499 -775 511 -741
rect 691 -775 703 -741
rect 883 -775 895 -741
rect -845 -781 -787 -775
rect -653 -781 -595 -775
rect -461 -781 -403 -775
rect -269 -781 -211 -775
rect -77 -781 -19 -775
rect 115 -781 173 -775
rect 307 -781 365 -775
rect 499 -781 557 -775
rect 691 -781 749 -775
rect 883 -781 941 -775
rect -845 -849 -787 -843
rect -653 -849 -595 -843
rect -461 -849 -403 -843
rect -269 -849 -211 -843
rect -77 -849 -19 -843
rect 115 -849 173 -843
rect 307 -849 365 -843
rect 499 -849 557 -843
rect 691 -849 749 -843
rect 883 -849 941 -843
rect -845 -883 -833 -849
rect -653 -883 -641 -849
rect -461 -883 -449 -849
rect -269 -883 -257 -849
rect -77 -883 -65 -849
rect 115 -883 127 -849
rect 307 -883 319 -849
rect 499 -883 511 -849
rect 691 -883 703 -849
rect 883 -883 895 -849
rect -845 -889 -787 -883
rect -653 -889 -595 -883
rect -461 -889 -403 -883
rect -269 -889 -211 -883
rect -77 -889 -19 -883
rect 115 -889 173 -883
rect 307 -889 365 -883
rect 499 -889 557 -883
rect 691 -889 749 -883
rect 883 -889 941 -883
rect -941 -1147 -883 -1141
rect -749 -1147 -691 -1141
rect -557 -1147 -499 -1141
rect -365 -1147 -307 -1141
rect -173 -1147 -115 -1141
rect 19 -1147 77 -1141
rect 211 -1147 269 -1141
rect 403 -1147 461 -1141
rect 595 -1147 653 -1141
rect 787 -1147 845 -1141
rect -941 -1181 -929 -1147
rect -749 -1181 -737 -1147
rect -557 -1181 -545 -1147
rect -365 -1181 -353 -1147
rect -173 -1181 -161 -1147
rect 19 -1181 31 -1147
rect 211 -1181 223 -1147
rect 403 -1181 415 -1147
rect 595 -1181 607 -1147
rect 787 -1181 799 -1147
rect -941 -1187 -883 -1181
rect -749 -1187 -691 -1181
rect -557 -1187 -499 -1181
rect -365 -1187 -307 -1181
rect -173 -1187 -115 -1181
rect 19 -1187 77 -1181
rect 211 -1187 269 -1181
rect 403 -1187 461 -1181
rect 595 -1187 653 -1181
rect 787 -1187 845 -1181
rect -941 -1255 -883 -1249
rect -749 -1255 -691 -1249
rect -557 -1255 -499 -1249
rect -365 -1255 -307 -1249
rect -173 -1255 -115 -1249
rect 19 -1255 77 -1249
rect 211 -1255 269 -1249
rect 403 -1255 461 -1249
rect 595 -1255 653 -1249
rect 787 -1255 845 -1249
rect -941 -1289 -929 -1255
rect -749 -1289 -737 -1255
rect -557 -1289 -545 -1255
rect -365 -1289 -353 -1255
rect -173 -1289 -161 -1255
rect 19 -1289 31 -1255
rect 211 -1289 223 -1255
rect 403 -1289 415 -1255
rect 595 -1289 607 -1255
rect 787 -1289 799 -1255
rect -941 -1295 -883 -1289
rect -749 -1295 -691 -1289
rect -557 -1295 -499 -1289
rect -365 -1295 -307 -1289
rect -173 -1295 -115 -1289
rect 19 -1295 77 -1289
rect 211 -1295 269 -1289
rect 403 -1295 461 -1289
rect 595 -1295 653 -1289
rect 787 -1295 845 -1289
rect -845 -1553 -787 -1547
rect -653 -1553 -595 -1547
rect -461 -1553 -403 -1547
rect -269 -1553 -211 -1547
rect -77 -1553 -19 -1547
rect 115 -1553 173 -1547
rect 307 -1553 365 -1547
rect 499 -1553 557 -1547
rect 691 -1553 749 -1547
rect 883 -1553 941 -1547
rect -845 -1587 -833 -1553
rect -653 -1587 -641 -1553
rect -461 -1587 -449 -1553
rect -269 -1587 -257 -1553
rect -77 -1587 -65 -1553
rect 115 -1587 127 -1553
rect 307 -1587 319 -1553
rect 499 -1587 511 -1553
rect 691 -1587 703 -1553
rect 883 -1587 895 -1553
rect -845 -1593 -787 -1587
rect -653 -1593 -595 -1587
rect -461 -1593 -403 -1587
rect -269 -1593 -211 -1587
rect -77 -1593 -19 -1587
rect 115 -1593 173 -1587
rect 307 -1593 365 -1587
rect 499 -1593 557 -1587
rect 691 -1593 749 -1587
rect 883 -1593 941 -1587
rect -845 -1661 -787 -1655
rect -653 -1661 -595 -1655
rect -461 -1661 -403 -1655
rect -269 -1661 -211 -1655
rect -77 -1661 -19 -1655
rect 115 -1661 173 -1655
rect 307 -1661 365 -1655
rect 499 -1661 557 -1655
rect 691 -1661 749 -1655
rect 883 -1661 941 -1655
rect -845 -1695 -833 -1661
rect -653 -1695 -641 -1661
rect -461 -1695 -449 -1661
rect -269 -1695 -257 -1661
rect -77 -1695 -65 -1661
rect 115 -1695 127 -1661
rect 307 -1695 319 -1661
rect 499 -1695 511 -1661
rect 691 -1695 703 -1661
rect 883 -1695 895 -1661
rect -845 -1701 -787 -1695
rect -653 -1701 -595 -1695
rect -461 -1701 -403 -1695
rect -269 -1701 -211 -1695
rect -77 -1701 -19 -1695
rect 115 -1701 173 -1695
rect 307 -1701 365 -1695
rect 499 -1701 557 -1695
rect 691 -1701 749 -1695
rect 883 -1701 941 -1695
rect -941 -1959 -883 -1953
rect -749 -1959 -691 -1953
rect -557 -1959 -499 -1953
rect -365 -1959 -307 -1953
rect -173 -1959 -115 -1953
rect 19 -1959 77 -1953
rect 211 -1959 269 -1953
rect 403 -1959 461 -1953
rect 595 -1959 653 -1953
rect 787 -1959 845 -1953
rect -941 -1993 -929 -1959
rect -749 -1993 -737 -1959
rect -557 -1993 -545 -1959
rect -365 -1993 -353 -1959
rect -173 -1993 -161 -1959
rect 19 -1993 31 -1959
rect 211 -1993 223 -1959
rect 403 -1993 415 -1959
rect 595 -1993 607 -1959
rect 787 -1993 799 -1959
rect -941 -1999 -883 -1993
rect -749 -1999 -691 -1993
rect -557 -1999 -499 -1993
rect -365 -1999 -307 -1993
rect -173 -1999 -115 -1993
rect 19 -1999 77 -1993
rect 211 -1999 269 -1993
rect 403 -1999 461 -1993
rect 595 -1999 653 -1993
rect 787 -1999 845 -1993
<< nwell >>
rect -1127 -2131 1127 2131
<< pmos >>
rect -927 1742 -897 1912
rect -831 1742 -801 1912
rect -735 1742 -705 1912
rect -639 1742 -609 1912
rect -543 1742 -513 1912
rect -447 1742 -417 1912
rect -351 1742 -321 1912
rect -255 1742 -225 1912
rect -159 1742 -129 1912
rect -63 1742 -33 1912
rect 33 1742 63 1912
rect 129 1742 159 1912
rect 225 1742 255 1912
rect 321 1742 351 1912
rect 417 1742 447 1912
rect 513 1742 543 1912
rect 609 1742 639 1912
rect 705 1742 735 1912
rect 801 1742 831 1912
rect 897 1742 927 1912
rect -927 1336 -897 1506
rect -831 1336 -801 1506
rect -735 1336 -705 1506
rect -639 1336 -609 1506
rect -543 1336 -513 1506
rect -447 1336 -417 1506
rect -351 1336 -321 1506
rect -255 1336 -225 1506
rect -159 1336 -129 1506
rect -63 1336 -33 1506
rect 33 1336 63 1506
rect 129 1336 159 1506
rect 225 1336 255 1506
rect 321 1336 351 1506
rect 417 1336 447 1506
rect 513 1336 543 1506
rect 609 1336 639 1506
rect 705 1336 735 1506
rect 801 1336 831 1506
rect 897 1336 927 1506
rect -927 930 -897 1100
rect -831 930 -801 1100
rect -735 930 -705 1100
rect -639 930 -609 1100
rect -543 930 -513 1100
rect -447 930 -417 1100
rect -351 930 -321 1100
rect -255 930 -225 1100
rect -159 930 -129 1100
rect -63 930 -33 1100
rect 33 930 63 1100
rect 129 930 159 1100
rect 225 930 255 1100
rect 321 930 351 1100
rect 417 930 447 1100
rect 513 930 543 1100
rect 609 930 639 1100
rect 705 930 735 1100
rect 801 930 831 1100
rect 897 930 927 1100
rect -927 524 -897 694
rect -831 524 -801 694
rect -735 524 -705 694
rect -639 524 -609 694
rect -543 524 -513 694
rect -447 524 -417 694
rect -351 524 -321 694
rect -255 524 -225 694
rect -159 524 -129 694
rect -63 524 -33 694
rect 33 524 63 694
rect 129 524 159 694
rect 225 524 255 694
rect 321 524 351 694
rect 417 524 447 694
rect 513 524 543 694
rect 609 524 639 694
rect 705 524 735 694
rect 801 524 831 694
rect 897 524 927 694
rect -927 118 -897 288
rect -831 118 -801 288
rect -735 118 -705 288
rect -639 118 -609 288
rect -543 118 -513 288
rect -447 118 -417 288
rect -351 118 -321 288
rect -255 118 -225 288
rect -159 118 -129 288
rect -63 118 -33 288
rect 33 118 63 288
rect 129 118 159 288
rect 225 118 255 288
rect 321 118 351 288
rect 417 118 447 288
rect 513 118 543 288
rect 609 118 639 288
rect 705 118 735 288
rect 801 118 831 288
rect 897 118 927 288
rect -927 -288 -897 -118
rect -831 -288 -801 -118
rect -735 -288 -705 -118
rect -639 -288 -609 -118
rect -543 -288 -513 -118
rect -447 -288 -417 -118
rect -351 -288 -321 -118
rect -255 -288 -225 -118
rect -159 -288 -129 -118
rect -63 -288 -33 -118
rect 33 -288 63 -118
rect 129 -288 159 -118
rect 225 -288 255 -118
rect 321 -288 351 -118
rect 417 -288 447 -118
rect 513 -288 543 -118
rect 609 -288 639 -118
rect 705 -288 735 -118
rect 801 -288 831 -118
rect 897 -288 927 -118
rect -927 -694 -897 -524
rect -831 -694 -801 -524
rect -735 -694 -705 -524
rect -639 -694 -609 -524
rect -543 -694 -513 -524
rect -447 -694 -417 -524
rect -351 -694 -321 -524
rect -255 -694 -225 -524
rect -159 -694 -129 -524
rect -63 -694 -33 -524
rect 33 -694 63 -524
rect 129 -694 159 -524
rect 225 -694 255 -524
rect 321 -694 351 -524
rect 417 -694 447 -524
rect 513 -694 543 -524
rect 609 -694 639 -524
rect 705 -694 735 -524
rect 801 -694 831 -524
rect 897 -694 927 -524
rect -927 -1100 -897 -930
rect -831 -1100 -801 -930
rect -735 -1100 -705 -930
rect -639 -1100 -609 -930
rect -543 -1100 -513 -930
rect -447 -1100 -417 -930
rect -351 -1100 -321 -930
rect -255 -1100 -225 -930
rect -159 -1100 -129 -930
rect -63 -1100 -33 -930
rect 33 -1100 63 -930
rect 129 -1100 159 -930
rect 225 -1100 255 -930
rect 321 -1100 351 -930
rect 417 -1100 447 -930
rect 513 -1100 543 -930
rect 609 -1100 639 -930
rect 705 -1100 735 -930
rect 801 -1100 831 -930
rect 897 -1100 927 -930
rect -927 -1506 -897 -1336
rect -831 -1506 -801 -1336
rect -735 -1506 -705 -1336
rect -639 -1506 -609 -1336
rect -543 -1506 -513 -1336
rect -447 -1506 -417 -1336
rect -351 -1506 -321 -1336
rect -255 -1506 -225 -1336
rect -159 -1506 -129 -1336
rect -63 -1506 -33 -1336
rect 33 -1506 63 -1336
rect 129 -1506 159 -1336
rect 225 -1506 255 -1336
rect 321 -1506 351 -1336
rect 417 -1506 447 -1336
rect 513 -1506 543 -1336
rect 609 -1506 639 -1336
rect 705 -1506 735 -1336
rect 801 -1506 831 -1336
rect 897 -1506 927 -1336
rect -927 -1912 -897 -1742
rect -831 -1912 -801 -1742
rect -735 -1912 -705 -1742
rect -639 -1912 -609 -1742
rect -543 -1912 -513 -1742
rect -447 -1912 -417 -1742
rect -351 -1912 -321 -1742
rect -255 -1912 -225 -1742
rect -159 -1912 -129 -1742
rect -63 -1912 -33 -1742
rect 33 -1912 63 -1742
rect 129 -1912 159 -1742
rect 225 -1912 255 -1742
rect 321 -1912 351 -1742
rect 417 -1912 447 -1742
rect 513 -1912 543 -1742
rect 609 -1912 639 -1742
rect 705 -1912 735 -1742
rect 801 -1912 831 -1742
rect 897 -1912 927 -1742
<< pdiff >>
rect -989 1900 -927 1912
rect -989 1754 -977 1900
rect -943 1754 -927 1900
rect -989 1742 -927 1754
rect -897 1900 -831 1912
rect -897 1754 -881 1900
rect -847 1754 -831 1900
rect -897 1742 -831 1754
rect -801 1900 -735 1912
rect -801 1754 -785 1900
rect -751 1754 -735 1900
rect -801 1742 -735 1754
rect -705 1900 -639 1912
rect -705 1754 -689 1900
rect -655 1754 -639 1900
rect -705 1742 -639 1754
rect -609 1900 -543 1912
rect -609 1754 -593 1900
rect -559 1754 -543 1900
rect -609 1742 -543 1754
rect -513 1900 -447 1912
rect -513 1754 -497 1900
rect -463 1754 -447 1900
rect -513 1742 -447 1754
rect -417 1900 -351 1912
rect -417 1754 -401 1900
rect -367 1754 -351 1900
rect -417 1742 -351 1754
rect -321 1900 -255 1912
rect -321 1754 -305 1900
rect -271 1754 -255 1900
rect -321 1742 -255 1754
rect -225 1900 -159 1912
rect -225 1754 -209 1900
rect -175 1754 -159 1900
rect -225 1742 -159 1754
rect -129 1900 -63 1912
rect -129 1754 -113 1900
rect -79 1754 -63 1900
rect -129 1742 -63 1754
rect -33 1900 33 1912
rect -33 1754 -17 1900
rect 17 1754 33 1900
rect -33 1742 33 1754
rect 63 1900 129 1912
rect 63 1754 79 1900
rect 113 1754 129 1900
rect 63 1742 129 1754
rect 159 1900 225 1912
rect 159 1754 175 1900
rect 209 1754 225 1900
rect 159 1742 225 1754
rect 255 1900 321 1912
rect 255 1754 271 1900
rect 305 1754 321 1900
rect 255 1742 321 1754
rect 351 1900 417 1912
rect 351 1754 367 1900
rect 401 1754 417 1900
rect 351 1742 417 1754
rect 447 1900 513 1912
rect 447 1754 463 1900
rect 497 1754 513 1900
rect 447 1742 513 1754
rect 543 1900 609 1912
rect 543 1754 559 1900
rect 593 1754 609 1900
rect 543 1742 609 1754
rect 639 1900 705 1912
rect 639 1754 655 1900
rect 689 1754 705 1900
rect 639 1742 705 1754
rect 735 1900 801 1912
rect 735 1754 751 1900
rect 785 1754 801 1900
rect 735 1742 801 1754
rect 831 1900 897 1912
rect 831 1754 847 1900
rect 881 1754 897 1900
rect 831 1742 897 1754
rect 927 1900 989 1912
rect 927 1754 943 1900
rect 977 1754 989 1900
rect 927 1742 989 1754
rect -989 1494 -927 1506
rect -989 1348 -977 1494
rect -943 1348 -927 1494
rect -989 1336 -927 1348
rect -897 1494 -831 1506
rect -897 1348 -881 1494
rect -847 1348 -831 1494
rect -897 1336 -831 1348
rect -801 1494 -735 1506
rect -801 1348 -785 1494
rect -751 1348 -735 1494
rect -801 1336 -735 1348
rect -705 1494 -639 1506
rect -705 1348 -689 1494
rect -655 1348 -639 1494
rect -705 1336 -639 1348
rect -609 1494 -543 1506
rect -609 1348 -593 1494
rect -559 1348 -543 1494
rect -609 1336 -543 1348
rect -513 1494 -447 1506
rect -513 1348 -497 1494
rect -463 1348 -447 1494
rect -513 1336 -447 1348
rect -417 1494 -351 1506
rect -417 1348 -401 1494
rect -367 1348 -351 1494
rect -417 1336 -351 1348
rect -321 1494 -255 1506
rect -321 1348 -305 1494
rect -271 1348 -255 1494
rect -321 1336 -255 1348
rect -225 1494 -159 1506
rect -225 1348 -209 1494
rect -175 1348 -159 1494
rect -225 1336 -159 1348
rect -129 1494 -63 1506
rect -129 1348 -113 1494
rect -79 1348 -63 1494
rect -129 1336 -63 1348
rect -33 1494 33 1506
rect -33 1348 -17 1494
rect 17 1348 33 1494
rect -33 1336 33 1348
rect 63 1494 129 1506
rect 63 1348 79 1494
rect 113 1348 129 1494
rect 63 1336 129 1348
rect 159 1494 225 1506
rect 159 1348 175 1494
rect 209 1348 225 1494
rect 159 1336 225 1348
rect 255 1494 321 1506
rect 255 1348 271 1494
rect 305 1348 321 1494
rect 255 1336 321 1348
rect 351 1494 417 1506
rect 351 1348 367 1494
rect 401 1348 417 1494
rect 351 1336 417 1348
rect 447 1494 513 1506
rect 447 1348 463 1494
rect 497 1348 513 1494
rect 447 1336 513 1348
rect 543 1494 609 1506
rect 543 1348 559 1494
rect 593 1348 609 1494
rect 543 1336 609 1348
rect 639 1494 705 1506
rect 639 1348 655 1494
rect 689 1348 705 1494
rect 639 1336 705 1348
rect 735 1494 801 1506
rect 735 1348 751 1494
rect 785 1348 801 1494
rect 735 1336 801 1348
rect 831 1494 897 1506
rect 831 1348 847 1494
rect 881 1348 897 1494
rect 831 1336 897 1348
rect 927 1494 989 1506
rect 927 1348 943 1494
rect 977 1348 989 1494
rect 927 1336 989 1348
rect -989 1088 -927 1100
rect -989 942 -977 1088
rect -943 942 -927 1088
rect -989 930 -927 942
rect -897 1088 -831 1100
rect -897 942 -881 1088
rect -847 942 -831 1088
rect -897 930 -831 942
rect -801 1088 -735 1100
rect -801 942 -785 1088
rect -751 942 -735 1088
rect -801 930 -735 942
rect -705 1088 -639 1100
rect -705 942 -689 1088
rect -655 942 -639 1088
rect -705 930 -639 942
rect -609 1088 -543 1100
rect -609 942 -593 1088
rect -559 942 -543 1088
rect -609 930 -543 942
rect -513 1088 -447 1100
rect -513 942 -497 1088
rect -463 942 -447 1088
rect -513 930 -447 942
rect -417 1088 -351 1100
rect -417 942 -401 1088
rect -367 942 -351 1088
rect -417 930 -351 942
rect -321 1088 -255 1100
rect -321 942 -305 1088
rect -271 942 -255 1088
rect -321 930 -255 942
rect -225 1088 -159 1100
rect -225 942 -209 1088
rect -175 942 -159 1088
rect -225 930 -159 942
rect -129 1088 -63 1100
rect -129 942 -113 1088
rect -79 942 -63 1088
rect -129 930 -63 942
rect -33 1088 33 1100
rect -33 942 -17 1088
rect 17 942 33 1088
rect -33 930 33 942
rect 63 1088 129 1100
rect 63 942 79 1088
rect 113 942 129 1088
rect 63 930 129 942
rect 159 1088 225 1100
rect 159 942 175 1088
rect 209 942 225 1088
rect 159 930 225 942
rect 255 1088 321 1100
rect 255 942 271 1088
rect 305 942 321 1088
rect 255 930 321 942
rect 351 1088 417 1100
rect 351 942 367 1088
rect 401 942 417 1088
rect 351 930 417 942
rect 447 1088 513 1100
rect 447 942 463 1088
rect 497 942 513 1088
rect 447 930 513 942
rect 543 1088 609 1100
rect 543 942 559 1088
rect 593 942 609 1088
rect 543 930 609 942
rect 639 1088 705 1100
rect 639 942 655 1088
rect 689 942 705 1088
rect 639 930 705 942
rect 735 1088 801 1100
rect 735 942 751 1088
rect 785 942 801 1088
rect 735 930 801 942
rect 831 1088 897 1100
rect 831 942 847 1088
rect 881 942 897 1088
rect 831 930 897 942
rect 927 1088 989 1100
rect 927 942 943 1088
rect 977 942 989 1088
rect 927 930 989 942
rect -989 682 -927 694
rect -989 536 -977 682
rect -943 536 -927 682
rect -989 524 -927 536
rect -897 682 -831 694
rect -897 536 -881 682
rect -847 536 -831 682
rect -897 524 -831 536
rect -801 682 -735 694
rect -801 536 -785 682
rect -751 536 -735 682
rect -801 524 -735 536
rect -705 682 -639 694
rect -705 536 -689 682
rect -655 536 -639 682
rect -705 524 -639 536
rect -609 682 -543 694
rect -609 536 -593 682
rect -559 536 -543 682
rect -609 524 -543 536
rect -513 682 -447 694
rect -513 536 -497 682
rect -463 536 -447 682
rect -513 524 -447 536
rect -417 682 -351 694
rect -417 536 -401 682
rect -367 536 -351 682
rect -417 524 -351 536
rect -321 682 -255 694
rect -321 536 -305 682
rect -271 536 -255 682
rect -321 524 -255 536
rect -225 682 -159 694
rect -225 536 -209 682
rect -175 536 -159 682
rect -225 524 -159 536
rect -129 682 -63 694
rect -129 536 -113 682
rect -79 536 -63 682
rect -129 524 -63 536
rect -33 682 33 694
rect -33 536 -17 682
rect 17 536 33 682
rect -33 524 33 536
rect 63 682 129 694
rect 63 536 79 682
rect 113 536 129 682
rect 63 524 129 536
rect 159 682 225 694
rect 159 536 175 682
rect 209 536 225 682
rect 159 524 225 536
rect 255 682 321 694
rect 255 536 271 682
rect 305 536 321 682
rect 255 524 321 536
rect 351 682 417 694
rect 351 536 367 682
rect 401 536 417 682
rect 351 524 417 536
rect 447 682 513 694
rect 447 536 463 682
rect 497 536 513 682
rect 447 524 513 536
rect 543 682 609 694
rect 543 536 559 682
rect 593 536 609 682
rect 543 524 609 536
rect 639 682 705 694
rect 639 536 655 682
rect 689 536 705 682
rect 639 524 705 536
rect 735 682 801 694
rect 735 536 751 682
rect 785 536 801 682
rect 735 524 801 536
rect 831 682 897 694
rect 831 536 847 682
rect 881 536 897 682
rect 831 524 897 536
rect 927 682 989 694
rect 927 536 943 682
rect 977 536 989 682
rect 927 524 989 536
rect -989 276 -927 288
rect -989 130 -977 276
rect -943 130 -927 276
rect -989 118 -927 130
rect -897 276 -831 288
rect -897 130 -881 276
rect -847 130 -831 276
rect -897 118 -831 130
rect -801 276 -735 288
rect -801 130 -785 276
rect -751 130 -735 276
rect -801 118 -735 130
rect -705 276 -639 288
rect -705 130 -689 276
rect -655 130 -639 276
rect -705 118 -639 130
rect -609 276 -543 288
rect -609 130 -593 276
rect -559 130 -543 276
rect -609 118 -543 130
rect -513 276 -447 288
rect -513 130 -497 276
rect -463 130 -447 276
rect -513 118 -447 130
rect -417 276 -351 288
rect -417 130 -401 276
rect -367 130 -351 276
rect -417 118 -351 130
rect -321 276 -255 288
rect -321 130 -305 276
rect -271 130 -255 276
rect -321 118 -255 130
rect -225 276 -159 288
rect -225 130 -209 276
rect -175 130 -159 276
rect -225 118 -159 130
rect -129 276 -63 288
rect -129 130 -113 276
rect -79 130 -63 276
rect -129 118 -63 130
rect -33 276 33 288
rect -33 130 -17 276
rect 17 130 33 276
rect -33 118 33 130
rect 63 276 129 288
rect 63 130 79 276
rect 113 130 129 276
rect 63 118 129 130
rect 159 276 225 288
rect 159 130 175 276
rect 209 130 225 276
rect 159 118 225 130
rect 255 276 321 288
rect 255 130 271 276
rect 305 130 321 276
rect 255 118 321 130
rect 351 276 417 288
rect 351 130 367 276
rect 401 130 417 276
rect 351 118 417 130
rect 447 276 513 288
rect 447 130 463 276
rect 497 130 513 276
rect 447 118 513 130
rect 543 276 609 288
rect 543 130 559 276
rect 593 130 609 276
rect 543 118 609 130
rect 639 276 705 288
rect 639 130 655 276
rect 689 130 705 276
rect 639 118 705 130
rect 735 276 801 288
rect 735 130 751 276
rect 785 130 801 276
rect 735 118 801 130
rect 831 276 897 288
rect 831 130 847 276
rect 881 130 897 276
rect 831 118 897 130
rect 927 276 989 288
rect 927 130 943 276
rect 977 130 989 276
rect 927 118 989 130
rect -989 -130 -927 -118
rect -989 -276 -977 -130
rect -943 -276 -927 -130
rect -989 -288 -927 -276
rect -897 -130 -831 -118
rect -897 -276 -881 -130
rect -847 -276 -831 -130
rect -897 -288 -831 -276
rect -801 -130 -735 -118
rect -801 -276 -785 -130
rect -751 -276 -735 -130
rect -801 -288 -735 -276
rect -705 -130 -639 -118
rect -705 -276 -689 -130
rect -655 -276 -639 -130
rect -705 -288 -639 -276
rect -609 -130 -543 -118
rect -609 -276 -593 -130
rect -559 -276 -543 -130
rect -609 -288 -543 -276
rect -513 -130 -447 -118
rect -513 -276 -497 -130
rect -463 -276 -447 -130
rect -513 -288 -447 -276
rect -417 -130 -351 -118
rect -417 -276 -401 -130
rect -367 -276 -351 -130
rect -417 -288 -351 -276
rect -321 -130 -255 -118
rect -321 -276 -305 -130
rect -271 -276 -255 -130
rect -321 -288 -255 -276
rect -225 -130 -159 -118
rect -225 -276 -209 -130
rect -175 -276 -159 -130
rect -225 -288 -159 -276
rect -129 -130 -63 -118
rect -129 -276 -113 -130
rect -79 -276 -63 -130
rect -129 -288 -63 -276
rect -33 -130 33 -118
rect -33 -276 -17 -130
rect 17 -276 33 -130
rect -33 -288 33 -276
rect 63 -130 129 -118
rect 63 -276 79 -130
rect 113 -276 129 -130
rect 63 -288 129 -276
rect 159 -130 225 -118
rect 159 -276 175 -130
rect 209 -276 225 -130
rect 159 -288 225 -276
rect 255 -130 321 -118
rect 255 -276 271 -130
rect 305 -276 321 -130
rect 255 -288 321 -276
rect 351 -130 417 -118
rect 351 -276 367 -130
rect 401 -276 417 -130
rect 351 -288 417 -276
rect 447 -130 513 -118
rect 447 -276 463 -130
rect 497 -276 513 -130
rect 447 -288 513 -276
rect 543 -130 609 -118
rect 543 -276 559 -130
rect 593 -276 609 -130
rect 543 -288 609 -276
rect 639 -130 705 -118
rect 639 -276 655 -130
rect 689 -276 705 -130
rect 639 -288 705 -276
rect 735 -130 801 -118
rect 735 -276 751 -130
rect 785 -276 801 -130
rect 735 -288 801 -276
rect 831 -130 897 -118
rect 831 -276 847 -130
rect 881 -276 897 -130
rect 831 -288 897 -276
rect 927 -130 989 -118
rect 927 -276 943 -130
rect 977 -276 989 -130
rect 927 -288 989 -276
rect -989 -536 -927 -524
rect -989 -682 -977 -536
rect -943 -682 -927 -536
rect -989 -694 -927 -682
rect -897 -536 -831 -524
rect -897 -682 -881 -536
rect -847 -682 -831 -536
rect -897 -694 -831 -682
rect -801 -536 -735 -524
rect -801 -682 -785 -536
rect -751 -682 -735 -536
rect -801 -694 -735 -682
rect -705 -536 -639 -524
rect -705 -682 -689 -536
rect -655 -682 -639 -536
rect -705 -694 -639 -682
rect -609 -536 -543 -524
rect -609 -682 -593 -536
rect -559 -682 -543 -536
rect -609 -694 -543 -682
rect -513 -536 -447 -524
rect -513 -682 -497 -536
rect -463 -682 -447 -536
rect -513 -694 -447 -682
rect -417 -536 -351 -524
rect -417 -682 -401 -536
rect -367 -682 -351 -536
rect -417 -694 -351 -682
rect -321 -536 -255 -524
rect -321 -682 -305 -536
rect -271 -682 -255 -536
rect -321 -694 -255 -682
rect -225 -536 -159 -524
rect -225 -682 -209 -536
rect -175 -682 -159 -536
rect -225 -694 -159 -682
rect -129 -536 -63 -524
rect -129 -682 -113 -536
rect -79 -682 -63 -536
rect -129 -694 -63 -682
rect -33 -536 33 -524
rect -33 -682 -17 -536
rect 17 -682 33 -536
rect -33 -694 33 -682
rect 63 -536 129 -524
rect 63 -682 79 -536
rect 113 -682 129 -536
rect 63 -694 129 -682
rect 159 -536 225 -524
rect 159 -682 175 -536
rect 209 -682 225 -536
rect 159 -694 225 -682
rect 255 -536 321 -524
rect 255 -682 271 -536
rect 305 -682 321 -536
rect 255 -694 321 -682
rect 351 -536 417 -524
rect 351 -682 367 -536
rect 401 -682 417 -536
rect 351 -694 417 -682
rect 447 -536 513 -524
rect 447 -682 463 -536
rect 497 -682 513 -536
rect 447 -694 513 -682
rect 543 -536 609 -524
rect 543 -682 559 -536
rect 593 -682 609 -536
rect 543 -694 609 -682
rect 639 -536 705 -524
rect 639 -682 655 -536
rect 689 -682 705 -536
rect 639 -694 705 -682
rect 735 -536 801 -524
rect 735 -682 751 -536
rect 785 -682 801 -536
rect 735 -694 801 -682
rect 831 -536 897 -524
rect 831 -682 847 -536
rect 881 -682 897 -536
rect 831 -694 897 -682
rect 927 -536 989 -524
rect 927 -682 943 -536
rect 977 -682 989 -536
rect 927 -694 989 -682
rect -989 -942 -927 -930
rect -989 -1088 -977 -942
rect -943 -1088 -927 -942
rect -989 -1100 -927 -1088
rect -897 -942 -831 -930
rect -897 -1088 -881 -942
rect -847 -1088 -831 -942
rect -897 -1100 -831 -1088
rect -801 -942 -735 -930
rect -801 -1088 -785 -942
rect -751 -1088 -735 -942
rect -801 -1100 -735 -1088
rect -705 -942 -639 -930
rect -705 -1088 -689 -942
rect -655 -1088 -639 -942
rect -705 -1100 -639 -1088
rect -609 -942 -543 -930
rect -609 -1088 -593 -942
rect -559 -1088 -543 -942
rect -609 -1100 -543 -1088
rect -513 -942 -447 -930
rect -513 -1088 -497 -942
rect -463 -1088 -447 -942
rect -513 -1100 -447 -1088
rect -417 -942 -351 -930
rect -417 -1088 -401 -942
rect -367 -1088 -351 -942
rect -417 -1100 -351 -1088
rect -321 -942 -255 -930
rect -321 -1088 -305 -942
rect -271 -1088 -255 -942
rect -321 -1100 -255 -1088
rect -225 -942 -159 -930
rect -225 -1088 -209 -942
rect -175 -1088 -159 -942
rect -225 -1100 -159 -1088
rect -129 -942 -63 -930
rect -129 -1088 -113 -942
rect -79 -1088 -63 -942
rect -129 -1100 -63 -1088
rect -33 -942 33 -930
rect -33 -1088 -17 -942
rect 17 -1088 33 -942
rect -33 -1100 33 -1088
rect 63 -942 129 -930
rect 63 -1088 79 -942
rect 113 -1088 129 -942
rect 63 -1100 129 -1088
rect 159 -942 225 -930
rect 159 -1088 175 -942
rect 209 -1088 225 -942
rect 159 -1100 225 -1088
rect 255 -942 321 -930
rect 255 -1088 271 -942
rect 305 -1088 321 -942
rect 255 -1100 321 -1088
rect 351 -942 417 -930
rect 351 -1088 367 -942
rect 401 -1088 417 -942
rect 351 -1100 417 -1088
rect 447 -942 513 -930
rect 447 -1088 463 -942
rect 497 -1088 513 -942
rect 447 -1100 513 -1088
rect 543 -942 609 -930
rect 543 -1088 559 -942
rect 593 -1088 609 -942
rect 543 -1100 609 -1088
rect 639 -942 705 -930
rect 639 -1088 655 -942
rect 689 -1088 705 -942
rect 639 -1100 705 -1088
rect 735 -942 801 -930
rect 735 -1088 751 -942
rect 785 -1088 801 -942
rect 735 -1100 801 -1088
rect 831 -942 897 -930
rect 831 -1088 847 -942
rect 881 -1088 897 -942
rect 831 -1100 897 -1088
rect 927 -942 989 -930
rect 927 -1088 943 -942
rect 977 -1088 989 -942
rect 927 -1100 989 -1088
rect -989 -1348 -927 -1336
rect -989 -1494 -977 -1348
rect -943 -1494 -927 -1348
rect -989 -1506 -927 -1494
rect -897 -1348 -831 -1336
rect -897 -1494 -881 -1348
rect -847 -1494 -831 -1348
rect -897 -1506 -831 -1494
rect -801 -1348 -735 -1336
rect -801 -1494 -785 -1348
rect -751 -1494 -735 -1348
rect -801 -1506 -735 -1494
rect -705 -1348 -639 -1336
rect -705 -1494 -689 -1348
rect -655 -1494 -639 -1348
rect -705 -1506 -639 -1494
rect -609 -1348 -543 -1336
rect -609 -1494 -593 -1348
rect -559 -1494 -543 -1348
rect -609 -1506 -543 -1494
rect -513 -1348 -447 -1336
rect -513 -1494 -497 -1348
rect -463 -1494 -447 -1348
rect -513 -1506 -447 -1494
rect -417 -1348 -351 -1336
rect -417 -1494 -401 -1348
rect -367 -1494 -351 -1348
rect -417 -1506 -351 -1494
rect -321 -1348 -255 -1336
rect -321 -1494 -305 -1348
rect -271 -1494 -255 -1348
rect -321 -1506 -255 -1494
rect -225 -1348 -159 -1336
rect -225 -1494 -209 -1348
rect -175 -1494 -159 -1348
rect -225 -1506 -159 -1494
rect -129 -1348 -63 -1336
rect -129 -1494 -113 -1348
rect -79 -1494 -63 -1348
rect -129 -1506 -63 -1494
rect -33 -1348 33 -1336
rect -33 -1494 -17 -1348
rect 17 -1494 33 -1348
rect -33 -1506 33 -1494
rect 63 -1348 129 -1336
rect 63 -1494 79 -1348
rect 113 -1494 129 -1348
rect 63 -1506 129 -1494
rect 159 -1348 225 -1336
rect 159 -1494 175 -1348
rect 209 -1494 225 -1348
rect 159 -1506 225 -1494
rect 255 -1348 321 -1336
rect 255 -1494 271 -1348
rect 305 -1494 321 -1348
rect 255 -1506 321 -1494
rect 351 -1348 417 -1336
rect 351 -1494 367 -1348
rect 401 -1494 417 -1348
rect 351 -1506 417 -1494
rect 447 -1348 513 -1336
rect 447 -1494 463 -1348
rect 497 -1494 513 -1348
rect 447 -1506 513 -1494
rect 543 -1348 609 -1336
rect 543 -1494 559 -1348
rect 593 -1494 609 -1348
rect 543 -1506 609 -1494
rect 639 -1348 705 -1336
rect 639 -1494 655 -1348
rect 689 -1494 705 -1348
rect 639 -1506 705 -1494
rect 735 -1348 801 -1336
rect 735 -1494 751 -1348
rect 785 -1494 801 -1348
rect 735 -1506 801 -1494
rect 831 -1348 897 -1336
rect 831 -1494 847 -1348
rect 881 -1494 897 -1348
rect 831 -1506 897 -1494
rect 927 -1348 989 -1336
rect 927 -1494 943 -1348
rect 977 -1494 989 -1348
rect 927 -1506 989 -1494
rect -989 -1754 -927 -1742
rect -989 -1900 -977 -1754
rect -943 -1900 -927 -1754
rect -989 -1912 -927 -1900
rect -897 -1754 -831 -1742
rect -897 -1900 -881 -1754
rect -847 -1900 -831 -1754
rect -897 -1912 -831 -1900
rect -801 -1754 -735 -1742
rect -801 -1900 -785 -1754
rect -751 -1900 -735 -1754
rect -801 -1912 -735 -1900
rect -705 -1754 -639 -1742
rect -705 -1900 -689 -1754
rect -655 -1900 -639 -1754
rect -705 -1912 -639 -1900
rect -609 -1754 -543 -1742
rect -609 -1900 -593 -1754
rect -559 -1900 -543 -1754
rect -609 -1912 -543 -1900
rect -513 -1754 -447 -1742
rect -513 -1900 -497 -1754
rect -463 -1900 -447 -1754
rect -513 -1912 -447 -1900
rect -417 -1754 -351 -1742
rect -417 -1900 -401 -1754
rect -367 -1900 -351 -1754
rect -417 -1912 -351 -1900
rect -321 -1754 -255 -1742
rect -321 -1900 -305 -1754
rect -271 -1900 -255 -1754
rect -321 -1912 -255 -1900
rect -225 -1754 -159 -1742
rect -225 -1900 -209 -1754
rect -175 -1900 -159 -1754
rect -225 -1912 -159 -1900
rect -129 -1754 -63 -1742
rect -129 -1900 -113 -1754
rect -79 -1900 -63 -1754
rect -129 -1912 -63 -1900
rect -33 -1754 33 -1742
rect -33 -1900 -17 -1754
rect 17 -1900 33 -1754
rect -33 -1912 33 -1900
rect 63 -1754 129 -1742
rect 63 -1900 79 -1754
rect 113 -1900 129 -1754
rect 63 -1912 129 -1900
rect 159 -1754 225 -1742
rect 159 -1900 175 -1754
rect 209 -1900 225 -1754
rect 159 -1912 225 -1900
rect 255 -1754 321 -1742
rect 255 -1900 271 -1754
rect 305 -1900 321 -1754
rect 255 -1912 321 -1900
rect 351 -1754 417 -1742
rect 351 -1900 367 -1754
rect 401 -1900 417 -1754
rect 351 -1912 417 -1900
rect 447 -1754 513 -1742
rect 447 -1900 463 -1754
rect 497 -1900 513 -1754
rect 447 -1912 513 -1900
rect 543 -1754 609 -1742
rect 543 -1900 559 -1754
rect 593 -1900 609 -1754
rect 543 -1912 609 -1900
rect 639 -1754 705 -1742
rect 639 -1900 655 -1754
rect 689 -1900 705 -1754
rect 639 -1912 705 -1900
rect 735 -1754 801 -1742
rect 735 -1900 751 -1754
rect 785 -1900 801 -1754
rect 735 -1912 801 -1900
rect 831 -1754 897 -1742
rect 831 -1900 847 -1754
rect 881 -1900 897 -1754
rect 831 -1912 897 -1900
rect 927 -1754 989 -1742
rect 927 -1900 943 -1754
rect 977 -1900 989 -1754
rect 927 -1912 989 -1900
<< pdiffc >>
rect -977 1754 -943 1900
rect -881 1754 -847 1900
rect -785 1754 -751 1900
rect -689 1754 -655 1900
rect -593 1754 -559 1900
rect -497 1754 -463 1900
rect -401 1754 -367 1900
rect -305 1754 -271 1900
rect -209 1754 -175 1900
rect -113 1754 -79 1900
rect -17 1754 17 1900
rect 79 1754 113 1900
rect 175 1754 209 1900
rect 271 1754 305 1900
rect 367 1754 401 1900
rect 463 1754 497 1900
rect 559 1754 593 1900
rect 655 1754 689 1900
rect 751 1754 785 1900
rect 847 1754 881 1900
rect 943 1754 977 1900
rect -977 1348 -943 1494
rect -881 1348 -847 1494
rect -785 1348 -751 1494
rect -689 1348 -655 1494
rect -593 1348 -559 1494
rect -497 1348 -463 1494
rect -401 1348 -367 1494
rect -305 1348 -271 1494
rect -209 1348 -175 1494
rect -113 1348 -79 1494
rect -17 1348 17 1494
rect 79 1348 113 1494
rect 175 1348 209 1494
rect 271 1348 305 1494
rect 367 1348 401 1494
rect 463 1348 497 1494
rect 559 1348 593 1494
rect 655 1348 689 1494
rect 751 1348 785 1494
rect 847 1348 881 1494
rect 943 1348 977 1494
rect -977 942 -943 1088
rect -881 942 -847 1088
rect -785 942 -751 1088
rect -689 942 -655 1088
rect -593 942 -559 1088
rect -497 942 -463 1088
rect -401 942 -367 1088
rect -305 942 -271 1088
rect -209 942 -175 1088
rect -113 942 -79 1088
rect -17 942 17 1088
rect 79 942 113 1088
rect 175 942 209 1088
rect 271 942 305 1088
rect 367 942 401 1088
rect 463 942 497 1088
rect 559 942 593 1088
rect 655 942 689 1088
rect 751 942 785 1088
rect 847 942 881 1088
rect 943 942 977 1088
rect -977 536 -943 682
rect -881 536 -847 682
rect -785 536 -751 682
rect -689 536 -655 682
rect -593 536 -559 682
rect -497 536 -463 682
rect -401 536 -367 682
rect -305 536 -271 682
rect -209 536 -175 682
rect -113 536 -79 682
rect -17 536 17 682
rect 79 536 113 682
rect 175 536 209 682
rect 271 536 305 682
rect 367 536 401 682
rect 463 536 497 682
rect 559 536 593 682
rect 655 536 689 682
rect 751 536 785 682
rect 847 536 881 682
rect 943 536 977 682
rect -977 130 -943 276
rect -881 130 -847 276
rect -785 130 -751 276
rect -689 130 -655 276
rect -593 130 -559 276
rect -497 130 -463 276
rect -401 130 -367 276
rect -305 130 -271 276
rect -209 130 -175 276
rect -113 130 -79 276
rect -17 130 17 276
rect 79 130 113 276
rect 175 130 209 276
rect 271 130 305 276
rect 367 130 401 276
rect 463 130 497 276
rect 559 130 593 276
rect 655 130 689 276
rect 751 130 785 276
rect 847 130 881 276
rect 943 130 977 276
rect -977 -276 -943 -130
rect -881 -276 -847 -130
rect -785 -276 -751 -130
rect -689 -276 -655 -130
rect -593 -276 -559 -130
rect -497 -276 -463 -130
rect -401 -276 -367 -130
rect -305 -276 -271 -130
rect -209 -276 -175 -130
rect -113 -276 -79 -130
rect -17 -276 17 -130
rect 79 -276 113 -130
rect 175 -276 209 -130
rect 271 -276 305 -130
rect 367 -276 401 -130
rect 463 -276 497 -130
rect 559 -276 593 -130
rect 655 -276 689 -130
rect 751 -276 785 -130
rect 847 -276 881 -130
rect 943 -276 977 -130
rect -977 -682 -943 -536
rect -881 -682 -847 -536
rect -785 -682 -751 -536
rect -689 -682 -655 -536
rect -593 -682 -559 -536
rect -497 -682 -463 -536
rect -401 -682 -367 -536
rect -305 -682 -271 -536
rect -209 -682 -175 -536
rect -113 -682 -79 -536
rect -17 -682 17 -536
rect 79 -682 113 -536
rect 175 -682 209 -536
rect 271 -682 305 -536
rect 367 -682 401 -536
rect 463 -682 497 -536
rect 559 -682 593 -536
rect 655 -682 689 -536
rect 751 -682 785 -536
rect 847 -682 881 -536
rect 943 -682 977 -536
rect -977 -1088 -943 -942
rect -881 -1088 -847 -942
rect -785 -1088 -751 -942
rect -689 -1088 -655 -942
rect -593 -1088 -559 -942
rect -497 -1088 -463 -942
rect -401 -1088 -367 -942
rect -305 -1088 -271 -942
rect -209 -1088 -175 -942
rect -113 -1088 -79 -942
rect -17 -1088 17 -942
rect 79 -1088 113 -942
rect 175 -1088 209 -942
rect 271 -1088 305 -942
rect 367 -1088 401 -942
rect 463 -1088 497 -942
rect 559 -1088 593 -942
rect 655 -1088 689 -942
rect 751 -1088 785 -942
rect 847 -1088 881 -942
rect 943 -1088 977 -942
rect -977 -1494 -943 -1348
rect -881 -1494 -847 -1348
rect -785 -1494 -751 -1348
rect -689 -1494 -655 -1348
rect -593 -1494 -559 -1348
rect -497 -1494 -463 -1348
rect -401 -1494 -367 -1348
rect -305 -1494 -271 -1348
rect -209 -1494 -175 -1348
rect -113 -1494 -79 -1348
rect -17 -1494 17 -1348
rect 79 -1494 113 -1348
rect 175 -1494 209 -1348
rect 271 -1494 305 -1348
rect 367 -1494 401 -1348
rect 463 -1494 497 -1348
rect 559 -1494 593 -1348
rect 655 -1494 689 -1348
rect 751 -1494 785 -1348
rect 847 -1494 881 -1348
rect 943 -1494 977 -1348
rect -977 -1900 -943 -1754
rect -881 -1900 -847 -1754
rect -785 -1900 -751 -1754
rect -689 -1900 -655 -1754
rect -593 -1900 -559 -1754
rect -497 -1900 -463 -1754
rect -401 -1900 -367 -1754
rect -305 -1900 -271 -1754
rect -209 -1900 -175 -1754
rect -113 -1900 -79 -1754
rect -17 -1900 17 -1754
rect 79 -1900 113 -1754
rect 175 -1900 209 -1754
rect 271 -1900 305 -1754
rect 367 -1900 401 -1754
rect 463 -1900 497 -1754
rect 559 -1900 593 -1754
rect 655 -1900 689 -1754
rect 751 -1900 785 -1754
rect 847 -1900 881 -1754
rect 943 -1900 977 -1754
<< nsubdiff >>
rect -1091 2061 -995 2095
rect 995 2061 1091 2095
rect -1091 1999 -1057 2061
rect 1057 1999 1091 2061
rect -1091 -2061 -1057 -1999
rect 1057 -2061 1091 -1999
rect -1091 -2095 -995 -2061
rect 995 -2095 1091 -2061
<< nsubdiffcont >>
rect -995 2061 995 2095
rect -1091 -1999 -1057 1999
rect 1057 -1999 1091 1999
rect -995 -2095 995 -2061
<< poly >>
rect -945 1993 -879 2009
rect -945 1959 -929 1993
rect -895 1959 -879 1993
rect -945 1943 -879 1959
rect -753 1993 -687 2009
rect -753 1959 -737 1993
rect -703 1959 -687 1993
rect -753 1943 -687 1959
rect -561 1993 -495 2009
rect -561 1959 -545 1993
rect -511 1959 -495 1993
rect -561 1943 -495 1959
rect -369 1993 -303 2009
rect -369 1959 -353 1993
rect -319 1959 -303 1993
rect -369 1943 -303 1959
rect -177 1993 -111 2009
rect -177 1959 -161 1993
rect -127 1959 -111 1993
rect -177 1943 -111 1959
rect 15 1993 81 2009
rect 15 1959 31 1993
rect 65 1959 81 1993
rect 15 1943 81 1959
rect 207 1993 273 2009
rect 207 1959 223 1993
rect 257 1959 273 1993
rect 207 1943 273 1959
rect 399 1993 465 2009
rect 399 1959 415 1993
rect 449 1959 465 1993
rect 399 1943 465 1959
rect 591 1993 657 2009
rect 591 1959 607 1993
rect 641 1959 657 1993
rect 591 1943 657 1959
rect 783 1993 849 2009
rect 783 1959 799 1993
rect 833 1959 849 1993
rect 783 1943 849 1959
rect -927 1912 -897 1943
rect -831 1912 -801 1938
rect -735 1912 -705 1943
rect -639 1912 -609 1938
rect -543 1912 -513 1943
rect -447 1912 -417 1938
rect -351 1912 -321 1943
rect -255 1912 -225 1938
rect -159 1912 -129 1943
rect -63 1912 -33 1938
rect 33 1912 63 1943
rect 129 1912 159 1938
rect 225 1912 255 1943
rect 321 1912 351 1938
rect 417 1912 447 1943
rect 513 1912 543 1938
rect 609 1912 639 1943
rect 705 1912 735 1938
rect 801 1912 831 1943
rect 897 1912 927 1938
rect -927 1716 -897 1742
rect -831 1711 -801 1742
rect -735 1716 -705 1742
rect -639 1711 -609 1742
rect -543 1716 -513 1742
rect -447 1711 -417 1742
rect -351 1716 -321 1742
rect -255 1711 -225 1742
rect -159 1716 -129 1742
rect -63 1711 -33 1742
rect 33 1716 63 1742
rect 129 1711 159 1742
rect 225 1716 255 1742
rect 321 1711 351 1742
rect 417 1716 447 1742
rect 513 1711 543 1742
rect 609 1716 639 1742
rect 705 1711 735 1742
rect 801 1716 831 1742
rect 897 1711 927 1742
rect -849 1695 -783 1711
rect -849 1661 -833 1695
rect -799 1661 -783 1695
rect -849 1645 -783 1661
rect -657 1695 -591 1711
rect -657 1661 -641 1695
rect -607 1661 -591 1695
rect -657 1645 -591 1661
rect -465 1695 -399 1711
rect -465 1661 -449 1695
rect -415 1661 -399 1695
rect -465 1645 -399 1661
rect -273 1695 -207 1711
rect -273 1661 -257 1695
rect -223 1661 -207 1695
rect -273 1645 -207 1661
rect -81 1695 -15 1711
rect -81 1661 -65 1695
rect -31 1661 -15 1695
rect -81 1645 -15 1661
rect 111 1695 177 1711
rect 111 1661 127 1695
rect 161 1661 177 1695
rect 111 1645 177 1661
rect 303 1695 369 1711
rect 303 1661 319 1695
rect 353 1661 369 1695
rect 303 1645 369 1661
rect 495 1695 561 1711
rect 495 1661 511 1695
rect 545 1661 561 1695
rect 495 1645 561 1661
rect 687 1695 753 1711
rect 687 1661 703 1695
rect 737 1661 753 1695
rect 687 1645 753 1661
rect 879 1695 945 1711
rect 879 1661 895 1695
rect 929 1661 945 1695
rect 879 1645 945 1661
rect -849 1587 -783 1603
rect -849 1553 -833 1587
rect -799 1553 -783 1587
rect -849 1537 -783 1553
rect -657 1587 -591 1603
rect -657 1553 -641 1587
rect -607 1553 -591 1587
rect -657 1537 -591 1553
rect -465 1587 -399 1603
rect -465 1553 -449 1587
rect -415 1553 -399 1587
rect -465 1537 -399 1553
rect -273 1587 -207 1603
rect -273 1553 -257 1587
rect -223 1553 -207 1587
rect -273 1537 -207 1553
rect -81 1587 -15 1603
rect -81 1553 -65 1587
rect -31 1553 -15 1587
rect -81 1537 -15 1553
rect 111 1587 177 1603
rect 111 1553 127 1587
rect 161 1553 177 1587
rect 111 1537 177 1553
rect 303 1587 369 1603
rect 303 1553 319 1587
rect 353 1553 369 1587
rect 303 1537 369 1553
rect 495 1587 561 1603
rect 495 1553 511 1587
rect 545 1553 561 1587
rect 495 1537 561 1553
rect 687 1587 753 1603
rect 687 1553 703 1587
rect 737 1553 753 1587
rect 687 1537 753 1553
rect 879 1587 945 1603
rect 879 1553 895 1587
rect 929 1553 945 1587
rect 879 1537 945 1553
rect -927 1506 -897 1532
rect -831 1506 -801 1537
rect -735 1506 -705 1532
rect -639 1506 -609 1537
rect -543 1506 -513 1532
rect -447 1506 -417 1537
rect -351 1506 -321 1532
rect -255 1506 -225 1537
rect -159 1506 -129 1532
rect -63 1506 -33 1537
rect 33 1506 63 1532
rect 129 1506 159 1537
rect 225 1506 255 1532
rect 321 1506 351 1537
rect 417 1506 447 1532
rect 513 1506 543 1537
rect 609 1506 639 1532
rect 705 1506 735 1537
rect 801 1506 831 1532
rect 897 1506 927 1537
rect -927 1305 -897 1336
rect -831 1310 -801 1336
rect -735 1305 -705 1336
rect -639 1310 -609 1336
rect -543 1305 -513 1336
rect -447 1310 -417 1336
rect -351 1305 -321 1336
rect -255 1310 -225 1336
rect -159 1305 -129 1336
rect -63 1310 -33 1336
rect 33 1305 63 1336
rect 129 1310 159 1336
rect 225 1305 255 1336
rect 321 1310 351 1336
rect 417 1305 447 1336
rect 513 1310 543 1336
rect 609 1305 639 1336
rect 705 1310 735 1336
rect 801 1305 831 1336
rect 897 1310 927 1336
rect -945 1289 -879 1305
rect -945 1255 -929 1289
rect -895 1255 -879 1289
rect -945 1239 -879 1255
rect -753 1289 -687 1305
rect -753 1255 -737 1289
rect -703 1255 -687 1289
rect -753 1239 -687 1255
rect -561 1289 -495 1305
rect -561 1255 -545 1289
rect -511 1255 -495 1289
rect -561 1239 -495 1255
rect -369 1289 -303 1305
rect -369 1255 -353 1289
rect -319 1255 -303 1289
rect -369 1239 -303 1255
rect -177 1289 -111 1305
rect -177 1255 -161 1289
rect -127 1255 -111 1289
rect -177 1239 -111 1255
rect 15 1289 81 1305
rect 15 1255 31 1289
rect 65 1255 81 1289
rect 15 1239 81 1255
rect 207 1289 273 1305
rect 207 1255 223 1289
rect 257 1255 273 1289
rect 207 1239 273 1255
rect 399 1289 465 1305
rect 399 1255 415 1289
rect 449 1255 465 1289
rect 399 1239 465 1255
rect 591 1289 657 1305
rect 591 1255 607 1289
rect 641 1255 657 1289
rect 591 1239 657 1255
rect 783 1289 849 1305
rect 783 1255 799 1289
rect 833 1255 849 1289
rect 783 1239 849 1255
rect -945 1181 -879 1197
rect -945 1147 -929 1181
rect -895 1147 -879 1181
rect -945 1131 -879 1147
rect -753 1181 -687 1197
rect -753 1147 -737 1181
rect -703 1147 -687 1181
rect -753 1131 -687 1147
rect -561 1181 -495 1197
rect -561 1147 -545 1181
rect -511 1147 -495 1181
rect -561 1131 -495 1147
rect -369 1181 -303 1197
rect -369 1147 -353 1181
rect -319 1147 -303 1181
rect -369 1131 -303 1147
rect -177 1181 -111 1197
rect -177 1147 -161 1181
rect -127 1147 -111 1181
rect -177 1131 -111 1147
rect 15 1181 81 1197
rect 15 1147 31 1181
rect 65 1147 81 1181
rect 15 1131 81 1147
rect 207 1181 273 1197
rect 207 1147 223 1181
rect 257 1147 273 1181
rect 207 1131 273 1147
rect 399 1181 465 1197
rect 399 1147 415 1181
rect 449 1147 465 1181
rect 399 1131 465 1147
rect 591 1181 657 1197
rect 591 1147 607 1181
rect 641 1147 657 1181
rect 591 1131 657 1147
rect 783 1181 849 1197
rect 783 1147 799 1181
rect 833 1147 849 1181
rect 783 1131 849 1147
rect -927 1100 -897 1131
rect -831 1100 -801 1126
rect -735 1100 -705 1131
rect -639 1100 -609 1126
rect -543 1100 -513 1131
rect -447 1100 -417 1126
rect -351 1100 -321 1131
rect -255 1100 -225 1126
rect -159 1100 -129 1131
rect -63 1100 -33 1126
rect 33 1100 63 1131
rect 129 1100 159 1126
rect 225 1100 255 1131
rect 321 1100 351 1126
rect 417 1100 447 1131
rect 513 1100 543 1126
rect 609 1100 639 1131
rect 705 1100 735 1126
rect 801 1100 831 1131
rect 897 1100 927 1126
rect -927 904 -897 930
rect -831 899 -801 930
rect -735 904 -705 930
rect -639 899 -609 930
rect -543 904 -513 930
rect -447 899 -417 930
rect -351 904 -321 930
rect -255 899 -225 930
rect -159 904 -129 930
rect -63 899 -33 930
rect 33 904 63 930
rect 129 899 159 930
rect 225 904 255 930
rect 321 899 351 930
rect 417 904 447 930
rect 513 899 543 930
rect 609 904 639 930
rect 705 899 735 930
rect 801 904 831 930
rect 897 899 927 930
rect -849 883 -783 899
rect -849 849 -833 883
rect -799 849 -783 883
rect -849 833 -783 849
rect -657 883 -591 899
rect -657 849 -641 883
rect -607 849 -591 883
rect -657 833 -591 849
rect -465 883 -399 899
rect -465 849 -449 883
rect -415 849 -399 883
rect -465 833 -399 849
rect -273 883 -207 899
rect -273 849 -257 883
rect -223 849 -207 883
rect -273 833 -207 849
rect -81 883 -15 899
rect -81 849 -65 883
rect -31 849 -15 883
rect -81 833 -15 849
rect 111 883 177 899
rect 111 849 127 883
rect 161 849 177 883
rect 111 833 177 849
rect 303 883 369 899
rect 303 849 319 883
rect 353 849 369 883
rect 303 833 369 849
rect 495 883 561 899
rect 495 849 511 883
rect 545 849 561 883
rect 495 833 561 849
rect 687 883 753 899
rect 687 849 703 883
rect 737 849 753 883
rect 687 833 753 849
rect 879 883 945 899
rect 879 849 895 883
rect 929 849 945 883
rect 879 833 945 849
rect -849 775 -783 791
rect -849 741 -833 775
rect -799 741 -783 775
rect -849 725 -783 741
rect -657 775 -591 791
rect -657 741 -641 775
rect -607 741 -591 775
rect -657 725 -591 741
rect -465 775 -399 791
rect -465 741 -449 775
rect -415 741 -399 775
rect -465 725 -399 741
rect -273 775 -207 791
rect -273 741 -257 775
rect -223 741 -207 775
rect -273 725 -207 741
rect -81 775 -15 791
rect -81 741 -65 775
rect -31 741 -15 775
rect -81 725 -15 741
rect 111 775 177 791
rect 111 741 127 775
rect 161 741 177 775
rect 111 725 177 741
rect 303 775 369 791
rect 303 741 319 775
rect 353 741 369 775
rect 303 725 369 741
rect 495 775 561 791
rect 495 741 511 775
rect 545 741 561 775
rect 495 725 561 741
rect 687 775 753 791
rect 687 741 703 775
rect 737 741 753 775
rect 687 725 753 741
rect 879 775 945 791
rect 879 741 895 775
rect 929 741 945 775
rect 879 725 945 741
rect -927 694 -897 720
rect -831 694 -801 725
rect -735 694 -705 720
rect -639 694 -609 725
rect -543 694 -513 720
rect -447 694 -417 725
rect -351 694 -321 720
rect -255 694 -225 725
rect -159 694 -129 720
rect -63 694 -33 725
rect 33 694 63 720
rect 129 694 159 725
rect 225 694 255 720
rect 321 694 351 725
rect 417 694 447 720
rect 513 694 543 725
rect 609 694 639 720
rect 705 694 735 725
rect 801 694 831 720
rect 897 694 927 725
rect -927 493 -897 524
rect -831 498 -801 524
rect -735 493 -705 524
rect -639 498 -609 524
rect -543 493 -513 524
rect -447 498 -417 524
rect -351 493 -321 524
rect -255 498 -225 524
rect -159 493 -129 524
rect -63 498 -33 524
rect 33 493 63 524
rect 129 498 159 524
rect 225 493 255 524
rect 321 498 351 524
rect 417 493 447 524
rect 513 498 543 524
rect 609 493 639 524
rect 705 498 735 524
rect 801 493 831 524
rect 897 498 927 524
rect -945 477 -879 493
rect -945 443 -929 477
rect -895 443 -879 477
rect -945 427 -879 443
rect -753 477 -687 493
rect -753 443 -737 477
rect -703 443 -687 477
rect -753 427 -687 443
rect -561 477 -495 493
rect -561 443 -545 477
rect -511 443 -495 477
rect -561 427 -495 443
rect -369 477 -303 493
rect -369 443 -353 477
rect -319 443 -303 477
rect -369 427 -303 443
rect -177 477 -111 493
rect -177 443 -161 477
rect -127 443 -111 477
rect -177 427 -111 443
rect 15 477 81 493
rect 15 443 31 477
rect 65 443 81 477
rect 15 427 81 443
rect 207 477 273 493
rect 207 443 223 477
rect 257 443 273 477
rect 207 427 273 443
rect 399 477 465 493
rect 399 443 415 477
rect 449 443 465 477
rect 399 427 465 443
rect 591 477 657 493
rect 591 443 607 477
rect 641 443 657 477
rect 591 427 657 443
rect 783 477 849 493
rect 783 443 799 477
rect 833 443 849 477
rect 783 427 849 443
rect -945 369 -879 385
rect -945 335 -929 369
rect -895 335 -879 369
rect -945 319 -879 335
rect -753 369 -687 385
rect -753 335 -737 369
rect -703 335 -687 369
rect -753 319 -687 335
rect -561 369 -495 385
rect -561 335 -545 369
rect -511 335 -495 369
rect -561 319 -495 335
rect -369 369 -303 385
rect -369 335 -353 369
rect -319 335 -303 369
rect -369 319 -303 335
rect -177 369 -111 385
rect -177 335 -161 369
rect -127 335 -111 369
rect -177 319 -111 335
rect 15 369 81 385
rect 15 335 31 369
rect 65 335 81 369
rect 15 319 81 335
rect 207 369 273 385
rect 207 335 223 369
rect 257 335 273 369
rect 207 319 273 335
rect 399 369 465 385
rect 399 335 415 369
rect 449 335 465 369
rect 399 319 465 335
rect 591 369 657 385
rect 591 335 607 369
rect 641 335 657 369
rect 591 319 657 335
rect 783 369 849 385
rect 783 335 799 369
rect 833 335 849 369
rect 783 319 849 335
rect -927 288 -897 319
rect -831 288 -801 314
rect -735 288 -705 319
rect -639 288 -609 314
rect -543 288 -513 319
rect -447 288 -417 314
rect -351 288 -321 319
rect -255 288 -225 314
rect -159 288 -129 319
rect -63 288 -33 314
rect 33 288 63 319
rect 129 288 159 314
rect 225 288 255 319
rect 321 288 351 314
rect 417 288 447 319
rect 513 288 543 314
rect 609 288 639 319
rect 705 288 735 314
rect 801 288 831 319
rect 897 288 927 314
rect -927 92 -897 118
rect -831 87 -801 118
rect -735 92 -705 118
rect -639 87 -609 118
rect -543 92 -513 118
rect -447 87 -417 118
rect -351 92 -321 118
rect -255 87 -225 118
rect -159 92 -129 118
rect -63 87 -33 118
rect 33 92 63 118
rect 129 87 159 118
rect 225 92 255 118
rect 321 87 351 118
rect 417 92 447 118
rect 513 87 543 118
rect 609 92 639 118
rect 705 87 735 118
rect 801 92 831 118
rect 897 87 927 118
rect -849 71 -783 87
rect -849 37 -833 71
rect -799 37 -783 71
rect -849 21 -783 37
rect -657 71 -591 87
rect -657 37 -641 71
rect -607 37 -591 71
rect -657 21 -591 37
rect -465 71 -399 87
rect -465 37 -449 71
rect -415 37 -399 71
rect -465 21 -399 37
rect -273 71 -207 87
rect -273 37 -257 71
rect -223 37 -207 71
rect -273 21 -207 37
rect -81 71 -15 87
rect -81 37 -65 71
rect -31 37 -15 71
rect -81 21 -15 37
rect 111 71 177 87
rect 111 37 127 71
rect 161 37 177 71
rect 111 21 177 37
rect 303 71 369 87
rect 303 37 319 71
rect 353 37 369 71
rect 303 21 369 37
rect 495 71 561 87
rect 495 37 511 71
rect 545 37 561 71
rect 495 21 561 37
rect 687 71 753 87
rect 687 37 703 71
rect 737 37 753 71
rect 687 21 753 37
rect 879 71 945 87
rect 879 37 895 71
rect 929 37 945 71
rect 879 21 945 37
rect -849 -37 -783 -21
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -849 -87 -783 -71
rect -657 -37 -591 -21
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -657 -87 -591 -71
rect -465 -37 -399 -21
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -465 -87 -399 -71
rect -273 -37 -207 -21
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -273 -87 -207 -71
rect -81 -37 -15 -21
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect -81 -87 -15 -71
rect 111 -37 177 -21
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 111 -87 177 -71
rect 303 -37 369 -21
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 303 -87 369 -71
rect 495 -37 561 -21
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 495 -87 561 -71
rect 687 -37 753 -21
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 687 -87 753 -71
rect 879 -37 945 -21
rect 879 -71 895 -37
rect 929 -71 945 -37
rect 879 -87 945 -71
rect -927 -118 -897 -92
rect -831 -118 -801 -87
rect -735 -118 -705 -92
rect -639 -118 -609 -87
rect -543 -118 -513 -92
rect -447 -118 -417 -87
rect -351 -118 -321 -92
rect -255 -118 -225 -87
rect -159 -118 -129 -92
rect -63 -118 -33 -87
rect 33 -118 63 -92
rect 129 -118 159 -87
rect 225 -118 255 -92
rect 321 -118 351 -87
rect 417 -118 447 -92
rect 513 -118 543 -87
rect 609 -118 639 -92
rect 705 -118 735 -87
rect 801 -118 831 -92
rect 897 -118 927 -87
rect -927 -319 -897 -288
rect -831 -314 -801 -288
rect -735 -319 -705 -288
rect -639 -314 -609 -288
rect -543 -319 -513 -288
rect -447 -314 -417 -288
rect -351 -319 -321 -288
rect -255 -314 -225 -288
rect -159 -319 -129 -288
rect -63 -314 -33 -288
rect 33 -319 63 -288
rect 129 -314 159 -288
rect 225 -319 255 -288
rect 321 -314 351 -288
rect 417 -319 447 -288
rect 513 -314 543 -288
rect 609 -319 639 -288
rect 705 -314 735 -288
rect 801 -319 831 -288
rect 897 -314 927 -288
rect -945 -335 -879 -319
rect -945 -369 -929 -335
rect -895 -369 -879 -335
rect -945 -385 -879 -369
rect -753 -335 -687 -319
rect -753 -369 -737 -335
rect -703 -369 -687 -335
rect -753 -385 -687 -369
rect -561 -335 -495 -319
rect -561 -369 -545 -335
rect -511 -369 -495 -335
rect -561 -385 -495 -369
rect -369 -335 -303 -319
rect -369 -369 -353 -335
rect -319 -369 -303 -335
rect -369 -385 -303 -369
rect -177 -335 -111 -319
rect -177 -369 -161 -335
rect -127 -369 -111 -335
rect -177 -385 -111 -369
rect 15 -335 81 -319
rect 15 -369 31 -335
rect 65 -369 81 -335
rect 15 -385 81 -369
rect 207 -335 273 -319
rect 207 -369 223 -335
rect 257 -369 273 -335
rect 207 -385 273 -369
rect 399 -335 465 -319
rect 399 -369 415 -335
rect 449 -369 465 -335
rect 399 -385 465 -369
rect 591 -335 657 -319
rect 591 -369 607 -335
rect 641 -369 657 -335
rect 591 -385 657 -369
rect 783 -335 849 -319
rect 783 -369 799 -335
rect 833 -369 849 -335
rect 783 -385 849 -369
rect -945 -443 -879 -427
rect -945 -477 -929 -443
rect -895 -477 -879 -443
rect -945 -493 -879 -477
rect -753 -443 -687 -427
rect -753 -477 -737 -443
rect -703 -477 -687 -443
rect -753 -493 -687 -477
rect -561 -443 -495 -427
rect -561 -477 -545 -443
rect -511 -477 -495 -443
rect -561 -493 -495 -477
rect -369 -443 -303 -427
rect -369 -477 -353 -443
rect -319 -477 -303 -443
rect -369 -493 -303 -477
rect -177 -443 -111 -427
rect -177 -477 -161 -443
rect -127 -477 -111 -443
rect -177 -493 -111 -477
rect 15 -443 81 -427
rect 15 -477 31 -443
rect 65 -477 81 -443
rect 15 -493 81 -477
rect 207 -443 273 -427
rect 207 -477 223 -443
rect 257 -477 273 -443
rect 207 -493 273 -477
rect 399 -443 465 -427
rect 399 -477 415 -443
rect 449 -477 465 -443
rect 399 -493 465 -477
rect 591 -443 657 -427
rect 591 -477 607 -443
rect 641 -477 657 -443
rect 591 -493 657 -477
rect 783 -443 849 -427
rect 783 -477 799 -443
rect 833 -477 849 -443
rect 783 -493 849 -477
rect -927 -524 -897 -493
rect -831 -524 -801 -498
rect -735 -524 -705 -493
rect -639 -524 -609 -498
rect -543 -524 -513 -493
rect -447 -524 -417 -498
rect -351 -524 -321 -493
rect -255 -524 -225 -498
rect -159 -524 -129 -493
rect -63 -524 -33 -498
rect 33 -524 63 -493
rect 129 -524 159 -498
rect 225 -524 255 -493
rect 321 -524 351 -498
rect 417 -524 447 -493
rect 513 -524 543 -498
rect 609 -524 639 -493
rect 705 -524 735 -498
rect 801 -524 831 -493
rect 897 -524 927 -498
rect -927 -720 -897 -694
rect -831 -725 -801 -694
rect -735 -720 -705 -694
rect -639 -725 -609 -694
rect -543 -720 -513 -694
rect -447 -725 -417 -694
rect -351 -720 -321 -694
rect -255 -725 -225 -694
rect -159 -720 -129 -694
rect -63 -725 -33 -694
rect 33 -720 63 -694
rect 129 -725 159 -694
rect 225 -720 255 -694
rect 321 -725 351 -694
rect 417 -720 447 -694
rect 513 -725 543 -694
rect 609 -720 639 -694
rect 705 -725 735 -694
rect 801 -720 831 -694
rect 897 -725 927 -694
rect -849 -741 -783 -725
rect -849 -775 -833 -741
rect -799 -775 -783 -741
rect -849 -791 -783 -775
rect -657 -741 -591 -725
rect -657 -775 -641 -741
rect -607 -775 -591 -741
rect -657 -791 -591 -775
rect -465 -741 -399 -725
rect -465 -775 -449 -741
rect -415 -775 -399 -741
rect -465 -791 -399 -775
rect -273 -741 -207 -725
rect -273 -775 -257 -741
rect -223 -775 -207 -741
rect -273 -791 -207 -775
rect -81 -741 -15 -725
rect -81 -775 -65 -741
rect -31 -775 -15 -741
rect -81 -791 -15 -775
rect 111 -741 177 -725
rect 111 -775 127 -741
rect 161 -775 177 -741
rect 111 -791 177 -775
rect 303 -741 369 -725
rect 303 -775 319 -741
rect 353 -775 369 -741
rect 303 -791 369 -775
rect 495 -741 561 -725
rect 495 -775 511 -741
rect 545 -775 561 -741
rect 495 -791 561 -775
rect 687 -741 753 -725
rect 687 -775 703 -741
rect 737 -775 753 -741
rect 687 -791 753 -775
rect 879 -741 945 -725
rect 879 -775 895 -741
rect 929 -775 945 -741
rect 879 -791 945 -775
rect -849 -849 -783 -833
rect -849 -883 -833 -849
rect -799 -883 -783 -849
rect -849 -899 -783 -883
rect -657 -849 -591 -833
rect -657 -883 -641 -849
rect -607 -883 -591 -849
rect -657 -899 -591 -883
rect -465 -849 -399 -833
rect -465 -883 -449 -849
rect -415 -883 -399 -849
rect -465 -899 -399 -883
rect -273 -849 -207 -833
rect -273 -883 -257 -849
rect -223 -883 -207 -849
rect -273 -899 -207 -883
rect -81 -849 -15 -833
rect -81 -883 -65 -849
rect -31 -883 -15 -849
rect -81 -899 -15 -883
rect 111 -849 177 -833
rect 111 -883 127 -849
rect 161 -883 177 -849
rect 111 -899 177 -883
rect 303 -849 369 -833
rect 303 -883 319 -849
rect 353 -883 369 -849
rect 303 -899 369 -883
rect 495 -849 561 -833
rect 495 -883 511 -849
rect 545 -883 561 -849
rect 495 -899 561 -883
rect 687 -849 753 -833
rect 687 -883 703 -849
rect 737 -883 753 -849
rect 687 -899 753 -883
rect 879 -849 945 -833
rect 879 -883 895 -849
rect 929 -883 945 -849
rect 879 -899 945 -883
rect -927 -930 -897 -904
rect -831 -930 -801 -899
rect -735 -930 -705 -904
rect -639 -930 -609 -899
rect -543 -930 -513 -904
rect -447 -930 -417 -899
rect -351 -930 -321 -904
rect -255 -930 -225 -899
rect -159 -930 -129 -904
rect -63 -930 -33 -899
rect 33 -930 63 -904
rect 129 -930 159 -899
rect 225 -930 255 -904
rect 321 -930 351 -899
rect 417 -930 447 -904
rect 513 -930 543 -899
rect 609 -930 639 -904
rect 705 -930 735 -899
rect 801 -930 831 -904
rect 897 -930 927 -899
rect -927 -1131 -897 -1100
rect -831 -1126 -801 -1100
rect -735 -1131 -705 -1100
rect -639 -1126 -609 -1100
rect -543 -1131 -513 -1100
rect -447 -1126 -417 -1100
rect -351 -1131 -321 -1100
rect -255 -1126 -225 -1100
rect -159 -1131 -129 -1100
rect -63 -1126 -33 -1100
rect 33 -1131 63 -1100
rect 129 -1126 159 -1100
rect 225 -1131 255 -1100
rect 321 -1126 351 -1100
rect 417 -1131 447 -1100
rect 513 -1126 543 -1100
rect 609 -1131 639 -1100
rect 705 -1126 735 -1100
rect 801 -1131 831 -1100
rect 897 -1126 927 -1100
rect -945 -1147 -879 -1131
rect -945 -1181 -929 -1147
rect -895 -1181 -879 -1147
rect -945 -1197 -879 -1181
rect -753 -1147 -687 -1131
rect -753 -1181 -737 -1147
rect -703 -1181 -687 -1147
rect -753 -1197 -687 -1181
rect -561 -1147 -495 -1131
rect -561 -1181 -545 -1147
rect -511 -1181 -495 -1147
rect -561 -1197 -495 -1181
rect -369 -1147 -303 -1131
rect -369 -1181 -353 -1147
rect -319 -1181 -303 -1147
rect -369 -1197 -303 -1181
rect -177 -1147 -111 -1131
rect -177 -1181 -161 -1147
rect -127 -1181 -111 -1147
rect -177 -1197 -111 -1181
rect 15 -1147 81 -1131
rect 15 -1181 31 -1147
rect 65 -1181 81 -1147
rect 15 -1197 81 -1181
rect 207 -1147 273 -1131
rect 207 -1181 223 -1147
rect 257 -1181 273 -1147
rect 207 -1197 273 -1181
rect 399 -1147 465 -1131
rect 399 -1181 415 -1147
rect 449 -1181 465 -1147
rect 399 -1197 465 -1181
rect 591 -1147 657 -1131
rect 591 -1181 607 -1147
rect 641 -1181 657 -1147
rect 591 -1197 657 -1181
rect 783 -1147 849 -1131
rect 783 -1181 799 -1147
rect 833 -1181 849 -1147
rect 783 -1197 849 -1181
rect -945 -1255 -879 -1239
rect -945 -1289 -929 -1255
rect -895 -1289 -879 -1255
rect -945 -1305 -879 -1289
rect -753 -1255 -687 -1239
rect -753 -1289 -737 -1255
rect -703 -1289 -687 -1255
rect -753 -1305 -687 -1289
rect -561 -1255 -495 -1239
rect -561 -1289 -545 -1255
rect -511 -1289 -495 -1255
rect -561 -1305 -495 -1289
rect -369 -1255 -303 -1239
rect -369 -1289 -353 -1255
rect -319 -1289 -303 -1255
rect -369 -1305 -303 -1289
rect -177 -1255 -111 -1239
rect -177 -1289 -161 -1255
rect -127 -1289 -111 -1255
rect -177 -1305 -111 -1289
rect 15 -1255 81 -1239
rect 15 -1289 31 -1255
rect 65 -1289 81 -1255
rect 15 -1305 81 -1289
rect 207 -1255 273 -1239
rect 207 -1289 223 -1255
rect 257 -1289 273 -1255
rect 207 -1305 273 -1289
rect 399 -1255 465 -1239
rect 399 -1289 415 -1255
rect 449 -1289 465 -1255
rect 399 -1305 465 -1289
rect 591 -1255 657 -1239
rect 591 -1289 607 -1255
rect 641 -1289 657 -1255
rect 591 -1305 657 -1289
rect 783 -1255 849 -1239
rect 783 -1289 799 -1255
rect 833 -1289 849 -1255
rect 783 -1305 849 -1289
rect -927 -1336 -897 -1305
rect -831 -1336 -801 -1310
rect -735 -1336 -705 -1305
rect -639 -1336 -609 -1310
rect -543 -1336 -513 -1305
rect -447 -1336 -417 -1310
rect -351 -1336 -321 -1305
rect -255 -1336 -225 -1310
rect -159 -1336 -129 -1305
rect -63 -1336 -33 -1310
rect 33 -1336 63 -1305
rect 129 -1336 159 -1310
rect 225 -1336 255 -1305
rect 321 -1336 351 -1310
rect 417 -1336 447 -1305
rect 513 -1336 543 -1310
rect 609 -1336 639 -1305
rect 705 -1336 735 -1310
rect 801 -1336 831 -1305
rect 897 -1336 927 -1310
rect -927 -1532 -897 -1506
rect -831 -1537 -801 -1506
rect -735 -1532 -705 -1506
rect -639 -1537 -609 -1506
rect -543 -1532 -513 -1506
rect -447 -1537 -417 -1506
rect -351 -1532 -321 -1506
rect -255 -1537 -225 -1506
rect -159 -1532 -129 -1506
rect -63 -1537 -33 -1506
rect 33 -1532 63 -1506
rect 129 -1537 159 -1506
rect 225 -1532 255 -1506
rect 321 -1537 351 -1506
rect 417 -1532 447 -1506
rect 513 -1537 543 -1506
rect 609 -1532 639 -1506
rect 705 -1537 735 -1506
rect 801 -1532 831 -1506
rect 897 -1537 927 -1506
rect -849 -1553 -783 -1537
rect -849 -1587 -833 -1553
rect -799 -1587 -783 -1553
rect -849 -1603 -783 -1587
rect -657 -1553 -591 -1537
rect -657 -1587 -641 -1553
rect -607 -1587 -591 -1553
rect -657 -1603 -591 -1587
rect -465 -1553 -399 -1537
rect -465 -1587 -449 -1553
rect -415 -1587 -399 -1553
rect -465 -1603 -399 -1587
rect -273 -1553 -207 -1537
rect -273 -1587 -257 -1553
rect -223 -1587 -207 -1553
rect -273 -1603 -207 -1587
rect -81 -1553 -15 -1537
rect -81 -1587 -65 -1553
rect -31 -1587 -15 -1553
rect -81 -1603 -15 -1587
rect 111 -1553 177 -1537
rect 111 -1587 127 -1553
rect 161 -1587 177 -1553
rect 111 -1603 177 -1587
rect 303 -1553 369 -1537
rect 303 -1587 319 -1553
rect 353 -1587 369 -1553
rect 303 -1603 369 -1587
rect 495 -1553 561 -1537
rect 495 -1587 511 -1553
rect 545 -1587 561 -1553
rect 495 -1603 561 -1587
rect 687 -1553 753 -1537
rect 687 -1587 703 -1553
rect 737 -1587 753 -1553
rect 687 -1603 753 -1587
rect 879 -1553 945 -1537
rect 879 -1587 895 -1553
rect 929 -1587 945 -1553
rect 879 -1603 945 -1587
rect -849 -1661 -783 -1645
rect -849 -1695 -833 -1661
rect -799 -1695 -783 -1661
rect -849 -1711 -783 -1695
rect -657 -1661 -591 -1645
rect -657 -1695 -641 -1661
rect -607 -1695 -591 -1661
rect -657 -1711 -591 -1695
rect -465 -1661 -399 -1645
rect -465 -1695 -449 -1661
rect -415 -1695 -399 -1661
rect -465 -1711 -399 -1695
rect -273 -1661 -207 -1645
rect -273 -1695 -257 -1661
rect -223 -1695 -207 -1661
rect -273 -1711 -207 -1695
rect -81 -1661 -15 -1645
rect -81 -1695 -65 -1661
rect -31 -1695 -15 -1661
rect -81 -1711 -15 -1695
rect 111 -1661 177 -1645
rect 111 -1695 127 -1661
rect 161 -1695 177 -1661
rect 111 -1711 177 -1695
rect 303 -1661 369 -1645
rect 303 -1695 319 -1661
rect 353 -1695 369 -1661
rect 303 -1711 369 -1695
rect 495 -1661 561 -1645
rect 495 -1695 511 -1661
rect 545 -1695 561 -1661
rect 495 -1711 561 -1695
rect 687 -1661 753 -1645
rect 687 -1695 703 -1661
rect 737 -1695 753 -1661
rect 687 -1711 753 -1695
rect 879 -1661 945 -1645
rect 879 -1695 895 -1661
rect 929 -1695 945 -1661
rect 879 -1711 945 -1695
rect -927 -1742 -897 -1716
rect -831 -1742 -801 -1711
rect -735 -1742 -705 -1716
rect -639 -1742 -609 -1711
rect -543 -1742 -513 -1716
rect -447 -1742 -417 -1711
rect -351 -1742 -321 -1716
rect -255 -1742 -225 -1711
rect -159 -1742 -129 -1716
rect -63 -1742 -33 -1711
rect 33 -1742 63 -1716
rect 129 -1742 159 -1711
rect 225 -1742 255 -1716
rect 321 -1742 351 -1711
rect 417 -1742 447 -1716
rect 513 -1742 543 -1711
rect 609 -1742 639 -1716
rect 705 -1742 735 -1711
rect 801 -1742 831 -1716
rect 897 -1742 927 -1711
rect -927 -1943 -897 -1912
rect -831 -1938 -801 -1912
rect -735 -1943 -705 -1912
rect -639 -1938 -609 -1912
rect -543 -1943 -513 -1912
rect -447 -1938 -417 -1912
rect -351 -1943 -321 -1912
rect -255 -1938 -225 -1912
rect -159 -1943 -129 -1912
rect -63 -1938 -33 -1912
rect 33 -1943 63 -1912
rect 129 -1938 159 -1912
rect 225 -1943 255 -1912
rect 321 -1938 351 -1912
rect 417 -1943 447 -1912
rect 513 -1938 543 -1912
rect 609 -1943 639 -1912
rect 705 -1938 735 -1912
rect 801 -1943 831 -1912
rect 897 -1938 927 -1912
rect -945 -1959 -879 -1943
rect -945 -1993 -929 -1959
rect -895 -1993 -879 -1959
rect -945 -2009 -879 -1993
rect -753 -1959 -687 -1943
rect -753 -1993 -737 -1959
rect -703 -1993 -687 -1959
rect -753 -2009 -687 -1993
rect -561 -1959 -495 -1943
rect -561 -1993 -545 -1959
rect -511 -1993 -495 -1959
rect -561 -2009 -495 -1993
rect -369 -1959 -303 -1943
rect -369 -1993 -353 -1959
rect -319 -1993 -303 -1959
rect -369 -2009 -303 -1993
rect -177 -1959 -111 -1943
rect -177 -1993 -161 -1959
rect -127 -1993 -111 -1959
rect -177 -2009 -111 -1993
rect 15 -1959 81 -1943
rect 15 -1993 31 -1959
rect 65 -1993 81 -1959
rect 15 -2009 81 -1993
rect 207 -1959 273 -1943
rect 207 -1993 223 -1959
rect 257 -1993 273 -1959
rect 207 -2009 273 -1993
rect 399 -1959 465 -1943
rect 399 -1993 415 -1959
rect 449 -1993 465 -1959
rect 399 -2009 465 -1993
rect 591 -1959 657 -1943
rect 591 -1993 607 -1959
rect 641 -1993 657 -1959
rect 591 -2009 657 -1993
rect 783 -1959 849 -1943
rect 783 -1993 799 -1959
rect 833 -1993 849 -1959
rect 783 -2009 849 -1993
<< polycont >>
rect -929 1959 -895 1993
rect -737 1959 -703 1993
rect -545 1959 -511 1993
rect -353 1959 -319 1993
rect -161 1959 -127 1993
rect 31 1959 65 1993
rect 223 1959 257 1993
rect 415 1959 449 1993
rect 607 1959 641 1993
rect 799 1959 833 1993
rect -833 1661 -799 1695
rect -641 1661 -607 1695
rect -449 1661 -415 1695
rect -257 1661 -223 1695
rect -65 1661 -31 1695
rect 127 1661 161 1695
rect 319 1661 353 1695
rect 511 1661 545 1695
rect 703 1661 737 1695
rect 895 1661 929 1695
rect -833 1553 -799 1587
rect -641 1553 -607 1587
rect -449 1553 -415 1587
rect -257 1553 -223 1587
rect -65 1553 -31 1587
rect 127 1553 161 1587
rect 319 1553 353 1587
rect 511 1553 545 1587
rect 703 1553 737 1587
rect 895 1553 929 1587
rect -929 1255 -895 1289
rect -737 1255 -703 1289
rect -545 1255 -511 1289
rect -353 1255 -319 1289
rect -161 1255 -127 1289
rect 31 1255 65 1289
rect 223 1255 257 1289
rect 415 1255 449 1289
rect 607 1255 641 1289
rect 799 1255 833 1289
rect -929 1147 -895 1181
rect -737 1147 -703 1181
rect -545 1147 -511 1181
rect -353 1147 -319 1181
rect -161 1147 -127 1181
rect 31 1147 65 1181
rect 223 1147 257 1181
rect 415 1147 449 1181
rect 607 1147 641 1181
rect 799 1147 833 1181
rect -833 849 -799 883
rect -641 849 -607 883
rect -449 849 -415 883
rect -257 849 -223 883
rect -65 849 -31 883
rect 127 849 161 883
rect 319 849 353 883
rect 511 849 545 883
rect 703 849 737 883
rect 895 849 929 883
rect -833 741 -799 775
rect -641 741 -607 775
rect -449 741 -415 775
rect -257 741 -223 775
rect -65 741 -31 775
rect 127 741 161 775
rect 319 741 353 775
rect 511 741 545 775
rect 703 741 737 775
rect 895 741 929 775
rect -929 443 -895 477
rect -737 443 -703 477
rect -545 443 -511 477
rect -353 443 -319 477
rect -161 443 -127 477
rect 31 443 65 477
rect 223 443 257 477
rect 415 443 449 477
rect 607 443 641 477
rect 799 443 833 477
rect -929 335 -895 369
rect -737 335 -703 369
rect -545 335 -511 369
rect -353 335 -319 369
rect -161 335 -127 369
rect 31 335 65 369
rect 223 335 257 369
rect 415 335 449 369
rect 607 335 641 369
rect 799 335 833 369
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -929 -369 -895 -335
rect -737 -369 -703 -335
rect -545 -369 -511 -335
rect -353 -369 -319 -335
rect -161 -369 -127 -335
rect 31 -369 65 -335
rect 223 -369 257 -335
rect 415 -369 449 -335
rect 607 -369 641 -335
rect 799 -369 833 -335
rect -929 -477 -895 -443
rect -737 -477 -703 -443
rect -545 -477 -511 -443
rect -353 -477 -319 -443
rect -161 -477 -127 -443
rect 31 -477 65 -443
rect 223 -477 257 -443
rect 415 -477 449 -443
rect 607 -477 641 -443
rect 799 -477 833 -443
rect -833 -775 -799 -741
rect -641 -775 -607 -741
rect -449 -775 -415 -741
rect -257 -775 -223 -741
rect -65 -775 -31 -741
rect 127 -775 161 -741
rect 319 -775 353 -741
rect 511 -775 545 -741
rect 703 -775 737 -741
rect 895 -775 929 -741
rect -833 -883 -799 -849
rect -641 -883 -607 -849
rect -449 -883 -415 -849
rect -257 -883 -223 -849
rect -65 -883 -31 -849
rect 127 -883 161 -849
rect 319 -883 353 -849
rect 511 -883 545 -849
rect 703 -883 737 -849
rect 895 -883 929 -849
rect -929 -1181 -895 -1147
rect -737 -1181 -703 -1147
rect -545 -1181 -511 -1147
rect -353 -1181 -319 -1147
rect -161 -1181 -127 -1147
rect 31 -1181 65 -1147
rect 223 -1181 257 -1147
rect 415 -1181 449 -1147
rect 607 -1181 641 -1147
rect 799 -1181 833 -1147
rect -929 -1289 -895 -1255
rect -737 -1289 -703 -1255
rect -545 -1289 -511 -1255
rect -353 -1289 -319 -1255
rect -161 -1289 -127 -1255
rect 31 -1289 65 -1255
rect 223 -1289 257 -1255
rect 415 -1289 449 -1255
rect 607 -1289 641 -1255
rect 799 -1289 833 -1255
rect -833 -1587 -799 -1553
rect -641 -1587 -607 -1553
rect -449 -1587 -415 -1553
rect -257 -1587 -223 -1553
rect -65 -1587 -31 -1553
rect 127 -1587 161 -1553
rect 319 -1587 353 -1553
rect 511 -1587 545 -1553
rect 703 -1587 737 -1553
rect 895 -1587 929 -1553
rect -833 -1695 -799 -1661
rect -641 -1695 -607 -1661
rect -449 -1695 -415 -1661
rect -257 -1695 -223 -1661
rect -65 -1695 -31 -1661
rect 127 -1695 161 -1661
rect 319 -1695 353 -1661
rect 511 -1695 545 -1661
rect 703 -1695 737 -1661
rect 895 -1695 929 -1661
rect -929 -1993 -895 -1959
rect -737 -1993 -703 -1959
rect -545 -1993 -511 -1959
rect -353 -1993 -319 -1959
rect -161 -1993 -127 -1959
rect 31 -1993 65 -1959
rect 223 -1993 257 -1959
rect 415 -1993 449 -1959
rect 607 -1993 641 -1959
rect 799 -1993 833 -1959
<< locali >>
rect -1091 2061 -995 2095
rect 995 2061 1091 2095
rect -1091 1999 -1057 2061
rect 1057 1999 1091 2061
rect -945 1959 -929 1993
rect -895 1959 -879 1993
rect -753 1959 -737 1993
rect -703 1959 -687 1993
rect -561 1959 -545 1993
rect -511 1959 -495 1993
rect -369 1959 -353 1993
rect -319 1959 -303 1993
rect -177 1959 -161 1993
rect -127 1959 -111 1993
rect 15 1959 31 1993
rect 65 1959 81 1993
rect 207 1959 223 1993
rect 257 1959 273 1993
rect 399 1959 415 1993
rect 449 1959 465 1993
rect 591 1959 607 1993
rect 641 1959 657 1993
rect 783 1959 799 1993
rect 833 1959 849 1993
rect -977 1900 -943 1916
rect -977 1738 -943 1754
rect -881 1900 -847 1916
rect -881 1738 -847 1754
rect -785 1900 -751 1916
rect -785 1738 -751 1754
rect -689 1900 -655 1916
rect -689 1738 -655 1754
rect -593 1900 -559 1916
rect -593 1738 -559 1754
rect -497 1900 -463 1916
rect -497 1738 -463 1754
rect -401 1900 -367 1916
rect -401 1738 -367 1754
rect -305 1900 -271 1916
rect -305 1738 -271 1754
rect -209 1900 -175 1916
rect -209 1738 -175 1754
rect -113 1900 -79 1916
rect -113 1738 -79 1754
rect -17 1900 17 1916
rect -17 1738 17 1754
rect 79 1900 113 1916
rect 79 1738 113 1754
rect 175 1900 209 1916
rect 175 1738 209 1754
rect 271 1900 305 1916
rect 271 1738 305 1754
rect 367 1900 401 1916
rect 367 1738 401 1754
rect 463 1900 497 1916
rect 463 1738 497 1754
rect 559 1900 593 1916
rect 559 1738 593 1754
rect 655 1900 689 1916
rect 655 1738 689 1754
rect 751 1900 785 1916
rect 751 1738 785 1754
rect 847 1900 881 1916
rect 847 1738 881 1754
rect 943 1900 977 1916
rect 943 1738 977 1754
rect -849 1661 -833 1695
rect -799 1661 -783 1695
rect -657 1661 -641 1695
rect -607 1661 -591 1695
rect -465 1661 -449 1695
rect -415 1661 -399 1695
rect -273 1661 -257 1695
rect -223 1661 -207 1695
rect -81 1661 -65 1695
rect -31 1661 -15 1695
rect 111 1661 127 1695
rect 161 1661 177 1695
rect 303 1661 319 1695
rect 353 1661 369 1695
rect 495 1661 511 1695
rect 545 1661 561 1695
rect 687 1661 703 1695
rect 737 1661 753 1695
rect 879 1661 895 1695
rect 929 1661 945 1695
rect -849 1553 -833 1587
rect -799 1553 -783 1587
rect -657 1553 -641 1587
rect -607 1553 -591 1587
rect -465 1553 -449 1587
rect -415 1553 -399 1587
rect -273 1553 -257 1587
rect -223 1553 -207 1587
rect -81 1553 -65 1587
rect -31 1553 -15 1587
rect 111 1553 127 1587
rect 161 1553 177 1587
rect 303 1553 319 1587
rect 353 1553 369 1587
rect 495 1553 511 1587
rect 545 1553 561 1587
rect 687 1553 703 1587
rect 737 1553 753 1587
rect 879 1553 895 1587
rect 929 1553 945 1587
rect -977 1494 -943 1510
rect -977 1332 -943 1348
rect -881 1494 -847 1510
rect -881 1332 -847 1348
rect -785 1494 -751 1510
rect -785 1332 -751 1348
rect -689 1494 -655 1510
rect -689 1332 -655 1348
rect -593 1494 -559 1510
rect -593 1332 -559 1348
rect -497 1494 -463 1510
rect -497 1332 -463 1348
rect -401 1494 -367 1510
rect -401 1332 -367 1348
rect -305 1494 -271 1510
rect -305 1332 -271 1348
rect -209 1494 -175 1510
rect -209 1332 -175 1348
rect -113 1494 -79 1510
rect -113 1332 -79 1348
rect -17 1494 17 1510
rect -17 1332 17 1348
rect 79 1494 113 1510
rect 79 1332 113 1348
rect 175 1494 209 1510
rect 175 1332 209 1348
rect 271 1494 305 1510
rect 271 1332 305 1348
rect 367 1494 401 1510
rect 367 1332 401 1348
rect 463 1494 497 1510
rect 463 1332 497 1348
rect 559 1494 593 1510
rect 559 1332 593 1348
rect 655 1494 689 1510
rect 655 1332 689 1348
rect 751 1494 785 1510
rect 751 1332 785 1348
rect 847 1494 881 1510
rect 847 1332 881 1348
rect 943 1494 977 1510
rect 943 1332 977 1348
rect -945 1255 -929 1289
rect -895 1255 -879 1289
rect -753 1255 -737 1289
rect -703 1255 -687 1289
rect -561 1255 -545 1289
rect -511 1255 -495 1289
rect -369 1255 -353 1289
rect -319 1255 -303 1289
rect -177 1255 -161 1289
rect -127 1255 -111 1289
rect 15 1255 31 1289
rect 65 1255 81 1289
rect 207 1255 223 1289
rect 257 1255 273 1289
rect 399 1255 415 1289
rect 449 1255 465 1289
rect 591 1255 607 1289
rect 641 1255 657 1289
rect 783 1255 799 1289
rect 833 1255 849 1289
rect -945 1147 -929 1181
rect -895 1147 -879 1181
rect -753 1147 -737 1181
rect -703 1147 -687 1181
rect -561 1147 -545 1181
rect -511 1147 -495 1181
rect -369 1147 -353 1181
rect -319 1147 -303 1181
rect -177 1147 -161 1181
rect -127 1147 -111 1181
rect 15 1147 31 1181
rect 65 1147 81 1181
rect 207 1147 223 1181
rect 257 1147 273 1181
rect 399 1147 415 1181
rect 449 1147 465 1181
rect 591 1147 607 1181
rect 641 1147 657 1181
rect 783 1147 799 1181
rect 833 1147 849 1181
rect -977 1088 -943 1104
rect -977 926 -943 942
rect -881 1088 -847 1104
rect -881 926 -847 942
rect -785 1088 -751 1104
rect -785 926 -751 942
rect -689 1088 -655 1104
rect -689 926 -655 942
rect -593 1088 -559 1104
rect -593 926 -559 942
rect -497 1088 -463 1104
rect -497 926 -463 942
rect -401 1088 -367 1104
rect -401 926 -367 942
rect -305 1088 -271 1104
rect -305 926 -271 942
rect -209 1088 -175 1104
rect -209 926 -175 942
rect -113 1088 -79 1104
rect -113 926 -79 942
rect -17 1088 17 1104
rect -17 926 17 942
rect 79 1088 113 1104
rect 79 926 113 942
rect 175 1088 209 1104
rect 175 926 209 942
rect 271 1088 305 1104
rect 271 926 305 942
rect 367 1088 401 1104
rect 367 926 401 942
rect 463 1088 497 1104
rect 463 926 497 942
rect 559 1088 593 1104
rect 559 926 593 942
rect 655 1088 689 1104
rect 655 926 689 942
rect 751 1088 785 1104
rect 751 926 785 942
rect 847 1088 881 1104
rect 847 926 881 942
rect 943 1088 977 1104
rect 943 926 977 942
rect -849 849 -833 883
rect -799 849 -783 883
rect -657 849 -641 883
rect -607 849 -591 883
rect -465 849 -449 883
rect -415 849 -399 883
rect -273 849 -257 883
rect -223 849 -207 883
rect -81 849 -65 883
rect -31 849 -15 883
rect 111 849 127 883
rect 161 849 177 883
rect 303 849 319 883
rect 353 849 369 883
rect 495 849 511 883
rect 545 849 561 883
rect 687 849 703 883
rect 737 849 753 883
rect 879 849 895 883
rect 929 849 945 883
rect -849 741 -833 775
rect -799 741 -783 775
rect -657 741 -641 775
rect -607 741 -591 775
rect -465 741 -449 775
rect -415 741 -399 775
rect -273 741 -257 775
rect -223 741 -207 775
rect -81 741 -65 775
rect -31 741 -15 775
rect 111 741 127 775
rect 161 741 177 775
rect 303 741 319 775
rect 353 741 369 775
rect 495 741 511 775
rect 545 741 561 775
rect 687 741 703 775
rect 737 741 753 775
rect 879 741 895 775
rect 929 741 945 775
rect -977 682 -943 698
rect -977 520 -943 536
rect -881 682 -847 698
rect -881 520 -847 536
rect -785 682 -751 698
rect -785 520 -751 536
rect -689 682 -655 698
rect -689 520 -655 536
rect -593 682 -559 698
rect -593 520 -559 536
rect -497 682 -463 698
rect -497 520 -463 536
rect -401 682 -367 698
rect -401 520 -367 536
rect -305 682 -271 698
rect -305 520 -271 536
rect -209 682 -175 698
rect -209 520 -175 536
rect -113 682 -79 698
rect -113 520 -79 536
rect -17 682 17 698
rect -17 520 17 536
rect 79 682 113 698
rect 79 520 113 536
rect 175 682 209 698
rect 175 520 209 536
rect 271 682 305 698
rect 271 520 305 536
rect 367 682 401 698
rect 367 520 401 536
rect 463 682 497 698
rect 463 520 497 536
rect 559 682 593 698
rect 559 520 593 536
rect 655 682 689 698
rect 655 520 689 536
rect 751 682 785 698
rect 751 520 785 536
rect 847 682 881 698
rect 847 520 881 536
rect 943 682 977 698
rect 943 520 977 536
rect -945 443 -929 477
rect -895 443 -879 477
rect -753 443 -737 477
rect -703 443 -687 477
rect -561 443 -545 477
rect -511 443 -495 477
rect -369 443 -353 477
rect -319 443 -303 477
rect -177 443 -161 477
rect -127 443 -111 477
rect 15 443 31 477
rect 65 443 81 477
rect 207 443 223 477
rect 257 443 273 477
rect 399 443 415 477
rect 449 443 465 477
rect 591 443 607 477
rect 641 443 657 477
rect 783 443 799 477
rect 833 443 849 477
rect -945 335 -929 369
rect -895 335 -879 369
rect -753 335 -737 369
rect -703 335 -687 369
rect -561 335 -545 369
rect -511 335 -495 369
rect -369 335 -353 369
rect -319 335 -303 369
rect -177 335 -161 369
rect -127 335 -111 369
rect 15 335 31 369
rect 65 335 81 369
rect 207 335 223 369
rect 257 335 273 369
rect 399 335 415 369
rect 449 335 465 369
rect 591 335 607 369
rect 641 335 657 369
rect 783 335 799 369
rect 833 335 849 369
rect -977 276 -943 292
rect -977 114 -943 130
rect -881 276 -847 292
rect -881 114 -847 130
rect -785 276 -751 292
rect -785 114 -751 130
rect -689 276 -655 292
rect -689 114 -655 130
rect -593 276 -559 292
rect -593 114 -559 130
rect -497 276 -463 292
rect -497 114 -463 130
rect -401 276 -367 292
rect -401 114 -367 130
rect -305 276 -271 292
rect -305 114 -271 130
rect -209 276 -175 292
rect -209 114 -175 130
rect -113 276 -79 292
rect -113 114 -79 130
rect -17 276 17 292
rect -17 114 17 130
rect 79 276 113 292
rect 79 114 113 130
rect 175 276 209 292
rect 175 114 209 130
rect 271 276 305 292
rect 271 114 305 130
rect 367 276 401 292
rect 367 114 401 130
rect 463 276 497 292
rect 463 114 497 130
rect 559 276 593 292
rect 559 114 593 130
rect 655 276 689 292
rect 655 114 689 130
rect 751 276 785 292
rect 751 114 785 130
rect 847 276 881 292
rect 847 114 881 130
rect 943 276 977 292
rect 943 114 977 130
rect -849 37 -833 71
rect -799 37 -783 71
rect -657 37 -641 71
rect -607 37 -591 71
rect -465 37 -449 71
rect -415 37 -399 71
rect -273 37 -257 71
rect -223 37 -207 71
rect -81 37 -65 71
rect -31 37 -15 71
rect 111 37 127 71
rect 161 37 177 71
rect 303 37 319 71
rect 353 37 369 71
rect 495 37 511 71
rect 545 37 561 71
rect 687 37 703 71
rect 737 37 753 71
rect 879 37 895 71
rect 929 37 945 71
rect -849 -71 -833 -37
rect -799 -71 -783 -37
rect -657 -71 -641 -37
rect -607 -71 -591 -37
rect -465 -71 -449 -37
rect -415 -71 -399 -37
rect -273 -71 -257 -37
rect -223 -71 -207 -37
rect -81 -71 -65 -37
rect -31 -71 -15 -37
rect 111 -71 127 -37
rect 161 -71 177 -37
rect 303 -71 319 -37
rect 353 -71 369 -37
rect 495 -71 511 -37
rect 545 -71 561 -37
rect 687 -71 703 -37
rect 737 -71 753 -37
rect 879 -71 895 -37
rect 929 -71 945 -37
rect -977 -130 -943 -114
rect -977 -292 -943 -276
rect -881 -130 -847 -114
rect -881 -292 -847 -276
rect -785 -130 -751 -114
rect -785 -292 -751 -276
rect -689 -130 -655 -114
rect -689 -292 -655 -276
rect -593 -130 -559 -114
rect -593 -292 -559 -276
rect -497 -130 -463 -114
rect -497 -292 -463 -276
rect -401 -130 -367 -114
rect -401 -292 -367 -276
rect -305 -130 -271 -114
rect -305 -292 -271 -276
rect -209 -130 -175 -114
rect -209 -292 -175 -276
rect -113 -130 -79 -114
rect -113 -292 -79 -276
rect -17 -130 17 -114
rect -17 -292 17 -276
rect 79 -130 113 -114
rect 79 -292 113 -276
rect 175 -130 209 -114
rect 175 -292 209 -276
rect 271 -130 305 -114
rect 271 -292 305 -276
rect 367 -130 401 -114
rect 367 -292 401 -276
rect 463 -130 497 -114
rect 463 -292 497 -276
rect 559 -130 593 -114
rect 559 -292 593 -276
rect 655 -130 689 -114
rect 655 -292 689 -276
rect 751 -130 785 -114
rect 751 -292 785 -276
rect 847 -130 881 -114
rect 847 -292 881 -276
rect 943 -130 977 -114
rect 943 -292 977 -276
rect -945 -369 -929 -335
rect -895 -369 -879 -335
rect -753 -369 -737 -335
rect -703 -369 -687 -335
rect -561 -369 -545 -335
rect -511 -369 -495 -335
rect -369 -369 -353 -335
rect -319 -369 -303 -335
rect -177 -369 -161 -335
rect -127 -369 -111 -335
rect 15 -369 31 -335
rect 65 -369 81 -335
rect 207 -369 223 -335
rect 257 -369 273 -335
rect 399 -369 415 -335
rect 449 -369 465 -335
rect 591 -369 607 -335
rect 641 -369 657 -335
rect 783 -369 799 -335
rect 833 -369 849 -335
rect -945 -477 -929 -443
rect -895 -477 -879 -443
rect -753 -477 -737 -443
rect -703 -477 -687 -443
rect -561 -477 -545 -443
rect -511 -477 -495 -443
rect -369 -477 -353 -443
rect -319 -477 -303 -443
rect -177 -477 -161 -443
rect -127 -477 -111 -443
rect 15 -477 31 -443
rect 65 -477 81 -443
rect 207 -477 223 -443
rect 257 -477 273 -443
rect 399 -477 415 -443
rect 449 -477 465 -443
rect 591 -477 607 -443
rect 641 -477 657 -443
rect 783 -477 799 -443
rect 833 -477 849 -443
rect -977 -536 -943 -520
rect -977 -698 -943 -682
rect -881 -536 -847 -520
rect -881 -698 -847 -682
rect -785 -536 -751 -520
rect -785 -698 -751 -682
rect -689 -536 -655 -520
rect -689 -698 -655 -682
rect -593 -536 -559 -520
rect -593 -698 -559 -682
rect -497 -536 -463 -520
rect -497 -698 -463 -682
rect -401 -536 -367 -520
rect -401 -698 -367 -682
rect -305 -536 -271 -520
rect -305 -698 -271 -682
rect -209 -536 -175 -520
rect -209 -698 -175 -682
rect -113 -536 -79 -520
rect -113 -698 -79 -682
rect -17 -536 17 -520
rect -17 -698 17 -682
rect 79 -536 113 -520
rect 79 -698 113 -682
rect 175 -536 209 -520
rect 175 -698 209 -682
rect 271 -536 305 -520
rect 271 -698 305 -682
rect 367 -536 401 -520
rect 367 -698 401 -682
rect 463 -536 497 -520
rect 463 -698 497 -682
rect 559 -536 593 -520
rect 559 -698 593 -682
rect 655 -536 689 -520
rect 655 -698 689 -682
rect 751 -536 785 -520
rect 751 -698 785 -682
rect 847 -536 881 -520
rect 847 -698 881 -682
rect 943 -536 977 -520
rect 943 -698 977 -682
rect -849 -775 -833 -741
rect -799 -775 -783 -741
rect -657 -775 -641 -741
rect -607 -775 -591 -741
rect -465 -775 -449 -741
rect -415 -775 -399 -741
rect -273 -775 -257 -741
rect -223 -775 -207 -741
rect -81 -775 -65 -741
rect -31 -775 -15 -741
rect 111 -775 127 -741
rect 161 -775 177 -741
rect 303 -775 319 -741
rect 353 -775 369 -741
rect 495 -775 511 -741
rect 545 -775 561 -741
rect 687 -775 703 -741
rect 737 -775 753 -741
rect 879 -775 895 -741
rect 929 -775 945 -741
rect -849 -883 -833 -849
rect -799 -883 -783 -849
rect -657 -883 -641 -849
rect -607 -883 -591 -849
rect -465 -883 -449 -849
rect -415 -883 -399 -849
rect -273 -883 -257 -849
rect -223 -883 -207 -849
rect -81 -883 -65 -849
rect -31 -883 -15 -849
rect 111 -883 127 -849
rect 161 -883 177 -849
rect 303 -883 319 -849
rect 353 -883 369 -849
rect 495 -883 511 -849
rect 545 -883 561 -849
rect 687 -883 703 -849
rect 737 -883 753 -849
rect 879 -883 895 -849
rect 929 -883 945 -849
rect -977 -942 -943 -926
rect -977 -1104 -943 -1088
rect -881 -942 -847 -926
rect -881 -1104 -847 -1088
rect -785 -942 -751 -926
rect -785 -1104 -751 -1088
rect -689 -942 -655 -926
rect -689 -1104 -655 -1088
rect -593 -942 -559 -926
rect -593 -1104 -559 -1088
rect -497 -942 -463 -926
rect -497 -1104 -463 -1088
rect -401 -942 -367 -926
rect -401 -1104 -367 -1088
rect -305 -942 -271 -926
rect -305 -1104 -271 -1088
rect -209 -942 -175 -926
rect -209 -1104 -175 -1088
rect -113 -942 -79 -926
rect -113 -1104 -79 -1088
rect -17 -942 17 -926
rect -17 -1104 17 -1088
rect 79 -942 113 -926
rect 79 -1104 113 -1088
rect 175 -942 209 -926
rect 175 -1104 209 -1088
rect 271 -942 305 -926
rect 271 -1104 305 -1088
rect 367 -942 401 -926
rect 367 -1104 401 -1088
rect 463 -942 497 -926
rect 463 -1104 497 -1088
rect 559 -942 593 -926
rect 559 -1104 593 -1088
rect 655 -942 689 -926
rect 655 -1104 689 -1088
rect 751 -942 785 -926
rect 751 -1104 785 -1088
rect 847 -942 881 -926
rect 847 -1104 881 -1088
rect 943 -942 977 -926
rect 943 -1104 977 -1088
rect -945 -1181 -929 -1147
rect -895 -1181 -879 -1147
rect -753 -1181 -737 -1147
rect -703 -1181 -687 -1147
rect -561 -1181 -545 -1147
rect -511 -1181 -495 -1147
rect -369 -1181 -353 -1147
rect -319 -1181 -303 -1147
rect -177 -1181 -161 -1147
rect -127 -1181 -111 -1147
rect 15 -1181 31 -1147
rect 65 -1181 81 -1147
rect 207 -1181 223 -1147
rect 257 -1181 273 -1147
rect 399 -1181 415 -1147
rect 449 -1181 465 -1147
rect 591 -1181 607 -1147
rect 641 -1181 657 -1147
rect 783 -1181 799 -1147
rect 833 -1181 849 -1147
rect -945 -1289 -929 -1255
rect -895 -1289 -879 -1255
rect -753 -1289 -737 -1255
rect -703 -1289 -687 -1255
rect -561 -1289 -545 -1255
rect -511 -1289 -495 -1255
rect -369 -1289 -353 -1255
rect -319 -1289 -303 -1255
rect -177 -1289 -161 -1255
rect -127 -1289 -111 -1255
rect 15 -1289 31 -1255
rect 65 -1289 81 -1255
rect 207 -1289 223 -1255
rect 257 -1289 273 -1255
rect 399 -1289 415 -1255
rect 449 -1289 465 -1255
rect 591 -1289 607 -1255
rect 641 -1289 657 -1255
rect 783 -1289 799 -1255
rect 833 -1289 849 -1255
rect -977 -1348 -943 -1332
rect -977 -1510 -943 -1494
rect -881 -1348 -847 -1332
rect -881 -1510 -847 -1494
rect -785 -1348 -751 -1332
rect -785 -1510 -751 -1494
rect -689 -1348 -655 -1332
rect -689 -1510 -655 -1494
rect -593 -1348 -559 -1332
rect -593 -1510 -559 -1494
rect -497 -1348 -463 -1332
rect -497 -1510 -463 -1494
rect -401 -1348 -367 -1332
rect -401 -1510 -367 -1494
rect -305 -1348 -271 -1332
rect -305 -1510 -271 -1494
rect -209 -1348 -175 -1332
rect -209 -1510 -175 -1494
rect -113 -1348 -79 -1332
rect -113 -1510 -79 -1494
rect -17 -1348 17 -1332
rect -17 -1510 17 -1494
rect 79 -1348 113 -1332
rect 79 -1510 113 -1494
rect 175 -1348 209 -1332
rect 175 -1510 209 -1494
rect 271 -1348 305 -1332
rect 271 -1510 305 -1494
rect 367 -1348 401 -1332
rect 367 -1510 401 -1494
rect 463 -1348 497 -1332
rect 463 -1510 497 -1494
rect 559 -1348 593 -1332
rect 559 -1510 593 -1494
rect 655 -1348 689 -1332
rect 655 -1510 689 -1494
rect 751 -1348 785 -1332
rect 751 -1510 785 -1494
rect 847 -1348 881 -1332
rect 847 -1510 881 -1494
rect 943 -1348 977 -1332
rect 943 -1510 977 -1494
rect -849 -1587 -833 -1553
rect -799 -1587 -783 -1553
rect -657 -1587 -641 -1553
rect -607 -1587 -591 -1553
rect -465 -1587 -449 -1553
rect -415 -1587 -399 -1553
rect -273 -1587 -257 -1553
rect -223 -1587 -207 -1553
rect -81 -1587 -65 -1553
rect -31 -1587 -15 -1553
rect 111 -1587 127 -1553
rect 161 -1587 177 -1553
rect 303 -1587 319 -1553
rect 353 -1587 369 -1553
rect 495 -1587 511 -1553
rect 545 -1587 561 -1553
rect 687 -1587 703 -1553
rect 737 -1587 753 -1553
rect 879 -1587 895 -1553
rect 929 -1587 945 -1553
rect -849 -1695 -833 -1661
rect -799 -1695 -783 -1661
rect -657 -1695 -641 -1661
rect -607 -1695 -591 -1661
rect -465 -1695 -449 -1661
rect -415 -1695 -399 -1661
rect -273 -1695 -257 -1661
rect -223 -1695 -207 -1661
rect -81 -1695 -65 -1661
rect -31 -1695 -15 -1661
rect 111 -1695 127 -1661
rect 161 -1695 177 -1661
rect 303 -1695 319 -1661
rect 353 -1695 369 -1661
rect 495 -1695 511 -1661
rect 545 -1695 561 -1661
rect 687 -1695 703 -1661
rect 737 -1695 753 -1661
rect 879 -1695 895 -1661
rect 929 -1695 945 -1661
rect -977 -1754 -943 -1738
rect -977 -1916 -943 -1900
rect -881 -1754 -847 -1738
rect -881 -1916 -847 -1900
rect -785 -1754 -751 -1738
rect -785 -1916 -751 -1900
rect -689 -1754 -655 -1738
rect -689 -1916 -655 -1900
rect -593 -1754 -559 -1738
rect -593 -1916 -559 -1900
rect -497 -1754 -463 -1738
rect -497 -1916 -463 -1900
rect -401 -1754 -367 -1738
rect -401 -1916 -367 -1900
rect -305 -1754 -271 -1738
rect -305 -1916 -271 -1900
rect -209 -1754 -175 -1738
rect -209 -1916 -175 -1900
rect -113 -1754 -79 -1738
rect -113 -1916 -79 -1900
rect -17 -1754 17 -1738
rect -17 -1916 17 -1900
rect 79 -1754 113 -1738
rect 79 -1916 113 -1900
rect 175 -1754 209 -1738
rect 175 -1916 209 -1900
rect 271 -1754 305 -1738
rect 271 -1916 305 -1900
rect 367 -1754 401 -1738
rect 367 -1916 401 -1900
rect 463 -1754 497 -1738
rect 463 -1916 497 -1900
rect 559 -1754 593 -1738
rect 559 -1916 593 -1900
rect 655 -1754 689 -1738
rect 655 -1916 689 -1900
rect 751 -1754 785 -1738
rect 751 -1916 785 -1900
rect 847 -1754 881 -1738
rect 847 -1916 881 -1900
rect 943 -1754 977 -1738
rect 943 -1916 977 -1900
rect -945 -1993 -929 -1959
rect -895 -1993 -879 -1959
rect -753 -1993 -737 -1959
rect -703 -1993 -687 -1959
rect -561 -1993 -545 -1959
rect -511 -1993 -495 -1959
rect -369 -1993 -353 -1959
rect -319 -1993 -303 -1959
rect -177 -1993 -161 -1959
rect -127 -1993 -111 -1959
rect 15 -1993 31 -1959
rect 65 -1993 81 -1959
rect 207 -1993 223 -1959
rect 257 -1993 273 -1959
rect 399 -1993 415 -1959
rect 449 -1993 465 -1959
rect 591 -1993 607 -1959
rect 641 -1993 657 -1959
rect 783 -1993 799 -1959
rect 833 -1993 849 -1959
rect -1091 -2061 -1057 -1999
rect 1057 -2061 1091 -1999
rect -1091 -2095 -995 -2061
rect 995 -2095 1091 -2061
<< viali >>
rect -929 1959 -895 1993
rect -737 1959 -703 1993
rect -545 1959 -511 1993
rect -353 1959 -319 1993
rect -161 1959 -127 1993
rect 31 1959 65 1993
rect 223 1959 257 1993
rect 415 1959 449 1993
rect 607 1959 641 1993
rect 799 1959 833 1993
rect -977 1754 -943 1900
rect -881 1754 -847 1900
rect -785 1754 -751 1900
rect -689 1754 -655 1900
rect -593 1754 -559 1900
rect -497 1754 -463 1900
rect -401 1754 -367 1900
rect -305 1754 -271 1900
rect -209 1754 -175 1900
rect -113 1754 -79 1900
rect -17 1754 17 1900
rect 79 1754 113 1900
rect 175 1754 209 1900
rect 271 1754 305 1900
rect 367 1754 401 1900
rect 463 1754 497 1900
rect 559 1754 593 1900
rect 655 1754 689 1900
rect 751 1754 785 1900
rect 847 1754 881 1900
rect 943 1754 977 1900
rect -833 1661 -799 1695
rect -641 1661 -607 1695
rect -449 1661 -415 1695
rect -257 1661 -223 1695
rect -65 1661 -31 1695
rect 127 1661 161 1695
rect 319 1661 353 1695
rect 511 1661 545 1695
rect 703 1661 737 1695
rect 895 1661 929 1695
rect -833 1553 -799 1587
rect -641 1553 -607 1587
rect -449 1553 -415 1587
rect -257 1553 -223 1587
rect -65 1553 -31 1587
rect 127 1553 161 1587
rect 319 1553 353 1587
rect 511 1553 545 1587
rect 703 1553 737 1587
rect 895 1553 929 1587
rect -977 1348 -943 1494
rect -881 1348 -847 1494
rect -785 1348 -751 1494
rect -689 1348 -655 1494
rect -593 1348 -559 1494
rect -497 1348 -463 1494
rect -401 1348 -367 1494
rect -305 1348 -271 1494
rect -209 1348 -175 1494
rect -113 1348 -79 1494
rect -17 1348 17 1494
rect 79 1348 113 1494
rect 175 1348 209 1494
rect 271 1348 305 1494
rect 367 1348 401 1494
rect 463 1348 497 1494
rect 559 1348 593 1494
rect 655 1348 689 1494
rect 751 1348 785 1494
rect 847 1348 881 1494
rect 943 1348 977 1494
rect -929 1255 -895 1289
rect -737 1255 -703 1289
rect -545 1255 -511 1289
rect -353 1255 -319 1289
rect -161 1255 -127 1289
rect 31 1255 65 1289
rect 223 1255 257 1289
rect 415 1255 449 1289
rect 607 1255 641 1289
rect 799 1255 833 1289
rect -929 1147 -895 1181
rect -737 1147 -703 1181
rect -545 1147 -511 1181
rect -353 1147 -319 1181
rect -161 1147 -127 1181
rect 31 1147 65 1181
rect 223 1147 257 1181
rect 415 1147 449 1181
rect 607 1147 641 1181
rect 799 1147 833 1181
rect -977 942 -943 1088
rect -881 942 -847 1088
rect -785 942 -751 1088
rect -689 942 -655 1088
rect -593 942 -559 1088
rect -497 942 -463 1088
rect -401 942 -367 1088
rect -305 942 -271 1088
rect -209 942 -175 1088
rect -113 942 -79 1088
rect -17 942 17 1088
rect 79 942 113 1088
rect 175 942 209 1088
rect 271 942 305 1088
rect 367 942 401 1088
rect 463 942 497 1088
rect 559 942 593 1088
rect 655 942 689 1088
rect 751 942 785 1088
rect 847 942 881 1088
rect 943 942 977 1088
rect -833 849 -799 883
rect -641 849 -607 883
rect -449 849 -415 883
rect -257 849 -223 883
rect -65 849 -31 883
rect 127 849 161 883
rect 319 849 353 883
rect 511 849 545 883
rect 703 849 737 883
rect 895 849 929 883
rect -833 741 -799 775
rect -641 741 -607 775
rect -449 741 -415 775
rect -257 741 -223 775
rect -65 741 -31 775
rect 127 741 161 775
rect 319 741 353 775
rect 511 741 545 775
rect 703 741 737 775
rect 895 741 929 775
rect -977 536 -943 682
rect -881 536 -847 682
rect -785 536 -751 682
rect -689 536 -655 682
rect -593 536 -559 682
rect -497 536 -463 682
rect -401 536 -367 682
rect -305 536 -271 682
rect -209 536 -175 682
rect -113 536 -79 682
rect -17 536 17 682
rect 79 536 113 682
rect 175 536 209 682
rect 271 536 305 682
rect 367 536 401 682
rect 463 536 497 682
rect 559 536 593 682
rect 655 536 689 682
rect 751 536 785 682
rect 847 536 881 682
rect 943 536 977 682
rect -929 443 -895 477
rect -737 443 -703 477
rect -545 443 -511 477
rect -353 443 -319 477
rect -161 443 -127 477
rect 31 443 65 477
rect 223 443 257 477
rect 415 443 449 477
rect 607 443 641 477
rect 799 443 833 477
rect -929 335 -895 369
rect -737 335 -703 369
rect -545 335 -511 369
rect -353 335 -319 369
rect -161 335 -127 369
rect 31 335 65 369
rect 223 335 257 369
rect 415 335 449 369
rect 607 335 641 369
rect 799 335 833 369
rect -977 130 -943 276
rect -881 130 -847 276
rect -785 130 -751 276
rect -689 130 -655 276
rect -593 130 -559 276
rect -497 130 -463 276
rect -401 130 -367 276
rect -305 130 -271 276
rect -209 130 -175 276
rect -113 130 -79 276
rect -17 130 17 276
rect 79 130 113 276
rect 175 130 209 276
rect 271 130 305 276
rect 367 130 401 276
rect 463 130 497 276
rect 559 130 593 276
rect 655 130 689 276
rect 751 130 785 276
rect 847 130 881 276
rect 943 130 977 276
rect -833 37 -799 71
rect -641 37 -607 71
rect -449 37 -415 71
rect -257 37 -223 71
rect -65 37 -31 71
rect 127 37 161 71
rect 319 37 353 71
rect 511 37 545 71
rect 703 37 737 71
rect 895 37 929 71
rect -833 -71 -799 -37
rect -641 -71 -607 -37
rect -449 -71 -415 -37
rect -257 -71 -223 -37
rect -65 -71 -31 -37
rect 127 -71 161 -37
rect 319 -71 353 -37
rect 511 -71 545 -37
rect 703 -71 737 -37
rect 895 -71 929 -37
rect -977 -276 -943 -130
rect -881 -276 -847 -130
rect -785 -276 -751 -130
rect -689 -276 -655 -130
rect -593 -276 -559 -130
rect -497 -276 -463 -130
rect -401 -276 -367 -130
rect -305 -276 -271 -130
rect -209 -276 -175 -130
rect -113 -276 -79 -130
rect -17 -276 17 -130
rect 79 -276 113 -130
rect 175 -276 209 -130
rect 271 -276 305 -130
rect 367 -276 401 -130
rect 463 -276 497 -130
rect 559 -276 593 -130
rect 655 -276 689 -130
rect 751 -276 785 -130
rect 847 -276 881 -130
rect 943 -276 977 -130
rect -929 -369 -895 -335
rect -737 -369 -703 -335
rect -545 -369 -511 -335
rect -353 -369 -319 -335
rect -161 -369 -127 -335
rect 31 -369 65 -335
rect 223 -369 257 -335
rect 415 -369 449 -335
rect 607 -369 641 -335
rect 799 -369 833 -335
rect -929 -477 -895 -443
rect -737 -477 -703 -443
rect -545 -477 -511 -443
rect -353 -477 -319 -443
rect -161 -477 -127 -443
rect 31 -477 65 -443
rect 223 -477 257 -443
rect 415 -477 449 -443
rect 607 -477 641 -443
rect 799 -477 833 -443
rect -977 -682 -943 -536
rect -881 -682 -847 -536
rect -785 -682 -751 -536
rect -689 -682 -655 -536
rect -593 -682 -559 -536
rect -497 -682 -463 -536
rect -401 -682 -367 -536
rect -305 -682 -271 -536
rect -209 -682 -175 -536
rect -113 -682 -79 -536
rect -17 -682 17 -536
rect 79 -682 113 -536
rect 175 -682 209 -536
rect 271 -682 305 -536
rect 367 -682 401 -536
rect 463 -682 497 -536
rect 559 -682 593 -536
rect 655 -682 689 -536
rect 751 -682 785 -536
rect 847 -682 881 -536
rect 943 -682 977 -536
rect -833 -775 -799 -741
rect -641 -775 -607 -741
rect -449 -775 -415 -741
rect -257 -775 -223 -741
rect -65 -775 -31 -741
rect 127 -775 161 -741
rect 319 -775 353 -741
rect 511 -775 545 -741
rect 703 -775 737 -741
rect 895 -775 929 -741
rect -833 -883 -799 -849
rect -641 -883 -607 -849
rect -449 -883 -415 -849
rect -257 -883 -223 -849
rect -65 -883 -31 -849
rect 127 -883 161 -849
rect 319 -883 353 -849
rect 511 -883 545 -849
rect 703 -883 737 -849
rect 895 -883 929 -849
rect -977 -1088 -943 -942
rect -881 -1088 -847 -942
rect -785 -1088 -751 -942
rect -689 -1088 -655 -942
rect -593 -1088 -559 -942
rect -497 -1088 -463 -942
rect -401 -1088 -367 -942
rect -305 -1088 -271 -942
rect -209 -1088 -175 -942
rect -113 -1088 -79 -942
rect -17 -1088 17 -942
rect 79 -1088 113 -942
rect 175 -1088 209 -942
rect 271 -1088 305 -942
rect 367 -1088 401 -942
rect 463 -1088 497 -942
rect 559 -1088 593 -942
rect 655 -1088 689 -942
rect 751 -1088 785 -942
rect 847 -1088 881 -942
rect 943 -1088 977 -942
rect -929 -1181 -895 -1147
rect -737 -1181 -703 -1147
rect -545 -1181 -511 -1147
rect -353 -1181 -319 -1147
rect -161 -1181 -127 -1147
rect 31 -1181 65 -1147
rect 223 -1181 257 -1147
rect 415 -1181 449 -1147
rect 607 -1181 641 -1147
rect 799 -1181 833 -1147
rect -929 -1289 -895 -1255
rect -737 -1289 -703 -1255
rect -545 -1289 -511 -1255
rect -353 -1289 -319 -1255
rect -161 -1289 -127 -1255
rect 31 -1289 65 -1255
rect 223 -1289 257 -1255
rect 415 -1289 449 -1255
rect 607 -1289 641 -1255
rect 799 -1289 833 -1255
rect -977 -1494 -943 -1348
rect -881 -1494 -847 -1348
rect -785 -1494 -751 -1348
rect -689 -1494 -655 -1348
rect -593 -1494 -559 -1348
rect -497 -1494 -463 -1348
rect -401 -1494 -367 -1348
rect -305 -1494 -271 -1348
rect -209 -1494 -175 -1348
rect -113 -1494 -79 -1348
rect -17 -1494 17 -1348
rect 79 -1494 113 -1348
rect 175 -1494 209 -1348
rect 271 -1494 305 -1348
rect 367 -1494 401 -1348
rect 463 -1494 497 -1348
rect 559 -1494 593 -1348
rect 655 -1494 689 -1348
rect 751 -1494 785 -1348
rect 847 -1494 881 -1348
rect 943 -1494 977 -1348
rect -833 -1587 -799 -1553
rect -641 -1587 -607 -1553
rect -449 -1587 -415 -1553
rect -257 -1587 -223 -1553
rect -65 -1587 -31 -1553
rect 127 -1587 161 -1553
rect 319 -1587 353 -1553
rect 511 -1587 545 -1553
rect 703 -1587 737 -1553
rect 895 -1587 929 -1553
rect -833 -1695 -799 -1661
rect -641 -1695 -607 -1661
rect -449 -1695 -415 -1661
rect -257 -1695 -223 -1661
rect -65 -1695 -31 -1661
rect 127 -1695 161 -1661
rect 319 -1695 353 -1661
rect 511 -1695 545 -1661
rect 703 -1695 737 -1661
rect 895 -1695 929 -1661
rect -977 -1900 -943 -1754
rect -881 -1900 -847 -1754
rect -785 -1900 -751 -1754
rect -689 -1900 -655 -1754
rect -593 -1900 -559 -1754
rect -497 -1900 -463 -1754
rect -401 -1900 -367 -1754
rect -305 -1900 -271 -1754
rect -209 -1900 -175 -1754
rect -113 -1900 -79 -1754
rect -17 -1900 17 -1754
rect 79 -1900 113 -1754
rect 175 -1900 209 -1754
rect 271 -1900 305 -1754
rect 367 -1900 401 -1754
rect 463 -1900 497 -1754
rect 559 -1900 593 -1754
rect 655 -1900 689 -1754
rect 751 -1900 785 -1754
rect 847 -1900 881 -1754
rect 943 -1900 977 -1754
rect -929 -1993 -895 -1959
rect -737 -1993 -703 -1959
rect -545 -1993 -511 -1959
rect -353 -1993 -319 -1959
rect -161 -1993 -127 -1959
rect 31 -1993 65 -1959
rect 223 -1993 257 -1959
rect 415 -1993 449 -1959
rect 607 -1993 641 -1959
rect 799 -1993 833 -1959
<< metal1 >>
rect -941 1993 -883 1999
rect -941 1959 -929 1993
rect -895 1959 -883 1993
rect -941 1953 -883 1959
rect -749 1993 -691 1999
rect -749 1959 -737 1993
rect -703 1959 -691 1993
rect -749 1953 -691 1959
rect -557 1993 -499 1999
rect -557 1959 -545 1993
rect -511 1959 -499 1993
rect -557 1953 -499 1959
rect -365 1993 -307 1999
rect -365 1959 -353 1993
rect -319 1959 -307 1993
rect -365 1953 -307 1959
rect -173 1993 -115 1999
rect -173 1959 -161 1993
rect -127 1959 -115 1993
rect -173 1953 -115 1959
rect 19 1993 77 1999
rect 19 1959 31 1993
rect 65 1959 77 1993
rect 19 1953 77 1959
rect 211 1993 269 1999
rect 211 1959 223 1993
rect 257 1959 269 1993
rect 211 1953 269 1959
rect 403 1993 461 1999
rect 403 1959 415 1993
rect 449 1959 461 1993
rect 403 1953 461 1959
rect 595 1993 653 1999
rect 595 1959 607 1993
rect 641 1959 653 1993
rect 595 1953 653 1959
rect 787 1993 845 1999
rect 787 1959 799 1993
rect 833 1959 845 1993
rect 787 1953 845 1959
rect -983 1900 -937 1912
rect -983 1754 -977 1900
rect -943 1754 -937 1900
rect -983 1742 -937 1754
rect -887 1900 -841 1912
rect -887 1754 -881 1900
rect -847 1754 -841 1900
rect -887 1742 -841 1754
rect -791 1900 -745 1912
rect -791 1754 -785 1900
rect -751 1754 -745 1900
rect -791 1742 -745 1754
rect -695 1900 -649 1912
rect -695 1754 -689 1900
rect -655 1754 -649 1900
rect -695 1742 -649 1754
rect -599 1900 -553 1912
rect -599 1754 -593 1900
rect -559 1754 -553 1900
rect -599 1742 -553 1754
rect -503 1900 -457 1912
rect -503 1754 -497 1900
rect -463 1754 -457 1900
rect -503 1742 -457 1754
rect -407 1900 -361 1912
rect -407 1754 -401 1900
rect -367 1754 -361 1900
rect -407 1742 -361 1754
rect -311 1900 -265 1912
rect -311 1754 -305 1900
rect -271 1754 -265 1900
rect -311 1742 -265 1754
rect -215 1900 -169 1912
rect -215 1754 -209 1900
rect -175 1754 -169 1900
rect -215 1742 -169 1754
rect -119 1900 -73 1912
rect -119 1754 -113 1900
rect -79 1754 -73 1900
rect -119 1742 -73 1754
rect -23 1900 23 1912
rect -23 1754 -17 1900
rect 17 1754 23 1900
rect -23 1742 23 1754
rect 73 1900 119 1912
rect 73 1754 79 1900
rect 113 1754 119 1900
rect 73 1742 119 1754
rect 169 1900 215 1912
rect 169 1754 175 1900
rect 209 1754 215 1900
rect 169 1742 215 1754
rect 265 1900 311 1912
rect 265 1754 271 1900
rect 305 1754 311 1900
rect 265 1742 311 1754
rect 361 1900 407 1912
rect 361 1754 367 1900
rect 401 1754 407 1900
rect 361 1742 407 1754
rect 457 1900 503 1912
rect 457 1754 463 1900
rect 497 1754 503 1900
rect 457 1742 503 1754
rect 553 1900 599 1912
rect 553 1754 559 1900
rect 593 1754 599 1900
rect 553 1742 599 1754
rect 649 1900 695 1912
rect 649 1754 655 1900
rect 689 1754 695 1900
rect 649 1742 695 1754
rect 745 1900 791 1912
rect 745 1754 751 1900
rect 785 1754 791 1900
rect 745 1742 791 1754
rect 841 1900 887 1912
rect 841 1754 847 1900
rect 881 1754 887 1900
rect 841 1742 887 1754
rect 937 1900 983 1912
rect 937 1754 943 1900
rect 977 1754 983 1900
rect 937 1742 983 1754
rect -845 1695 -787 1701
rect -845 1661 -833 1695
rect -799 1661 -787 1695
rect -845 1655 -787 1661
rect -653 1695 -595 1701
rect -653 1661 -641 1695
rect -607 1661 -595 1695
rect -653 1655 -595 1661
rect -461 1695 -403 1701
rect -461 1661 -449 1695
rect -415 1661 -403 1695
rect -461 1655 -403 1661
rect -269 1695 -211 1701
rect -269 1661 -257 1695
rect -223 1661 -211 1695
rect -269 1655 -211 1661
rect -77 1695 -19 1701
rect -77 1661 -65 1695
rect -31 1661 -19 1695
rect -77 1655 -19 1661
rect 115 1695 173 1701
rect 115 1661 127 1695
rect 161 1661 173 1695
rect 115 1655 173 1661
rect 307 1695 365 1701
rect 307 1661 319 1695
rect 353 1661 365 1695
rect 307 1655 365 1661
rect 499 1695 557 1701
rect 499 1661 511 1695
rect 545 1661 557 1695
rect 499 1655 557 1661
rect 691 1695 749 1701
rect 691 1661 703 1695
rect 737 1661 749 1695
rect 691 1655 749 1661
rect 883 1695 941 1701
rect 883 1661 895 1695
rect 929 1661 941 1695
rect 883 1655 941 1661
rect -845 1587 -787 1593
rect -845 1553 -833 1587
rect -799 1553 -787 1587
rect -845 1547 -787 1553
rect -653 1587 -595 1593
rect -653 1553 -641 1587
rect -607 1553 -595 1587
rect -653 1547 -595 1553
rect -461 1587 -403 1593
rect -461 1553 -449 1587
rect -415 1553 -403 1587
rect -461 1547 -403 1553
rect -269 1587 -211 1593
rect -269 1553 -257 1587
rect -223 1553 -211 1587
rect -269 1547 -211 1553
rect -77 1587 -19 1593
rect -77 1553 -65 1587
rect -31 1553 -19 1587
rect -77 1547 -19 1553
rect 115 1587 173 1593
rect 115 1553 127 1587
rect 161 1553 173 1587
rect 115 1547 173 1553
rect 307 1587 365 1593
rect 307 1553 319 1587
rect 353 1553 365 1587
rect 307 1547 365 1553
rect 499 1587 557 1593
rect 499 1553 511 1587
rect 545 1553 557 1587
rect 499 1547 557 1553
rect 691 1587 749 1593
rect 691 1553 703 1587
rect 737 1553 749 1587
rect 691 1547 749 1553
rect 883 1587 941 1593
rect 883 1553 895 1587
rect 929 1553 941 1587
rect 883 1547 941 1553
rect -983 1494 -937 1506
rect -983 1348 -977 1494
rect -943 1348 -937 1494
rect -983 1336 -937 1348
rect -887 1494 -841 1506
rect -887 1348 -881 1494
rect -847 1348 -841 1494
rect -887 1336 -841 1348
rect -791 1494 -745 1506
rect -791 1348 -785 1494
rect -751 1348 -745 1494
rect -791 1336 -745 1348
rect -695 1494 -649 1506
rect -695 1348 -689 1494
rect -655 1348 -649 1494
rect -695 1336 -649 1348
rect -599 1494 -553 1506
rect -599 1348 -593 1494
rect -559 1348 -553 1494
rect -599 1336 -553 1348
rect -503 1494 -457 1506
rect -503 1348 -497 1494
rect -463 1348 -457 1494
rect -503 1336 -457 1348
rect -407 1494 -361 1506
rect -407 1348 -401 1494
rect -367 1348 -361 1494
rect -407 1336 -361 1348
rect -311 1494 -265 1506
rect -311 1348 -305 1494
rect -271 1348 -265 1494
rect -311 1336 -265 1348
rect -215 1494 -169 1506
rect -215 1348 -209 1494
rect -175 1348 -169 1494
rect -215 1336 -169 1348
rect -119 1494 -73 1506
rect -119 1348 -113 1494
rect -79 1348 -73 1494
rect -119 1336 -73 1348
rect -23 1494 23 1506
rect -23 1348 -17 1494
rect 17 1348 23 1494
rect -23 1336 23 1348
rect 73 1494 119 1506
rect 73 1348 79 1494
rect 113 1348 119 1494
rect 73 1336 119 1348
rect 169 1494 215 1506
rect 169 1348 175 1494
rect 209 1348 215 1494
rect 169 1336 215 1348
rect 265 1494 311 1506
rect 265 1348 271 1494
rect 305 1348 311 1494
rect 265 1336 311 1348
rect 361 1494 407 1506
rect 361 1348 367 1494
rect 401 1348 407 1494
rect 361 1336 407 1348
rect 457 1494 503 1506
rect 457 1348 463 1494
rect 497 1348 503 1494
rect 457 1336 503 1348
rect 553 1494 599 1506
rect 553 1348 559 1494
rect 593 1348 599 1494
rect 553 1336 599 1348
rect 649 1494 695 1506
rect 649 1348 655 1494
rect 689 1348 695 1494
rect 649 1336 695 1348
rect 745 1494 791 1506
rect 745 1348 751 1494
rect 785 1348 791 1494
rect 745 1336 791 1348
rect 841 1494 887 1506
rect 841 1348 847 1494
rect 881 1348 887 1494
rect 841 1336 887 1348
rect 937 1494 983 1506
rect 937 1348 943 1494
rect 977 1348 983 1494
rect 937 1336 983 1348
rect -941 1289 -883 1295
rect -941 1255 -929 1289
rect -895 1255 -883 1289
rect -941 1249 -883 1255
rect -749 1289 -691 1295
rect -749 1255 -737 1289
rect -703 1255 -691 1289
rect -749 1249 -691 1255
rect -557 1289 -499 1295
rect -557 1255 -545 1289
rect -511 1255 -499 1289
rect -557 1249 -499 1255
rect -365 1289 -307 1295
rect -365 1255 -353 1289
rect -319 1255 -307 1289
rect -365 1249 -307 1255
rect -173 1289 -115 1295
rect -173 1255 -161 1289
rect -127 1255 -115 1289
rect -173 1249 -115 1255
rect 19 1289 77 1295
rect 19 1255 31 1289
rect 65 1255 77 1289
rect 19 1249 77 1255
rect 211 1289 269 1295
rect 211 1255 223 1289
rect 257 1255 269 1289
rect 211 1249 269 1255
rect 403 1289 461 1295
rect 403 1255 415 1289
rect 449 1255 461 1289
rect 403 1249 461 1255
rect 595 1289 653 1295
rect 595 1255 607 1289
rect 641 1255 653 1289
rect 595 1249 653 1255
rect 787 1289 845 1295
rect 787 1255 799 1289
rect 833 1255 845 1289
rect 787 1249 845 1255
rect -941 1181 -883 1187
rect -941 1147 -929 1181
rect -895 1147 -883 1181
rect -941 1141 -883 1147
rect -749 1181 -691 1187
rect -749 1147 -737 1181
rect -703 1147 -691 1181
rect -749 1141 -691 1147
rect -557 1181 -499 1187
rect -557 1147 -545 1181
rect -511 1147 -499 1181
rect -557 1141 -499 1147
rect -365 1181 -307 1187
rect -365 1147 -353 1181
rect -319 1147 -307 1181
rect -365 1141 -307 1147
rect -173 1181 -115 1187
rect -173 1147 -161 1181
rect -127 1147 -115 1181
rect -173 1141 -115 1147
rect 19 1181 77 1187
rect 19 1147 31 1181
rect 65 1147 77 1181
rect 19 1141 77 1147
rect 211 1181 269 1187
rect 211 1147 223 1181
rect 257 1147 269 1181
rect 211 1141 269 1147
rect 403 1181 461 1187
rect 403 1147 415 1181
rect 449 1147 461 1181
rect 403 1141 461 1147
rect 595 1181 653 1187
rect 595 1147 607 1181
rect 641 1147 653 1181
rect 595 1141 653 1147
rect 787 1181 845 1187
rect 787 1147 799 1181
rect 833 1147 845 1181
rect 787 1141 845 1147
rect -983 1088 -937 1100
rect -983 942 -977 1088
rect -943 942 -937 1088
rect -983 930 -937 942
rect -887 1088 -841 1100
rect -887 942 -881 1088
rect -847 942 -841 1088
rect -887 930 -841 942
rect -791 1088 -745 1100
rect -791 942 -785 1088
rect -751 942 -745 1088
rect -791 930 -745 942
rect -695 1088 -649 1100
rect -695 942 -689 1088
rect -655 942 -649 1088
rect -695 930 -649 942
rect -599 1088 -553 1100
rect -599 942 -593 1088
rect -559 942 -553 1088
rect -599 930 -553 942
rect -503 1088 -457 1100
rect -503 942 -497 1088
rect -463 942 -457 1088
rect -503 930 -457 942
rect -407 1088 -361 1100
rect -407 942 -401 1088
rect -367 942 -361 1088
rect -407 930 -361 942
rect -311 1088 -265 1100
rect -311 942 -305 1088
rect -271 942 -265 1088
rect -311 930 -265 942
rect -215 1088 -169 1100
rect -215 942 -209 1088
rect -175 942 -169 1088
rect -215 930 -169 942
rect -119 1088 -73 1100
rect -119 942 -113 1088
rect -79 942 -73 1088
rect -119 930 -73 942
rect -23 1088 23 1100
rect -23 942 -17 1088
rect 17 942 23 1088
rect -23 930 23 942
rect 73 1088 119 1100
rect 73 942 79 1088
rect 113 942 119 1088
rect 73 930 119 942
rect 169 1088 215 1100
rect 169 942 175 1088
rect 209 942 215 1088
rect 169 930 215 942
rect 265 1088 311 1100
rect 265 942 271 1088
rect 305 942 311 1088
rect 265 930 311 942
rect 361 1088 407 1100
rect 361 942 367 1088
rect 401 942 407 1088
rect 361 930 407 942
rect 457 1088 503 1100
rect 457 942 463 1088
rect 497 942 503 1088
rect 457 930 503 942
rect 553 1088 599 1100
rect 553 942 559 1088
rect 593 942 599 1088
rect 553 930 599 942
rect 649 1088 695 1100
rect 649 942 655 1088
rect 689 942 695 1088
rect 649 930 695 942
rect 745 1088 791 1100
rect 745 942 751 1088
rect 785 942 791 1088
rect 745 930 791 942
rect 841 1088 887 1100
rect 841 942 847 1088
rect 881 942 887 1088
rect 841 930 887 942
rect 937 1088 983 1100
rect 937 942 943 1088
rect 977 942 983 1088
rect 937 930 983 942
rect -845 883 -787 889
rect -845 849 -833 883
rect -799 849 -787 883
rect -845 843 -787 849
rect -653 883 -595 889
rect -653 849 -641 883
rect -607 849 -595 883
rect -653 843 -595 849
rect -461 883 -403 889
rect -461 849 -449 883
rect -415 849 -403 883
rect -461 843 -403 849
rect -269 883 -211 889
rect -269 849 -257 883
rect -223 849 -211 883
rect -269 843 -211 849
rect -77 883 -19 889
rect -77 849 -65 883
rect -31 849 -19 883
rect -77 843 -19 849
rect 115 883 173 889
rect 115 849 127 883
rect 161 849 173 883
rect 115 843 173 849
rect 307 883 365 889
rect 307 849 319 883
rect 353 849 365 883
rect 307 843 365 849
rect 499 883 557 889
rect 499 849 511 883
rect 545 849 557 883
rect 499 843 557 849
rect 691 883 749 889
rect 691 849 703 883
rect 737 849 749 883
rect 691 843 749 849
rect 883 883 941 889
rect 883 849 895 883
rect 929 849 941 883
rect 883 843 941 849
rect -845 775 -787 781
rect -845 741 -833 775
rect -799 741 -787 775
rect -845 735 -787 741
rect -653 775 -595 781
rect -653 741 -641 775
rect -607 741 -595 775
rect -653 735 -595 741
rect -461 775 -403 781
rect -461 741 -449 775
rect -415 741 -403 775
rect -461 735 -403 741
rect -269 775 -211 781
rect -269 741 -257 775
rect -223 741 -211 775
rect -269 735 -211 741
rect -77 775 -19 781
rect -77 741 -65 775
rect -31 741 -19 775
rect -77 735 -19 741
rect 115 775 173 781
rect 115 741 127 775
rect 161 741 173 775
rect 115 735 173 741
rect 307 775 365 781
rect 307 741 319 775
rect 353 741 365 775
rect 307 735 365 741
rect 499 775 557 781
rect 499 741 511 775
rect 545 741 557 775
rect 499 735 557 741
rect 691 775 749 781
rect 691 741 703 775
rect 737 741 749 775
rect 691 735 749 741
rect 883 775 941 781
rect 883 741 895 775
rect 929 741 941 775
rect 883 735 941 741
rect -983 682 -937 694
rect -983 536 -977 682
rect -943 536 -937 682
rect -983 524 -937 536
rect -887 682 -841 694
rect -887 536 -881 682
rect -847 536 -841 682
rect -887 524 -841 536
rect -791 682 -745 694
rect -791 536 -785 682
rect -751 536 -745 682
rect -791 524 -745 536
rect -695 682 -649 694
rect -695 536 -689 682
rect -655 536 -649 682
rect -695 524 -649 536
rect -599 682 -553 694
rect -599 536 -593 682
rect -559 536 -553 682
rect -599 524 -553 536
rect -503 682 -457 694
rect -503 536 -497 682
rect -463 536 -457 682
rect -503 524 -457 536
rect -407 682 -361 694
rect -407 536 -401 682
rect -367 536 -361 682
rect -407 524 -361 536
rect -311 682 -265 694
rect -311 536 -305 682
rect -271 536 -265 682
rect -311 524 -265 536
rect -215 682 -169 694
rect -215 536 -209 682
rect -175 536 -169 682
rect -215 524 -169 536
rect -119 682 -73 694
rect -119 536 -113 682
rect -79 536 -73 682
rect -119 524 -73 536
rect -23 682 23 694
rect -23 536 -17 682
rect 17 536 23 682
rect -23 524 23 536
rect 73 682 119 694
rect 73 536 79 682
rect 113 536 119 682
rect 73 524 119 536
rect 169 682 215 694
rect 169 536 175 682
rect 209 536 215 682
rect 169 524 215 536
rect 265 682 311 694
rect 265 536 271 682
rect 305 536 311 682
rect 265 524 311 536
rect 361 682 407 694
rect 361 536 367 682
rect 401 536 407 682
rect 361 524 407 536
rect 457 682 503 694
rect 457 536 463 682
rect 497 536 503 682
rect 457 524 503 536
rect 553 682 599 694
rect 553 536 559 682
rect 593 536 599 682
rect 553 524 599 536
rect 649 682 695 694
rect 649 536 655 682
rect 689 536 695 682
rect 649 524 695 536
rect 745 682 791 694
rect 745 536 751 682
rect 785 536 791 682
rect 745 524 791 536
rect 841 682 887 694
rect 841 536 847 682
rect 881 536 887 682
rect 841 524 887 536
rect 937 682 983 694
rect 937 536 943 682
rect 977 536 983 682
rect 937 524 983 536
rect -941 477 -883 483
rect -941 443 -929 477
rect -895 443 -883 477
rect -941 437 -883 443
rect -749 477 -691 483
rect -749 443 -737 477
rect -703 443 -691 477
rect -749 437 -691 443
rect -557 477 -499 483
rect -557 443 -545 477
rect -511 443 -499 477
rect -557 437 -499 443
rect -365 477 -307 483
rect -365 443 -353 477
rect -319 443 -307 477
rect -365 437 -307 443
rect -173 477 -115 483
rect -173 443 -161 477
rect -127 443 -115 477
rect -173 437 -115 443
rect 19 477 77 483
rect 19 443 31 477
rect 65 443 77 477
rect 19 437 77 443
rect 211 477 269 483
rect 211 443 223 477
rect 257 443 269 477
rect 211 437 269 443
rect 403 477 461 483
rect 403 443 415 477
rect 449 443 461 477
rect 403 437 461 443
rect 595 477 653 483
rect 595 443 607 477
rect 641 443 653 477
rect 595 437 653 443
rect 787 477 845 483
rect 787 443 799 477
rect 833 443 845 477
rect 787 437 845 443
rect -941 369 -883 375
rect -941 335 -929 369
rect -895 335 -883 369
rect -941 329 -883 335
rect -749 369 -691 375
rect -749 335 -737 369
rect -703 335 -691 369
rect -749 329 -691 335
rect -557 369 -499 375
rect -557 335 -545 369
rect -511 335 -499 369
rect -557 329 -499 335
rect -365 369 -307 375
rect -365 335 -353 369
rect -319 335 -307 369
rect -365 329 -307 335
rect -173 369 -115 375
rect -173 335 -161 369
rect -127 335 -115 369
rect -173 329 -115 335
rect 19 369 77 375
rect 19 335 31 369
rect 65 335 77 369
rect 19 329 77 335
rect 211 369 269 375
rect 211 335 223 369
rect 257 335 269 369
rect 211 329 269 335
rect 403 369 461 375
rect 403 335 415 369
rect 449 335 461 369
rect 403 329 461 335
rect 595 369 653 375
rect 595 335 607 369
rect 641 335 653 369
rect 595 329 653 335
rect 787 369 845 375
rect 787 335 799 369
rect 833 335 845 369
rect 787 329 845 335
rect -983 276 -937 288
rect -983 130 -977 276
rect -943 130 -937 276
rect -983 118 -937 130
rect -887 276 -841 288
rect -887 130 -881 276
rect -847 130 -841 276
rect -887 118 -841 130
rect -791 276 -745 288
rect -791 130 -785 276
rect -751 130 -745 276
rect -791 118 -745 130
rect -695 276 -649 288
rect -695 130 -689 276
rect -655 130 -649 276
rect -695 118 -649 130
rect -599 276 -553 288
rect -599 130 -593 276
rect -559 130 -553 276
rect -599 118 -553 130
rect -503 276 -457 288
rect -503 130 -497 276
rect -463 130 -457 276
rect -503 118 -457 130
rect -407 276 -361 288
rect -407 130 -401 276
rect -367 130 -361 276
rect -407 118 -361 130
rect -311 276 -265 288
rect -311 130 -305 276
rect -271 130 -265 276
rect -311 118 -265 130
rect -215 276 -169 288
rect -215 130 -209 276
rect -175 130 -169 276
rect -215 118 -169 130
rect -119 276 -73 288
rect -119 130 -113 276
rect -79 130 -73 276
rect -119 118 -73 130
rect -23 276 23 288
rect -23 130 -17 276
rect 17 130 23 276
rect -23 118 23 130
rect 73 276 119 288
rect 73 130 79 276
rect 113 130 119 276
rect 73 118 119 130
rect 169 276 215 288
rect 169 130 175 276
rect 209 130 215 276
rect 169 118 215 130
rect 265 276 311 288
rect 265 130 271 276
rect 305 130 311 276
rect 265 118 311 130
rect 361 276 407 288
rect 361 130 367 276
rect 401 130 407 276
rect 361 118 407 130
rect 457 276 503 288
rect 457 130 463 276
rect 497 130 503 276
rect 457 118 503 130
rect 553 276 599 288
rect 553 130 559 276
rect 593 130 599 276
rect 553 118 599 130
rect 649 276 695 288
rect 649 130 655 276
rect 689 130 695 276
rect 649 118 695 130
rect 745 276 791 288
rect 745 130 751 276
rect 785 130 791 276
rect 745 118 791 130
rect 841 276 887 288
rect 841 130 847 276
rect 881 130 887 276
rect 841 118 887 130
rect 937 276 983 288
rect 937 130 943 276
rect 977 130 983 276
rect 937 118 983 130
rect -845 71 -787 77
rect -845 37 -833 71
rect -799 37 -787 71
rect -845 31 -787 37
rect -653 71 -595 77
rect -653 37 -641 71
rect -607 37 -595 71
rect -653 31 -595 37
rect -461 71 -403 77
rect -461 37 -449 71
rect -415 37 -403 71
rect -461 31 -403 37
rect -269 71 -211 77
rect -269 37 -257 71
rect -223 37 -211 71
rect -269 31 -211 37
rect -77 71 -19 77
rect -77 37 -65 71
rect -31 37 -19 71
rect -77 31 -19 37
rect 115 71 173 77
rect 115 37 127 71
rect 161 37 173 71
rect 115 31 173 37
rect 307 71 365 77
rect 307 37 319 71
rect 353 37 365 71
rect 307 31 365 37
rect 499 71 557 77
rect 499 37 511 71
rect 545 37 557 71
rect 499 31 557 37
rect 691 71 749 77
rect 691 37 703 71
rect 737 37 749 71
rect 691 31 749 37
rect 883 71 941 77
rect 883 37 895 71
rect 929 37 941 71
rect 883 31 941 37
rect -845 -37 -787 -31
rect -845 -71 -833 -37
rect -799 -71 -787 -37
rect -845 -77 -787 -71
rect -653 -37 -595 -31
rect -653 -71 -641 -37
rect -607 -71 -595 -37
rect -653 -77 -595 -71
rect -461 -37 -403 -31
rect -461 -71 -449 -37
rect -415 -71 -403 -37
rect -461 -77 -403 -71
rect -269 -37 -211 -31
rect -269 -71 -257 -37
rect -223 -71 -211 -37
rect -269 -77 -211 -71
rect -77 -37 -19 -31
rect -77 -71 -65 -37
rect -31 -71 -19 -37
rect -77 -77 -19 -71
rect 115 -37 173 -31
rect 115 -71 127 -37
rect 161 -71 173 -37
rect 115 -77 173 -71
rect 307 -37 365 -31
rect 307 -71 319 -37
rect 353 -71 365 -37
rect 307 -77 365 -71
rect 499 -37 557 -31
rect 499 -71 511 -37
rect 545 -71 557 -37
rect 499 -77 557 -71
rect 691 -37 749 -31
rect 691 -71 703 -37
rect 737 -71 749 -37
rect 691 -77 749 -71
rect 883 -37 941 -31
rect 883 -71 895 -37
rect 929 -71 941 -37
rect 883 -77 941 -71
rect -983 -130 -937 -118
rect -983 -276 -977 -130
rect -943 -276 -937 -130
rect -983 -288 -937 -276
rect -887 -130 -841 -118
rect -887 -276 -881 -130
rect -847 -276 -841 -130
rect -887 -288 -841 -276
rect -791 -130 -745 -118
rect -791 -276 -785 -130
rect -751 -276 -745 -130
rect -791 -288 -745 -276
rect -695 -130 -649 -118
rect -695 -276 -689 -130
rect -655 -276 -649 -130
rect -695 -288 -649 -276
rect -599 -130 -553 -118
rect -599 -276 -593 -130
rect -559 -276 -553 -130
rect -599 -288 -553 -276
rect -503 -130 -457 -118
rect -503 -276 -497 -130
rect -463 -276 -457 -130
rect -503 -288 -457 -276
rect -407 -130 -361 -118
rect -407 -276 -401 -130
rect -367 -276 -361 -130
rect -407 -288 -361 -276
rect -311 -130 -265 -118
rect -311 -276 -305 -130
rect -271 -276 -265 -130
rect -311 -288 -265 -276
rect -215 -130 -169 -118
rect -215 -276 -209 -130
rect -175 -276 -169 -130
rect -215 -288 -169 -276
rect -119 -130 -73 -118
rect -119 -276 -113 -130
rect -79 -276 -73 -130
rect -119 -288 -73 -276
rect -23 -130 23 -118
rect -23 -276 -17 -130
rect 17 -276 23 -130
rect -23 -288 23 -276
rect 73 -130 119 -118
rect 73 -276 79 -130
rect 113 -276 119 -130
rect 73 -288 119 -276
rect 169 -130 215 -118
rect 169 -276 175 -130
rect 209 -276 215 -130
rect 169 -288 215 -276
rect 265 -130 311 -118
rect 265 -276 271 -130
rect 305 -276 311 -130
rect 265 -288 311 -276
rect 361 -130 407 -118
rect 361 -276 367 -130
rect 401 -276 407 -130
rect 361 -288 407 -276
rect 457 -130 503 -118
rect 457 -276 463 -130
rect 497 -276 503 -130
rect 457 -288 503 -276
rect 553 -130 599 -118
rect 553 -276 559 -130
rect 593 -276 599 -130
rect 553 -288 599 -276
rect 649 -130 695 -118
rect 649 -276 655 -130
rect 689 -276 695 -130
rect 649 -288 695 -276
rect 745 -130 791 -118
rect 745 -276 751 -130
rect 785 -276 791 -130
rect 745 -288 791 -276
rect 841 -130 887 -118
rect 841 -276 847 -130
rect 881 -276 887 -130
rect 841 -288 887 -276
rect 937 -130 983 -118
rect 937 -276 943 -130
rect 977 -276 983 -130
rect 937 -288 983 -276
rect -941 -335 -883 -329
rect -941 -369 -929 -335
rect -895 -369 -883 -335
rect -941 -375 -883 -369
rect -749 -335 -691 -329
rect -749 -369 -737 -335
rect -703 -369 -691 -335
rect -749 -375 -691 -369
rect -557 -335 -499 -329
rect -557 -369 -545 -335
rect -511 -369 -499 -335
rect -557 -375 -499 -369
rect -365 -335 -307 -329
rect -365 -369 -353 -335
rect -319 -369 -307 -335
rect -365 -375 -307 -369
rect -173 -335 -115 -329
rect -173 -369 -161 -335
rect -127 -369 -115 -335
rect -173 -375 -115 -369
rect 19 -335 77 -329
rect 19 -369 31 -335
rect 65 -369 77 -335
rect 19 -375 77 -369
rect 211 -335 269 -329
rect 211 -369 223 -335
rect 257 -369 269 -335
rect 211 -375 269 -369
rect 403 -335 461 -329
rect 403 -369 415 -335
rect 449 -369 461 -335
rect 403 -375 461 -369
rect 595 -335 653 -329
rect 595 -369 607 -335
rect 641 -369 653 -335
rect 595 -375 653 -369
rect 787 -335 845 -329
rect 787 -369 799 -335
rect 833 -369 845 -335
rect 787 -375 845 -369
rect -941 -443 -883 -437
rect -941 -477 -929 -443
rect -895 -477 -883 -443
rect -941 -483 -883 -477
rect -749 -443 -691 -437
rect -749 -477 -737 -443
rect -703 -477 -691 -443
rect -749 -483 -691 -477
rect -557 -443 -499 -437
rect -557 -477 -545 -443
rect -511 -477 -499 -443
rect -557 -483 -499 -477
rect -365 -443 -307 -437
rect -365 -477 -353 -443
rect -319 -477 -307 -443
rect -365 -483 -307 -477
rect -173 -443 -115 -437
rect -173 -477 -161 -443
rect -127 -477 -115 -443
rect -173 -483 -115 -477
rect 19 -443 77 -437
rect 19 -477 31 -443
rect 65 -477 77 -443
rect 19 -483 77 -477
rect 211 -443 269 -437
rect 211 -477 223 -443
rect 257 -477 269 -443
rect 211 -483 269 -477
rect 403 -443 461 -437
rect 403 -477 415 -443
rect 449 -477 461 -443
rect 403 -483 461 -477
rect 595 -443 653 -437
rect 595 -477 607 -443
rect 641 -477 653 -443
rect 595 -483 653 -477
rect 787 -443 845 -437
rect 787 -477 799 -443
rect 833 -477 845 -443
rect 787 -483 845 -477
rect -983 -536 -937 -524
rect -983 -682 -977 -536
rect -943 -682 -937 -536
rect -983 -694 -937 -682
rect -887 -536 -841 -524
rect -887 -682 -881 -536
rect -847 -682 -841 -536
rect -887 -694 -841 -682
rect -791 -536 -745 -524
rect -791 -682 -785 -536
rect -751 -682 -745 -536
rect -791 -694 -745 -682
rect -695 -536 -649 -524
rect -695 -682 -689 -536
rect -655 -682 -649 -536
rect -695 -694 -649 -682
rect -599 -536 -553 -524
rect -599 -682 -593 -536
rect -559 -682 -553 -536
rect -599 -694 -553 -682
rect -503 -536 -457 -524
rect -503 -682 -497 -536
rect -463 -682 -457 -536
rect -503 -694 -457 -682
rect -407 -536 -361 -524
rect -407 -682 -401 -536
rect -367 -682 -361 -536
rect -407 -694 -361 -682
rect -311 -536 -265 -524
rect -311 -682 -305 -536
rect -271 -682 -265 -536
rect -311 -694 -265 -682
rect -215 -536 -169 -524
rect -215 -682 -209 -536
rect -175 -682 -169 -536
rect -215 -694 -169 -682
rect -119 -536 -73 -524
rect -119 -682 -113 -536
rect -79 -682 -73 -536
rect -119 -694 -73 -682
rect -23 -536 23 -524
rect -23 -682 -17 -536
rect 17 -682 23 -536
rect -23 -694 23 -682
rect 73 -536 119 -524
rect 73 -682 79 -536
rect 113 -682 119 -536
rect 73 -694 119 -682
rect 169 -536 215 -524
rect 169 -682 175 -536
rect 209 -682 215 -536
rect 169 -694 215 -682
rect 265 -536 311 -524
rect 265 -682 271 -536
rect 305 -682 311 -536
rect 265 -694 311 -682
rect 361 -536 407 -524
rect 361 -682 367 -536
rect 401 -682 407 -536
rect 361 -694 407 -682
rect 457 -536 503 -524
rect 457 -682 463 -536
rect 497 -682 503 -536
rect 457 -694 503 -682
rect 553 -536 599 -524
rect 553 -682 559 -536
rect 593 -682 599 -536
rect 553 -694 599 -682
rect 649 -536 695 -524
rect 649 -682 655 -536
rect 689 -682 695 -536
rect 649 -694 695 -682
rect 745 -536 791 -524
rect 745 -682 751 -536
rect 785 -682 791 -536
rect 745 -694 791 -682
rect 841 -536 887 -524
rect 841 -682 847 -536
rect 881 -682 887 -536
rect 841 -694 887 -682
rect 937 -536 983 -524
rect 937 -682 943 -536
rect 977 -682 983 -536
rect 937 -694 983 -682
rect -845 -741 -787 -735
rect -845 -775 -833 -741
rect -799 -775 -787 -741
rect -845 -781 -787 -775
rect -653 -741 -595 -735
rect -653 -775 -641 -741
rect -607 -775 -595 -741
rect -653 -781 -595 -775
rect -461 -741 -403 -735
rect -461 -775 -449 -741
rect -415 -775 -403 -741
rect -461 -781 -403 -775
rect -269 -741 -211 -735
rect -269 -775 -257 -741
rect -223 -775 -211 -741
rect -269 -781 -211 -775
rect -77 -741 -19 -735
rect -77 -775 -65 -741
rect -31 -775 -19 -741
rect -77 -781 -19 -775
rect 115 -741 173 -735
rect 115 -775 127 -741
rect 161 -775 173 -741
rect 115 -781 173 -775
rect 307 -741 365 -735
rect 307 -775 319 -741
rect 353 -775 365 -741
rect 307 -781 365 -775
rect 499 -741 557 -735
rect 499 -775 511 -741
rect 545 -775 557 -741
rect 499 -781 557 -775
rect 691 -741 749 -735
rect 691 -775 703 -741
rect 737 -775 749 -741
rect 691 -781 749 -775
rect 883 -741 941 -735
rect 883 -775 895 -741
rect 929 -775 941 -741
rect 883 -781 941 -775
rect -845 -849 -787 -843
rect -845 -883 -833 -849
rect -799 -883 -787 -849
rect -845 -889 -787 -883
rect -653 -849 -595 -843
rect -653 -883 -641 -849
rect -607 -883 -595 -849
rect -653 -889 -595 -883
rect -461 -849 -403 -843
rect -461 -883 -449 -849
rect -415 -883 -403 -849
rect -461 -889 -403 -883
rect -269 -849 -211 -843
rect -269 -883 -257 -849
rect -223 -883 -211 -849
rect -269 -889 -211 -883
rect -77 -849 -19 -843
rect -77 -883 -65 -849
rect -31 -883 -19 -849
rect -77 -889 -19 -883
rect 115 -849 173 -843
rect 115 -883 127 -849
rect 161 -883 173 -849
rect 115 -889 173 -883
rect 307 -849 365 -843
rect 307 -883 319 -849
rect 353 -883 365 -849
rect 307 -889 365 -883
rect 499 -849 557 -843
rect 499 -883 511 -849
rect 545 -883 557 -849
rect 499 -889 557 -883
rect 691 -849 749 -843
rect 691 -883 703 -849
rect 737 -883 749 -849
rect 691 -889 749 -883
rect 883 -849 941 -843
rect 883 -883 895 -849
rect 929 -883 941 -849
rect 883 -889 941 -883
rect -983 -942 -937 -930
rect -983 -1088 -977 -942
rect -943 -1088 -937 -942
rect -983 -1100 -937 -1088
rect -887 -942 -841 -930
rect -887 -1088 -881 -942
rect -847 -1088 -841 -942
rect -887 -1100 -841 -1088
rect -791 -942 -745 -930
rect -791 -1088 -785 -942
rect -751 -1088 -745 -942
rect -791 -1100 -745 -1088
rect -695 -942 -649 -930
rect -695 -1088 -689 -942
rect -655 -1088 -649 -942
rect -695 -1100 -649 -1088
rect -599 -942 -553 -930
rect -599 -1088 -593 -942
rect -559 -1088 -553 -942
rect -599 -1100 -553 -1088
rect -503 -942 -457 -930
rect -503 -1088 -497 -942
rect -463 -1088 -457 -942
rect -503 -1100 -457 -1088
rect -407 -942 -361 -930
rect -407 -1088 -401 -942
rect -367 -1088 -361 -942
rect -407 -1100 -361 -1088
rect -311 -942 -265 -930
rect -311 -1088 -305 -942
rect -271 -1088 -265 -942
rect -311 -1100 -265 -1088
rect -215 -942 -169 -930
rect -215 -1088 -209 -942
rect -175 -1088 -169 -942
rect -215 -1100 -169 -1088
rect -119 -942 -73 -930
rect -119 -1088 -113 -942
rect -79 -1088 -73 -942
rect -119 -1100 -73 -1088
rect -23 -942 23 -930
rect -23 -1088 -17 -942
rect 17 -1088 23 -942
rect -23 -1100 23 -1088
rect 73 -942 119 -930
rect 73 -1088 79 -942
rect 113 -1088 119 -942
rect 73 -1100 119 -1088
rect 169 -942 215 -930
rect 169 -1088 175 -942
rect 209 -1088 215 -942
rect 169 -1100 215 -1088
rect 265 -942 311 -930
rect 265 -1088 271 -942
rect 305 -1088 311 -942
rect 265 -1100 311 -1088
rect 361 -942 407 -930
rect 361 -1088 367 -942
rect 401 -1088 407 -942
rect 361 -1100 407 -1088
rect 457 -942 503 -930
rect 457 -1088 463 -942
rect 497 -1088 503 -942
rect 457 -1100 503 -1088
rect 553 -942 599 -930
rect 553 -1088 559 -942
rect 593 -1088 599 -942
rect 553 -1100 599 -1088
rect 649 -942 695 -930
rect 649 -1088 655 -942
rect 689 -1088 695 -942
rect 649 -1100 695 -1088
rect 745 -942 791 -930
rect 745 -1088 751 -942
rect 785 -1088 791 -942
rect 745 -1100 791 -1088
rect 841 -942 887 -930
rect 841 -1088 847 -942
rect 881 -1088 887 -942
rect 841 -1100 887 -1088
rect 937 -942 983 -930
rect 937 -1088 943 -942
rect 977 -1088 983 -942
rect 937 -1100 983 -1088
rect -941 -1147 -883 -1141
rect -941 -1181 -929 -1147
rect -895 -1181 -883 -1147
rect -941 -1187 -883 -1181
rect -749 -1147 -691 -1141
rect -749 -1181 -737 -1147
rect -703 -1181 -691 -1147
rect -749 -1187 -691 -1181
rect -557 -1147 -499 -1141
rect -557 -1181 -545 -1147
rect -511 -1181 -499 -1147
rect -557 -1187 -499 -1181
rect -365 -1147 -307 -1141
rect -365 -1181 -353 -1147
rect -319 -1181 -307 -1147
rect -365 -1187 -307 -1181
rect -173 -1147 -115 -1141
rect -173 -1181 -161 -1147
rect -127 -1181 -115 -1147
rect -173 -1187 -115 -1181
rect 19 -1147 77 -1141
rect 19 -1181 31 -1147
rect 65 -1181 77 -1147
rect 19 -1187 77 -1181
rect 211 -1147 269 -1141
rect 211 -1181 223 -1147
rect 257 -1181 269 -1147
rect 211 -1187 269 -1181
rect 403 -1147 461 -1141
rect 403 -1181 415 -1147
rect 449 -1181 461 -1147
rect 403 -1187 461 -1181
rect 595 -1147 653 -1141
rect 595 -1181 607 -1147
rect 641 -1181 653 -1147
rect 595 -1187 653 -1181
rect 787 -1147 845 -1141
rect 787 -1181 799 -1147
rect 833 -1181 845 -1147
rect 787 -1187 845 -1181
rect -941 -1255 -883 -1249
rect -941 -1289 -929 -1255
rect -895 -1289 -883 -1255
rect -941 -1295 -883 -1289
rect -749 -1255 -691 -1249
rect -749 -1289 -737 -1255
rect -703 -1289 -691 -1255
rect -749 -1295 -691 -1289
rect -557 -1255 -499 -1249
rect -557 -1289 -545 -1255
rect -511 -1289 -499 -1255
rect -557 -1295 -499 -1289
rect -365 -1255 -307 -1249
rect -365 -1289 -353 -1255
rect -319 -1289 -307 -1255
rect -365 -1295 -307 -1289
rect -173 -1255 -115 -1249
rect -173 -1289 -161 -1255
rect -127 -1289 -115 -1255
rect -173 -1295 -115 -1289
rect 19 -1255 77 -1249
rect 19 -1289 31 -1255
rect 65 -1289 77 -1255
rect 19 -1295 77 -1289
rect 211 -1255 269 -1249
rect 211 -1289 223 -1255
rect 257 -1289 269 -1255
rect 211 -1295 269 -1289
rect 403 -1255 461 -1249
rect 403 -1289 415 -1255
rect 449 -1289 461 -1255
rect 403 -1295 461 -1289
rect 595 -1255 653 -1249
rect 595 -1289 607 -1255
rect 641 -1289 653 -1255
rect 595 -1295 653 -1289
rect 787 -1255 845 -1249
rect 787 -1289 799 -1255
rect 833 -1289 845 -1255
rect 787 -1295 845 -1289
rect -983 -1348 -937 -1336
rect -983 -1494 -977 -1348
rect -943 -1494 -937 -1348
rect -983 -1506 -937 -1494
rect -887 -1348 -841 -1336
rect -887 -1494 -881 -1348
rect -847 -1494 -841 -1348
rect -887 -1506 -841 -1494
rect -791 -1348 -745 -1336
rect -791 -1494 -785 -1348
rect -751 -1494 -745 -1348
rect -791 -1506 -745 -1494
rect -695 -1348 -649 -1336
rect -695 -1494 -689 -1348
rect -655 -1494 -649 -1348
rect -695 -1506 -649 -1494
rect -599 -1348 -553 -1336
rect -599 -1494 -593 -1348
rect -559 -1494 -553 -1348
rect -599 -1506 -553 -1494
rect -503 -1348 -457 -1336
rect -503 -1494 -497 -1348
rect -463 -1494 -457 -1348
rect -503 -1506 -457 -1494
rect -407 -1348 -361 -1336
rect -407 -1494 -401 -1348
rect -367 -1494 -361 -1348
rect -407 -1506 -361 -1494
rect -311 -1348 -265 -1336
rect -311 -1494 -305 -1348
rect -271 -1494 -265 -1348
rect -311 -1506 -265 -1494
rect -215 -1348 -169 -1336
rect -215 -1494 -209 -1348
rect -175 -1494 -169 -1348
rect -215 -1506 -169 -1494
rect -119 -1348 -73 -1336
rect -119 -1494 -113 -1348
rect -79 -1494 -73 -1348
rect -119 -1506 -73 -1494
rect -23 -1348 23 -1336
rect -23 -1494 -17 -1348
rect 17 -1494 23 -1348
rect -23 -1506 23 -1494
rect 73 -1348 119 -1336
rect 73 -1494 79 -1348
rect 113 -1494 119 -1348
rect 73 -1506 119 -1494
rect 169 -1348 215 -1336
rect 169 -1494 175 -1348
rect 209 -1494 215 -1348
rect 169 -1506 215 -1494
rect 265 -1348 311 -1336
rect 265 -1494 271 -1348
rect 305 -1494 311 -1348
rect 265 -1506 311 -1494
rect 361 -1348 407 -1336
rect 361 -1494 367 -1348
rect 401 -1494 407 -1348
rect 361 -1506 407 -1494
rect 457 -1348 503 -1336
rect 457 -1494 463 -1348
rect 497 -1494 503 -1348
rect 457 -1506 503 -1494
rect 553 -1348 599 -1336
rect 553 -1494 559 -1348
rect 593 -1494 599 -1348
rect 553 -1506 599 -1494
rect 649 -1348 695 -1336
rect 649 -1494 655 -1348
rect 689 -1494 695 -1348
rect 649 -1506 695 -1494
rect 745 -1348 791 -1336
rect 745 -1494 751 -1348
rect 785 -1494 791 -1348
rect 745 -1506 791 -1494
rect 841 -1348 887 -1336
rect 841 -1494 847 -1348
rect 881 -1494 887 -1348
rect 841 -1506 887 -1494
rect 937 -1348 983 -1336
rect 937 -1494 943 -1348
rect 977 -1494 983 -1348
rect 937 -1506 983 -1494
rect -845 -1553 -787 -1547
rect -845 -1587 -833 -1553
rect -799 -1587 -787 -1553
rect -845 -1593 -787 -1587
rect -653 -1553 -595 -1547
rect -653 -1587 -641 -1553
rect -607 -1587 -595 -1553
rect -653 -1593 -595 -1587
rect -461 -1553 -403 -1547
rect -461 -1587 -449 -1553
rect -415 -1587 -403 -1553
rect -461 -1593 -403 -1587
rect -269 -1553 -211 -1547
rect -269 -1587 -257 -1553
rect -223 -1587 -211 -1553
rect -269 -1593 -211 -1587
rect -77 -1553 -19 -1547
rect -77 -1587 -65 -1553
rect -31 -1587 -19 -1553
rect -77 -1593 -19 -1587
rect 115 -1553 173 -1547
rect 115 -1587 127 -1553
rect 161 -1587 173 -1553
rect 115 -1593 173 -1587
rect 307 -1553 365 -1547
rect 307 -1587 319 -1553
rect 353 -1587 365 -1553
rect 307 -1593 365 -1587
rect 499 -1553 557 -1547
rect 499 -1587 511 -1553
rect 545 -1587 557 -1553
rect 499 -1593 557 -1587
rect 691 -1553 749 -1547
rect 691 -1587 703 -1553
rect 737 -1587 749 -1553
rect 691 -1593 749 -1587
rect 883 -1553 941 -1547
rect 883 -1587 895 -1553
rect 929 -1587 941 -1553
rect 883 -1593 941 -1587
rect -845 -1661 -787 -1655
rect -845 -1695 -833 -1661
rect -799 -1695 -787 -1661
rect -845 -1701 -787 -1695
rect -653 -1661 -595 -1655
rect -653 -1695 -641 -1661
rect -607 -1695 -595 -1661
rect -653 -1701 -595 -1695
rect -461 -1661 -403 -1655
rect -461 -1695 -449 -1661
rect -415 -1695 -403 -1661
rect -461 -1701 -403 -1695
rect -269 -1661 -211 -1655
rect -269 -1695 -257 -1661
rect -223 -1695 -211 -1661
rect -269 -1701 -211 -1695
rect -77 -1661 -19 -1655
rect -77 -1695 -65 -1661
rect -31 -1695 -19 -1661
rect -77 -1701 -19 -1695
rect 115 -1661 173 -1655
rect 115 -1695 127 -1661
rect 161 -1695 173 -1661
rect 115 -1701 173 -1695
rect 307 -1661 365 -1655
rect 307 -1695 319 -1661
rect 353 -1695 365 -1661
rect 307 -1701 365 -1695
rect 499 -1661 557 -1655
rect 499 -1695 511 -1661
rect 545 -1695 557 -1661
rect 499 -1701 557 -1695
rect 691 -1661 749 -1655
rect 691 -1695 703 -1661
rect 737 -1695 749 -1661
rect 691 -1701 749 -1695
rect 883 -1661 941 -1655
rect 883 -1695 895 -1661
rect 929 -1695 941 -1661
rect 883 -1701 941 -1695
rect -983 -1754 -937 -1742
rect -983 -1900 -977 -1754
rect -943 -1900 -937 -1754
rect -983 -1912 -937 -1900
rect -887 -1754 -841 -1742
rect -887 -1900 -881 -1754
rect -847 -1900 -841 -1754
rect -887 -1912 -841 -1900
rect -791 -1754 -745 -1742
rect -791 -1900 -785 -1754
rect -751 -1900 -745 -1754
rect -791 -1912 -745 -1900
rect -695 -1754 -649 -1742
rect -695 -1900 -689 -1754
rect -655 -1900 -649 -1754
rect -695 -1912 -649 -1900
rect -599 -1754 -553 -1742
rect -599 -1900 -593 -1754
rect -559 -1900 -553 -1754
rect -599 -1912 -553 -1900
rect -503 -1754 -457 -1742
rect -503 -1900 -497 -1754
rect -463 -1900 -457 -1754
rect -503 -1912 -457 -1900
rect -407 -1754 -361 -1742
rect -407 -1900 -401 -1754
rect -367 -1900 -361 -1754
rect -407 -1912 -361 -1900
rect -311 -1754 -265 -1742
rect -311 -1900 -305 -1754
rect -271 -1900 -265 -1754
rect -311 -1912 -265 -1900
rect -215 -1754 -169 -1742
rect -215 -1900 -209 -1754
rect -175 -1900 -169 -1754
rect -215 -1912 -169 -1900
rect -119 -1754 -73 -1742
rect -119 -1900 -113 -1754
rect -79 -1900 -73 -1754
rect -119 -1912 -73 -1900
rect -23 -1754 23 -1742
rect -23 -1900 -17 -1754
rect 17 -1900 23 -1754
rect -23 -1912 23 -1900
rect 73 -1754 119 -1742
rect 73 -1900 79 -1754
rect 113 -1900 119 -1754
rect 73 -1912 119 -1900
rect 169 -1754 215 -1742
rect 169 -1900 175 -1754
rect 209 -1900 215 -1754
rect 169 -1912 215 -1900
rect 265 -1754 311 -1742
rect 265 -1900 271 -1754
rect 305 -1900 311 -1754
rect 265 -1912 311 -1900
rect 361 -1754 407 -1742
rect 361 -1900 367 -1754
rect 401 -1900 407 -1754
rect 361 -1912 407 -1900
rect 457 -1754 503 -1742
rect 457 -1900 463 -1754
rect 497 -1900 503 -1754
rect 457 -1912 503 -1900
rect 553 -1754 599 -1742
rect 553 -1900 559 -1754
rect 593 -1900 599 -1754
rect 553 -1912 599 -1900
rect 649 -1754 695 -1742
rect 649 -1900 655 -1754
rect 689 -1900 695 -1754
rect 649 -1912 695 -1900
rect 745 -1754 791 -1742
rect 745 -1900 751 -1754
rect 785 -1900 791 -1754
rect 745 -1912 791 -1900
rect 841 -1754 887 -1742
rect 841 -1900 847 -1754
rect 881 -1900 887 -1754
rect 841 -1912 887 -1900
rect 937 -1754 983 -1742
rect 937 -1900 943 -1754
rect 977 -1900 983 -1754
rect 937 -1912 983 -1900
rect -941 -1959 -883 -1953
rect -941 -1993 -929 -1959
rect -895 -1993 -883 -1959
rect -941 -1999 -883 -1993
rect -749 -1959 -691 -1953
rect -749 -1993 -737 -1959
rect -703 -1993 -691 -1959
rect -749 -1999 -691 -1993
rect -557 -1959 -499 -1953
rect -557 -1993 -545 -1959
rect -511 -1993 -499 -1959
rect -557 -1999 -499 -1993
rect -365 -1959 -307 -1953
rect -365 -1993 -353 -1959
rect -319 -1993 -307 -1959
rect -365 -1999 -307 -1993
rect -173 -1959 -115 -1953
rect -173 -1993 -161 -1959
rect -127 -1993 -115 -1959
rect -173 -1999 -115 -1993
rect 19 -1959 77 -1953
rect 19 -1993 31 -1959
rect 65 -1993 77 -1959
rect 19 -1999 77 -1993
rect 211 -1959 269 -1953
rect 211 -1993 223 -1959
rect 257 -1993 269 -1959
rect 211 -1999 269 -1993
rect 403 -1959 461 -1953
rect 403 -1993 415 -1959
rect 449 -1993 461 -1959
rect 403 -1999 461 -1993
rect 595 -1959 653 -1953
rect 595 -1993 607 -1959
rect 641 -1993 653 -1959
rect 595 -1999 653 -1993
rect 787 -1959 845 -1953
rect 787 -1993 799 -1959
rect 833 -1993 845 -1959
rect 787 -1999 845 -1993
<< properties >>
string FIXED_BBOX -1074 -2078 1074 2078
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.85 l 0.15 m 10 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
