magic
tech sky130A
magscale 1 2
timestamp 1669661075
<< poly >>
rect 94 792 272 822
rect 224 -80 266 56
rect 172 -108 270 -80
rect 172 -156 196 -108
rect 246 -156 270 -108
rect 172 -186 270 -156
rect 174 -992 272 -964
rect 174 -1040 198 -992
rect 248 -1040 272 -992
rect 174 -1070 272 -1040
rect 224 -1234 270 -1070
<< polycont >>
rect 196 -156 246 -108
rect 198 -1040 248 -992
<< locali >>
rect 180 -104 258 -92
rect 180 -160 192 -104
rect 248 -160 258 -104
rect 180 -174 258 -160
rect 182 -988 260 -976
rect 182 -1044 194 -988
rect 250 -1044 260 -988
rect 182 -1058 260 -1044
<< viali >>
rect 192 -108 248 -104
rect 192 -156 196 -108
rect 196 -156 246 -108
rect 246 -156 248 -108
rect 192 -160 248 -156
rect 194 -992 250 -988
rect 194 -1040 198 -992
rect 198 -1040 248 -992
rect 248 -1040 250 -992
rect 194 -1044 250 -1040
rect 158 -2242 212 -2192
<< metal1 >>
rect 176 -98 262 -88
rect 172 -104 262 -98
rect 172 -152 192 -104
rect 176 -160 192 -152
rect 248 -150 262 -104
rect 248 -160 268 -150
rect 176 -178 268 -160
rect 224 -972 268 -178
rect 178 -974 268 -972
rect 178 -982 264 -974
rect 174 -988 264 -982
rect 174 -1036 194 -988
rect 178 -1044 194 -1036
rect 250 -1044 264 -988
rect 178 -1062 264 -1044
rect 296 -1258 324 78
rect 172 -2176 202 -1920
rect 144 -2192 226 -2176
rect 144 -2242 158 -2192
rect 212 -2242 226 -2192
rect 144 -2256 226 -2242
use sky130_fd_pr__nfet_01v8_E8KW6F  sky130_fd_pr__nfet_01v8_E8KW6F_0
timestamp 1667954557
transform 1 0 246 0 1 -1588
box -88 -376 88 376
use sky130_fd_pr__pfet_01v8_JJT9EJ  sky130_fd_pr__pfet_01v8_JJT9EJ_0
timestamp 1669522153
transform 1 0 183 0 1 418
box -183 -412 183 412
<< end >>
