magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect 30 1005 88 1011
rect 30 971 42 1005
rect 30 965 88 971
<< nwell >>
rect -183 -1058 183 1024
<< pmos >>
rect -89 -996 -29 924
rect 29 -996 89 924
<< pdiff >>
rect -147 899 -89 924
rect -147 865 -135 899
rect -101 865 -89 899
rect -147 831 -89 865
rect -147 797 -135 831
rect -101 797 -89 831
rect -147 763 -89 797
rect -147 729 -135 763
rect -101 729 -89 763
rect -147 695 -89 729
rect -147 661 -135 695
rect -101 661 -89 695
rect -147 627 -89 661
rect -147 593 -135 627
rect -101 593 -89 627
rect -147 559 -89 593
rect -147 525 -135 559
rect -101 525 -89 559
rect -147 491 -89 525
rect -147 457 -135 491
rect -101 457 -89 491
rect -147 423 -89 457
rect -147 389 -135 423
rect -101 389 -89 423
rect -147 355 -89 389
rect -147 321 -135 355
rect -101 321 -89 355
rect -147 287 -89 321
rect -147 253 -135 287
rect -101 253 -89 287
rect -147 219 -89 253
rect -147 185 -135 219
rect -101 185 -89 219
rect -147 151 -89 185
rect -147 117 -135 151
rect -101 117 -89 151
rect -147 83 -89 117
rect -147 49 -135 83
rect -101 49 -89 83
rect -147 15 -89 49
rect -147 -19 -135 15
rect -101 -19 -89 15
rect -147 -53 -89 -19
rect -147 -87 -135 -53
rect -101 -87 -89 -53
rect -147 -121 -89 -87
rect -147 -155 -135 -121
rect -101 -155 -89 -121
rect -147 -189 -89 -155
rect -147 -223 -135 -189
rect -101 -223 -89 -189
rect -147 -257 -89 -223
rect -147 -291 -135 -257
rect -101 -291 -89 -257
rect -147 -325 -89 -291
rect -147 -359 -135 -325
rect -101 -359 -89 -325
rect -147 -393 -89 -359
rect -147 -427 -135 -393
rect -101 -427 -89 -393
rect -147 -461 -89 -427
rect -147 -495 -135 -461
rect -101 -495 -89 -461
rect -147 -529 -89 -495
rect -147 -563 -135 -529
rect -101 -563 -89 -529
rect -147 -597 -89 -563
rect -147 -631 -135 -597
rect -101 -631 -89 -597
rect -147 -665 -89 -631
rect -147 -699 -135 -665
rect -101 -699 -89 -665
rect -147 -733 -89 -699
rect -147 -767 -135 -733
rect -101 -767 -89 -733
rect -147 -801 -89 -767
rect -147 -835 -135 -801
rect -101 -835 -89 -801
rect -147 -869 -89 -835
rect -147 -903 -135 -869
rect -101 -903 -89 -869
rect -147 -937 -89 -903
rect -147 -971 -135 -937
rect -101 -971 -89 -937
rect -147 -996 -89 -971
rect -29 899 29 924
rect -29 865 -17 899
rect 17 865 29 899
rect -29 831 29 865
rect -29 797 -17 831
rect 17 797 29 831
rect -29 763 29 797
rect -29 729 -17 763
rect 17 729 29 763
rect -29 695 29 729
rect -29 661 -17 695
rect 17 661 29 695
rect -29 627 29 661
rect -29 593 -17 627
rect 17 593 29 627
rect -29 559 29 593
rect -29 525 -17 559
rect 17 525 29 559
rect -29 491 29 525
rect -29 457 -17 491
rect 17 457 29 491
rect -29 423 29 457
rect -29 389 -17 423
rect 17 389 29 423
rect -29 355 29 389
rect -29 321 -17 355
rect 17 321 29 355
rect -29 287 29 321
rect -29 253 -17 287
rect 17 253 29 287
rect -29 219 29 253
rect -29 185 -17 219
rect 17 185 29 219
rect -29 151 29 185
rect -29 117 -17 151
rect 17 117 29 151
rect -29 83 29 117
rect -29 49 -17 83
rect 17 49 29 83
rect -29 15 29 49
rect -29 -19 -17 15
rect 17 -19 29 15
rect -29 -53 29 -19
rect -29 -87 -17 -53
rect 17 -87 29 -53
rect -29 -121 29 -87
rect -29 -155 -17 -121
rect 17 -155 29 -121
rect -29 -189 29 -155
rect -29 -223 -17 -189
rect 17 -223 29 -189
rect -29 -257 29 -223
rect -29 -291 -17 -257
rect 17 -291 29 -257
rect -29 -325 29 -291
rect -29 -359 -17 -325
rect 17 -359 29 -325
rect -29 -393 29 -359
rect -29 -427 -17 -393
rect 17 -427 29 -393
rect -29 -461 29 -427
rect -29 -495 -17 -461
rect 17 -495 29 -461
rect -29 -529 29 -495
rect -29 -563 -17 -529
rect 17 -563 29 -529
rect -29 -597 29 -563
rect -29 -631 -17 -597
rect 17 -631 29 -597
rect -29 -665 29 -631
rect -29 -699 -17 -665
rect 17 -699 29 -665
rect -29 -733 29 -699
rect -29 -767 -17 -733
rect 17 -767 29 -733
rect -29 -801 29 -767
rect -29 -835 -17 -801
rect 17 -835 29 -801
rect -29 -869 29 -835
rect -29 -903 -17 -869
rect 17 -903 29 -869
rect -29 -937 29 -903
rect -29 -971 -17 -937
rect 17 -971 29 -937
rect -29 -996 29 -971
rect 89 899 147 924
rect 89 865 101 899
rect 135 865 147 899
rect 89 831 147 865
rect 89 797 101 831
rect 135 797 147 831
rect 89 763 147 797
rect 89 729 101 763
rect 135 729 147 763
rect 89 695 147 729
rect 89 661 101 695
rect 135 661 147 695
rect 89 627 147 661
rect 89 593 101 627
rect 135 593 147 627
rect 89 559 147 593
rect 89 525 101 559
rect 135 525 147 559
rect 89 491 147 525
rect 89 457 101 491
rect 135 457 147 491
rect 89 423 147 457
rect 89 389 101 423
rect 135 389 147 423
rect 89 355 147 389
rect 89 321 101 355
rect 135 321 147 355
rect 89 287 147 321
rect 89 253 101 287
rect 135 253 147 287
rect 89 219 147 253
rect 89 185 101 219
rect 135 185 147 219
rect 89 151 147 185
rect 89 117 101 151
rect 135 117 147 151
rect 89 83 147 117
rect 89 49 101 83
rect 135 49 147 83
rect 89 15 147 49
rect 89 -19 101 15
rect 135 -19 147 15
rect 89 -53 147 -19
rect 89 -87 101 -53
rect 135 -87 147 -53
rect 89 -121 147 -87
rect 89 -155 101 -121
rect 135 -155 147 -121
rect 89 -189 147 -155
rect 89 -223 101 -189
rect 135 -223 147 -189
rect 89 -257 147 -223
rect 89 -291 101 -257
rect 135 -291 147 -257
rect 89 -325 147 -291
rect 89 -359 101 -325
rect 135 -359 147 -325
rect 89 -393 147 -359
rect 89 -427 101 -393
rect 135 -427 147 -393
rect 89 -461 147 -427
rect 89 -495 101 -461
rect 135 -495 147 -461
rect 89 -529 147 -495
rect 89 -563 101 -529
rect 135 -563 147 -529
rect 89 -597 147 -563
rect 89 -631 101 -597
rect 135 -631 147 -597
rect 89 -665 147 -631
rect 89 -699 101 -665
rect 135 -699 147 -665
rect 89 -733 147 -699
rect 89 -767 101 -733
rect 135 -767 147 -733
rect 89 -801 147 -767
rect 89 -835 101 -801
rect 135 -835 147 -801
rect 89 -869 147 -835
rect 89 -903 101 -869
rect 135 -903 147 -869
rect 89 -937 147 -903
rect 89 -971 101 -937
rect 135 -971 147 -937
rect 89 -996 147 -971
<< pdiffc >>
rect -135 865 -101 899
rect -135 797 -101 831
rect -135 729 -101 763
rect -135 661 -101 695
rect -135 593 -101 627
rect -135 525 -101 559
rect -135 457 -101 491
rect -135 389 -101 423
rect -135 321 -101 355
rect -135 253 -101 287
rect -135 185 -101 219
rect -135 117 -101 151
rect -135 49 -101 83
rect -135 -19 -101 15
rect -135 -87 -101 -53
rect -135 -155 -101 -121
rect -135 -223 -101 -189
rect -135 -291 -101 -257
rect -135 -359 -101 -325
rect -135 -427 -101 -393
rect -135 -495 -101 -461
rect -135 -563 -101 -529
rect -135 -631 -101 -597
rect -135 -699 -101 -665
rect -135 -767 -101 -733
rect -135 -835 -101 -801
rect -135 -903 -101 -869
rect -135 -971 -101 -937
rect -17 865 17 899
rect -17 797 17 831
rect -17 729 17 763
rect -17 661 17 695
rect -17 593 17 627
rect -17 525 17 559
rect -17 457 17 491
rect -17 389 17 423
rect -17 321 17 355
rect -17 253 17 287
rect -17 185 17 219
rect -17 117 17 151
rect -17 49 17 83
rect -17 -19 17 15
rect -17 -87 17 -53
rect -17 -155 17 -121
rect -17 -223 17 -189
rect -17 -291 17 -257
rect -17 -359 17 -325
rect -17 -427 17 -393
rect -17 -495 17 -461
rect -17 -563 17 -529
rect -17 -631 17 -597
rect -17 -699 17 -665
rect -17 -767 17 -733
rect -17 -835 17 -801
rect -17 -903 17 -869
rect -17 -971 17 -937
rect 101 865 135 899
rect 101 797 135 831
rect 101 729 135 763
rect 101 661 135 695
rect 101 593 135 627
rect 101 525 135 559
rect 101 457 135 491
rect 101 389 135 423
rect 101 321 135 355
rect 101 253 135 287
rect 101 185 135 219
rect 101 117 135 151
rect 101 49 135 83
rect 101 -19 135 15
rect 101 -87 135 -53
rect 101 -155 135 -121
rect 101 -223 135 -189
rect 101 -291 135 -257
rect 101 -359 135 -325
rect 101 -427 135 -393
rect 101 -495 135 -461
rect 101 -563 135 -529
rect 101 -631 135 -597
rect 101 -699 135 -665
rect 101 -767 135 -733
rect 101 -835 135 -801
rect 101 -903 135 -869
rect 101 -971 135 -937
<< poly >>
rect -89 1005 92 1021
rect -89 971 42 1005
rect 76 971 92 1005
rect -89 955 92 971
rect -89 924 -29 955
rect 29 924 89 955
rect -89 -1018 -29 -996
rect 29 -1018 89 -996
rect -89 -1054 89 -1018
<< polycont >>
rect 42 971 76 1005
<< locali >>
rect 26 971 42 1005
rect 76 971 92 1005
rect -135 899 -101 928
rect -135 831 -101 847
rect -135 763 -101 775
rect -135 695 -101 703
rect -135 627 -101 631
rect -135 521 -101 525
rect -135 449 -101 457
rect -135 377 -101 389
rect -135 305 -101 321
rect -135 233 -101 253
rect -135 161 -101 185
rect -135 89 -101 117
rect -135 17 -101 49
rect -135 -53 -101 -19
rect -135 -121 -101 -89
rect -135 -189 -101 -161
rect -135 -257 -101 -233
rect -135 -325 -101 -305
rect -135 -393 -101 -377
rect -135 -461 -101 -449
rect -135 -529 -101 -521
rect -135 -597 -101 -593
rect -135 -703 -101 -699
rect -135 -775 -101 -767
rect -135 -847 -101 -835
rect -135 -919 -101 -903
rect -135 -1000 -101 -971
rect -17 899 17 928
rect -17 831 17 847
rect -17 763 17 775
rect -17 695 17 703
rect -17 627 17 631
rect -17 521 17 525
rect -17 449 17 457
rect -17 377 17 389
rect -17 305 17 321
rect -17 233 17 253
rect -17 161 17 185
rect -17 89 17 117
rect -17 17 17 49
rect -17 -53 17 -19
rect -17 -121 17 -89
rect -17 -189 17 -161
rect -17 -257 17 -233
rect -17 -325 17 -305
rect -17 -393 17 -377
rect -17 -461 17 -449
rect -17 -529 17 -521
rect -17 -597 17 -593
rect -17 -703 17 -699
rect -17 -775 17 -767
rect -17 -847 17 -835
rect -17 -919 17 -903
rect -17 -1000 17 -971
rect 101 899 135 928
rect 101 831 135 847
rect 101 763 135 775
rect 101 695 135 703
rect 101 627 135 631
rect 101 521 135 525
rect 101 449 135 457
rect 101 377 135 389
rect 101 305 135 321
rect 101 233 135 253
rect 101 161 135 185
rect 101 89 135 117
rect 101 17 135 49
rect 101 -53 135 -19
rect 101 -121 135 -89
rect 101 -189 135 -161
rect 101 -257 135 -233
rect 101 -325 135 -305
rect 101 -393 135 -377
rect 101 -461 135 -449
rect 101 -529 135 -521
rect 101 -597 135 -593
rect 101 -703 135 -699
rect 101 -775 135 -767
rect 101 -847 135 -835
rect 101 -919 135 -903
rect 101 -1000 135 -971
<< viali >>
rect 42 971 76 1005
rect -135 865 -101 881
rect -135 847 -101 865
rect -135 797 -101 809
rect -135 775 -101 797
rect -135 729 -101 737
rect -135 703 -101 729
rect -135 661 -101 665
rect -135 631 -101 661
rect -135 559 -101 593
rect -135 491 -101 521
rect -135 487 -101 491
rect -135 423 -101 449
rect -135 415 -101 423
rect -135 355 -101 377
rect -135 343 -101 355
rect -135 287 -101 305
rect -135 271 -101 287
rect -135 219 -101 233
rect -135 199 -101 219
rect -135 151 -101 161
rect -135 127 -101 151
rect -135 83 -101 89
rect -135 55 -101 83
rect -135 15 -101 17
rect -135 -17 -101 15
rect -135 -87 -101 -55
rect -135 -89 -101 -87
rect -135 -155 -101 -127
rect -135 -161 -101 -155
rect -135 -223 -101 -199
rect -135 -233 -101 -223
rect -135 -291 -101 -271
rect -135 -305 -101 -291
rect -135 -359 -101 -343
rect -135 -377 -101 -359
rect -135 -427 -101 -415
rect -135 -449 -101 -427
rect -135 -495 -101 -487
rect -135 -521 -101 -495
rect -135 -563 -101 -559
rect -135 -593 -101 -563
rect -135 -665 -101 -631
rect -135 -733 -101 -703
rect -135 -737 -101 -733
rect -135 -801 -101 -775
rect -135 -809 -101 -801
rect -135 -869 -101 -847
rect -135 -881 -101 -869
rect -135 -937 -101 -919
rect -135 -953 -101 -937
rect -17 865 17 881
rect -17 847 17 865
rect -17 797 17 809
rect -17 775 17 797
rect -17 729 17 737
rect -17 703 17 729
rect -17 661 17 665
rect -17 631 17 661
rect -17 559 17 593
rect -17 491 17 521
rect -17 487 17 491
rect -17 423 17 449
rect -17 415 17 423
rect -17 355 17 377
rect -17 343 17 355
rect -17 287 17 305
rect -17 271 17 287
rect -17 219 17 233
rect -17 199 17 219
rect -17 151 17 161
rect -17 127 17 151
rect -17 83 17 89
rect -17 55 17 83
rect -17 15 17 17
rect -17 -17 17 15
rect -17 -87 17 -55
rect -17 -89 17 -87
rect -17 -155 17 -127
rect -17 -161 17 -155
rect -17 -223 17 -199
rect -17 -233 17 -223
rect -17 -291 17 -271
rect -17 -305 17 -291
rect -17 -359 17 -343
rect -17 -377 17 -359
rect -17 -427 17 -415
rect -17 -449 17 -427
rect -17 -495 17 -487
rect -17 -521 17 -495
rect -17 -563 17 -559
rect -17 -593 17 -563
rect -17 -665 17 -631
rect -17 -733 17 -703
rect -17 -737 17 -733
rect -17 -801 17 -775
rect -17 -809 17 -801
rect -17 -869 17 -847
rect -17 -881 17 -869
rect -17 -937 17 -919
rect -17 -953 17 -937
rect 101 865 135 881
rect 101 847 135 865
rect 101 797 135 809
rect 101 775 135 797
rect 101 729 135 737
rect 101 703 135 729
rect 101 661 135 665
rect 101 631 135 661
rect 101 559 135 593
rect 101 491 135 521
rect 101 487 135 491
rect 101 423 135 449
rect 101 415 135 423
rect 101 355 135 377
rect 101 343 135 355
rect 101 287 135 305
rect 101 271 135 287
rect 101 219 135 233
rect 101 199 135 219
rect 101 151 135 161
rect 101 127 135 151
rect 101 83 135 89
rect 101 55 135 83
rect 101 15 135 17
rect 101 -17 135 15
rect 101 -87 135 -55
rect 101 -89 135 -87
rect 101 -155 135 -127
rect 101 -161 135 -155
rect 101 -223 135 -199
rect 101 -233 135 -223
rect 101 -291 135 -271
rect 101 -305 135 -291
rect 101 -359 135 -343
rect 101 -377 135 -359
rect 101 -427 135 -415
rect 101 -449 135 -427
rect 101 -495 135 -487
rect 101 -521 135 -495
rect 101 -563 135 -559
rect 101 -593 135 -563
rect 101 -665 135 -631
rect 101 -733 135 -703
rect 101 -737 135 -733
rect 101 -801 135 -775
rect 101 -809 135 -801
rect 101 -869 135 -847
rect 101 -881 135 -869
rect 101 -937 135 -919
rect 101 -953 135 -937
<< metal1 >>
rect 30 1005 88 1011
rect 30 971 42 1005
rect 76 971 88 1005
rect 30 965 88 971
rect -141 881 -95 924
rect -141 847 -135 881
rect -101 847 -95 881
rect -141 809 -95 847
rect -141 775 -135 809
rect -101 775 -95 809
rect -141 737 -95 775
rect -141 703 -135 737
rect -101 703 -95 737
rect -141 665 -95 703
rect -141 631 -135 665
rect -101 631 -95 665
rect -141 593 -95 631
rect -141 559 -135 593
rect -101 559 -95 593
rect -141 521 -95 559
rect -141 487 -135 521
rect -101 487 -95 521
rect -141 449 -95 487
rect -141 415 -135 449
rect -101 415 -95 449
rect -141 377 -95 415
rect -141 343 -135 377
rect -101 343 -95 377
rect -141 305 -95 343
rect -141 271 -135 305
rect -101 271 -95 305
rect -141 233 -95 271
rect -141 199 -135 233
rect -101 199 -95 233
rect -141 161 -95 199
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -199 -95 -161
rect -141 -233 -135 -199
rect -101 -233 -95 -199
rect -141 -271 -95 -233
rect -141 -305 -135 -271
rect -101 -305 -95 -271
rect -141 -343 -95 -305
rect -141 -377 -135 -343
rect -101 -377 -95 -343
rect -141 -415 -95 -377
rect -141 -449 -135 -415
rect -101 -449 -95 -415
rect -141 -487 -95 -449
rect -141 -521 -135 -487
rect -101 -521 -95 -487
rect -141 -559 -95 -521
rect -141 -593 -135 -559
rect -101 -593 -95 -559
rect -141 -631 -95 -593
rect -141 -665 -135 -631
rect -101 -665 -95 -631
rect -141 -703 -95 -665
rect -141 -737 -135 -703
rect -101 -737 -95 -703
rect -141 -775 -95 -737
rect -141 -809 -135 -775
rect -101 -809 -95 -775
rect -141 -847 -95 -809
rect -141 -881 -135 -847
rect -101 -881 -95 -847
rect -141 -919 -95 -881
rect -141 -953 -135 -919
rect -101 -953 -95 -919
rect -141 -996 -95 -953
rect -23 881 23 924
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -919 23 -881
rect -23 -953 -17 -919
rect 17 -953 23 -919
rect -23 -996 23 -953
rect 95 881 141 924
rect 95 847 101 881
rect 135 847 141 881
rect 95 809 141 847
rect 95 775 101 809
rect 135 775 141 809
rect 95 737 141 775
rect 95 703 101 737
rect 135 703 141 737
rect 95 665 141 703
rect 95 631 101 665
rect 135 631 141 665
rect 95 593 141 631
rect 95 559 101 593
rect 135 559 141 593
rect 95 521 141 559
rect 95 487 101 521
rect 135 487 141 521
rect 95 449 141 487
rect 95 415 101 449
rect 135 415 141 449
rect 95 377 141 415
rect 95 343 101 377
rect 135 343 141 377
rect 95 305 141 343
rect 95 271 101 305
rect 135 271 141 305
rect 95 233 141 271
rect 95 199 101 233
rect 135 199 141 233
rect 95 161 141 199
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -199 141 -161
rect 95 -233 101 -199
rect 135 -233 141 -199
rect 95 -271 141 -233
rect 95 -305 101 -271
rect 135 -305 141 -271
rect 95 -343 141 -305
rect 95 -377 101 -343
rect 135 -377 141 -343
rect 95 -415 141 -377
rect 95 -449 101 -415
rect 135 -449 141 -415
rect 95 -487 141 -449
rect 95 -521 101 -487
rect 135 -521 141 -487
rect 95 -559 141 -521
rect 95 -593 101 -559
rect 135 -593 141 -559
rect 95 -631 141 -593
rect 95 -665 101 -631
rect 135 -665 141 -631
rect 95 -703 141 -665
rect 95 -737 101 -703
rect 135 -737 141 -703
rect 95 -775 141 -737
rect 95 -809 101 -775
rect 135 -809 141 -775
rect 95 -847 141 -809
rect 95 -881 101 -847
rect 135 -881 141 -847
rect 95 -919 141 -881
rect 95 -953 101 -919
rect 135 -953 141 -919
rect 95 -996 141 -953
<< end >>
