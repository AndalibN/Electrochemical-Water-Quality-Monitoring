magic
tech sky130A
timestamp 1667316071
<< nmos >>
rect -104 -500 -54 500
rect -25 -500 25 500
rect 54 -500 104 500
<< ndiff >>
rect -133 494 -104 500
rect -133 -494 -127 494
rect -110 -494 -104 494
rect -133 -500 -104 -494
rect -54 494 -25 500
rect -54 -494 -48 494
rect -31 -494 -25 494
rect -54 -500 -25 -494
rect 25 494 54 500
rect 25 -494 31 494
rect 48 -494 54 494
rect 25 -500 54 -494
rect 104 494 133 500
rect 104 -494 110 494
rect 127 -494 133 494
rect 104 -500 133 -494
<< ndiffc >>
rect -127 -494 -110 494
rect -48 -494 -31 494
rect 31 -494 48 494
rect 110 -494 127 494
<< poly >>
rect -104 536 -54 544
rect -104 519 -96 536
rect -62 519 -54 536
rect -104 500 -54 519
rect -25 536 25 544
rect -25 519 -17 536
rect 17 519 25 536
rect -25 500 25 519
rect 54 536 104 544
rect 54 519 62 536
rect 96 519 104 536
rect 54 500 104 519
rect -104 -519 -54 -500
rect -104 -536 -96 -519
rect -62 -536 -54 -519
rect -104 -544 -54 -536
rect -25 -519 25 -500
rect -25 -536 -17 -519
rect 17 -536 25 -519
rect -25 -544 25 -536
rect 54 -519 104 -500
rect 54 -536 62 -519
rect 96 -536 104 -519
rect 54 -544 104 -536
<< polycont >>
rect -96 519 -62 536
rect -17 519 17 536
rect 62 519 96 536
rect -96 -536 -62 -519
rect -17 -536 17 -519
rect 62 -536 96 -519
<< locali >>
rect -104 519 -96 536
rect -62 519 -54 536
rect -25 519 -17 536
rect 17 519 25 536
rect 54 519 62 536
rect 96 519 104 536
rect -127 494 -110 502
rect -127 -502 -110 -494
rect -48 494 -31 502
rect -48 -502 -31 -494
rect 31 494 48 502
rect 31 -502 48 -494
rect 110 494 127 502
rect 110 -502 127 -494
rect -104 -536 -96 -519
rect -62 -536 -54 -519
rect -25 -536 -17 -519
rect 17 -536 25 -519
rect 54 -536 62 -519
rect 96 -536 104 -519
<< viali >>
rect -96 519 -62 536
rect -17 519 17 536
rect 62 519 96 536
rect -127 -494 -110 494
rect -48 -494 -31 494
rect 31 -494 48 494
rect 110 -494 127 494
rect -96 -536 -62 -519
rect -17 -536 17 -519
rect 62 -536 96 -519
<< metal1 >>
rect -102 536 -56 539
rect -102 519 -96 536
rect -62 519 -56 536
rect -102 516 -56 519
rect -23 536 23 539
rect -23 519 -17 536
rect 17 519 23 536
rect -23 516 23 519
rect 56 536 102 539
rect 56 519 62 536
rect 96 519 102 536
rect 56 516 102 519
rect -130 494 -107 500
rect -130 -494 -127 494
rect -110 -494 -107 494
rect -130 -500 -107 -494
rect -51 494 -28 500
rect -51 -494 -48 494
rect -31 -494 -28 494
rect -51 -500 -28 -494
rect 28 494 51 500
rect 28 -494 31 494
rect 48 -494 51 494
rect 28 -500 51 -494
rect 107 494 130 500
rect 107 -494 110 494
rect 127 -494 130 494
rect 107 -500 130 -494
rect -102 -519 -56 -516
rect -102 -536 -96 -519
rect -62 -536 -56 -519
rect -102 -539 -56 -536
rect -23 -519 23 -516
rect -23 -536 -17 -519
rect 17 -536 23 -519
rect -23 -539 23 -536
rect 56 -519 102 -516
rect 56 -536 62 -519
rect 96 -536 102 -519
rect 56 -539 102 -536
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
