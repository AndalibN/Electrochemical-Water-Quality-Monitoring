magic
tech sky130A
magscale 1 2
timestamp 1668714113
<< metal3 >>
rect -1509 1422 -10 1450
rect -1509 78 -94 1422
rect -30 78 -10 1422
rect -1509 50 -10 78
rect 110 1422 1609 1450
rect 110 78 1525 1422
rect 1589 78 1609 1422
rect 110 50 1609 78
rect -1509 -78 -10 -50
rect -1509 -1422 -94 -78
rect -30 -1422 -10 -78
rect -1509 -1450 -10 -1422
rect 110 -78 1609 -50
rect 110 -1422 1525 -78
rect 1589 -1422 1609 -78
rect 110 -1450 1609 -1422
<< via3 >>
rect -94 78 -30 1422
rect 1525 78 1589 1422
rect -94 -1422 -30 -78
rect 1525 -1422 1589 -78
<< mimcap >>
rect -1409 1310 -209 1350
rect -1409 190 -1369 1310
rect -249 190 -209 1310
rect -1409 150 -209 190
rect 210 1310 1410 1350
rect 210 190 250 1310
rect 1370 190 1410 1310
rect 210 150 1410 190
rect -1409 -190 -209 -150
rect -1409 -1310 -1369 -190
rect -249 -1310 -209 -190
rect -1409 -1350 -209 -1310
rect 210 -190 1410 -150
rect 210 -1310 250 -190
rect 1370 -1310 1410 -190
rect 210 -1350 1410 -1310
<< mimcapcontact >>
rect -1369 190 -249 1310
rect 250 190 1370 1310
rect -1369 -1310 -249 -190
rect 250 -1310 1370 -190
<< metal4 >>
rect -861 1311 -757 1500
rect -141 1438 -37 1500
rect -141 1422 -14 1438
rect -1370 1310 -248 1311
rect -1370 190 -1369 1310
rect -249 190 -248 1310
rect -1370 189 -248 190
rect -861 -189 -757 189
rect -141 78 -94 1422
rect -30 78 -14 1422
rect 758 1311 862 1500
rect 1478 1438 1582 1500
rect 1478 1422 1605 1438
rect 249 1310 1371 1311
rect 249 190 250 1310
rect 1370 190 1371 1310
rect 249 189 1371 190
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -1370 -190 -248 -189
rect -1370 -1310 -1369 -190
rect -249 -1310 -248 -190
rect -1370 -1311 -248 -1310
rect -861 -1500 -757 -1311
rect -141 -1422 -94 -78
rect -30 -1422 -14 -78
rect 758 -189 862 189
rect 1478 78 1525 1422
rect 1589 78 1605 1422
rect 1478 62 1605 78
rect 1478 -62 1582 62
rect 1478 -78 1605 -62
rect 249 -190 1371 -189
rect 249 -1310 250 -190
rect 1370 -1310 1371 -190
rect 249 -1311 1371 -1310
rect -141 -1438 -14 -1422
rect -141 -1500 -37 -1438
rect 758 -1500 862 -1311
rect 1478 -1422 1525 -78
rect 1589 -1422 1605 -78
rect 1478 -1438 1605 -1422
rect 1478 -1500 1582 -1438
<< properties >>
string FIXED_BBOX 10 50 1410 1450
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 6 l 6 val 76.56 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
