magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -183 -412 183 412
<< pmos >>
rect -89 -350 -29 350
rect 29 -350 89 350
<< pdiff >>
rect -147 323 -89 350
rect -147 289 -135 323
rect -101 289 -89 323
rect -147 255 -89 289
rect -147 221 -135 255
rect -101 221 -89 255
rect -147 187 -89 221
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -221 -89 -187
rect -147 -255 -135 -221
rect -101 -255 -89 -221
rect -147 -289 -89 -255
rect -147 -323 -135 -289
rect -101 -323 -89 -289
rect -147 -350 -89 -323
rect -29 323 29 350
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -350 29 -323
rect 89 323 147 350
rect 89 289 101 323
rect 135 289 147 323
rect 89 255 147 289
rect 89 221 101 255
rect 135 221 147 255
rect 89 187 147 221
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -221 147 -187
rect 89 -255 101 -221
rect 135 -255 147 -221
rect 89 -289 147 -255
rect 89 -323 101 -289
rect 135 -323 147 -289
rect 89 -350 147 -323
<< pdiffc >>
rect -135 289 -101 323
rect -135 221 -101 255
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -135 -255 -101 -221
rect -135 -323 -101 -289
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect 101 289 135 323
rect 101 221 135 255
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 101 -255 135 -221
rect 101 -323 135 -289
<< poly >>
rect -89 350 -29 376
rect 29 350 89 376
rect -89 -376 -29 -350
rect 29 -376 89 -350
<< locali >>
rect -135 323 -101 354
rect -135 255 -101 271
rect -135 187 -101 199
rect -135 119 -101 127
rect -135 51 -101 55
rect -135 -55 -101 -51
rect -135 -127 -101 -119
rect -135 -199 -101 -187
rect -135 -271 -101 -255
rect -135 -354 -101 -323
rect -17 323 17 354
rect -17 255 17 271
rect -17 187 17 199
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -199 17 -187
rect -17 -271 17 -255
rect -17 -354 17 -323
rect 101 323 135 354
rect 101 255 135 271
rect 101 187 135 199
rect 101 119 135 127
rect 101 51 135 55
rect 101 -55 135 -51
rect 101 -127 135 -119
rect 101 -199 135 -187
rect 101 -271 135 -255
rect 101 -354 135 -323
<< viali >>
rect -135 289 -101 305
rect -135 271 -101 289
rect -135 221 -101 233
rect -135 199 -101 221
rect -135 153 -101 161
rect -135 127 -101 153
rect -135 85 -101 89
rect -135 55 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -55
rect -135 -89 -101 -85
rect -135 -153 -101 -127
rect -135 -161 -101 -153
rect -135 -221 -101 -199
rect -135 -233 -101 -221
rect -135 -289 -101 -271
rect -135 -305 -101 -289
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect 101 289 135 305
rect 101 271 135 289
rect 101 221 135 233
rect 101 199 135 221
rect 101 153 135 161
rect 101 127 135 153
rect 101 85 135 89
rect 101 55 135 85
rect 101 -17 135 17
rect 101 -85 135 -55
rect 101 -89 135 -85
rect 101 -153 135 -127
rect 101 -161 135 -153
rect 101 -221 135 -199
rect 101 -233 135 -221
rect 101 -289 135 -271
rect 101 -305 135 -289
<< metal1 >>
rect -141 305 -95 350
rect -141 271 -135 305
rect -101 271 -95 305
rect -141 233 -95 271
rect -141 199 -135 233
rect -101 199 -95 233
rect -141 161 -95 199
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -199 -95 -161
rect -141 -233 -135 -199
rect -101 -233 -95 -199
rect -141 -271 -95 -233
rect -141 -305 -135 -271
rect -101 -305 -95 -271
rect -141 -350 -95 -305
rect -23 305 23 350
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -350 23 -305
rect 95 305 141 350
rect 95 271 101 305
rect 135 271 141 305
rect 95 233 141 271
rect 95 199 101 233
rect 135 199 141 233
rect 95 161 141 199
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -199 141 -161
rect 95 -233 101 -199
rect 135 -233 141 -199
rect 95 -271 141 -233
rect 95 -305 101 -271
rect 135 -305 141 -271
rect 95 -350 141 -305
<< end >>
