magic
tech sky130A
magscale 1 2
timestamp 1666801420
<< error_p >>
rect -32 4011 32 4017
rect -32 3977 -20 4011
rect -32 3971 32 3977
rect -32 2095 32 2101
rect -32 2061 -20 2095
rect -32 2055 32 2061
rect -32 1987 32 1993
rect -32 1953 -20 1987
rect -32 1947 32 1953
rect -32 71 32 77
rect -32 37 -20 71
rect -32 31 32 37
rect -32 -37 32 -31
rect -32 -71 -20 -37
rect -32 -77 32 -71
rect -32 -1953 32 -1947
rect -32 -1987 -20 -1953
rect -32 -1993 32 -1987
rect -32 -2061 32 -2055
rect -32 -2095 -20 -2061
rect -32 -2101 32 -2095
rect -32 -3977 32 -3971
rect -32 -4011 -20 -3977
rect -32 -4017 32 -4011
<< pwell >>
rect -232 -4149 232 4149
<< nmos >>
rect -36 2133 36 3939
rect -36 109 36 1915
rect -36 -1915 36 -109
rect -36 -3939 36 -2133
<< ndiff >>
rect -94 3927 -36 3939
rect -94 2145 -82 3927
rect -48 2145 -36 3927
rect -94 2133 -36 2145
rect 36 3927 94 3939
rect 36 2145 48 3927
rect 82 2145 94 3927
rect 36 2133 94 2145
rect -94 1903 -36 1915
rect -94 121 -82 1903
rect -48 121 -36 1903
rect -94 109 -36 121
rect 36 1903 94 1915
rect 36 121 48 1903
rect 82 121 94 1903
rect 36 109 94 121
rect -94 -121 -36 -109
rect -94 -1903 -82 -121
rect -48 -1903 -36 -121
rect -94 -1915 -36 -1903
rect 36 -121 94 -109
rect 36 -1903 48 -121
rect 82 -1903 94 -121
rect 36 -1915 94 -1903
rect -94 -2145 -36 -2133
rect -94 -3927 -82 -2145
rect -48 -3927 -36 -2145
rect -94 -3939 -36 -3927
rect 36 -2145 94 -2133
rect 36 -3927 48 -2145
rect 82 -3927 94 -2145
rect 36 -3939 94 -3927
<< ndiffc >>
rect -82 2145 -48 3927
rect 48 2145 82 3927
rect -82 121 -48 1903
rect 48 121 82 1903
rect -82 -1903 -48 -121
rect 48 -1903 82 -121
rect -82 -3927 -48 -2145
rect 48 -3927 82 -2145
<< psubdiff >>
rect -196 4079 -100 4113
rect 100 4079 196 4113
rect -196 4017 -162 4079
rect 162 4017 196 4079
rect -196 -4079 -162 -4017
rect 162 -4079 196 -4017
rect -196 -4113 -100 -4079
rect 100 -4113 196 -4079
<< psubdiffcont >>
rect -100 4079 100 4113
rect -196 -4017 -162 4017
rect 162 -4017 196 4017
rect -100 -4113 100 -4079
<< poly >>
rect -36 4011 36 4027
rect -36 3977 -20 4011
rect 20 3977 36 4011
rect -36 3939 36 3977
rect -36 2095 36 2133
rect -36 2061 -20 2095
rect 20 2061 36 2095
rect -36 2045 36 2061
rect -36 1987 36 2003
rect -36 1953 -20 1987
rect 20 1953 36 1987
rect -36 1915 36 1953
rect -36 71 36 109
rect -36 37 -20 71
rect 20 37 36 71
rect -36 21 36 37
rect -36 -37 36 -21
rect -36 -71 -20 -37
rect 20 -71 36 -37
rect -36 -109 36 -71
rect -36 -1953 36 -1915
rect -36 -1987 -20 -1953
rect 20 -1987 36 -1953
rect -36 -2003 36 -1987
rect -36 -2061 36 -2045
rect -36 -2095 -20 -2061
rect 20 -2095 36 -2061
rect -36 -2133 36 -2095
rect -36 -3977 36 -3939
rect -36 -4011 -20 -3977
rect 20 -4011 36 -3977
rect -36 -4027 36 -4011
<< polycont >>
rect -20 3977 20 4011
rect -20 2061 20 2095
rect -20 1953 20 1987
rect -20 37 20 71
rect -20 -71 20 -37
rect -20 -1987 20 -1953
rect -20 -2095 20 -2061
rect -20 -4011 20 -3977
<< locali >>
rect -196 4079 -100 4113
rect 100 4079 196 4113
rect -196 4017 -162 4079
rect 162 4017 196 4079
rect -36 3977 -20 4011
rect 20 3977 36 4011
rect -82 3927 -48 3943
rect -82 2129 -48 2145
rect 48 3927 82 3943
rect 48 2129 82 2145
rect -36 2061 -20 2095
rect 20 2061 36 2095
rect -36 1953 -20 1987
rect 20 1953 36 1987
rect -82 1903 -48 1919
rect -82 105 -48 121
rect 48 1903 82 1919
rect 48 105 82 121
rect -36 37 -20 71
rect 20 37 36 71
rect -36 -71 -20 -37
rect 20 -71 36 -37
rect -82 -121 -48 -105
rect -82 -1919 -48 -1903
rect 48 -121 82 -105
rect 48 -1919 82 -1903
rect -36 -1987 -20 -1953
rect 20 -1987 36 -1953
rect -36 -2095 -20 -2061
rect 20 -2095 36 -2061
rect -82 -2145 -48 -2129
rect -82 -3943 -48 -3927
rect 48 -2145 82 -2129
rect 48 -3943 82 -3927
rect -36 -4011 -20 -3977
rect 20 -4011 36 -3977
rect -196 -4079 -162 -4017
rect 162 -4079 196 -4017
rect -196 -4113 -100 -4079
rect 100 -4113 196 -4079
<< viali >>
rect -20 3977 20 4011
rect -82 2145 -48 3927
rect 48 2145 82 3927
rect -20 2061 20 2095
rect -20 1953 20 1987
rect -82 121 -48 1903
rect 48 121 82 1903
rect -20 37 20 71
rect -20 -71 20 -37
rect -82 -1903 -48 -121
rect 48 -1903 82 -121
rect -20 -1987 20 -1953
rect -20 -2095 20 -2061
rect -82 -3927 -48 -2145
rect 48 -3927 82 -2145
rect -20 -4011 20 -3977
<< metal1 >>
rect -32 4011 32 4017
rect -32 3977 -20 4011
rect 20 3977 32 4011
rect -32 3971 32 3977
rect -88 3927 -42 3939
rect -88 2145 -82 3927
rect -48 2145 -42 3927
rect -88 2133 -42 2145
rect 42 3927 88 3939
rect 42 2145 48 3927
rect 82 2145 88 3927
rect 42 2133 88 2145
rect -32 2095 32 2101
rect -32 2061 -20 2095
rect 20 2061 32 2095
rect -32 2055 32 2061
rect -32 1987 32 1993
rect -32 1953 -20 1987
rect 20 1953 32 1987
rect -32 1947 32 1953
rect -88 1903 -42 1915
rect -88 121 -82 1903
rect -48 121 -42 1903
rect -88 109 -42 121
rect 42 1903 88 1915
rect 42 121 48 1903
rect 82 121 88 1903
rect 42 109 88 121
rect -32 71 32 77
rect -32 37 -20 71
rect 20 37 32 71
rect -32 31 32 37
rect -32 -37 32 -31
rect -32 -71 -20 -37
rect 20 -71 32 -37
rect -32 -77 32 -71
rect -88 -121 -42 -109
rect -88 -1903 -82 -121
rect -48 -1903 -42 -121
rect -88 -1915 -42 -1903
rect 42 -121 88 -109
rect 42 -1903 48 -121
rect 82 -1903 88 -121
rect 42 -1915 88 -1903
rect -32 -1953 32 -1947
rect -32 -1987 -20 -1953
rect 20 -1987 32 -1953
rect -32 -1993 32 -1987
rect -32 -2061 32 -2055
rect -32 -2095 -20 -2061
rect 20 -2095 32 -2061
rect -32 -2101 32 -2095
rect -88 -2145 -42 -2133
rect -88 -3927 -82 -2145
rect -48 -3927 -42 -2145
rect -88 -3939 -42 -3927
rect 42 -2145 88 -2133
rect 42 -3927 48 -2145
rect 82 -3927 88 -2145
rect 42 -3939 88 -3927
rect -32 -3977 32 -3971
rect -32 -4011 -20 -3977
rect 20 -4011 32 -3977
rect -32 -4017 32 -4011
<< properties >>
string FIXED_BBOX -179 -4096 179 4096
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 9.028 l 0.361 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
