magic
tech sky130A
magscale 1 2
timestamp 1668114367
<< psubdiff >>
rect -10835 6139 -10678 6144
rect -9376 6139 -9219 6144
rect -10841 6120 -10817 6139
rect -9220 6120 -9196 6139
rect -10841 5954 -10835 6120
rect -9219 5954 -9196 6120
rect -3582 5300 -3524 5310
rect -4802 5234 -4778 5300
rect -3524 5234 -3500 5300
rect -10859 -141 -10835 -21
rect -9200 -141 -9176 -21
rect -10835 -165 -10678 -141
rect -9376 -165 -9219 -141
rect 16371 409 16762 433
rect -4818 -484 -4794 -418
rect -3500 -484 -3476 -418
rect -4770 -500 -4712 -484
rect -3582 -490 -3524 -484
rect 16371 -550 16762 -526
rect 11594 -950 11650 -942
rect 12386 -950 12442 -942
rect 11568 -1012 11592 -950
rect 12428 -966 12452 -950
rect 12442 -1012 12452 -966
rect 11562 -2658 11586 -2600
rect 12442 -2650 12464 -2600
rect 12440 -2658 12464 -2650
rect 11594 -2674 11650 -2658
rect 12386 -2674 12442 -2658
<< psubdiffcont >>
rect -10817 6120 -9220 6139
rect -10835 5954 -9219 6120
rect -10835 -21 -10678 5954
rect -9376 -21 -9219 5954
rect -4778 5234 -3524 5300
rect -10835 -141 -9200 -21
rect -4770 -418 -4712 5234
rect -3582 -418 -3524 5234
rect -4794 -484 -3500 -418
rect 16371 -526 16762 409
rect 11592 -966 12428 -950
rect 11592 -1012 12442 -966
rect 11594 -2600 11650 -1012
rect 12386 -2600 12442 -1012
rect 11586 -2650 12442 -2600
rect 11586 -2658 12440 -2650
<< locali >>
rect -10833 6136 -10817 6139
rect -10835 6120 -10817 6136
rect -9220 6120 -9204 6139
rect -9219 5954 -9204 6120
rect -9380 5178 -9376 5240
rect -3582 5300 -3524 5302
rect -4794 5240 -4778 5300
rect -9219 5234 -4778 5240
rect -3524 5234 -3508 5300
rect -9219 5178 -4770 5234
rect -10851 -141 -10835 -21
rect -9200 -141 -9184 -21
rect -10835 -157 -10678 -141
rect -9376 -157 -9219 -141
rect -3584 5074 -3582 5196
rect 4920 5196 5102 5197
rect -3524 5074 5102 5196
rect -4810 -484 -4794 -418
rect -3500 -484 -3484 -418
rect -4770 -492 -4712 -484
rect 4920 -1358 5102 5074
rect 15860 66 16249 499
rect 16371 409 16762 425
rect 15542 -680 15931 -247
rect 16371 -542 16762 -526
rect 11576 -1012 11592 -950
rect 12428 -966 12444 -950
rect 12442 -1012 12444 -966
rect 4920 -1460 11594 -1358
rect 11570 -2658 11586 -2600
rect 12442 -2650 12456 -2600
rect 12440 -2658 12456 -2650
rect 11594 -2666 11650 -2658
rect 12386 -2666 12442 -2658
<< viali >>
rect 11884 -2646 11918 -2610
<< metal1 >>
rect 12160 15706 12274 15718
rect 12160 15616 12174 15706
rect 12264 15616 12274 15706
rect 12160 15136 12274 15616
rect 12014 14972 12274 15136
rect 12014 14388 12188 14972
rect 11994 7232 12194 14388
rect 20136 7232 23624 7236
rect 11994 6964 23624 7232
rect 11994 5860 12194 6964
rect 11994 5842 12190 5860
rect 11266 5836 12190 5842
rect 9442 5832 12190 5836
rect 5786 5828 12190 5832
rect 3948 5824 12190 5828
rect 318 5822 12190 5824
rect -3232 5820 12190 5822
rect -5082 5818 12190 5820
rect -8278 5814 -7116 5816
rect -6022 5814 12190 5818
rect -9428 5810 12190 5814
rect -9632 5808 12190 5810
rect -9840 5792 12190 5808
rect -9840 5786 11310 5792
rect -9840 5782 9472 5786
rect -9840 5778 5816 5782
rect -9840 5774 3996 5778
rect -9840 5772 454 5774
rect -9840 5770 -5996 5772
rect -5082 5770 -3214 5772
rect -9840 5768 -9628 5770
rect -9428 5768 -8266 5770
rect -7158 5768 -5996 5770
rect -9840 5582 -9810 5768
rect -10078 5542 -9810 5582
rect -10192 148 -10158 5364
rect -10078 396 -10044 5542
rect -9888 5395 -9859 5542
rect 19960 5486 23624 6964
rect 4138 5476 11300 5478
rect 18103 5476 23624 5486
rect 4138 5467 23624 5476
rect -3183 5462 23624 5467
rect -4229 5458 23624 5462
rect -5264 5454 23624 5458
rect -6319 5452 23624 5454
rect -7377 5448 23624 5452
rect -8432 5446 23624 5448
rect -9502 5444 23624 5446
rect -9810 5419 23624 5444
rect -9810 5411 18284 5419
rect -9810 5407 -4184 5411
rect -3183 5410 18284 5411
rect -3183 5409 5970 5410
rect 11122 5408 18284 5410
rect -9810 5403 -5239 5407
rect -9810 5401 -6297 5403
rect -9810 5397 -7352 5401
rect -9810 5396 -8422 5397
rect -9502 5395 -8422 5396
rect -9888 5367 -9855 5395
rect -9883 5366 -9855 5367
rect -9883 5364 -9826 5366
rect -9964 148 -9930 5364
rect -9883 5333 -9816 5364
rect -9850 396 -9816 5333
rect -9736 148 -9702 5348
rect -7498 5074 -6336 5076
rect -5242 5074 -4238 5078
rect -8648 5070 -4238 5074
rect -8852 5068 -4238 5070
rect -9060 5032 -4238 5068
rect -9060 5030 -5216 5032
rect -9060 5028 -8848 5030
rect -8648 5028 -7486 5030
rect -6378 5028 -5216 5030
rect -9060 2670 -9030 5028
rect -9060 2644 -9028 2670
rect -9058 148 -9028 2644
rect -10420 120 -9028 148
rect -10420 114 -9032 120
rect -10420 112 -9702 114
rect -4580 -342 -4546 5032
rect -4386 -264 -4352 4739
rect -4272 -229 -4238 5032
rect -3967 4922 -3857 4924
rect -3967 4903 -3924 4922
rect -3968 4892 -3924 4903
rect -4158 4863 -3924 4892
rect -3865 4863 -3857 4922
rect -4158 4859 -3857 4863
rect -4158 -264 -4124 4859
rect -3967 4858 -3857 4859
rect -2972 4832 -2706 4834
rect -2972 4830 -2518 4832
rect -3748 4828 -2518 4830
rect -3748 4824 -2498 4828
rect -4004 4780 -2498 4824
rect -4004 4776 -2962 4780
rect -2856 4778 -2590 4780
rect -4004 4770 -3738 4776
rect -4386 -300 -4124 -264
rect -4158 -301 -4124 -300
rect -4044 -342 -4010 4739
rect -3930 3167 -3896 4739
rect -3022 3167 -2636 3168
rect -3930 3160 -2636 3167
rect -3930 3054 -2736 3160
rect -2646 3054 -2636 3160
rect -3930 3052 -2636 3054
rect -3930 -229 -3896 3052
rect -2556 2962 -2498 4780
rect 19960 4184 23624 5419
rect -2556 2956 -2496 2962
rect -2554 810 -2496 2956
rect -3294 790 -2496 810
rect -3302 674 -2496 790
rect 15544 734 15612 738
rect -3302 664 -2504 674
rect 10688 664 15612 734
rect -3302 -150 -3240 664
rect -3328 -166 -3088 -150
rect -3328 -272 -3188 -166
rect -3098 -272 -3088 -166
rect -3328 -286 -3088 -272
rect -4580 -370 -3980 -342
rect -4580 -372 -4546 -370
rect 10688 -682 10752 664
rect 15542 437 15612 664
rect 12541 378 12794 383
rect 12541 318 12814 378
rect 12541 171 12612 318
rect 10688 -766 10762 -682
rect 10692 -818 10762 -766
rect 12540 -770 12611 -637
rect 12015 -818 12612 -770
rect 10689 -822 12612 -818
rect 12782 -821 12814 318
rect 10689 -869 12089 -822
rect 12540 -825 12611 -822
rect 11942 -1060 12008 -1059
rect 12044 -1060 12089 -869
rect 11942 -1092 12121 -1060
rect 11942 -1093 12008 -1092
rect 11883 -2576 11917 -1127
rect 12001 -1176 12035 -1127
rect 12090 -1176 12121 -1092
rect 12001 -1214 12121 -1176
rect 12778 -1114 12894 -821
rect 16178 -884 16248 -592
rect 19960 -884 20376 4184
rect 12778 -1204 12780 -1114
rect 12886 -1204 12894 -1114
rect 16174 -1152 20396 -884
rect 16178 -1160 16248 -1152
rect 12778 -1214 12894 -1204
rect 12001 -2469 12035 -1214
rect 12090 -1215 12121 -1214
rect 11882 -2596 11917 -2576
rect 11882 -2604 11930 -2596
rect 11874 -2610 11930 -2604
rect 11874 -2646 11884 -2610
rect 11918 -2646 11930 -2610
rect 11874 -2650 11930 -2646
rect 11876 -2652 11930 -2650
rect 11882 -2658 11930 -2652
rect 11609 -2985 11742 -2980
rect 11882 -2985 11917 -2658
rect 11609 -3004 11917 -2985
rect 11169 -3006 11917 -3004
rect 11169 -3112 11179 -3006
rect 11269 -3016 11917 -3006
rect 11269 -3022 11742 -3016
rect 11269 -3112 11639 -3022
rect 11169 -3120 11639 -3112
rect -12830 -12434 -12666 -11710
rect -11458 -12434 -9328 -12386
rect -12830 -12608 -9328 -12434
rect -12830 -12616 -10162 -12608
rect -12670 -12994 -10162 -12616
rect -11458 -13222 -10162 -12994
rect -9446 -13222 -9328 -12608
rect -11458 -13408 -9328 -13222
<< via1 >>
rect 12174 15616 12264 15706
rect -3924 4863 -3865 4922
rect -2736 3054 -2646 3160
rect -3188 -272 -3098 -166
rect 12780 -1204 12886 -1114
rect 11179 -3112 11269 -3006
rect -10162 -13222 -9446 -12608
<< metal2 >>
rect 12222 18274 12376 18290
rect 12222 18150 12232 18274
rect 12366 18150 12376 18274
rect 12222 17998 12376 18150
rect 12224 15718 12376 17998
rect 12160 15706 12376 15718
rect 12160 15616 12174 15706
rect 12264 15616 12376 15706
rect 12160 15602 12376 15616
rect -3929 4922 -3859 4936
rect -3929 4863 -3924 4922
rect -3865 4863 -3859 4922
rect -3929 4767 -3859 4863
rect -3930 4751 -3859 4767
rect -3930 4739 -3896 4751
rect -2752 3160 -2080 3176
rect -2752 3054 -2736 3160
rect -2646 3156 -2080 3160
rect -2646 3056 -2172 3156
rect -2090 3056 -2080 3156
rect -2646 3054 -2080 3056
rect -2752 3042 -2080 3054
rect -3204 -166 -2532 -150
rect -3204 -272 -3188 -166
rect -3098 -170 -2532 -166
rect -3098 -270 -2624 -170
rect -2542 -270 -2532 -170
rect -3098 -272 -2532 -270
rect -3204 -284 -2532 -272
rect 12768 -1114 12902 -1098
rect 12768 -1204 12780 -1114
rect 12886 -1204 12902 -1114
rect 12768 -1678 12902 -1204
rect 12768 -1760 12782 -1678
rect 12882 -1760 12902 -1678
rect 12768 -1770 12902 -1760
rect 10613 -3006 11285 -2994
rect 10613 -3008 11179 -3006
rect 10613 -3108 10623 -3008
rect 10705 -3108 11179 -3008
rect 10613 -3112 11179 -3108
rect 11269 -3112 11285 -3006
rect 10613 -3128 11285 -3112
rect -10334 -12472 -8220 -12300
rect -10334 -12608 -7008 -12472
rect -10334 -13222 -10162 -12608
rect -9446 -12692 -7008 -12608
rect -9446 -13222 -7724 -12692
rect -10334 -13290 -7724 -13222
rect -7060 -13290 -7008 -12692
rect -10334 -13442 -7008 -13290
rect -10334 -13630 -8220 -13442
<< via2 >>
rect 12232 18150 12366 18274
rect -2172 3056 -2090 3156
rect -2624 -270 -2542 -170
rect 12782 -1760 12882 -1678
rect 10623 -3108 10705 -3008
rect -7724 -13290 -7060 -12692
<< metal3 >>
rect 12222 18812 12376 18822
rect 12222 18690 12234 18812
rect 12362 18690 12376 18812
rect 12222 18274 12376 18690
rect 12222 18150 12232 18274
rect 12366 18150 12376 18274
rect 12222 18138 12376 18150
rect -2188 3156 -1704 3170
rect -2188 3056 -2172 3156
rect -2090 3148 -1704 3156
rect -2090 3056 -1792 3148
rect -2188 3048 -1792 3056
rect -1710 3048 -1704 3148
rect -2188 3042 -1704 3048
rect -2640 -170 -2156 -156
rect -2640 -270 -2624 -170
rect -2542 -178 -2156 -170
rect -2542 -270 -2244 -178
rect -2640 -278 -2244 -270
rect -2162 -278 -2156 -178
rect -2640 -284 -2156 -278
rect 12768 -1678 12896 -1662
rect 12768 -1760 12782 -1678
rect 12882 -1760 12896 -1678
rect 12768 -2058 12896 -1760
rect 12768 -2140 12774 -2058
rect 12874 -2140 12896 -2058
rect 12768 -2146 12896 -2140
rect 10237 -3000 10721 -2994
rect 10237 -3100 10243 -3000
rect 10325 -3008 10721 -3000
rect 10325 -3100 10623 -3008
rect 10237 -3108 10623 -3100
rect 10705 -3108 10721 -3008
rect 10237 -3122 10721 -3108
rect -7862 -12692 -5372 -12540
rect -7862 -13290 -7724 -12692
rect -7060 -12710 -5372 -12692
rect -7060 -13290 -6156 -12710
rect -5474 -13290 -5372 -12710
rect -7862 -13494 -5372 -13290
<< via3 >>
rect 12234 18690 12362 18812
rect -1792 3048 -1710 3148
rect -2244 -278 -2162 -178
rect 12774 -2140 12874 -2058
rect 10243 -3100 10325 -3000
rect -6156 -13290 -5474 -12710
<< metal4 >>
rect -14426 108220 -10732 108236
rect -74552 105142 -10732 108220
rect -74524 38474 -73976 105142
rect -14426 95268 -10732 105142
rect -14426 95062 -10530 95268
rect -14426 92162 -14028 95062
rect -10978 92162 -10530 95062
rect -14426 91956 -10530 92162
rect -14426 91564 -10732 91956
rect -74524 38414 -43004 38474
rect -74524 37878 -42740 38414
rect -43256 14624 -42740 37878
rect -2422 37134 948 37444
rect -2422 34974 -1756 37134
rect 700 34974 948 37134
rect -2422 34644 948 34974
rect -3326 31444 574 31449
rect -3326 29194 3120 31444
rect -3326 29034 3122 29194
rect -3326 29025 574 29034
rect -3319 28424 -1362 29025
rect -3319 27093 -3158 28424
rect -1463 27093 -1362 28424
rect -3319 26992 -1362 27093
rect 1258 26950 3122 29034
rect 9000 26950 9318 26958
rect 1258 26352 9318 26950
rect 9000 23118 9318 26352
rect 16060 23290 16738 23780
rect 16030 23286 16738 23290
rect 13764 23162 16738 23286
rect 13764 23160 16210 23162
rect 8958 23036 12366 23118
rect 8958 22928 9068 23036
rect 10130 22892 10234 23036
rect 11300 22920 11402 23036
rect 12192 23034 12366 23036
rect 4708 19556 5026 19562
rect 8448 19556 8558 19696
rect 4708 19482 8558 19556
rect 9622 19482 9732 19704
rect 10790 19482 10900 19698
rect 4708 19396 10900 19482
rect 12224 19462 12366 23034
rect 13764 22928 13868 23160
rect 14936 22928 15038 23160
rect 16106 22928 16210 23160
rect 13332 19718 13358 19722
rect 13252 19462 13362 19716
rect 14422 19462 14532 19704
rect 15596 19462 15700 19708
rect 12224 19458 15700 19462
rect 4708 19018 5026 19396
rect 8448 19392 10900 19396
rect 12222 19336 15700 19458
rect 12222 19334 13246 19336
rect 12222 19240 12376 19334
rect 4708 18934 12372 19018
rect 4708 18812 12376 18934
rect 4708 18690 12234 18812
rect 12362 18690 12376 18812
rect 4708 18678 12376 18690
rect 4708 15760 5026 18678
rect 12222 18670 12376 18678
rect 4708 15750 5036 15760
rect 4698 14624 5036 15750
rect -43258 14026 5036 14624
rect -43258 14016 4970 14026
rect 119418 12528 121128 12672
rect 118990 11886 121128 12528
rect 118276 11748 122126 11886
rect 127318 11748 127974 21024
rect 118276 10604 127974 11748
rect 118276 10602 119986 10604
rect 117062 10030 119986 10602
rect 116204 9962 119986 10030
rect 120416 10510 127974 10604
rect 120416 10320 127556 10510
rect 120416 9962 122126 10320
rect 116204 8678 118772 9962
rect 116204 8308 117914 8678
rect 114922 8106 117914 8308
rect 114922 7702 116632 8106
rect 113890 6562 116632 7702
rect 112572 6384 116632 6562
rect 112572 4816 115600 6384
rect 112572 4568 114282 4816
rect 111788 3676 114282 4568
rect -1804 3148 -1643 3158
rect -1804 3048 -1792 3148
rect -1710 3048 -1643 3148
rect -1804 3038 -1643 3048
rect -1803 2938 -1647 3038
rect 1404 2982 1685 3201
rect 598 2940 1685 2982
rect 596 2938 1685 2940
rect -2053 2911 1685 2938
rect -2053 2849 659 2911
rect -1482 2770 -1378 2849
rect -464 2771 -360 2849
rect 544 2771 659 2849
rect -1923 -168 -1813 -44
rect -2256 -172 -1813 -168
rect -903 -172 -799 -47
rect 116 -172 220 -47
rect -2256 -178 686 -172
rect -2256 -278 -2244 -178
rect -2162 -278 686 -178
rect -2256 -288 686 -278
rect -1840 -608 -1503 -288
rect -7700 -769 -1503 -608
rect -7700 -1431 -7640 -769
rect -6676 -1431 -1503 -769
rect -7700 -1552 -1503 -1431
rect -1840 -1553 -1503 -1552
rect 1404 -3215 1685 2911
rect 111788 2466 113498 3676
rect 109830 1682 113498 2466
rect 109830 -1844 112642 1682
rect 12764 -2058 12884 -2046
rect 12764 -2140 12774 -2058
rect 12874 -2140 12884 -2058
rect 12764 -2249 12884 -2140
rect 12752 -2519 12939 -2249
rect 12698 -2665 12939 -2519
rect 3171 -2978 5778 -2970
rect 3171 -2990 10134 -2978
rect 3171 -3000 10337 -2990
rect 3171 -3057 10243 -3000
rect -4398 -4109 1711 -3215
rect 3171 -3425 3243 -3057
rect 3561 -3100 10243 -3057
rect 10325 -3100 10337 -3000
rect 3561 -3110 10337 -3100
rect 3561 -3165 10134 -3110
rect 12698 -3127 12914 -2665
rect 105234 -3126 112642 -1844
rect 3561 -3425 5778 -3165
rect 3171 -3483 5778 -3425
rect -4398 -6488 -3094 -4109
rect -20648 -6606 -3094 -6488
rect -21348 -9656 -3094 -6606
rect -21348 -9692 -3122 -9656
rect -21348 -11652 -19660 -9692
rect 12347 -11292 12982 -3127
rect 105234 -10052 110862 -3126
rect 12347 -11697 12401 -11292
rect 12941 -11697 12982 -11292
rect 12347 -11751 12982 -11697
rect -6292 -12692 -3718 -12590
rect -6292 -12710 -4384 -12692
rect -6292 -13290 -6156 -12710
rect -5474 -13256 -4384 -12710
rect -3754 -13256 -3718 -12692
rect 57958 -12742 110862 -10052
rect 3806 -12852 4130 -12825
rect 57958 -12852 105602 -12742
rect -5474 -13290 -3718 -13256
rect 3755 -12870 105602 -12852
rect 3755 -13273 59016 -12870
rect 3755 -13290 58709 -13273
rect -6292 -13442 -3718 -13290
rect 3806 -14863 4130 -13290
rect 3806 -14876 9858 -14863
rect 3433 -14978 9858 -14876
rect 3433 -14990 9891 -14978
rect 4266 -15282 4369 -14990
rect 6109 -15281 6213 -14990
rect 7947 -15280 8051 -14990
rect 9787 -15281 9891 -14990
rect 3447 -22395 3538 -22151
rect 3440 -22399 3897 -22395
rect 5291 -22399 5382 -22151
rect 7127 -22399 7218 -22152
rect 8960 -22399 9051 -22152
rect 3440 -22533 9924 -22399
rect 5005 -23084 5301 -22533
rect 4768 -23822 5588 -23084
<< via4 >>
rect -14028 92162 -10978 95062
rect -1756 34974 700 37134
rect -3158 27093 -1463 28424
rect -7640 -1431 -6676 -769
rect 3243 -3425 3561 -3057
rect 12401 -11697 12941 -11292
rect -4384 -13256 -3754 -12692
<< metal5 >>
rect -14216 95062 -10604 95120
rect -14216 92162 -14028 95062
rect -10978 92162 -10604 95062
rect -14216 80710 -10604 92162
rect -2376 78208 662 78210
rect 1106 78208 4698 81418
rect -5366 78204 4698 78208
rect -8312 78182 4698 78204
rect -8386 76612 4698 78182
rect -8386 76610 -2328 76612
rect 634 76610 4698 76612
rect -8386 76606 -5274 76610
rect -8386 75000 -5332 76606
rect 1106 76598 4698 76610
rect -8386 69974 -5330 75000
rect -8284 69964 -5330 69974
rect -1892 39558 890 67140
rect -1880 37134 860 39558
rect -1880 34974 -1756 37134
rect 700 34974 860 37134
rect -1880 34800 860 34974
rect -38928 -695 -6516 -611
rect -69916 -769 -6516 -695
rect -69916 -1431 -7640 -769
rect -6676 -1431 -6516 -769
rect -69916 -1590 -6516 -1431
rect -69916 -1674 -38628 -1590
rect -68712 -28661 -67840 -1674
rect 3192 -3057 3605 -2971
rect 3192 -3425 3243 -3057
rect 3561 -3425 3605 -3057
rect 3192 -5356 3605 -3425
rect 3192 -8176 6555 -5356
rect 3192 -8829 3605 -8176
rect 217 -9405 3605 -8829
rect 219 -12637 973 -9405
rect 3192 -9407 3605 -9405
rect 1748 -11292 12999 -11213
rect 1748 -11383 12401 -11292
rect -4502 -12692 973 -12637
rect -4502 -13256 -4384 -12692
rect -3754 -13256 973 -12692
rect -4502 -13260 973 -13256
rect 1662 -11697 12401 -11383
rect 12941 -11697 12999 -11292
rect 1662 -11769 12999 -11697
rect -4502 -13391 908 -13260
rect 1662 -28336 2090 -11769
rect 68184 -27520 68988 -25318
rect 62230 -28162 68988 -27520
rect 119854 -27752 121030 -27712
rect 119402 -28162 121030 -27752
rect 62230 -28336 121030 -28162
rect -34584 -28361 121030 -28336
rect -38928 -28661 121030 -28361
rect -68712 -29560 121030 -28661
rect -68078 -29561 121030 -29560
rect -68078 -29567 -34519 -29561
rect -68078 -29640 -36790 -29567
rect 62230 -29694 121030 -29561
rect 62230 -29742 68940 -29694
rect 119854 -29704 121030 -29694
use LG  LG_0
timestamp 1668113732
transform -1 0 117890 0 1 55546
box -81282 -83494 47246 55400
use LS  LS_0
timestamp 1668104415
transform 1 0 -18930 0 1 -2358
box -34810 -19320 6180 -3320
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC1
timestamp 1667951165
transform 1 0 9723 0 1 21290
box -1711 -1620 1710 1640
use sky130_fd_pr__cap_mim_m3_1_FLZ2GZ  XC3
timestamp 1667951165
transform 1 0 6250 0 1 -18718
box -3568 -3440 3668 3440
use sky130_fd_pr__cap_mim_m3_1_HYGCGT  XC4
timestamp 1667951165
transform 1 0 14527 0 1 21308
box -1711 -1620 1710 1640
use sky130_fd_pr__nfet_01v8_TAQE79  XM2
timestamp 1668019001
transform 1 0 -9947 0 1 2880
box -257 -2568 257 2568
use sky130_fd_pr__nfet_01v8_PAV6Y8  XM3
timestamp 1668017392
transform 1 0 11959 0 1 -1798
box -88 -755 88 755
use ind1p2n  ind1p2n_0
timestamp 1667951165
transform -1 0 -40100 0 -1 13436
box -39200 -37500 -3800 -2500
use ind2p69  ind2p69_0
timestamp 1667951165
transform -1 0 -60784 0 -1 57164
box -53200 -45000 5400 5000
use ind2p69  ind2p69_1
timestamp 1667951165
transform 1 0 51308 0 -1 54230
box -53200 -45000 5400 5000
use sky130_fd_pr__cap_mim_m3_1_LJH8TW  sky130_fd_pr__cap_mim_m3_1_LJH8TW_1
timestamp 1667951165
transform 1 0 -801 0 1 1362
box -1489 -1410 1488 1410
use sky130_fd_pr__nfet_01v8_TAQE79  sky130_fd_pr__nfet_01v8_TAQE79_0
timestamp 1668019001
transform 1 0 -4141 0 1 2255
box -257 -2568 257 2568
use sky130_fd_pr__res_xhigh_po_0p35_BZ5JJG  sky130_fd_pr__res_xhigh_po_0p35_BZ5JJG_0
timestamp 1667951165
transform -1 0 15895 0 -1 -91
box -355 -589 355 589
use sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ  sky130_fd_pr__res_xhigh_po_0p35_NE8FRQ_0
timestamp 1667951165
transform -1 0 12576 0 1 -217
box -37 -502 37 502
<< labels >>
rlabel metal4 16310 23440 16548 23660 1 RFOUT
port 1 n
rlabel metal4 4768 -23822 5588 -23084 1 RFIN
port 2 n
rlabel metal5 3996 -7994 6312 -5678 1 GND
port 3 n
rlabel metal1 20408 4420 23150 6956 1 VDD
port 4 n
<< properties >>
string LEFview true
<< end >>
