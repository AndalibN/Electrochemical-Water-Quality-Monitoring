magic
tech sky130A
timestamp 1667254537
<< nmos >>
rect -25 -5000 25 5000
<< ndiff >>
rect -54 4994 -25 5000
rect -54 -4994 -48 4994
rect -31 -4994 -25 4994
rect -54 -5000 -25 -4994
rect 25 4994 54 5000
rect 25 -4994 31 4994
rect 48 -4994 54 4994
rect 25 -5000 54 -4994
<< ndiffc >>
rect -48 -4994 -31 4994
rect 31 -4994 48 4994
<< poly >>
rect -25 5036 25 5044
rect -25 5019 -17 5036
rect 17 5019 25 5036
rect -25 5000 25 5019
rect -25 -5019 25 -5000
rect -25 -5036 -17 -5019
rect 17 -5036 25 -5019
rect -25 -5044 25 -5036
<< polycont >>
rect -17 5019 17 5036
rect -17 -5036 17 -5019
<< locali >>
rect -25 5019 -17 5036
rect 17 5019 25 5036
rect -48 4994 -31 5002
rect -48 -5002 -31 -4994
rect 31 4994 48 5002
rect 31 -5002 48 -4994
rect -25 -5036 -17 -5019
rect 17 -5036 25 -5019
<< viali >>
rect -17 5019 17 5036
rect -48 -4994 -31 4994
rect 31 -4994 48 4994
rect -17 -5036 17 -5019
<< metal1 >>
rect -23 5036 23 5039
rect -23 5019 -17 5036
rect 17 5019 23 5036
rect -23 5016 23 5019
rect -51 4994 -28 5000
rect -51 -4994 -48 4994
rect -31 -4994 -28 4994
rect -51 -5000 -28 -4994
rect 28 4994 51 5000
rect 28 -4994 31 4994
rect 48 -4994 51 4994
rect 28 -5000 51 -4994
rect -23 -5019 23 -5016
rect -23 -5036 -17 -5019
rect 17 -5036 23 -5019
rect -23 -5039 23 -5036
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 100.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
