magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< nwell >>
rect -223 -5100 223 5100
<< pmos >>
rect -129 -5000 -29 5000
rect 29 -5000 129 5000
<< pdiff >>
rect -187 4988 -129 5000
rect -187 -4988 -175 4988
rect -141 -4988 -129 4988
rect -187 -5000 -129 -4988
rect -29 4988 29 5000
rect -29 -4988 -17 4988
rect 17 -4988 29 4988
rect -29 -5000 29 -4988
rect 129 4988 187 5000
rect 129 -4988 141 4988
rect 175 -4988 187 4988
rect 129 -5000 187 -4988
<< pdiffc >>
rect -175 -4988 -141 4988
rect -17 -4988 17 4988
rect 141 -4988 175 4988
<< poly >>
rect -129 5081 -29 5097
rect -129 5047 -113 5081
rect -45 5047 -29 5081
rect -129 5000 -29 5047
rect 29 5081 129 5097
rect 29 5047 45 5081
rect 113 5047 129 5081
rect 29 5000 129 5047
rect -129 -5047 -29 -5000
rect -129 -5081 -113 -5047
rect -45 -5081 -29 -5047
rect -129 -5097 -29 -5081
rect 29 -5047 129 -5000
rect 29 -5081 45 -5047
rect 113 -5081 129 -5047
rect 29 -5097 129 -5081
<< polycont >>
rect -113 5047 -45 5081
rect 45 5047 113 5081
rect -113 -5081 -45 -5047
rect 45 -5081 113 -5047
<< locali >>
rect -129 5047 -113 5081
rect -45 5047 -29 5081
rect 29 5047 45 5081
rect 113 5047 129 5081
rect -175 4988 -141 5004
rect -175 -5004 -141 -4988
rect -17 4988 17 5004
rect -17 -5004 17 -4988
rect 141 4988 175 5004
rect 141 -5004 175 -4988
rect -129 -5081 -113 -5047
rect -45 -5081 -29 -5047
rect 29 -5081 45 -5047
rect 113 -5081 129 -5047
<< viali >>
rect -113 5047 -45 5081
rect 45 5047 113 5081
rect -175 -4988 -141 4988
rect -17 -4988 17 4988
rect 141 -4988 175 4988
rect -113 -5081 -45 -5047
rect 45 -5081 113 -5047
<< metal1 >>
rect -125 5081 -33 5087
rect -125 5047 -113 5081
rect -45 5047 -33 5081
rect -125 5041 -33 5047
rect 33 5081 125 5087
rect 33 5047 45 5081
rect 113 5047 125 5081
rect 33 5041 125 5047
rect -181 4988 -135 5000
rect -181 -4988 -175 4988
rect -141 -4988 -135 4988
rect -181 -5000 -135 -4988
rect -23 4988 23 5000
rect -23 -4988 -17 4988
rect 17 -4988 23 4988
rect -23 -5000 23 -4988
rect 135 4988 181 5000
rect 135 -4988 141 4988
rect 175 -4988 181 4988
rect 135 -5000 181 -4988
rect -125 -5047 -33 -5041
rect -125 -5081 -113 -5047
rect -45 -5081 -33 -5047
rect -125 -5087 -33 -5081
rect 33 -5047 125 -5041
rect 33 -5081 45 -5047
rect 113 -5081 125 -5047
rect 33 -5087 125 -5081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 50.0 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
