magic
tech sky130A
magscale 1 2
timestamp 1666102132
<< pwell >>
rect -246 -1319 246 1319
<< nmos >>
rect -50 109 50 1109
rect -50 -1109 50 -109
<< ndiff >>
rect -108 1097 -50 1109
rect -108 121 -96 1097
rect -62 121 -50 1097
rect -108 109 -50 121
rect 50 1097 108 1109
rect 50 121 62 1097
rect 96 121 108 1097
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -1097 -96 -121
rect -62 -1097 -50 -121
rect -108 -1109 -50 -1097
rect 50 -121 108 -109
rect 50 -1097 62 -121
rect 96 -1097 108 -121
rect 50 -1109 108 -1097
<< ndiffc >>
rect -96 121 -62 1097
rect 62 121 96 1097
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
<< psubdiff >>
rect -210 1249 -114 1283
rect 114 1249 210 1283
rect -210 1187 -176 1249
rect 176 1187 210 1249
rect -210 -1249 -176 -1187
rect 176 -1249 210 -1187
rect -210 -1283 -114 -1249
rect 114 -1283 210 -1249
<< psubdiffcont >>
rect -114 1249 114 1283
rect -210 -1187 -176 1187
rect 176 -1187 210 1187
rect -114 -1283 114 -1249
<< poly >>
rect -50 1181 50 1197
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -50 1109 50 1147
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -1147 50 -1109
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1197 50 -1181
<< polycont >>
rect -34 1147 34 1181
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1181 34 -1147
<< locali >>
rect -210 1249 -114 1283
rect 114 1249 210 1283
rect -210 1187 -176 1249
rect 176 1187 210 1249
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -96 1097 -62 1113
rect -96 105 -62 121
rect 62 1097 96 1113
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -1113 -62 -1097
rect 62 -121 96 -105
rect 62 -1113 96 -1097
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -210 -1249 -176 -1187
rect 176 -1249 210 -1187
rect -210 -1283 -114 -1249
rect 114 -1283 210 -1249
<< viali >>
rect -34 1147 34 1181
rect -96 121 -62 1097
rect 62 121 96 1097
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -34 -1181 34 -1147
<< metal1 >>
rect -46 1181 46 1187
rect -46 1147 -34 1181
rect 34 1147 46 1181
rect -46 1141 46 1147
rect -102 1097 -56 1109
rect -102 121 -96 1097
rect -62 121 -56 1097
rect -102 109 -56 121
rect 56 1097 102 1109
rect 56 121 62 1097
rect 96 121 102 1097
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -1097 -96 -121
rect -62 -1097 -56 -121
rect -102 -1109 -56 -1097
rect 56 -121 102 -109
rect 56 -1097 62 -121
rect 96 -1097 102 -121
rect 56 -1109 102 -1097
rect -46 -1147 46 -1141
rect -46 -1181 -34 -1147
rect 34 -1181 46 -1147
rect -46 -1187 46 -1181
<< properties >>
string FIXED_BBOX -193 -1266 193 1266
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
