magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -184 -544 184 578
<< pmos >>
rect -90 -444 90 516
<< pdiff >>
rect -148 495 -90 516
rect -148 461 -136 495
rect -102 461 -90 495
rect -148 427 -90 461
rect -148 393 -136 427
rect -102 393 -90 427
rect -148 359 -90 393
rect -148 325 -136 359
rect -102 325 -90 359
rect -148 291 -90 325
rect -148 257 -136 291
rect -102 257 -90 291
rect -148 223 -90 257
rect -148 189 -136 223
rect -102 189 -90 223
rect -148 155 -90 189
rect -148 121 -136 155
rect -102 121 -90 155
rect -148 87 -90 121
rect -148 53 -136 87
rect -102 53 -90 87
rect -148 19 -90 53
rect -148 -15 -136 19
rect -102 -15 -90 19
rect -148 -49 -90 -15
rect -148 -83 -136 -49
rect -102 -83 -90 -49
rect -148 -117 -90 -83
rect -148 -151 -136 -117
rect -102 -151 -90 -117
rect -148 -185 -90 -151
rect -148 -219 -136 -185
rect -102 -219 -90 -185
rect -148 -253 -90 -219
rect -148 -287 -136 -253
rect -102 -287 -90 -253
rect -148 -321 -90 -287
rect -148 -355 -136 -321
rect -102 -355 -90 -321
rect -148 -389 -90 -355
rect -148 -423 -136 -389
rect -102 -423 -90 -389
rect -148 -444 -90 -423
rect 90 495 148 516
rect 90 461 102 495
rect 136 461 148 495
rect 90 427 148 461
rect 90 393 102 427
rect 136 393 148 427
rect 90 359 148 393
rect 90 325 102 359
rect 136 325 148 359
rect 90 291 148 325
rect 90 257 102 291
rect 136 257 148 291
rect 90 223 148 257
rect 90 189 102 223
rect 136 189 148 223
rect 90 155 148 189
rect 90 121 102 155
rect 136 121 148 155
rect 90 87 148 121
rect 90 53 102 87
rect 136 53 148 87
rect 90 19 148 53
rect 90 -15 102 19
rect 136 -15 148 19
rect 90 -49 148 -15
rect 90 -83 102 -49
rect 136 -83 148 -49
rect 90 -117 148 -83
rect 90 -151 102 -117
rect 136 -151 148 -117
rect 90 -185 148 -151
rect 90 -219 102 -185
rect 136 -219 148 -185
rect 90 -253 148 -219
rect 90 -287 102 -253
rect 136 -287 148 -253
rect 90 -321 148 -287
rect 90 -355 102 -321
rect 136 -355 148 -321
rect 90 -389 148 -355
rect 90 -423 102 -389
rect 136 -423 148 -389
rect 90 -444 148 -423
<< pdiffc >>
rect -136 461 -102 495
rect -136 393 -102 427
rect -136 325 -102 359
rect -136 257 -102 291
rect -136 189 -102 223
rect -136 121 -102 155
rect -136 53 -102 87
rect -136 -15 -102 19
rect -136 -83 -102 -49
rect -136 -151 -102 -117
rect -136 -219 -102 -185
rect -136 -287 -102 -253
rect -136 -355 -102 -321
rect -136 -423 -102 -389
rect 102 461 136 495
rect 102 393 136 427
rect 102 325 136 359
rect 102 257 136 291
rect 102 189 136 223
rect 102 121 136 155
rect 102 53 136 87
rect 102 -15 136 19
rect 102 -83 136 -49
rect 102 -151 136 -117
rect 102 -219 136 -185
rect 102 -287 136 -253
rect 102 -355 136 -321
rect 102 -423 136 -389
<< poly >>
rect -90 516 90 542
rect -90 -491 90 -444
rect -90 -525 -51 -491
rect -17 -525 17 -491
rect 51 -525 90 -491
rect -90 -541 90 -525
<< polycont >>
rect -51 -525 -17 -491
rect 17 -525 51 -491
<< locali >>
rect -136 495 -102 520
rect -136 427 -102 451
rect -136 359 -102 379
rect -136 291 -102 307
rect -136 223 -102 235
rect -136 155 -102 163
rect -136 87 -102 91
rect -136 -19 -102 -15
rect -136 -91 -102 -83
rect -136 -163 -102 -151
rect -136 -235 -102 -219
rect -136 -307 -102 -287
rect -136 -379 -102 -355
rect -136 -448 -102 -423
rect 102 495 136 520
rect 102 427 136 451
rect 102 359 136 379
rect 102 291 136 307
rect 102 223 136 235
rect 102 155 136 163
rect 102 87 136 91
rect 102 -19 136 -15
rect 102 -91 136 -83
rect 102 -163 136 -151
rect 102 -235 136 -219
rect 102 -307 136 -287
rect 102 -379 136 -355
rect 102 -448 136 -423
rect -90 -525 -53 -491
rect -17 -525 17 -491
rect 53 -525 90 -491
<< viali >>
rect -136 461 -102 485
rect -136 451 -102 461
rect -136 393 -102 413
rect -136 379 -102 393
rect -136 325 -102 341
rect -136 307 -102 325
rect -136 257 -102 269
rect -136 235 -102 257
rect -136 189 -102 197
rect -136 163 -102 189
rect -136 121 -102 125
rect -136 91 -102 121
rect -136 19 -102 53
rect -136 -49 -102 -19
rect -136 -53 -102 -49
rect -136 -117 -102 -91
rect -136 -125 -102 -117
rect -136 -185 -102 -163
rect -136 -197 -102 -185
rect -136 -253 -102 -235
rect -136 -269 -102 -253
rect -136 -321 -102 -307
rect -136 -341 -102 -321
rect -136 -389 -102 -379
rect -136 -413 -102 -389
rect 102 461 136 485
rect 102 451 136 461
rect 102 393 136 413
rect 102 379 136 393
rect 102 325 136 341
rect 102 307 136 325
rect 102 257 136 269
rect 102 235 136 257
rect 102 189 136 197
rect 102 163 136 189
rect 102 121 136 125
rect 102 91 136 121
rect 102 19 136 53
rect 102 -49 136 -19
rect 102 -53 136 -49
rect 102 -117 136 -91
rect 102 -125 136 -117
rect 102 -185 136 -163
rect 102 -197 136 -185
rect 102 -253 136 -235
rect 102 -269 136 -253
rect 102 -321 136 -307
rect 102 -341 136 -321
rect 102 -389 136 -379
rect 102 -413 136 -389
rect -53 -525 -51 -491
rect -51 -525 -19 -491
rect 19 -525 51 -491
rect 51 -525 53 -491
<< metal1 >>
rect -142 485 -96 516
rect -142 451 -136 485
rect -102 451 -96 485
rect -142 413 -96 451
rect -142 379 -136 413
rect -102 379 -96 413
rect -142 341 -96 379
rect -142 307 -136 341
rect -102 307 -96 341
rect -142 269 -96 307
rect -142 235 -136 269
rect -102 235 -96 269
rect -142 197 -96 235
rect -142 163 -136 197
rect -102 163 -96 197
rect -142 125 -96 163
rect -142 91 -136 125
rect -102 91 -96 125
rect -142 53 -96 91
rect -142 19 -136 53
rect -102 19 -96 53
rect -142 -19 -96 19
rect -142 -53 -136 -19
rect -102 -53 -96 -19
rect -142 -91 -96 -53
rect -142 -125 -136 -91
rect -102 -125 -96 -91
rect -142 -163 -96 -125
rect -142 -197 -136 -163
rect -102 -197 -96 -163
rect -142 -235 -96 -197
rect -142 -269 -136 -235
rect -102 -269 -96 -235
rect -142 -307 -96 -269
rect -142 -341 -136 -307
rect -102 -341 -96 -307
rect -142 -379 -96 -341
rect -142 -413 -136 -379
rect -102 -413 -96 -379
rect -142 -444 -96 -413
rect 96 485 142 516
rect 96 451 102 485
rect 136 451 142 485
rect 96 413 142 451
rect 96 379 102 413
rect 136 379 142 413
rect 96 341 142 379
rect 96 307 102 341
rect 136 307 142 341
rect 96 269 142 307
rect 96 235 102 269
rect 136 235 142 269
rect 96 197 142 235
rect 96 163 102 197
rect 136 163 142 197
rect 96 125 142 163
rect 96 91 102 125
rect 136 91 142 125
rect 96 53 142 91
rect 96 19 102 53
rect 136 19 142 53
rect 96 -19 142 19
rect 96 -53 102 -19
rect 136 -53 142 -19
rect 96 -91 142 -53
rect 96 -125 102 -91
rect 136 -125 142 -91
rect 96 -163 142 -125
rect 96 -197 102 -163
rect 136 -197 142 -163
rect 96 -235 142 -197
rect 96 -269 102 -235
rect 136 -269 142 -235
rect 96 -307 142 -269
rect 96 -341 102 -307
rect 136 -341 142 -307
rect 96 -379 142 -341
rect 96 -413 102 -379
rect 136 -413 142 -379
rect 96 -444 142 -413
rect -86 -491 86 -485
rect -86 -525 -53 -491
rect -19 -525 19 -491
rect 53 -525 86 -491
rect -86 -531 86 -525
<< end >>
