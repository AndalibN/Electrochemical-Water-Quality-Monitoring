magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -570 -202 2756 990
rect -54 -204 2756 -202
rect 606 -208 1874 -204
<< pwell >>
rect 2104 -266 2306 -264
rect -428 -286 -220 -272
rect -446 -364 -220 -286
rect -446 -1198 -234 -364
rect -8 -370 230 -284
rect 1036 -288 1516 -286
rect 12 -1198 122 -370
rect 464 -374 1896 -288
rect 524 -406 1896 -374
rect 2104 -380 2756 -266
rect 524 -1028 1848 -406
rect 524 -1198 646 -1028
rect 1126 -1198 1248 -1028
rect 1700 -1198 1848 -1028
rect 2128 -1198 2232 -380
rect 2460 -390 2756 -380
rect 2520 -1198 2698 -390
rect -446 -1396 2704 -1198
<< nmos >>
rect 794 -1002 854 -402
rect 912 -1002 972 -402
rect 1386 -1002 1446 -402
rect 1504 -1002 1564 -402
<< pmos >>
rect 678 58 738 658
rect 796 58 856 658
rect 914 58 974 658
rect 1032 58 1092 658
rect 1270 58 1330 658
rect 1388 58 1448 658
rect 1506 58 1566 658
rect 1624 58 1684 658
<< ndiff >>
rect 736 -447 794 -402
rect 736 -481 748 -447
rect 782 -481 794 -447
rect 736 -515 794 -481
rect 736 -549 748 -515
rect 782 -549 794 -515
rect 736 -583 794 -549
rect 736 -617 748 -583
rect 782 -617 794 -583
rect 736 -651 794 -617
rect 736 -685 748 -651
rect 782 -685 794 -651
rect 736 -719 794 -685
rect 736 -753 748 -719
rect 782 -753 794 -719
rect 736 -787 794 -753
rect 736 -821 748 -787
rect 782 -821 794 -787
rect 736 -855 794 -821
rect 736 -889 748 -855
rect 782 -889 794 -855
rect 736 -923 794 -889
rect 736 -957 748 -923
rect 782 -957 794 -923
rect 736 -1002 794 -957
rect 854 -447 912 -402
rect 854 -481 866 -447
rect 900 -481 912 -447
rect 854 -515 912 -481
rect 854 -549 866 -515
rect 900 -549 912 -515
rect 854 -583 912 -549
rect 854 -617 866 -583
rect 900 -617 912 -583
rect 854 -651 912 -617
rect 854 -685 866 -651
rect 900 -685 912 -651
rect 854 -719 912 -685
rect 854 -753 866 -719
rect 900 -753 912 -719
rect 854 -787 912 -753
rect 854 -821 866 -787
rect 900 -821 912 -787
rect 854 -855 912 -821
rect 854 -889 866 -855
rect 900 -889 912 -855
rect 854 -923 912 -889
rect 854 -957 866 -923
rect 900 -957 912 -923
rect 854 -1002 912 -957
rect 972 -447 1030 -402
rect 972 -481 984 -447
rect 1018 -481 1030 -447
rect 972 -515 1030 -481
rect 972 -549 984 -515
rect 1018 -549 1030 -515
rect 972 -583 1030 -549
rect 972 -617 984 -583
rect 1018 -617 1030 -583
rect 972 -651 1030 -617
rect 972 -685 984 -651
rect 1018 -685 1030 -651
rect 972 -719 1030 -685
rect 972 -753 984 -719
rect 1018 -753 1030 -719
rect 972 -787 1030 -753
rect 972 -821 984 -787
rect 1018 -821 1030 -787
rect 972 -855 1030 -821
rect 972 -889 984 -855
rect 1018 -889 1030 -855
rect 972 -923 1030 -889
rect 972 -957 984 -923
rect 1018 -957 1030 -923
rect 972 -1002 1030 -957
rect 1328 -447 1386 -402
rect 1328 -481 1340 -447
rect 1374 -481 1386 -447
rect 1328 -515 1386 -481
rect 1328 -549 1340 -515
rect 1374 -549 1386 -515
rect 1328 -583 1386 -549
rect 1328 -617 1340 -583
rect 1374 -617 1386 -583
rect 1328 -651 1386 -617
rect 1328 -685 1340 -651
rect 1374 -685 1386 -651
rect 1328 -719 1386 -685
rect 1328 -753 1340 -719
rect 1374 -753 1386 -719
rect 1328 -787 1386 -753
rect 1328 -821 1340 -787
rect 1374 -821 1386 -787
rect 1328 -855 1386 -821
rect 1328 -889 1340 -855
rect 1374 -889 1386 -855
rect 1328 -923 1386 -889
rect 1328 -957 1340 -923
rect 1374 -957 1386 -923
rect 1328 -1002 1386 -957
rect 1446 -447 1504 -402
rect 1446 -481 1458 -447
rect 1492 -481 1504 -447
rect 1446 -515 1504 -481
rect 1446 -549 1458 -515
rect 1492 -549 1504 -515
rect 1446 -583 1504 -549
rect 1446 -617 1458 -583
rect 1492 -617 1504 -583
rect 1446 -651 1504 -617
rect 1446 -685 1458 -651
rect 1492 -685 1504 -651
rect 1446 -719 1504 -685
rect 1446 -753 1458 -719
rect 1492 -753 1504 -719
rect 1446 -787 1504 -753
rect 1446 -821 1458 -787
rect 1492 -821 1504 -787
rect 1446 -855 1504 -821
rect 1446 -889 1458 -855
rect 1492 -889 1504 -855
rect 1446 -923 1504 -889
rect 1446 -957 1458 -923
rect 1492 -957 1504 -923
rect 1446 -1002 1504 -957
rect 1564 -447 1622 -402
rect 1564 -481 1576 -447
rect 1610 -481 1622 -447
rect 1564 -515 1622 -481
rect 1564 -549 1576 -515
rect 1610 -549 1622 -515
rect 1564 -583 1622 -549
rect 1564 -617 1576 -583
rect 1610 -617 1622 -583
rect 1564 -651 1622 -617
rect 1564 -685 1576 -651
rect 1610 -685 1622 -651
rect 1564 -719 1622 -685
rect 1564 -753 1576 -719
rect 1610 -753 1622 -719
rect 1564 -787 1622 -753
rect 1564 -821 1576 -787
rect 1610 -821 1622 -787
rect 1564 -855 1622 -821
rect 1564 -889 1576 -855
rect 1610 -889 1622 -855
rect 1564 -923 1622 -889
rect 1564 -957 1576 -923
rect 1610 -957 1622 -923
rect 1564 -1002 1622 -957
<< pdiff >>
rect 620 613 678 658
rect 620 579 632 613
rect 666 579 678 613
rect 620 545 678 579
rect 620 511 632 545
rect 666 511 678 545
rect 620 477 678 511
rect 620 443 632 477
rect 666 443 678 477
rect 620 409 678 443
rect 620 375 632 409
rect 666 375 678 409
rect 620 341 678 375
rect 620 307 632 341
rect 666 307 678 341
rect 620 273 678 307
rect 620 239 632 273
rect 666 239 678 273
rect 620 205 678 239
rect 620 171 632 205
rect 666 171 678 205
rect 620 137 678 171
rect 620 103 632 137
rect 666 103 678 137
rect 620 58 678 103
rect 738 613 796 658
rect 738 579 750 613
rect 784 579 796 613
rect 738 545 796 579
rect 738 511 750 545
rect 784 511 796 545
rect 738 477 796 511
rect 738 443 750 477
rect 784 443 796 477
rect 738 409 796 443
rect 738 375 750 409
rect 784 375 796 409
rect 738 341 796 375
rect 738 307 750 341
rect 784 307 796 341
rect 738 273 796 307
rect 738 239 750 273
rect 784 239 796 273
rect 738 205 796 239
rect 738 171 750 205
rect 784 171 796 205
rect 738 137 796 171
rect 738 103 750 137
rect 784 103 796 137
rect 738 58 796 103
rect 856 613 914 658
rect 856 579 868 613
rect 902 579 914 613
rect 856 545 914 579
rect 856 511 868 545
rect 902 511 914 545
rect 856 477 914 511
rect 856 443 868 477
rect 902 443 914 477
rect 856 409 914 443
rect 856 375 868 409
rect 902 375 914 409
rect 856 341 914 375
rect 856 307 868 341
rect 902 307 914 341
rect 856 273 914 307
rect 856 239 868 273
rect 902 239 914 273
rect 856 205 914 239
rect 856 171 868 205
rect 902 171 914 205
rect 856 137 914 171
rect 856 103 868 137
rect 902 103 914 137
rect 856 58 914 103
rect 974 613 1032 658
rect 974 579 986 613
rect 1020 579 1032 613
rect 974 545 1032 579
rect 974 511 986 545
rect 1020 511 1032 545
rect 974 477 1032 511
rect 974 443 986 477
rect 1020 443 1032 477
rect 974 409 1032 443
rect 974 375 986 409
rect 1020 375 1032 409
rect 974 341 1032 375
rect 974 307 986 341
rect 1020 307 1032 341
rect 974 273 1032 307
rect 974 239 986 273
rect 1020 239 1032 273
rect 974 205 1032 239
rect 974 171 986 205
rect 1020 171 1032 205
rect 974 137 1032 171
rect 974 103 986 137
rect 1020 103 1032 137
rect 974 58 1032 103
rect 1092 613 1150 658
rect 1092 579 1104 613
rect 1138 579 1150 613
rect 1092 545 1150 579
rect 1092 511 1104 545
rect 1138 511 1150 545
rect 1092 477 1150 511
rect 1092 443 1104 477
rect 1138 443 1150 477
rect 1092 409 1150 443
rect 1092 375 1104 409
rect 1138 375 1150 409
rect 1092 341 1150 375
rect 1092 307 1104 341
rect 1138 307 1150 341
rect 1092 273 1150 307
rect 1092 239 1104 273
rect 1138 239 1150 273
rect 1092 205 1150 239
rect 1092 171 1104 205
rect 1138 171 1150 205
rect 1092 137 1150 171
rect 1092 103 1104 137
rect 1138 103 1150 137
rect 1092 58 1150 103
rect 1212 613 1270 658
rect 1212 579 1224 613
rect 1258 579 1270 613
rect 1212 545 1270 579
rect 1212 511 1224 545
rect 1258 511 1270 545
rect 1212 477 1270 511
rect 1212 443 1224 477
rect 1258 443 1270 477
rect 1212 409 1270 443
rect 1212 375 1224 409
rect 1258 375 1270 409
rect 1212 341 1270 375
rect 1212 307 1224 341
rect 1258 307 1270 341
rect 1212 273 1270 307
rect 1212 239 1224 273
rect 1258 239 1270 273
rect 1212 205 1270 239
rect 1212 171 1224 205
rect 1258 171 1270 205
rect 1212 137 1270 171
rect 1212 103 1224 137
rect 1258 103 1270 137
rect 1212 58 1270 103
rect 1330 613 1388 658
rect 1330 579 1342 613
rect 1376 579 1388 613
rect 1330 545 1388 579
rect 1330 511 1342 545
rect 1376 511 1388 545
rect 1330 477 1388 511
rect 1330 443 1342 477
rect 1376 443 1388 477
rect 1330 409 1388 443
rect 1330 375 1342 409
rect 1376 375 1388 409
rect 1330 341 1388 375
rect 1330 307 1342 341
rect 1376 307 1388 341
rect 1330 273 1388 307
rect 1330 239 1342 273
rect 1376 239 1388 273
rect 1330 205 1388 239
rect 1330 171 1342 205
rect 1376 171 1388 205
rect 1330 137 1388 171
rect 1330 103 1342 137
rect 1376 103 1388 137
rect 1330 58 1388 103
rect 1448 613 1506 658
rect 1448 579 1460 613
rect 1494 579 1506 613
rect 1448 545 1506 579
rect 1448 511 1460 545
rect 1494 511 1506 545
rect 1448 477 1506 511
rect 1448 443 1460 477
rect 1494 443 1506 477
rect 1448 409 1506 443
rect 1448 375 1460 409
rect 1494 375 1506 409
rect 1448 341 1506 375
rect 1448 307 1460 341
rect 1494 307 1506 341
rect 1448 273 1506 307
rect 1448 239 1460 273
rect 1494 239 1506 273
rect 1448 205 1506 239
rect 1448 171 1460 205
rect 1494 171 1506 205
rect 1448 137 1506 171
rect 1448 103 1460 137
rect 1494 103 1506 137
rect 1448 58 1506 103
rect 1566 613 1624 658
rect 1566 579 1578 613
rect 1612 579 1624 613
rect 1566 545 1624 579
rect 1566 511 1578 545
rect 1612 511 1624 545
rect 1566 477 1624 511
rect 1566 443 1578 477
rect 1612 443 1624 477
rect 1566 409 1624 443
rect 1566 375 1578 409
rect 1612 375 1624 409
rect 1566 341 1624 375
rect 1566 307 1578 341
rect 1612 307 1624 341
rect 1566 273 1624 307
rect 1566 239 1578 273
rect 1612 239 1624 273
rect 1566 205 1624 239
rect 1566 171 1578 205
rect 1612 171 1624 205
rect 1566 137 1624 171
rect 1566 103 1578 137
rect 1612 103 1624 137
rect 1566 58 1624 103
rect 1684 613 1742 658
rect 1684 579 1696 613
rect 1730 579 1742 613
rect 1684 545 1742 579
rect 1684 511 1696 545
rect 1730 511 1742 545
rect 1684 477 1742 511
rect 1684 443 1696 477
rect 1730 443 1742 477
rect 1684 409 1742 443
rect 1684 375 1696 409
rect 1730 375 1742 409
rect 1684 341 1742 375
rect 1684 307 1696 341
rect 1730 307 1742 341
rect 1684 273 1742 307
rect 1684 239 1696 273
rect 1730 239 1742 273
rect 1684 205 1742 239
rect 1684 171 1696 205
rect 1730 171 1742 205
rect 1684 137 1742 171
rect 1684 103 1696 137
rect 1730 103 1742 137
rect 1684 58 1742 103
<< ndiffc >>
rect 748 -481 782 -447
rect 748 -549 782 -515
rect 748 -617 782 -583
rect 748 -685 782 -651
rect 748 -753 782 -719
rect 748 -821 782 -787
rect 748 -889 782 -855
rect 748 -957 782 -923
rect 866 -481 900 -447
rect 866 -549 900 -515
rect 866 -617 900 -583
rect 866 -685 900 -651
rect 866 -753 900 -719
rect 866 -821 900 -787
rect 866 -889 900 -855
rect 866 -957 900 -923
rect 984 -481 1018 -447
rect 984 -549 1018 -515
rect 984 -617 1018 -583
rect 984 -685 1018 -651
rect 984 -753 1018 -719
rect 984 -821 1018 -787
rect 984 -889 1018 -855
rect 984 -957 1018 -923
rect 1340 -481 1374 -447
rect 1340 -549 1374 -515
rect 1340 -617 1374 -583
rect 1340 -685 1374 -651
rect 1340 -753 1374 -719
rect 1340 -821 1374 -787
rect 1340 -889 1374 -855
rect 1340 -957 1374 -923
rect 1458 -481 1492 -447
rect 1458 -549 1492 -515
rect 1458 -617 1492 -583
rect 1458 -685 1492 -651
rect 1458 -753 1492 -719
rect 1458 -821 1492 -787
rect 1458 -889 1492 -855
rect 1458 -957 1492 -923
rect 1576 -481 1610 -447
rect 1576 -549 1610 -515
rect 1576 -617 1610 -583
rect 1576 -685 1610 -651
rect 1576 -753 1610 -719
rect 1576 -821 1610 -787
rect 1576 -889 1610 -855
rect 1576 -957 1610 -923
<< pdiffc >>
rect 632 579 666 613
rect 632 511 666 545
rect 632 443 666 477
rect 632 375 666 409
rect 632 307 666 341
rect 632 239 666 273
rect 632 171 666 205
rect 632 103 666 137
rect 750 579 784 613
rect 750 511 784 545
rect 750 443 784 477
rect 750 375 784 409
rect 750 307 784 341
rect 750 239 784 273
rect 750 171 784 205
rect 750 103 784 137
rect 868 579 902 613
rect 868 511 902 545
rect 868 443 902 477
rect 868 375 902 409
rect 868 307 902 341
rect 868 239 902 273
rect 868 171 902 205
rect 868 103 902 137
rect 986 579 1020 613
rect 986 511 1020 545
rect 986 443 1020 477
rect 986 375 1020 409
rect 986 307 1020 341
rect 986 239 1020 273
rect 986 171 1020 205
rect 986 103 1020 137
rect 1104 579 1138 613
rect 1104 511 1138 545
rect 1104 443 1138 477
rect 1104 375 1138 409
rect 1104 307 1138 341
rect 1104 239 1138 273
rect 1104 171 1138 205
rect 1104 103 1138 137
rect 1224 579 1258 613
rect 1224 511 1258 545
rect 1224 443 1258 477
rect 1224 375 1258 409
rect 1224 307 1258 341
rect 1224 239 1258 273
rect 1224 171 1258 205
rect 1224 103 1258 137
rect 1342 579 1376 613
rect 1342 511 1376 545
rect 1342 443 1376 477
rect 1342 375 1376 409
rect 1342 307 1376 341
rect 1342 239 1376 273
rect 1342 171 1376 205
rect 1342 103 1376 137
rect 1460 579 1494 613
rect 1460 511 1494 545
rect 1460 443 1494 477
rect 1460 375 1494 409
rect 1460 307 1494 341
rect 1460 239 1494 273
rect 1460 171 1494 205
rect 1460 103 1494 137
rect 1578 579 1612 613
rect 1578 511 1612 545
rect 1578 443 1612 477
rect 1578 375 1612 409
rect 1578 307 1612 341
rect 1578 239 1612 273
rect 1578 171 1612 205
rect 1578 103 1612 137
rect 1696 579 1730 613
rect 1696 511 1730 545
rect 1696 443 1730 477
rect 1696 375 1730 409
rect 1696 307 1730 341
rect 1696 239 1730 273
rect 1696 171 1730 205
rect 1696 103 1730 137
<< psubdiff >>
rect -402 -304 -246 -298
rect -402 -312 -319 -304
rect -420 -338 -319 -312
rect -285 -338 -246 -304
rect -420 -372 -260 -338
rect 18 -344 58 -310
rect 92 -344 126 -310
rect 160 -344 204 -310
rect -420 -1290 -387 -372
rect -285 -1224 -260 -372
rect 38 -398 96 -344
rect 490 -348 568 -314
rect 602 -348 661 -314
rect 695 -348 729 -314
rect 763 -348 797 -314
rect 831 -348 862 -314
rect 38 -432 50 -398
rect 84 -432 96 -398
rect 38 -466 96 -432
rect 38 -500 50 -466
rect 84 -500 96 -466
rect 38 -534 96 -500
rect 38 -568 50 -534
rect 84 -568 96 -534
rect 38 -602 96 -568
rect 38 -636 50 -602
rect 84 -636 96 -602
rect 38 -670 96 -636
rect 38 -704 50 -670
rect 84 -704 96 -670
rect 38 -738 96 -704
rect 38 -772 50 -738
rect 84 -772 96 -738
rect 38 -806 96 -772
rect 38 -840 50 -806
rect 84 -840 96 -806
rect 38 -874 96 -840
rect 38 -908 50 -874
rect 84 -908 96 -874
rect 38 -942 96 -908
rect 38 -976 50 -942
rect 84 -976 96 -942
rect 38 -1010 96 -976
rect 38 -1044 50 -1010
rect 84 -1044 96 -1010
rect 550 -382 620 -348
rect 1062 -346 1170 -312
rect 1204 -346 1276 -312
rect 1310 -346 1344 -312
rect 1378 -346 1412 -312
rect 1446 -346 1490 -312
rect 550 -416 568 -382
rect 602 -416 620 -382
rect 1152 -382 1222 -346
rect 1686 -330 1870 -314
rect 1686 -364 1757 -330
rect 1791 -364 1870 -330
rect 550 -450 620 -416
rect 550 -484 568 -450
rect 602 -484 620 -450
rect 550 -518 620 -484
rect 550 -552 568 -518
rect 602 -552 620 -518
rect 550 -586 620 -552
rect 550 -620 568 -586
rect 602 -620 620 -586
rect 550 -654 620 -620
rect 550 -688 568 -654
rect 602 -688 620 -654
rect 550 -722 620 -688
rect 550 -756 568 -722
rect 602 -756 620 -722
rect 550 -790 620 -756
rect 550 -824 568 -790
rect 602 -824 620 -790
rect 550 -858 620 -824
rect 550 -892 568 -858
rect 602 -892 620 -858
rect 550 -926 620 -892
rect 550 -960 568 -926
rect 602 -960 620 -926
rect 550 -994 620 -960
rect 38 -1088 96 -1044
rect 550 -1028 568 -994
rect 602 -1028 620 -994
rect 1152 -416 1170 -382
rect 1204 -416 1222 -382
rect 1686 -380 1870 -364
rect 2130 -305 2280 -290
rect 2130 -339 2163 -305
rect 2197 -339 2280 -305
rect 2130 -354 2280 -339
rect 1152 -450 1222 -416
rect 1152 -484 1170 -450
rect 1204 -484 1222 -450
rect 1152 -518 1222 -484
rect 1152 -552 1170 -518
rect 1204 -552 1222 -518
rect 1152 -586 1222 -552
rect 1152 -620 1170 -586
rect 1204 -620 1222 -586
rect 1152 -654 1222 -620
rect 1152 -688 1170 -654
rect 1204 -688 1222 -654
rect 1152 -722 1222 -688
rect 1152 -756 1170 -722
rect 1204 -756 1222 -722
rect 1152 -790 1222 -756
rect 1152 -824 1170 -790
rect 1204 -824 1222 -790
rect 1152 -858 1222 -824
rect 1152 -892 1170 -858
rect 1204 -892 1222 -858
rect 1152 -926 1222 -892
rect 1152 -960 1170 -926
rect 1204 -960 1222 -926
rect 1152 -994 1222 -960
rect 1152 -1028 1170 -994
rect 1204 -1028 1222 -994
rect 1726 -445 1822 -380
rect 1726 -479 1757 -445
rect 1791 -479 1822 -445
rect 1726 -513 1822 -479
rect 1726 -547 1757 -513
rect 1791 -547 1822 -513
rect 1726 -581 1822 -547
rect 1726 -615 1757 -581
rect 1791 -615 1822 -581
rect 1726 -649 1822 -615
rect 1726 -683 1757 -649
rect 1791 -683 1822 -649
rect 1726 -717 1822 -683
rect 1726 -751 1757 -717
rect 1791 -751 1822 -717
rect 1726 -785 1822 -751
rect 1726 -819 1757 -785
rect 1791 -819 1822 -785
rect 1726 -853 1822 -819
rect 1726 -887 1757 -853
rect 1791 -887 1822 -853
rect 1726 -921 1822 -887
rect 1726 -955 1757 -921
rect 1791 -955 1822 -921
rect 1726 -989 1822 -955
rect 1726 -1023 1757 -989
rect 1791 -1023 1822 -989
rect 550 -1052 620 -1028
rect 1152 -1054 1222 -1028
rect 1726 -1057 1822 -1023
rect 1726 -1091 1757 -1057
rect 1791 -1091 1822 -1057
rect 1726 -1125 1822 -1091
rect 1726 -1159 1757 -1125
rect 1791 -1159 1822 -1125
rect 1726 -1224 1822 -1159
rect 2154 -398 2206 -354
rect 2486 -304 2730 -292
rect 2486 -338 2605 -304
rect 2639 -338 2730 -304
rect 2486 -364 2730 -338
rect 2546 -372 2672 -364
rect 2154 -432 2163 -398
rect 2197 -432 2206 -398
rect 2154 -466 2206 -432
rect 2154 -500 2163 -466
rect 2197 -500 2206 -466
rect 2154 -534 2206 -500
rect 2154 -568 2163 -534
rect 2197 -568 2206 -534
rect 2154 -602 2206 -568
rect 2154 -636 2163 -602
rect 2197 -636 2206 -602
rect 2154 -670 2206 -636
rect 2154 -704 2163 -670
rect 2197 -704 2206 -670
rect 2154 -738 2206 -704
rect 2154 -772 2163 -738
rect 2197 -772 2206 -738
rect 2154 -806 2206 -772
rect 2154 -840 2163 -806
rect 2197 -840 2206 -806
rect 2154 -874 2206 -840
rect 2154 -908 2163 -874
rect 2197 -908 2206 -874
rect 2154 -942 2206 -908
rect 2154 -976 2163 -942
rect 2197 -976 2206 -942
rect 2154 -1010 2206 -976
rect 2154 -1044 2163 -1010
rect 2197 -1044 2206 -1010
rect 2154 -1078 2206 -1044
rect 2154 -1112 2163 -1078
rect 2197 -1112 2206 -1078
rect 2154 -1146 2206 -1112
rect 2154 -1180 2163 -1146
rect 2197 -1180 2206 -1146
rect 2154 -1224 2206 -1180
rect 2546 -406 2605 -372
rect 2639 -406 2672 -372
rect 2546 -440 2672 -406
rect 2546 -474 2605 -440
rect 2639 -474 2672 -440
rect 2546 -508 2672 -474
rect 2546 -542 2605 -508
rect 2639 -542 2672 -508
rect 2546 -576 2672 -542
rect 2546 -610 2605 -576
rect 2639 -610 2672 -576
rect 2546 -644 2672 -610
rect 2546 -678 2605 -644
rect 2639 -678 2672 -644
rect 2546 -712 2672 -678
rect 2546 -746 2605 -712
rect 2639 -746 2672 -712
rect 2546 -780 2672 -746
rect 2546 -814 2605 -780
rect 2639 -814 2672 -780
rect 2546 -848 2672 -814
rect 2546 -882 2605 -848
rect 2639 -882 2672 -848
rect 2546 -916 2672 -882
rect 2546 -950 2605 -916
rect 2639 -950 2672 -916
rect 2546 -984 2672 -950
rect 2546 -1018 2605 -984
rect 2639 -1018 2672 -984
rect 2546 -1052 2672 -1018
rect 2546 -1086 2605 -1052
rect 2639 -1086 2672 -1052
rect 2546 -1120 2672 -1086
rect 2546 -1154 2605 -1120
rect 2639 -1154 2672 -1120
rect 2546 -1188 2672 -1154
rect 2546 -1222 2605 -1188
rect 2639 -1222 2672 -1188
rect 2546 -1224 2672 -1222
rect -285 -1256 2678 -1224
rect -420 -1358 -319 -1290
rect 2639 -1358 2678 -1256
rect -420 -1370 2678 -1358
<< nsubdiff >>
rect -332 935 2584 952
rect -332 901 -243 935
rect -209 901 -175 935
rect -141 901 -107 935
rect -73 901 -39 935
rect -5 901 29 935
rect 63 901 97 935
rect 131 901 165 935
rect 199 901 233 935
rect 267 901 301 935
rect 335 901 369 935
rect 403 901 437 935
rect 471 901 505 935
rect 539 901 573 935
rect 607 901 641 935
rect 675 901 709 935
rect 743 901 777 935
rect 811 901 845 935
rect 879 901 913 935
rect 947 901 981 935
rect 1015 901 1049 935
rect 1083 901 1117 935
rect 1151 901 1185 935
rect 1219 901 1253 935
rect 1287 901 1321 935
rect 1355 901 1389 935
rect 1423 901 1457 935
rect 1491 901 1525 935
rect 1559 901 1593 935
rect 1627 901 1661 935
rect 1695 901 1729 935
rect 1763 901 1797 935
rect 1831 901 1865 935
rect 1899 901 1933 935
rect 1967 901 2001 935
rect 2035 901 2069 935
rect 2103 901 2137 935
rect 2171 901 2205 935
rect 2239 901 2273 935
rect 2307 901 2341 935
rect 2375 901 2409 935
rect 2443 901 2584 935
rect -332 860 2584 901
rect -332 823 -256 860
rect -332 789 -313 823
rect -279 789 -256 823
rect -332 755 -256 789
rect -332 721 -313 755
rect -279 721 -256 755
rect -332 687 -256 721
rect -332 653 -313 687
rect -279 653 -256 687
rect -332 619 -256 653
rect 2500 779 2584 860
rect 2500 745 2523 779
rect 2557 745 2584 779
rect 2500 711 2584 745
rect 2500 677 2523 711
rect 2557 677 2584 711
rect -332 585 -313 619
rect -279 585 -256 619
rect -332 551 -256 585
rect -332 517 -313 551
rect -279 517 -256 551
rect -332 483 -256 517
rect -332 449 -313 483
rect -279 449 -256 483
rect -332 415 -256 449
rect -332 381 -313 415
rect -279 381 -256 415
rect -332 347 -256 381
rect -332 313 -313 347
rect -279 313 -256 347
rect -332 279 -256 313
rect -332 245 -313 279
rect -279 245 -256 279
rect -332 211 -256 245
rect -332 177 -313 211
rect -279 177 -256 211
rect -332 143 -256 177
rect -332 109 -313 143
rect -279 109 -256 143
rect -332 75 -256 109
rect -332 41 -313 75
rect -279 41 -256 75
rect -332 -58 -256 41
rect 2500 643 2584 677
rect 2500 609 2523 643
rect 2557 609 2584 643
rect 2500 575 2584 609
rect 2500 541 2523 575
rect 2557 541 2584 575
rect 2500 507 2584 541
rect 2500 473 2523 507
rect 2557 473 2584 507
rect 2500 439 2584 473
rect 2500 405 2523 439
rect 2557 405 2584 439
rect 2500 371 2584 405
rect 2500 337 2523 371
rect 2557 337 2584 371
rect 2500 303 2584 337
rect 2500 269 2523 303
rect 2557 269 2584 303
rect 2500 235 2584 269
rect 2500 201 2523 235
rect 2557 201 2584 235
rect 2500 167 2584 201
rect 2500 133 2523 167
rect 2557 133 2584 167
rect 2500 99 2584 133
rect 2500 65 2523 99
rect 2557 65 2584 99
rect -332 -60 -74 -58
rect -332 -70 316 -60
rect -332 -104 -278 -70
rect -244 -104 -210 -70
rect -176 -104 -142 -70
rect -108 -71 316 -70
rect -108 -104 -33 -71
rect -332 -105 -33 -104
rect 1 -105 35 -71
rect 69 -105 103 -71
rect 137 -105 171 -71
rect 205 -105 239 -71
rect 273 -105 316 -71
rect -332 -122 316 -105
rect 486 -67 876 -56
rect 486 -101 527 -67
rect 561 -101 595 -67
rect 629 -101 663 -67
rect 697 -101 731 -67
rect 765 -101 799 -67
rect 833 -101 876 -67
rect 486 -118 876 -101
rect 1076 -69 1466 -58
rect 1076 -103 1117 -69
rect 1151 -103 1185 -69
rect 1219 -103 1253 -69
rect 1287 -103 1321 -69
rect 1355 -103 1389 -69
rect 1423 -103 1466 -69
rect 1076 -120 1466 -103
rect 2500 31 2584 65
rect 1640 -77 1964 -66
rect 1640 -111 1714 -77
rect 1748 -111 1782 -77
rect 1816 -111 1850 -77
rect 1884 -111 1964 -77
rect 1640 -124 1964 -111
rect 2096 -79 2322 -70
rect 2096 -113 2154 -79
rect 2188 -113 2222 -79
rect 2256 -113 2322 -79
rect 2096 -124 2322 -113
rect 2500 -3 2523 31
rect 2557 -3 2584 31
rect 2500 -134 2584 -3
<< psubdiffcont >>
rect -319 -338 -285 -304
rect 58 -344 92 -310
rect 126 -344 160 -310
rect -387 -1256 -285 -372
rect 568 -348 602 -314
rect 661 -348 695 -314
rect 729 -348 763 -314
rect 797 -348 831 -314
rect 50 -432 84 -398
rect 50 -500 84 -466
rect 50 -568 84 -534
rect 50 -636 84 -602
rect 50 -704 84 -670
rect 50 -772 84 -738
rect 50 -840 84 -806
rect 50 -908 84 -874
rect 50 -976 84 -942
rect 50 -1044 84 -1010
rect 1170 -346 1204 -312
rect 1276 -346 1310 -312
rect 1344 -346 1378 -312
rect 1412 -346 1446 -312
rect 568 -416 602 -382
rect 1757 -364 1791 -330
rect 568 -484 602 -450
rect 568 -552 602 -518
rect 568 -620 602 -586
rect 568 -688 602 -654
rect 568 -756 602 -722
rect 568 -824 602 -790
rect 568 -892 602 -858
rect 568 -960 602 -926
rect 568 -1028 602 -994
rect 1170 -416 1204 -382
rect 2163 -339 2197 -305
rect 1170 -484 1204 -450
rect 1170 -552 1204 -518
rect 1170 -620 1204 -586
rect 1170 -688 1204 -654
rect 1170 -756 1204 -722
rect 1170 -824 1204 -790
rect 1170 -892 1204 -858
rect 1170 -960 1204 -926
rect 1170 -1028 1204 -994
rect 1757 -479 1791 -445
rect 1757 -547 1791 -513
rect 1757 -615 1791 -581
rect 1757 -683 1791 -649
rect 1757 -751 1791 -717
rect 1757 -819 1791 -785
rect 1757 -887 1791 -853
rect 1757 -955 1791 -921
rect 1757 -1023 1791 -989
rect 1757 -1091 1791 -1057
rect 1757 -1159 1791 -1125
rect 2605 -338 2639 -304
rect 2163 -432 2197 -398
rect 2163 -500 2197 -466
rect 2163 -568 2197 -534
rect 2163 -636 2197 -602
rect 2163 -704 2197 -670
rect 2163 -772 2197 -738
rect 2163 -840 2197 -806
rect 2163 -908 2197 -874
rect 2163 -976 2197 -942
rect 2163 -1044 2197 -1010
rect 2163 -1112 2197 -1078
rect 2163 -1180 2197 -1146
rect 2605 -406 2639 -372
rect 2605 -474 2639 -440
rect 2605 -542 2639 -508
rect 2605 -610 2639 -576
rect 2605 -678 2639 -644
rect 2605 -746 2639 -712
rect 2605 -814 2639 -780
rect 2605 -882 2639 -848
rect 2605 -950 2639 -916
rect 2605 -1018 2639 -984
rect 2605 -1086 2639 -1052
rect 2605 -1154 2639 -1120
rect 2605 -1222 2639 -1188
rect -387 -1290 2639 -1256
rect -319 -1358 2639 -1290
<< nsubdiffcont >>
rect -243 901 -209 935
rect -175 901 -141 935
rect -107 901 -73 935
rect -39 901 -5 935
rect 29 901 63 935
rect 97 901 131 935
rect 165 901 199 935
rect 233 901 267 935
rect 301 901 335 935
rect 369 901 403 935
rect 437 901 471 935
rect 505 901 539 935
rect 573 901 607 935
rect 641 901 675 935
rect 709 901 743 935
rect 777 901 811 935
rect 845 901 879 935
rect 913 901 947 935
rect 981 901 1015 935
rect 1049 901 1083 935
rect 1117 901 1151 935
rect 1185 901 1219 935
rect 1253 901 1287 935
rect 1321 901 1355 935
rect 1389 901 1423 935
rect 1457 901 1491 935
rect 1525 901 1559 935
rect 1593 901 1627 935
rect 1661 901 1695 935
rect 1729 901 1763 935
rect 1797 901 1831 935
rect 1865 901 1899 935
rect 1933 901 1967 935
rect 2001 901 2035 935
rect 2069 901 2103 935
rect 2137 901 2171 935
rect 2205 901 2239 935
rect 2273 901 2307 935
rect 2341 901 2375 935
rect 2409 901 2443 935
rect -313 789 -279 823
rect -313 721 -279 755
rect -313 653 -279 687
rect 2523 745 2557 779
rect 2523 677 2557 711
rect -313 585 -279 619
rect -313 517 -279 551
rect -313 449 -279 483
rect -313 381 -279 415
rect -313 313 -279 347
rect -313 245 -279 279
rect -313 177 -279 211
rect -313 109 -279 143
rect -313 41 -279 75
rect 2523 609 2557 643
rect 2523 541 2557 575
rect 2523 473 2557 507
rect 2523 405 2557 439
rect 2523 337 2557 371
rect 2523 269 2557 303
rect 2523 201 2557 235
rect 2523 133 2557 167
rect 2523 65 2557 99
rect -278 -104 -244 -70
rect -210 -104 -176 -70
rect -142 -104 -108 -70
rect -33 -105 1 -71
rect 35 -105 69 -71
rect 103 -105 137 -71
rect 171 -105 205 -71
rect 239 -105 273 -71
rect 527 -101 561 -67
rect 595 -101 629 -67
rect 663 -101 697 -67
rect 731 -101 765 -67
rect 799 -101 833 -67
rect 1117 -103 1151 -69
rect 1185 -103 1219 -69
rect 1253 -103 1287 -69
rect 1321 -103 1355 -69
rect 1389 -103 1423 -69
rect 1714 -111 1748 -77
rect 1782 -111 1816 -77
rect 1850 -111 1884 -77
rect 2154 -113 2188 -79
rect 2222 -113 2256 -79
rect 2523 -3 2557 31
<< poly >>
rect 212 782 738 818
rect -130 708 154 744
rect -130 640 -84 708
rect 94 688 154 708
rect 212 686 272 782
rect 330 688 508 726
rect 678 658 738 782
rect 796 784 1330 818
rect 796 658 856 784
rect 914 684 1092 722
rect 914 658 974 684
rect 1032 658 1092 684
rect 1270 658 1330 784
rect 1868 790 2024 820
rect 1868 738 1902 790
rect 1986 736 2024 790
rect 2222 784 2378 814
rect 2222 736 2260 784
rect 2340 734 2378 784
rect 1506 684 1684 722
rect 1388 658 1448 684
rect 1506 658 1566 684
rect 1624 658 1684 684
rect -136 98 -76 140
rect -160 88 -76 98
rect -160 74 -78 88
rect -160 40 -137 74
rect -103 40 -78 74
rect -160 16 -78 40
rect 94 4 272 36
rect -638 -214 -506 -164
rect 214 -182 296 -160
rect 342 -182 376 50
rect 678 32 738 58
rect 796 32 856 58
rect 914 32 974 58
rect 1032 32 1092 58
rect 1270 32 1330 58
rect 1388 32 1448 58
rect 1506 32 1566 58
rect 1624 32 1684 58
rect 678 0 856 32
rect 214 -184 376 -182
rect -638 -215 -88 -214
rect -638 -249 -586 -215
rect -552 -232 -88 -215
rect 214 -218 237 -184
rect 271 -218 376 -184
rect 214 -222 376 -218
rect -552 -249 -86 -232
rect 214 -242 296 -222
rect -638 -258 -86 -249
rect -638 -298 -506 -258
rect -128 -368 -86 -258
rect 342 -374 376 -222
rect 626 -152 708 -146
rect 926 -152 960 32
rect 1270 0 1448 32
rect 1518 -148 1552 32
rect 626 -170 960 -152
rect 626 -204 649 -170
rect 683 -182 960 -170
rect 683 -204 708 -182
rect 626 -228 708 -204
rect -126 -1166 -88 -762
rect 926 -376 960 -182
rect 1236 -172 1552 -148
rect 1236 -206 1259 -172
rect 1293 -182 1552 -172
rect 1293 -206 1318 -182
rect 1236 -226 1318 -206
rect 794 -402 854 -376
rect 912 -402 972 -376
rect 1518 -376 1552 -182
rect 1754 -178 1836 -156
rect 1986 -178 2028 6
rect 1754 -180 2028 -178
rect 1754 -214 1777 -180
rect 1811 -210 2028 -180
rect 1811 -214 1836 -210
rect 1754 -238 1836 -214
rect 220 -1078 258 -1012
rect 1386 -402 1446 -376
rect 1504 -402 1564 -376
rect 1986 -380 2028 -210
rect 2170 -174 2252 -150
rect 2336 -174 2378 6
rect 2170 -208 2193 -174
rect 2227 -206 2378 -174
rect 2227 -208 2252 -206
rect 2170 -232 2252 -208
rect 794 -1028 854 -1002
rect 912 -1028 972 -1002
rect 1386 -1028 1446 -1002
rect 1504 -1028 1564 -1002
rect 806 -1078 840 -1028
rect 1400 -1078 1434 -1028
rect 220 -1110 1434 -1078
rect 220 -1166 254 -1110
rect -126 -1200 254 -1166
rect 2336 -384 2378 -206
<< polycont >>
rect -137 40 -103 74
rect -586 -249 -552 -215
rect 237 -218 271 -184
rect 649 -204 683 -170
rect 1259 -206 1293 -172
rect 1777 -214 1811 -180
rect 2193 -208 2227 -174
<< locali >>
rect -326 935 2578 948
rect -326 901 -243 935
rect -209 931 -175 935
rect -209 901 -182 931
rect -141 901 -107 935
rect -73 901 -39 935
rect -5 901 29 935
rect 63 901 97 935
rect 131 927 165 935
rect 131 901 163 927
rect 199 901 233 935
rect 267 901 301 935
rect 335 901 369 935
rect 403 901 437 935
rect 471 901 505 935
rect 539 901 573 935
rect 607 901 641 935
rect 675 901 709 935
rect 743 925 777 935
rect 743 901 747 925
rect 811 901 845 935
rect 879 901 913 935
rect 947 901 981 935
rect 1015 901 1049 935
rect 1083 901 1117 935
rect 1151 901 1185 935
rect 1219 901 1253 935
rect 1287 901 1321 935
rect 1355 925 1389 935
rect 1371 901 1389 925
rect 1423 901 1457 935
rect 1491 901 1525 935
rect 1559 901 1593 935
rect 1627 901 1661 935
rect 1695 901 1729 935
rect 1763 901 1797 935
rect 1831 901 1865 935
rect 1899 928 1933 935
rect 1899 901 1928 928
rect 1967 901 2001 935
rect 2035 901 2069 935
rect 2103 901 2137 935
rect 2171 901 2205 935
rect 2239 901 2273 935
rect 2307 934 2341 935
rect 2313 901 2341 934
rect 2375 901 2409 935
rect 2443 901 2578 935
rect -326 897 -182 901
rect -148 897 163 901
rect -326 893 163 897
rect 197 893 747 901
rect -326 891 747 893
rect 781 891 1337 901
rect 1371 894 1928 901
rect 1962 900 2279 901
rect 2313 900 2578 901
rect 1962 894 2578 900
rect 1371 891 2578 894
rect -326 874 2578 891
rect -326 823 -264 874
rect -326 789 -313 823
rect -279 789 -264 823
rect -326 755 -264 789
rect -326 721 -313 755
rect -279 721 -264 755
rect -326 687 -264 721
rect -326 653 -313 687
rect -279 653 -264 687
rect 2504 779 2578 874
rect 2504 745 2523 779
rect 2557 745 2578 779
rect 2504 711 2578 745
rect 2504 677 2523 711
rect 2557 677 2578 711
rect -326 619 -264 653
rect -326 585 -313 619
rect -279 585 -264 619
rect -326 551 -264 585
rect -326 517 -313 551
rect -279 517 -264 551
rect -326 483 -264 517
rect -326 449 -313 483
rect -279 449 -264 483
rect -326 415 -264 449
rect -326 381 -313 415
rect -279 381 -264 415
rect -326 347 -264 381
rect -326 313 -313 347
rect -279 313 -264 347
rect -326 279 -264 313
rect -326 245 -313 279
rect -279 245 -264 279
rect -326 211 -264 245
rect -326 177 -313 211
rect -279 177 -264 211
rect -326 143 -264 177
rect -326 109 -313 143
rect -279 109 -264 143
rect -326 75 -264 109
rect 632 627 666 662
rect 632 555 666 579
rect 632 483 666 511
rect 632 411 666 443
rect 632 341 666 375
rect 632 273 666 305
rect 632 205 666 233
rect 632 137 666 161
rect -326 41 -313 75
rect -279 41 -264 75
rect -326 -62 -264 41
rect -156 74 -82 94
rect -156 40 -138 74
rect -103 40 -82 74
rect 632 54 666 89
rect 750 627 784 662
rect 750 555 784 579
rect 750 483 784 511
rect 750 411 784 443
rect 750 341 784 375
rect 750 273 784 305
rect 750 205 784 233
rect 750 137 784 161
rect 750 54 784 89
rect 868 627 902 662
rect 868 555 902 579
rect 868 483 902 511
rect 868 411 902 443
rect 868 341 902 375
rect 868 273 902 305
rect 868 205 902 233
rect 868 137 902 161
rect 868 54 902 89
rect 986 627 1020 662
rect 986 555 1020 579
rect 986 483 1020 511
rect 986 411 1020 443
rect 986 341 1020 375
rect 986 273 1020 305
rect 986 205 1020 233
rect 986 137 1020 161
rect 986 54 1020 89
rect 1104 627 1138 662
rect 1104 555 1138 579
rect 1104 483 1138 511
rect 1104 411 1138 443
rect 1104 341 1138 375
rect 1104 273 1138 305
rect 1104 205 1138 233
rect 1104 137 1138 161
rect 1104 54 1138 89
rect 1224 627 1258 662
rect 1224 555 1258 579
rect 1224 483 1258 511
rect 1224 411 1258 443
rect 1224 341 1258 375
rect 1224 273 1258 305
rect 1224 205 1258 233
rect 1224 137 1258 161
rect 1224 54 1258 89
rect 1342 627 1376 662
rect 1342 555 1376 579
rect 1342 483 1376 511
rect 1342 411 1376 443
rect 1342 341 1376 375
rect 1342 273 1376 305
rect 1342 205 1376 233
rect 1342 137 1376 161
rect 1342 54 1376 89
rect 1460 627 1494 662
rect 1460 555 1494 579
rect 1460 483 1494 511
rect 1460 411 1494 443
rect 1460 341 1494 375
rect 1460 273 1494 305
rect 1460 205 1494 233
rect 1460 137 1494 161
rect 1460 54 1494 89
rect 1578 627 1612 662
rect 1578 555 1612 579
rect 1578 483 1612 511
rect 1578 411 1612 443
rect 1578 341 1612 375
rect 1578 273 1612 305
rect 1578 205 1612 233
rect 1578 137 1612 161
rect 1578 54 1612 89
rect 1696 627 1730 662
rect 1696 555 1730 579
rect 1696 483 1730 511
rect 1696 411 1730 443
rect 1696 341 1730 375
rect 1696 273 1730 305
rect 1696 205 1730 233
rect 1696 137 1730 161
rect 1696 54 1730 89
rect 2504 643 2578 677
rect 2504 609 2523 643
rect 2557 609 2578 643
rect 2504 575 2578 609
rect 2504 541 2523 575
rect 2557 541 2578 575
rect 2504 507 2578 541
rect 2504 473 2523 507
rect 2557 473 2578 507
rect 2504 439 2578 473
rect 2504 405 2523 439
rect 2557 405 2578 439
rect 2504 371 2578 405
rect 2504 337 2523 371
rect 2557 337 2578 371
rect 2504 303 2578 337
rect 2504 269 2523 303
rect 2557 269 2578 303
rect 2504 235 2578 269
rect 2504 201 2523 235
rect 2557 201 2578 235
rect 2504 167 2578 201
rect 2504 133 2523 167
rect 2557 133 2578 167
rect 2504 99 2578 133
rect 2504 65 2523 99
rect 2557 65 2578 99
rect -156 24 -82 40
rect 2504 31 2578 65
rect 2504 -3 2523 31
rect 2557 -3 2578 31
rect -326 -70 312 -62
rect -326 -104 -278 -70
rect -244 -104 -210 -70
rect -176 -104 -142 -70
rect -108 -71 312 -70
rect -108 -104 -33 -71
rect -326 -105 -33 -104
rect 1 -105 35 -71
rect 69 -105 103 -71
rect 137 -105 171 -71
rect 205 -105 239 -71
rect 273 -72 312 -71
rect -326 -106 268 -105
rect 302 -106 312 -72
rect -326 -116 312 -106
rect 488 -64 872 -58
rect 488 -98 500 -64
rect 534 -67 872 -64
rect 488 -101 527 -98
rect 561 -101 595 -67
rect 629 -101 663 -67
rect 697 -101 731 -67
rect 765 -101 799 -67
rect 833 -76 872 -67
rect 488 -110 827 -101
rect 861 -110 872 -76
rect 488 -114 872 -110
rect 1078 -68 1462 -60
rect 1078 -102 1091 -68
rect 1125 -69 1462 -68
rect 1078 -103 1117 -102
rect 1151 -103 1185 -69
rect 1219 -103 1253 -69
rect 1287 -103 1321 -69
rect 1355 -103 1389 -69
rect 1423 -74 1462 -69
rect 1662 -69 1700 -68
rect 1662 -72 1664 -69
rect 1078 -108 1414 -103
rect 1448 -108 1462 -74
rect 1078 -116 1462 -108
rect 1646 -103 1664 -72
rect 1698 -72 1700 -69
rect 2258 -70 2300 -66
rect 1698 -77 1958 -72
rect 2126 -74 2166 -70
rect 2258 -74 2262 -70
rect 1698 -103 1714 -77
rect 1646 -111 1714 -103
rect 1748 -111 1782 -77
rect 1816 -111 1850 -77
rect 1884 -96 1958 -77
rect 1884 -111 1891 -96
rect 1646 -116 1891 -111
rect -68 -118 312 -116
rect 1888 -130 1891 -116
rect 1925 -116 1958 -96
rect 2100 -108 2129 -74
rect 2163 -79 2262 -74
rect 2100 -113 2154 -108
rect 2188 -113 2222 -79
rect 2256 -104 2262 -79
rect 2296 -74 2300 -70
rect 2296 -104 2318 -74
rect 2256 -113 2318 -104
rect 1925 -130 1928 -116
rect 2100 -120 2318 -113
rect 2504 -130 2578 -3
rect -636 -212 -510 -168
rect -636 -246 -587 -212
rect -553 -215 -510 -212
rect -636 -249 -586 -246
rect -552 -249 -510 -215
rect 218 -184 292 -164
rect 218 -218 236 -184
rect 271 -218 292 -184
rect 218 -234 292 -218
rect 630 -170 704 -150
rect 630 -204 648 -170
rect 683 -204 704 -170
rect 630 -220 704 -204
rect 1240 -172 1314 -152
rect 1240 -206 1258 -172
rect 1293 -206 1314 -172
rect 1240 -222 1314 -206
rect 1758 -180 1832 -160
rect 1758 -214 1776 -180
rect 1811 -214 1832 -180
rect 1758 -230 1832 -214
rect 2174 -174 2248 -154
rect 2174 -208 2192 -174
rect 2227 -208 2248 -174
rect 2174 -224 2248 -208
rect -636 -294 -510 -249
rect -394 -304 -254 -298
rect -394 -320 -319 -304
rect -420 -338 -319 -320
rect -285 -338 -254 -304
rect 2138 -305 2272 -290
rect -420 -348 -260 -338
rect 26 -344 58 -310
rect 92 -344 126 -310
rect 160 -344 196 -310
rect -420 -372 -346 -348
rect -312 -372 -260 -348
rect -420 -1290 -387 -372
rect -285 -1224 -260 -372
rect 38 -357 96 -344
rect 498 -348 568 -314
rect 602 -348 661 -314
rect 695 -348 729 -314
rect 763 -348 797 -314
rect 831 -348 854 -314
rect 1070 -346 1170 -312
rect 1204 -346 1276 -312
rect 1310 -346 1344 -312
rect 1378 -346 1412 -312
rect 1446 -346 1482 -312
rect 1694 -330 1862 -314
rect 38 -391 50 -357
rect 84 -391 96 -357
rect 38 -398 96 -391
rect 38 -432 50 -398
rect 84 -432 96 -398
rect 38 -466 96 -432
rect 38 -500 50 -466
rect 84 -500 96 -466
rect 38 -534 96 -500
rect 38 -568 50 -534
rect 84 -568 96 -534
rect 38 -602 96 -568
rect 38 -636 50 -602
rect 84 -636 96 -602
rect 38 -670 96 -636
rect 38 -704 50 -670
rect 84 -704 96 -670
rect 38 -738 96 -704
rect 38 -772 50 -738
rect 84 -772 96 -738
rect 38 -806 96 -772
rect 38 -840 50 -806
rect 84 -840 96 -806
rect 38 -874 96 -840
rect 38 -908 50 -874
rect 84 -908 96 -874
rect 38 -942 96 -908
rect 38 -976 50 -942
rect 84 -976 96 -942
rect 38 -1010 96 -976
rect 38 -1044 50 -1010
rect 84 -1017 96 -1010
rect 38 -1051 52 -1044
rect 86 -1051 96 -1017
rect 550 -364 620 -348
rect 550 -398 565 -364
rect 599 -382 620 -364
rect 550 -416 568 -398
rect 602 -416 620 -382
rect 1152 -365 1222 -346
rect 1152 -382 1172 -365
rect 550 -450 620 -416
rect 550 -484 568 -450
rect 602 -484 620 -450
rect 550 -518 620 -484
rect 550 -552 568 -518
rect 602 -552 620 -518
rect 550 -586 620 -552
rect 550 -620 568 -586
rect 602 -620 620 -586
rect 550 -654 620 -620
rect 550 -688 568 -654
rect 602 -688 620 -654
rect 550 -722 620 -688
rect 550 -756 568 -722
rect 602 -756 620 -722
rect 550 -790 620 -756
rect 550 -824 568 -790
rect 602 -824 620 -790
rect 550 -858 620 -824
rect 550 -892 568 -858
rect 602 -892 620 -858
rect 550 -926 620 -892
rect 550 -960 568 -926
rect 602 -960 620 -926
rect 550 -974 620 -960
rect 550 -1028 568 -974
rect 602 -1028 620 -974
rect 748 -433 782 -398
rect 748 -505 782 -481
rect 748 -577 782 -549
rect 748 -649 782 -617
rect 748 -719 782 -685
rect 748 -787 782 -755
rect 748 -855 782 -827
rect 748 -923 782 -899
rect 748 -1006 782 -971
rect 866 -433 900 -398
rect 866 -505 900 -481
rect 866 -577 900 -549
rect 866 -649 900 -617
rect 866 -719 900 -685
rect 866 -787 900 -755
rect 866 -855 900 -827
rect 866 -923 900 -899
rect 866 -1006 900 -971
rect 984 -433 1018 -398
rect 984 -505 1018 -481
rect 984 -577 1018 -549
rect 984 -649 1018 -617
rect 984 -719 1018 -685
rect 984 -787 1018 -755
rect 984 -855 1018 -827
rect 984 -923 1018 -899
rect 984 -1006 1018 -971
rect 1152 -416 1170 -382
rect 1206 -399 1222 -365
rect 1694 -364 1757 -330
rect 1791 -364 1862 -330
rect 2138 -339 2163 -305
rect 2197 -306 2272 -305
rect 2197 -339 2230 -306
rect 2138 -340 2230 -339
rect 2264 -340 2272 -306
rect 2138 -354 2272 -340
rect 2494 -304 2722 -292
rect 2494 -309 2605 -304
rect 2494 -343 2509 -309
rect 2543 -338 2605 -309
rect 2639 -338 2722 -304
rect 2543 -343 2722 -338
rect 1694 -368 1862 -364
rect 1694 -380 1764 -368
rect 1204 -416 1222 -399
rect 1152 -450 1222 -416
rect 1152 -484 1170 -450
rect 1204 -484 1222 -450
rect 1152 -518 1222 -484
rect 1152 -552 1170 -518
rect 1204 -552 1222 -518
rect 1152 -586 1222 -552
rect 1152 -620 1170 -586
rect 1204 -620 1222 -586
rect 1152 -654 1222 -620
rect 1152 -688 1170 -654
rect 1204 -688 1222 -654
rect 1152 -722 1222 -688
rect 1152 -756 1170 -722
rect 1204 -756 1222 -722
rect 1152 -790 1222 -756
rect 1152 -824 1170 -790
rect 1204 -824 1222 -790
rect 1152 -858 1222 -824
rect 1152 -892 1170 -858
rect 1204 -892 1222 -858
rect 1152 -926 1222 -892
rect 1152 -960 1170 -926
rect 1204 -960 1222 -926
rect 1152 -976 1222 -960
rect 550 -1044 620 -1028
rect 1152 -1010 1169 -976
rect 1203 -994 1222 -976
rect 1152 -1028 1170 -1010
rect 1204 -1028 1222 -994
rect 1340 -433 1374 -398
rect 1340 -505 1374 -481
rect 1340 -577 1374 -549
rect 1340 -649 1374 -617
rect 1340 -719 1374 -685
rect 1340 -787 1374 -755
rect 1340 -855 1374 -827
rect 1340 -923 1374 -899
rect 1340 -1006 1374 -971
rect 1458 -433 1492 -398
rect 1458 -505 1492 -481
rect 1458 -577 1492 -549
rect 1458 -649 1492 -617
rect 1458 -719 1492 -685
rect 1458 -787 1492 -755
rect 1458 -855 1492 -827
rect 1458 -923 1492 -899
rect 1458 -1006 1492 -971
rect 1576 -433 1610 -398
rect 1576 -505 1610 -481
rect 1576 -577 1610 -549
rect 1576 -649 1610 -617
rect 1576 -719 1610 -685
rect 1576 -787 1610 -755
rect 1576 -855 1610 -827
rect 1576 -923 1610 -899
rect 1576 -1006 1610 -971
rect 1726 -402 1764 -380
rect 1798 -380 1862 -368
rect 1798 -402 1822 -380
rect 1726 -445 1822 -402
rect 1726 -479 1757 -445
rect 1791 -479 1822 -445
rect 1726 -513 1822 -479
rect 1726 -547 1757 -513
rect 1791 -547 1822 -513
rect 1726 -581 1822 -547
rect 1726 -615 1757 -581
rect 1791 -615 1822 -581
rect 1726 -649 1822 -615
rect 1726 -683 1757 -649
rect 1791 -683 1822 -649
rect 1726 -717 1822 -683
rect 1726 -751 1757 -717
rect 1791 -751 1822 -717
rect 1726 -785 1822 -751
rect 1726 -819 1757 -785
rect 1791 -819 1822 -785
rect 1726 -853 1822 -819
rect 1726 -887 1757 -853
rect 1791 -887 1822 -853
rect 1726 -921 1822 -887
rect 1726 -955 1757 -921
rect 1791 -955 1822 -921
rect 1726 -989 1822 -955
rect 1152 -1046 1222 -1028
rect 1726 -1023 1757 -989
rect 1791 -1023 1822 -989
rect 38 -1080 96 -1051
rect 1726 -1057 1822 -1023
rect 1726 -1091 1757 -1057
rect 1791 -1091 1822 -1057
rect 1726 -1125 1822 -1091
rect 1726 -1159 1757 -1125
rect 1791 -1159 1822 -1125
rect 1726 -1224 1822 -1159
rect 2154 -398 2206 -354
rect 2494 -364 2722 -343
rect 2154 -432 2163 -398
rect 2197 -432 2206 -398
rect 2154 -466 2206 -432
rect 2154 -500 2163 -466
rect 2197 -500 2206 -466
rect 2154 -534 2206 -500
rect 2154 -568 2163 -534
rect 2197 -568 2206 -534
rect 2154 -602 2206 -568
rect 2154 -636 2163 -602
rect 2197 -636 2206 -602
rect 2154 -670 2206 -636
rect 2154 -704 2163 -670
rect 2197 -704 2206 -670
rect 2154 -738 2206 -704
rect 2154 -772 2163 -738
rect 2197 -772 2206 -738
rect 2154 -806 2206 -772
rect 2154 -840 2163 -806
rect 2197 -840 2206 -806
rect 2154 -874 2206 -840
rect 2154 -908 2163 -874
rect 2197 -908 2206 -874
rect 2154 -942 2206 -908
rect 2154 -976 2163 -942
rect 2197 -976 2206 -942
rect 2154 -1010 2206 -976
rect 2154 -1044 2163 -1010
rect 2197 -1044 2206 -1010
rect 2154 -1078 2206 -1044
rect 2154 -1112 2163 -1078
rect 2197 -1112 2206 -1078
rect 2154 -1146 2206 -1112
rect 2154 -1180 2163 -1146
rect 2197 -1180 2206 -1146
rect 2154 -1224 2206 -1180
rect 2546 -372 2672 -364
rect 2546 -406 2605 -372
rect 2639 -406 2672 -372
rect 2546 -440 2672 -406
rect 2546 -474 2605 -440
rect 2639 -474 2672 -440
rect 2546 -508 2672 -474
rect 2546 -542 2605 -508
rect 2639 -542 2672 -508
rect 2546 -576 2672 -542
rect 2546 -610 2605 -576
rect 2639 -610 2672 -576
rect 2546 -644 2672 -610
rect 2546 -678 2605 -644
rect 2639 -678 2672 -644
rect 2546 -712 2672 -678
rect 2546 -746 2605 -712
rect 2639 -746 2672 -712
rect 2546 -780 2672 -746
rect 2546 -814 2605 -780
rect 2639 -814 2672 -780
rect 2546 -848 2672 -814
rect 2546 -882 2605 -848
rect 2639 -882 2672 -848
rect 2546 -916 2672 -882
rect 2546 -950 2605 -916
rect 2639 -950 2672 -916
rect 2546 -984 2672 -950
rect 2546 -1018 2605 -984
rect 2639 -1018 2672 -984
rect 2546 -1052 2672 -1018
rect 2546 -1086 2605 -1052
rect 2639 -1086 2672 -1052
rect 2546 -1120 2672 -1086
rect 2546 -1154 2605 -1120
rect 2639 -1154 2672 -1120
rect 2546 -1188 2672 -1154
rect 2546 -1222 2605 -1188
rect 2639 -1222 2672 -1188
rect 2546 -1224 2672 -1222
rect -285 -1237 2672 -1224
rect -285 -1255 53 -1237
rect -285 -1256 -181 -1255
rect -147 -1256 53 -1255
rect 87 -1256 2672 -1237
rect -420 -1358 -319 -1290
rect 2639 -1358 2670 -1256
rect -420 -1362 2670 -1358
rect -386 -1370 2670 -1362
<< viali >>
rect -182 901 -175 931
rect -175 901 -148 931
rect 163 901 165 927
rect 165 901 197 927
rect 747 901 777 925
rect 777 901 781 925
rect 1337 901 1355 925
rect 1355 901 1371 925
rect 1928 901 1933 928
rect 1933 901 1962 928
rect 2279 901 2307 934
rect 2307 901 2313 934
rect -182 897 -148 901
rect 163 893 197 901
rect 747 891 781 901
rect 1337 891 1371 901
rect 1928 894 1962 901
rect 2279 900 2313 901
rect 632 613 666 627
rect 632 593 666 613
rect 632 545 666 555
rect 632 521 666 545
rect 632 477 666 483
rect 632 449 666 477
rect 632 409 666 411
rect 632 377 666 409
rect 632 307 666 339
rect 632 305 666 307
rect 632 239 666 267
rect 632 233 666 239
rect 632 171 666 195
rect 632 161 666 171
rect 632 103 666 123
rect -138 40 -137 74
rect -137 40 -104 74
rect 632 89 666 103
rect 750 613 784 627
rect 750 593 784 613
rect 750 545 784 555
rect 750 521 784 545
rect 750 477 784 483
rect 750 449 784 477
rect 750 409 784 411
rect 750 377 784 409
rect 750 307 784 339
rect 750 305 784 307
rect 750 239 784 267
rect 750 233 784 239
rect 750 171 784 195
rect 750 161 784 171
rect 750 103 784 123
rect 750 89 784 103
rect 868 613 902 627
rect 868 593 902 613
rect 868 545 902 555
rect 868 521 902 545
rect 868 477 902 483
rect 868 449 902 477
rect 868 409 902 411
rect 868 377 902 409
rect 868 307 902 339
rect 868 305 902 307
rect 868 239 902 267
rect 868 233 902 239
rect 868 171 902 195
rect 868 161 902 171
rect 868 103 902 123
rect 868 89 902 103
rect 986 613 1020 627
rect 986 593 1020 613
rect 986 545 1020 555
rect 986 521 1020 545
rect 986 477 1020 483
rect 986 449 1020 477
rect 986 409 1020 411
rect 986 377 1020 409
rect 986 307 1020 339
rect 986 305 1020 307
rect 986 239 1020 267
rect 986 233 1020 239
rect 986 171 1020 195
rect 986 161 1020 171
rect 986 103 1020 123
rect 986 89 1020 103
rect 1104 613 1138 627
rect 1104 593 1138 613
rect 1104 545 1138 555
rect 1104 521 1138 545
rect 1104 477 1138 483
rect 1104 449 1138 477
rect 1104 409 1138 411
rect 1104 377 1138 409
rect 1104 307 1138 339
rect 1104 305 1138 307
rect 1104 239 1138 267
rect 1104 233 1138 239
rect 1104 171 1138 195
rect 1104 161 1138 171
rect 1104 103 1138 123
rect 1104 89 1138 103
rect 1224 613 1258 627
rect 1224 593 1258 613
rect 1224 545 1258 555
rect 1224 521 1258 545
rect 1224 477 1258 483
rect 1224 449 1258 477
rect 1224 409 1258 411
rect 1224 377 1258 409
rect 1224 307 1258 339
rect 1224 305 1258 307
rect 1224 239 1258 267
rect 1224 233 1258 239
rect 1224 171 1258 195
rect 1224 161 1258 171
rect 1224 103 1258 123
rect 1224 89 1258 103
rect 1342 613 1376 627
rect 1342 593 1376 613
rect 1342 545 1376 555
rect 1342 521 1376 545
rect 1342 477 1376 483
rect 1342 449 1376 477
rect 1342 409 1376 411
rect 1342 377 1376 409
rect 1342 307 1376 339
rect 1342 305 1376 307
rect 1342 239 1376 267
rect 1342 233 1376 239
rect 1342 171 1376 195
rect 1342 161 1376 171
rect 1342 103 1376 123
rect 1342 89 1376 103
rect 1460 613 1494 627
rect 1460 593 1494 613
rect 1460 545 1494 555
rect 1460 521 1494 545
rect 1460 477 1494 483
rect 1460 449 1494 477
rect 1460 409 1494 411
rect 1460 377 1494 409
rect 1460 307 1494 339
rect 1460 305 1494 307
rect 1460 239 1494 267
rect 1460 233 1494 239
rect 1460 171 1494 195
rect 1460 161 1494 171
rect 1460 103 1494 123
rect 1460 89 1494 103
rect 1578 613 1612 627
rect 1578 593 1612 613
rect 1578 545 1612 555
rect 1578 521 1612 545
rect 1578 477 1612 483
rect 1578 449 1612 477
rect 1578 409 1612 411
rect 1578 377 1612 409
rect 1578 307 1612 339
rect 1578 305 1612 307
rect 1578 239 1612 267
rect 1578 233 1612 239
rect 1578 171 1612 195
rect 1578 161 1612 171
rect 1578 103 1612 123
rect 1578 89 1612 103
rect 1696 613 1730 627
rect 1696 593 1730 613
rect 1696 545 1730 555
rect 1696 521 1730 545
rect 1696 477 1730 483
rect 1696 449 1730 477
rect 1696 409 1730 411
rect 1696 377 1730 409
rect 1696 307 1730 339
rect 1696 305 1730 307
rect 1696 239 1730 267
rect 1696 233 1730 239
rect 1696 171 1730 195
rect 1696 161 1730 171
rect 1696 103 1730 123
rect 1696 89 1730 103
rect 268 -105 273 -72
rect 273 -105 302 -72
rect 268 -106 302 -105
rect 500 -67 534 -64
rect 500 -98 527 -67
rect 527 -98 534 -67
rect 827 -101 833 -76
rect 833 -101 861 -76
rect 827 -110 861 -101
rect 1091 -69 1125 -68
rect 1091 -102 1117 -69
rect 1117 -102 1125 -69
rect 1414 -103 1423 -74
rect 1423 -103 1448 -74
rect 1414 -108 1448 -103
rect 1664 -103 1698 -69
rect 1891 -130 1925 -96
rect 2129 -79 2163 -74
rect 2129 -108 2154 -79
rect 2154 -108 2163 -79
rect 2262 -104 2296 -70
rect -587 -215 -553 -212
rect -587 -246 -586 -215
rect -586 -246 -553 -215
rect 236 -218 237 -184
rect 237 -218 270 -184
rect 648 -204 649 -170
rect 649 -204 682 -170
rect 1258 -206 1259 -172
rect 1259 -206 1292 -172
rect 1776 -214 1777 -180
rect 1777 -214 1810 -180
rect 2192 -208 2193 -174
rect 2193 -208 2226 -174
rect -346 -372 -312 -348
rect -346 -382 -312 -372
rect 50 -391 84 -357
rect 52 -1044 84 -1017
rect 84 -1044 86 -1017
rect 52 -1051 86 -1044
rect 565 -382 599 -364
rect 565 -398 568 -382
rect 568 -398 599 -382
rect 1172 -382 1206 -365
rect 568 -994 602 -974
rect 568 -1008 602 -994
rect 748 -447 782 -433
rect 748 -467 782 -447
rect 748 -515 782 -505
rect 748 -539 782 -515
rect 748 -583 782 -577
rect 748 -611 782 -583
rect 748 -651 782 -649
rect 748 -683 782 -651
rect 748 -753 782 -721
rect 748 -755 782 -753
rect 748 -821 782 -793
rect 748 -827 782 -821
rect 748 -889 782 -865
rect 748 -899 782 -889
rect 748 -957 782 -937
rect 748 -971 782 -957
rect 866 -447 900 -433
rect 866 -467 900 -447
rect 866 -515 900 -505
rect 866 -539 900 -515
rect 866 -583 900 -577
rect 866 -611 900 -583
rect 866 -651 900 -649
rect 866 -683 900 -651
rect 866 -753 900 -721
rect 866 -755 900 -753
rect 866 -821 900 -793
rect 866 -827 900 -821
rect 866 -889 900 -865
rect 866 -899 900 -889
rect 866 -957 900 -937
rect 866 -971 900 -957
rect 984 -447 1018 -433
rect 984 -467 1018 -447
rect 984 -515 1018 -505
rect 984 -539 1018 -515
rect 984 -583 1018 -577
rect 984 -611 1018 -583
rect 984 -651 1018 -649
rect 984 -683 1018 -651
rect 984 -753 1018 -721
rect 984 -755 1018 -753
rect 984 -821 1018 -793
rect 984 -827 1018 -821
rect 984 -889 1018 -865
rect 984 -899 1018 -889
rect 984 -957 1018 -937
rect 984 -971 1018 -957
rect 1172 -399 1204 -382
rect 1204 -399 1206 -382
rect 2230 -340 2264 -306
rect 2509 -343 2543 -309
rect 1169 -994 1203 -976
rect 1169 -1010 1170 -994
rect 1170 -1010 1203 -994
rect 1340 -447 1374 -433
rect 1340 -467 1374 -447
rect 1340 -515 1374 -505
rect 1340 -539 1374 -515
rect 1340 -583 1374 -577
rect 1340 -611 1374 -583
rect 1340 -651 1374 -649
rect 1340 -683 1374 -651
rect 1340 -753 1374 -721
rect 1340 -755 1374 -753
rect 1340 -821 1374 -793
rect 1340 -827 1374 -821
rect 1340 -889 1374 -865
rect 1340 -899 1374 -889
rect 1340 -957 1374 -937
rect 1340 -971 1374 -957
rect 1458 -447 1492 -433
rect 1458 -467 1492 -447
rect 1458 -515 1492 -505
rect 1458 -539 1492 -515
rect 1458 -583 1492 -577
rect 1458 -611 1492 -583
rect 1458 -651 1492 -649
rect 1458 -683 1492 -651
rect 1458 -753 1492 -721
rect 1458 -755 1492 -753
rect 1458 -821 1492 -793
rect 1458 -827 1492 -821
rect 1458 -889 1492 -865
rect 1458 -899 1492 -889
rect 1458 -957 1492 -937
rect 1458 -971 1492 -957
rect 1576 -447 1610 -433
rect 1576 -467 1610 -447
rect 1576 -515 1610 -505
rect 1576 -539 1610 -515
rect 1576 -583 1610 -577
rect 1576 -611 1610 -583
rect 1576 -651 1610 -649
rect 1576 -683 1610 -651
rect 1576 -753 1610 -721
rect 1576 -755 1610 -753
rect 1576 -821 1610 -793
rect 1576 -827 1610 -821
rect 1576 -889 1610 -865
rect 1576 -899 1610 -889
rect 1576 -957 1610 -937
rect 1576 -971 1610 -957
rect 1764 -402 1798 -368
rect -181 -1256 -147 -1255
rect 53 -1256 87 -1237
rect -181 -1289 -147 -1256
rect 53 -1271 87 -1256
rect 166 -1296 200 -1262
rect 563 -1293 597 -1259
rect 749 -1295 783 -1261
rect 1170 -1301 1204 -1267
rect 1336 -1296 1370 -1262
rect 1928 -1294 1962 -1260
rect 2278 -1297 2312 -1263
<< metal1 >>
rect -194 931 -136 946
rect -194 897 -182 931
rect -148 897 -136 931
rect -194 886 -136 897
rect 146 927 214 944
rect 146 893 163 927
rect 197 893 214 927
rect -178 620 -150 886
rect 146 882 214 893
rect 728 925 802 942
rect 728 891 747 925
rect 781 891 802 925
rect 150 880 212 882
rect 168 656 196 880
rect 728 878 802 891
rect 1318 940 1386 944
rect 1318 925 1390 940
rect 1318 891 1337 925
rect 1371 891 1390 925
rect 1318 878 1390 891
rect 1908 928 1980 946
rect 1908 894 1928 928
rect 1962 894 1980 928
rect 1908 882 1980 894
rect 2266 934 2330 940
rect 2266 900 2279 934
rect 2313 900 2330 934
rect 2266 888 2330 900
rect 1910 878 1980 882
rect 286 736 552 768
rect 286 660 318 736
rect 520 658 552 736
rect 750 658 784 878
rect 1318 876 1386 878
rect 870 732 1136 764
rect 870 658 902 732
rect 1104 658 1136 732
rect 1342 658 1374 876
rect 1462 732 1728 764
rect 1462 658 1494 732
rect 1696 658 1728 732
rect 1926 712 1966 878
rect 2110 810 2196 822
rect 2110 758 2127 810
rect 2179 758 2196 810
rect 2110 748 2196 758
rect 2166 700 2196 748
rect 2284 714 2314 888
rect 2404 812 2486 826
rect 2404 760 2413 812
rect 2465 760 2486 812
rect 2404 748 2486 760
rect 2404 698 2432 748
rect 626 627 672 658
rect 626 593 632 627
rect 666 593 672 627
rect 626 555 672 593
rect 626 521 632 555
rect 666 521 672 555
rect 626 483 672 521
rect 626 449 632 483
rect 666 449 672 483
rect 626 411 672 449
rect 626 377 632 411
rect 666 377 672 411
rect 626 339 672 377
rect 626 305 632 339
rect 666 305 672 339
rect 626 267 672 305
rect 626 233 632 267
rect 666 233 672 267
rect 626 195 672 233
rect 626 161 632 195
rect 666 161 672 195
rect -158 74 -80 98
rect -158 40 -138 74
rect -104 68 -80 74
rect -52 68 -22 148
rect 626 123 672 161
rect 626 89 632 123
rect 666 89 672 123
rect 404 78 408 80
rect 404 74 432 78
rect -104 40 -22 68
rect -158 36 -22 40
rect -158 18 -80 36
rect -808 -214 -700 -178
rect -628 -212 -512 -170
rect -628 -214 -587 -212
rect -808 -246 -587 -214
rect -553 -246 -512 -212
rect -808 -264 -512 -246
rect -808 -298 -700 -264
rect -628 -290 -512 -264
rect -362 -340 -290 -334
rect -362 -392 -354 -340
rect -302 -392 -290 -340
rect -362 -400 -290 -392
rect -52 -394 -22 36
rect 50 -4 80 70
rect 290 -4 320 68
rect 50 -32 320 -4
rect 252 -65 318 -60
rect 252 -117 259 -65
rect 311 -117 318 -65
rect 252 -126 318 -117
rect 404 -156 432 70
rect 626 58 672 89
rect 744 627 790 658
rect 744 593 750 627
rect 784 593 790 627
rect 744 555 790 593
rect 744 521 750 555
rect 784 521 790 555
rect 744 483 790 521
rect 744 449 750 483
rect 784 449 790 483
rect 744 411 790 449
rect 744 377 750 411
rect 784 377 790 411
rect 744 339 790 377
rect 744 305 750 339
rect 784 305 790 339
rect 744 267 790 305
rect 744 233 750 267
rect 784 233 790 267
rect 744 195 790 233
rect 744 161 750 195
rect 784 161 790 195
rect 744 123 790 161
rect 744 89 750 123
rect 784 89 790 123
rect 744 58 790 89
rect 862 627 908 658
rect 862 593 868 627
rect 902 593 908 627
rect 862 555 908 593
rect 862 521 868 555
rect 902 521 908 555
rect 862 483 908 521
rect 862 449 868 483
rect 902 449 908 483
rect 862 411 908 449
rect 862 377 868 411
rect 902 377 908 411
rect 862 339 908 377
rect 862 305 868 339
rect 902 305 908 339
rect 862 267 908 305
rect 862 233 868 267
rect 902 233 908 267
rect 862 195 908 233
rect 862 161 868 195
rect 902 161 908 195
rect 862 123 908 161
rect 862 89 868 123
rect 902 89 908 123
rect 862 58 908 89
rect 980 627 1026 658
rect 980 593 986 627
rect 1020 593 1026 627
rect 980 555 1026 593
rect 980 521 986 555
rect 1020 521 1026 555
rect 980 483 1026 521
rect 980 449 986 483
rect 1020 449 1026 483
rect 980 411 1026 449
rect 980 377 986 411
rect 1020 377 1026 411
rect 980 339 1026 377
rect 980 305 986 339
rect 1020 305 1026 339
rect 980 267 1026 305
rect 980 233 986 267
rect 1020 233 1026 267
rect 980 195 1026 233
rect 980 161 986 195
rect 1020 161 1026 195
rect 980 123 1026 161
rect 980 89 986 123
rect 1020 89 1026 123
rect 980 58 1026 89
rect 1098 627 1144 658
rect 1098 593 1104 627
rect 1138 593 1144 627
rect 1098 555 1144 593
rect 1098 521 1104 555
rect 1138 521 1144 555
rect 1098 483 1144 521
rect 1098 449 1104 483
rect 1138 449 1144 483
rect 1098 411 1144 449
rect 1098 377 1104 411
rect 1138 377 1144 411
rect 1098 339 1144 377
rect 1098 305 1104 339
rect 1138 305 1144 339
rect 1098 267 1144 305
rect 1098 233 1104 267
rect 1138 233 1144 267
rect 1098 195 1144 233
rect 1098 161 1104 195
rect 1138 161 1144 195
rect 1098 123 1144 161
rect 1098 89 1104 123
rect 1138 89 1144 123
rect 1098 58 1144 89
rect 1218 627 1264 658
rect 1218 593 1224 627
rect 1258 593 1264 627
rect 1218 555 1264 593
rect 1218 521 1224 555
rect 1258 521 1264 555
rect 1218 483 1264 521
rect 1218 449 1224 483
rect 1258 449 1264 483
rect 1218 411 1264 449
rect 1218 377 1224 411
rect 1258 377 1264 411
rect 1218 339 1264 377
rect 1218 305 1224 339
rect 1258 305 1264 339
rect 1218 267 1264 305
rect 1218 233 1224 267
rect 1258 233 1264 267
rect 1218 195 1264 233
rect 1218 161 1224 195
rect 1258 161 1264 195
rect 1218 123 1264 161
rect 1218 89 1224 123
rect 1258 89 1264 123
rect 1218 58 1264 89
rect 1336 627 1382 658
rect 1336 593 1342 627
rect 1376 593 1382 627
rect 1336 555 1382 593
rect 1336 521 1342 555
rect 1376 521 1382 555
rect 1336 483 1382 521
rect 1336 449 1342 483
rect 1376 449 1382 483
rect 1336 411 1382 449
rect 1336 377 1342 411
rect 1376 377 1382 411
rect 1336 339 1382 377
rect 1336 305 1342 339
rect 1376 305 1382 339
rect 1336 267 1382 305
rect 1336 233 1342 267
rect 1376 233 1382 267
rect 1336 195 1382 233
rect 1336 161 1342 195
rect 1376 161 1382 195
rect 1336 123 1382 161
rect 1336 89 1342 123
rect 1376 89 1382 123
rect 1336 58 1382 89
rect 1454 627 1500 658
rect 1454 593 1460 627
rect 1494 593 1500 627
rect 1454 555 1500 593
rect 1454 521 1460 555
rect 1494 521 1500 555
rect 1454 483 1500 521
rect 1454 449 1460 483
rect 1494 449 1500 483
rect 1454 411 1500 449
rect 1454 377 1460 411
rect 1494 377 1500 411
rect 1454 339 1500 377
rect 1454 305 1460 339
rect 1494 305 1500 339
rect 1454 267 1500 305
rect 1454 233 1460 267
rect 1494 233 1500 267
rect 1454 195 1500 233
rect 1454 161 1460 195
rect 1494 161 1500 195
rect 1454 123 1500 161
rect 1454 89 1460 123
rect 1494 89 1500 123
rect 1454 58 1500 89
rect 1572 627 1618 658
rect 1572 593 1578 627
rect 1612 593 1618 627
rect 1572 555 1618 593
rect 1572 521 1578 555
rect 1612 521 1618 555
rect 1572 483 1618 521
rect 1572 449 1578 483
rect 1612 449 1618 483
rect 1572 411 1618 449
rect 1572 377 1578 411
rect 1612 377 1618 411
rect 1572 339 1618 377
rect 1572 305 1578 339
rect 1612 305 1618 339
rect 1572 267 1618 305
rect 1572 233 1578 267
rect 1612 233 1618 267
rect 1572 195 1618 233
rect 1572 161 1578 195
rect 1612 161 1618 195
rect 1572 123 1618 161
rect 1572 89 1578 123
rect 1612 89 1618 123
rect 1572 58 1618 89
rect 1690 627 1736 658
rect 1690 593 1696 627
rect 1730 593 1736 627
rect 1690 555 1736 593
rect 1690 521 1696 555
rect 1730 521 1736 555
rect 1690 483 1736 521
rect 1690 449 1696 483
rect 1730 449 1736 483
rect 1690 411 1736 449
rect 1690 377 1696 411
rect 1730 377 1736 411
rect 1690 339 1736 377
rect 1690 305 1696 339
rect 1730 305 1736 339
rect 1690 267 1736 305
rect 1690 233 1696 267
rect 1730 233 1736 267
rect 1690 195 1736 233
rect 1690 161 1696 195
rect 1730 161 1736 195
rect 1690 123 1736 161
rect 1690 89 1696 123
rect 1730 89 1736 123
rect 1690 58 1736 89
rect 634 -8 664 58
rect 874 -8 904 58
rect 634 -36 904 -8
rect 486 -57 552 -52
rect 486 -109 493 -57
rect 545 -109 552 -57
rect 486 -118 552 -109
rect 810 -70 878 -64
rect 810 -122 818 -70
rect 870 -122 878 -70
rect 810 -132 878 -122
rect 628 -156 706 -146
rect 216 -175 294 -160
rect 216 -227 227 -175
rect 279 -227 294 -175
rect 216 -240 294 -227
rect 404 -170 706 -156
rect 404 -184 648 -170
rect 36 -347 98 -338
rect 36 -399 42 -347
rect 94 -399 98 -347
rect 36 -408 98 -399
rect 404 -402 432 -184
rect 628 -204 648 -184
rect 682 -204 706 -170
rect 628 -226 706 -204
rect 988 -154 1016 58
rect 1226 -8 1256 58
rect 1466 -8 1496 58
rect 1226 -36 1496 -8
rect 1076 -66 1148 -48
rect 1076 -118 1084 -66
rect 1136 -118 1148 -66
rect 1076 -124 1148 -118
rect 1396 -72 1466 -66
rect 1396 -124 1405 -72
rect 1457 -124 1466 -72
rect 1396 -130 1466 -124
rect 1238 -154 1316 -148
rect 988 -172 1316 -154
rect 988 -182 1258 -172
rect 552 -355 622 -346
rect 552 -407 558 -355
rect 610 -407 622 -355
rect 988 -402 1016 -182
rect 1238 -206 1258 -182
rect 1292 -206 1316 -172
rect 1238 -226 1316 -206
rect 1580 -178 1608 58
rect 1814 -26 1846 26
rect 2044 -26 2072 28
rect 1640 -63 1728 -48
rect 1814 -54 2072 -26
rect 1640 -115 1658 -63
rect 1710 -115 1728 -63
rect 1640 -124 1728 -115
rect 1872 -90 1942 -82
rect 1872 -142 1881 -90
rect 1933 -142 1942 -90
rect 1872 -148 1942 -142
rect 1756 -171 1834 -156
rect 1756 -178 1767 -171
rect 1580 -210 1767 -178
rect 1152 -357 1222 -346
rect 552 -418 622 -407
rect 742 -433 788 -402
rect 742 -467 748 -433
rect 782 -467 788 -433
rect 742 -505 788 -467
rect 742 -539 748 -505
rect 782 -539 788 -505
rect 742 -577 788 -539
rect 742 -611 748 -577
rect 782 -611 788 -577
rect 742 -649 788 -611
rect 742 -683 748 -649
rect 782 -683 788 -649
rect 742 -721 788 -683
rect -182 -1242 -146 -742
rect 742 -755 748 -721
rect 782 -755 788 -721
rect 742 -793 788 -755
rect 742 -827 748 -793
rect 782 -827 788 -793
rect 742 -865 788 -827
rect 742 -899 748 -865
rect 782 -899 788 -865
rect 742 -937 788 -899
rect 554 -964 616 -958
rect 38 -1006 96 -998
rect 38 -1058 42 -1006
rect 94 -1058 96 -1006
rect 38 -1066 96 -1058
rect 36 -1229 100 -1224
rect -200 -1255 -128 -1242
rect -200 -1289 -181 -1255
rect -147 -1289 -128 -1255
rect -200 -1306 -128 -1289
rect 36 -1281 42 -1229
rect 94 -1281 100 -1229
rect 164 -1252 202 -988
rect 554 -1016 558 -964
rect 610 -1016 616 -964
rect 742 -971 748 -937
rect 782 -971 788 -937
rect 742 -1002 788 -971
rect 860 -433 906 -402
rect 860 -467 866 -433
rect 900 -467 906 -433
rect 860 -505 906 -467
rect 860 -539 866 -505
rect 900 -539 906 -505
rect 860 -577 906 -539
rect 860 -611 866 -577
rect 900 -611 906 -577
rect 860 -649 906 -611
rect 860 -683 866 -649
rect 900 -683 906 -649
rect 860 -721 906 -683
rect 860 -755 866 -721
rect 900 -755 906 -721
rect 860 -793 906 -755
rect 860 -827 866 -793
rect 900 -827 906 -793
rect 860 -865 906 -827
rect 860 -899 866 -865
rect 900 -899 906 -865
rect 860 -937 906 -899
rect 860 -971 866 -937
rect 900 -971 906 -937
rect 860 -1002 906 -971
rect 978 -433 1024 -402
rect 1152 -409 1160 -357
rect 1212 -409 1222 -357
rect 1580 -402 1608 -210
rect 1756 -223 1767 -210
rect 1819 -223 1834 -171
rect 1756 -236 1834 -223
rect 2044 -178 2072 -54
rect 2106 -58 2180 -48
rect 2106 -110 2118 -58
rect 2170 -110 2180 -58
rect 2106 -122 2180 -110
rect 2244 -60 2318 -48
rect 2244 -112 2254 -60
rect 2306 -112 2318 -60
rect 2244 -120 2318 -112
rect 2172 -174 2250 -150
rect 2172 -178 2192 -174
rect 2044 -208 2192 -178
rect 2226 -208 2250 -174
rect 2044 -210 2250 -208
rect 1744 -361 1810 -354
rect 1152 -418 1222 -409
rect 978 -467 984 -433
rect 1018 -467 1024 -433
rect 978 -505 1024 -467
rect 978 -539 984 -505
rect 1018 -539 1024 -505
rect 978 -577 1024 -539
rect 978 -611 984 -577
rect 1018 -611 1024 -577
rect 978 -649 1024 -611
rect 978 -683 984 -649
rect 1018 -683 1024 -649
rect 978 -721 1024 -683
rect 978 -755 984 -721
rect 1018 -755 1024 -721
rect 978 -793 1024 -755
rect 978 -827 984 -793
rect 1018 -827 1024 -793
rect 978 -865 1024 -827
rect 978 -899 984 -865
rect 1018 -899 1024 -865
rect 978 -937 1024 -899
rect 978 -971 984 -937
rect 1018 -971 1024 -937
rect 1334 -433 1380 -402
rect 1334 -467 1340 -433
rect 1374 -467 1380 -433
rect 1334 -505 1380 -467
rect 1334 -539 1340 -505
rect 1374 -539 1380 -505
rect 1334 -577 1380 -539
rect 1334 -611 1340 -577
rect 1374 -611 1380 -577
rect 1334 -649 1380 -611
rect 1334 -683 1340 -649
rect 1374 -683 1380 -649
rect 1334 -721 1380 -683
rect 1334 -755 1340 -721
rect 1374 -755 1380 -721
rect 1334 -793 1380 -755
rect 1334 -827 1340 -793
rect 1374 -827 1380 -793
rect 1334 -865 1380 -827
rect 1334 -899 1340 -865
rect 1374 -899 1380 -865
rect 1334 -937 1380 -899
rect 978 -1002 1024 -971
rect 1154 -966 1218 -964
rect 554 -1022 616 -1016
rect 536 -1249 626 -1238
rect 752 -1248 780 -1002
rect 1154 -1018 1160 -966
rect 1212 -1018 1218 -966
rect 1334 -971 1340 -937
rect 1374 -971 1380 -937
rect 1334 -1002 1380 -971
rect 1452 -433 1498 -402
rect 1452 -467 1458 -433
rect 1492 -467 1498 -433
rect 1452 -505 1498 -467
rect 1452 -539 1458 -505
rect 1492 -539 1498 -505
rect 1452 -577 1498 -539
rect 1452 -611 1458 -577
rect 1492 -611 1498 -577
rect 1452 -649 1498 -611
rect 1452 -683 1458 -649
rect 1492 -683 1498 -649
rect 1452 -721 1498 -683
rect 1452 -755 1458 -721
rect 1492 -755 1498 -721
rect 1452 -793 1498 -755
rect 1452 -827 1458 -793
rect 1492 -827 1498 -793
rect 1452 -865 1498 -827
rect 1452 -899 1458 -865
rect 1492 -899 1498 -865
rect 1452 -937 1498 -899
rect 1452 -971 1458 -937
rect 1492 -971 1498 -937
rect 1452 -1002 1498 -971
rect 1570 -433 1616 -402
rect 1744 -413 1754 -361
rect 1806 -413 1810 -361
rect 1744 -424 1810 -413
rect 2044 -416 2072 -210
rect 2172 -230 2250 -210
rect 2404 -170 2434 22
rect 2694 -170 2776 -140
rect 2404 -202 2776 -170
rect 2216 -294 2280 -290
rect 2216 -346 2222 -294
rect 2274 -346 2280 -294
rect 2216 -354 2280 -346
rect 2404 -412 2434 -202
rect 2694 -226 2776 -202
rect 2486 -300 2556 -292
rect 2486 -352 2500 -300
rect 2552 -352 2556 -300
rect 2486 -364 2556 -352
rect 1570 -467 1576 -433
rect 1610 -467 1616 -433
rect 1570 -505 1616 -467
rect 1570 -539 1576 -505
rect 1610 -539 1616 -505
rect 1570 -577 1616 -539
rect 1570 -611 1576 -577
rect 1610 -611 1616 -577
rect 1570 -649 1616 -611
rect 1570 -683 1576 -649
rect 1610 -683 1616 -649
rect 1570 -721 1616 -683
rect 1570 -755 1576 -721
rect 1610 -755 1616 -721
rect 1570 -793 1616 -755
rect 1570 -827 1576 -793
rect 1610 -827 1616 -793
rect 1570 -865 1616 -827
rect 1570 -899 1576 -865
rect 1610 -899 1616 -865
rect 1570 -937 1616 -899
rect 1570 -971 1576 -937
rect 1610 -971 1616 -937
rect 1570 -1002 1616 -971
rect 1154 -1024 1218 -1018
rect 1340 -1244 1372 -1002
rect 36 -1292 100 -1281
rect 150 -1262 218 -1252
rect 150 -1296 166 -1262
rect 200 -1296 218 -1262
rect 150 -1310 218 -1296
rect 536 -1301 555 -1249
rect 607 -1301 626 -1249
rect 536 -1316 626 -1301
rect 734 -1261 800 -1248
rect 734 -1295 749 -1261
rect 783 -1295 800 -1261
rect 734 -1312 800 -1295
rect 1146 -1257 1230 -1246
rect 1146 -1309 1162 -1257
rect 1214 -1309 1230 -1257
rect 1146 -1320 1230 -1309
rect 1318 -1262 1390 -1244
rect 1932 -1246 1964 -1098
rect 1318 -1296 1336 -1262
rect 1370 -1296 1390 -1262
rect 1318 -1314 1390 -1296
rect 1910 -1260 1982 -1246
rect 2278 -1254 2316 -1102
rect 1910 -1294 1928 -1260
rect 1962 -1294 1982 -1260
rect 1910 -1310 1982 -1294
rect 2264 -1263 2328 -1254
rect 2264 -1297 2278 -1263
rect 2312 -1297 2328 -1263
rect 2264 -1310 2328 -1297
<< via1 >>
rect 2127 758 2179 810
rect 2413 760 2465 812
rect -354 -348 -302 -340
rect -354 -382 -346 -348
rect -346 -382 -312 -348
rect -312 -382 -302 -348
rect -354 -392 -302 -382
rect 259 -72 311 -65
rect 259 -106 268 -72
rect 268 -106 302 -72
rect 302 -106 311 -72
rect 259 -117 311 -106
rect 493 -64 545 -57
rect 493 -98 500 -64
rect 500 -98 534 -64
rect 534 -98 545 -64
rect 493 -109 545 -98
rect 818 -76 870 -70
rect 818 -110 827 -76
rect 827 -110 861 -76
rect 861 -110 870 -76
rect 818 -122 870 -110
rect 227 -184 279 -175
rect 227 -218 236 -184
rect 236 -218 270 -184
rect 270 -218 279 -184
rect 227 -227 279 -218
rect 42 -357 94 -347
rect 42 -391 50 -357
rect 50 -391 84 -357
rect 84 -391 94 -357
rect 42 -399 94 -391
rect 1084 -68 1136 -66
rect 1084 -102 1091 -68
rect 1091 -102 1125 -68
rect 1125 -102 1136 -68
rect 1084 -118 1136 -102
rect 1405 -74 1457 -72
rect 1405 -108 1414 -74
rect 1414 -108 1448 -74
rect 1448 -108 1457 -74
rect 1405 -124 1457 -108
rect 558 -364 610 -355
rect 558 -398 565 -364
rect 565 -398 599 -364
rect 599 -398 610 -364
rect 558 -407 610 -398
rect 1658 -69 1710 -63
rect 1658 -103 1664 -69
rect 1664 -103 1698 -69
rect 1698 -103 1710 -69
rect 1658 -115 1710 -103
rect 1881 -96 1933 -90
rect 1881 -130 1891 -96
rect 1891 -130 1925 -96
rect 1925 -130 1933 -96
rect 1881 -142 1933 -130
rect 1767 -180 1819 -171
rect 42 -1017 94 -1006
rect 42 -1051 52 -1017
rect 52 -1051 86 -1017
rect 86 -1051 94 -1017
rect 42 -1058 94 -1051
rect 42 -1237 94 -1229
rect 42 -1271 53 -1237
rect 53 -1271 87 -1237
rect 87 -1271 94 -1237
rect 42 -1281 94 -1271
rect 558 -974 610 -964
rect 558 -1008 568 -974
rect 568 -1008 602 -974
rect 602 -1008 610 -974
rect 558 -1016 610 -1008
rect 1160 -365 1212 -357
rect 1160 -399 1172 -365
rect 1172 -399 1206 -365
rect 1206 -399 1212 -365
rect 1160 -409 1212 -399
rect 1767 -214 1776 -180
rect 1776 -214 1810 -180
rect 1810 -214 1819 -180
rect 1767 -223 1819 -214
rect 2118 -74 2170 -58
rect 2118 -108 2129 -74
rect 2129 -108 2163 -74
rect 2163 -108 2170 -74
rect 2118 -110 2170 -108
rect 2254 -70 2306 -60
rect 2254 -104 2262 -70
rect 2262 -104 2296 -70
rect 2296 -104 2306 -70
rect 2254 -112 2306 -104
rect 1160 -976 1212 -966
rect 1160 -1010 1169 -976
rect 1169 -1010 1203 -976
rect 1203 -1010 1212 -976
rect 1160 -1018 1212 -1010
rect 1754 -368 1806 -361
rect 1754 -402 1764 -368
rect 1764 -402 1798 -368
rect 1798 -402 1806 -368
rect 1754 -413 1806 -402
rect 2222 -306 2274 -294
rect 2222 -340 2230 -306
rect 2230 -340 2264 -306
rect 2264 -340 2274 -306
rect 2222 -346 2274 -340
rect 2500 -309 2552 -300
rect 2500 -343 2509 -309
rect 2509 -343 2543 -309
rect 2543 -343 2552 -309
rect 2500 -352 2552 -343
rect 555 -1259 607 -1249
rect 555 -1293 563 -1259
rect 563 -1293 597 -1259
rect 597 -1293 607 -1259
rect 555 -1301 607 -1293
rect 1162 -1267 1214 -1257
rect 1162 -1301 1170 -1267
rect 1170 -1301 1204 -1267
rect 1204 -1301 1214 -1267
rect 1162 -1309 1214 -1301
<< metal2 >>
rect 2164 826 2432 854
rect 2164 824 2486 826
rect 2164 820 2196 824
rect 2110 810 2196 820
rect 2110 758 2127 810
rect 2179 758 2196 810
rect 2110 746 2196 758
rect 2404 812 2486 824
rect 2404 760 2413 812
rect 2465 760 2486 812
rect 2404 748 2486 760
rect 252 -65 318 -56
rect 252 -117 259 -65
rect 311 -74 318 -65
rect 486 -57 552 -52
rect 486 -74 493 -57
rect 311 -106 493 -74
rect 311 -117 318 -106
rect 252 -126 318 -117
rect 486 -109 493 -106
rect 545 -109 552 -57
rect 812 -64 876 -58
rect 486 -118 552 -109
rect 810 -70 878 -64
rect 1076 -66 1148 -52
rect 1640 -63 1728 -48
rect 1076 -70 1084 -66
rect 810 -122 818 -70
rect 870 -100 1084 -70
rect 870 -122 878 -100
rect 810 -132 878 -122
rect 1076 -118 1084 -100
rect 1136 -118 1148 -66
rect 1076 -128 1148 -118
rect 1396 -72 1466 -66
rect 1396 -124 1405 -72
rect 1457 -74 1466 -72
rect 1640 -74 1658 -63
rect 1457 -104 1658 -74
rect 1457 -124 1466 -104
rect 1640 -115 1658 -104
rect 1710 -115 1728 -63
rect 2106 -58 2180 -48
rect 2106 -82 2118 -58
rect 1640 -124 1728 -115
rect 1872 -90 2118 -82
rect 1396 -130 1466 -124
rect 1872 -142 1881 -90
rect 1933 -110 2118 -90
rect 2170 -110 2180 -58
rect 1933 -142 1942 -110
rect 2106 -122 2180 -110
rect 2244 -60 2318 -48
rect 2244 -112 2254 -60
rect 2306 -82 2318 -60
rect 2306 -110 2520 -82
rect 2306 -112 2318 -110
rect 2244 -120 2318 -112
rect 1872 -148 1942 -142
rect 214 -175 296 -160
rect 214 -184 227 -175
rect 154 -216 227 -184
rect 154 -272 186 -216
rect 214 -227 227 -216
rect 279 -227 296 -175
rect 214 -242 296 -227
rect 1754 -171 1836 -156
rect 1754 -223 1767 -171
rect 1819 -223 1836 -171
rect 1754 -238 1836 -223
rect 1780 -272 1812 -238
rect 154 -302 1812 -272
rect 2216 -294 2280 -290
rect 2216 -324 2222 -294
rect -338 -330 82 -324
rect 2202 -330 2222 -324
rect -338 -332 606 -330
rect 1170 -332 1210 -330
rect 1760 -332 2222 -330
rect -338 -334 2222 -332
rect -362 -340 2222 -334
rect -362 -392 -354 -340
rect -302 -346 2222 -340
rect 2274 -308 2280 -294
rect 2486 -300 2556 -292
rect 2486 -308 2500 -300
rect 2274 -336 2500 -308
rect 2274 -346 2280 -336
rect -302 -347 2280 -346
rect -302 -354 42 -347
rect -302 -392 -290 -354
rect -362 -398 -290 -392
rect -362 -400 -292 -398
rect 36 -399 42 -354
rect 94 -354 2280 -347
rect 2486 -352 2500 -336
rect 2552 -352 2556 -300
rect 94 -355 2230 -354
rect 94 -360 558 -355
rect 94 -399 98 -360
rect 36 -408 98 -399
rect 550 -407 558 -360
rect 610 -357 2230 -355
rect 610 -364 1160 -357
rect 610 -407 622 -364
rect 550 -418 622 -407
rect 1152 -409 1160 -364
rect 1212 -360 2230 -357
rect 1212 -409 1222 -360
rect 1152 -418 1222 -409
rect 1744 -361 1810 -360
rect 1744 -413 1754 -361
rect 1806 -413 1810 -361
rect 2486 -364 2556 -352
rect 1744 -424 1810 -413
rect 552 -964 618 -958
rect 38 -1006 96 -998
rect 38 -1058 42 -1006
rect 94 -1058 96 -1006
rect 552 -1016 558 -964
rect 610 -1016 618 -964
rect 552 -1024 618 -1016
rect 1152 -966 1220 -964
rect 1152 -1018 1160 -966
rect 1212 -1018 1220 -966
rect 38 -1066 96 -1058
rect 50 -1224 82 -1066
rect 36 -1229 100 -1224
rect 36 -1281 42 -1229
rect 94 -1281 100 -1229
rect 562 -1238 604 -1024
rect 1152 -1026 1220 -1018
rect 36 -1292 100 -1281
rect 536 -1249 626 -1238
rect 1168 -1244 1210 -1026
rect 536 -1301 555 -1249
rect 607 -1301 626 -1249
rect 536 -1316 626 -1301
rect 1144 -1257 1232 -1244
rect 1144 -1309 1162 -1257
rect 1214 -1309 1232 -1257
rect 1144 -1322 1232 -1309
use sky130_fd_pr__nfet_01v8_7R257D  sky130_fd_pr__nfet_01v8_7R257D_0
timestamp 1669522153
transform 1 0 -104 0 1 -572
box -114 -206 114 206
use sky130_fd_pr__nfet_01v8_M8KAMF  sky130_fd_pr__nfet_01v8_M8KAMF_0
timestamp 1669522153
transform 1 0 240 0 1 -698
box -114 -326 114 326
use sky130_fd_pr__nfet_01v8_N56T4C  sky130_fd_pr__nfet_01v8_N56T4C_0
timestamp 1669522153
transform 1 0 358 0 1 -698
box -114 -326 114 326
use sky130_fd_pr__nfet_01v8_ZU5QBV  sky130_fd_pr__nfet_01v8_ZU5QBV_0
timestamp 1669522153
transform 1 0 2008 0 1 -756
box -114 -376 114 376
use sky130_fd_pr__nfet_01v8_ZU5QBV  sky130_fd_pr__nfet_01v8_ZU5QBV_1
timestamp 1669522153
transform 1 0 2358 0 1 -758
box -114 -376 114 376
use sky130_fd_pr__pfet_01v8_EKD6RN  sky130_fd_pr__pfet_01v8_EKD6RN_0
timestamp 1669522153
transform 1 0 419 0 1 362
box -183 -362 183 362
use sky130_fd_pr__pfet_01v8_EKD6RN  sky130_fd_pr__pfet_01v8_EKD6RN_1
timestamp 1669522153
transform 1 0 183 0 1 362
box -183 -362 183 362
use sky130_fd_pr__pfet_01v8_GRHA7T  sky130_fd_pr__pfet_01v8_GRHA7T_0
timestamp 1669522153
transform 1 0 -106 0 1 382
box -124 -302 124 302
use sky130_fd_pr__pfet_01v8_JJT9EJ  sky130_fd_pr__pfet_01v8_JJT9EJ_0
timestamp 1669522153
transform 1 0 2299 0 1 366
box -183 -412 183 412
use sky130_fd_pr__pfet_01v8_JJT9EJ  sky130_fd_pr__pfet_01v8_JJT9EJ_1
timestamp 1669522153
transform 1 0 1947 0 1 366
box -183 -412 183 412
<< labels >>
rlabel locali s -382 -1322 2596 -1252 4 gnd
port 1 nsew
rlabel metal1 s -800 -278 -720 -194 4 In
port 2 nsew
rlabel metal1 s 2716 -212 2760 -152 4 Out
port 3 nsew
rlabel nwell s -232 894 2424 940 4 VDD
port 4 nsew
<< end >>
