magic
tech sky130A
magscale 1 2
timestamp 1667321908
<< nmoslvt >>
rect -270 60163 270 79963
rect -270 40145 270 59945
rect -270 20127 270 39927
rect -270 109 270 19909
rect -270 -19909 270 -109
rect -270 -39927 270 -20127
rect -270 -59945 270 -40145
rect -270 -79963 270 -60163
<< ndiff >>
rect -328 79951 -270 79963
rect -328 60175 -316 79951
rect -282 60175 -270 79951
rect -328 60163 -270 60175
rect 270 79951 328 79963
rect 270 60175 282 79951
rect 316 60175 328 79951
rect 270 60163 328 60175
rect -328 59933 -270 59945
rect -328 40157 -316 59933
rect -282 40157 -270 59933
rect -328 40145 -270 40157
rect 270 59933 328 59945
rect 270 40157 282 59933
rect 316 40157 328 59933
rect 270 40145 328 40157
rect -328 39915 -270 39927
rect -328 20139 -316 39915
rect -282 20139 -270 39915
rect -328 20127 -270 20139
rect 270 39915 328 39927
rect 270 20139 282 39915
rect 316 20139 328 39915
rect 270 20127 328 20139
rect -328 19897 -270 19909
rect -328 121 -316 19897
rect -282 121 -270 19897
rect -328 109 -270 121
rect 270 19897 328 19909
rect 270 121 282 19897
rect 316 121 328 19897
rect 270 109 328 121
rect -328 -121 -270 -109
rect -328 -19897 -316 -121
rect -282 -19897 -270 -121
rect -328 -19909 -270 -19897
rect 270 -121 328 -109
rect 270 -19897 282 -121
rect 316 -19897 328 -121
rect 270 -19909 328 -19897
rect -328 -20139 -270 -20127
rect -328 -39915 -316 -20139
rect -282 -39915 -270 -20139
rect -328 -39927 -270 -39915
rect 270 -20139 328 -20127
rect 270 -39915 282 -20139
rect 316 -39915 328 -20139
rect 270 -39927 328 -39915
rect -328 -40157 -270 -40145
rect -328 -59933 -316 -40157
rect -282 -59933 -270 -40157
rect -328 -59945 -270 -59933
rect 270 -40157 328 -40145
rect 270 -59933 282 -40157
rect 316 -59933 328 -40157
rect 270 -59945 328 -59933
rect -328 -60175 -270 -60163
rect -328 -79951 -316 -60175
rect -282 -79951 -270 -60175
rect -328 -79963 -270 -79951
rect 270 -60175 328 -60163
rect 270 -79951 282 -60175
rect 316 -79951 328 -60175
rect 270 -79963 328 -79951
<< ndiffc >>
rect -316 60175 -282 79951
rect 282 60175 316 79951
rect -316 40157 -282 59933
rect 282 40157 316 59933
rect -316 20139 -282 39915
rect 282 20139 316 39915
rect -316 121 -282 19897
rect 282 121 316 19897
rect -316 -19897 -282 -121
rect 282 -19897 316 -121
rect -316 -39915 -282 -20139
rect 282 -39915 316 -20139
rect -316 -59933 -282 -40157
rect 282 -59933 316 -40157
rect -316 -79951 -282 -60175
rect 282 -79951 316 -60175
<< poly >>
rect -270 80035 270 80051
rect -270 80001 -254 80035
rect 254 80001 270 80035
rect -270 79963 270 80001
rect -270 60125 270 60163
rect -270 60091 -254 60125
rect 254 60091 270 60125
rect -270 60075 270 60091
rect -270 60017 270 60033
rect -270 59983 -254 60017
rect 254 59983 270 60017
rect -270 59945 270 59983
rect -270 40107 270 40145
rect -270 40073 -254 40107
rect 254 40073 270 40107
rect -270 40057 270 40073
rect -270 39999 270 40015
rect -270 39965 -254 39999
rect 254 39965 270 39999
rect -270 39927 270 39965
rect -270 20089 270 20127
rect -270 20055 -254 20089
rect 254 20055 270 20089
rect -270 20039 270 20055
rect -270 19981 270 19997
rect -270 19947 -254 19981
rect 254 19947 270 19981
rect -270 19909 270 19947
rect -270 71 270 109
rect -270 37 -254 71
rect 254 37 270 71
rect -270 21 270 37
rect -270 -37 270 -21
rect -270 -71 -254 -37
rect 254 -71 270 -37
rect -270 -109 270 -71
rect -270 -19947 270 -19909
rect -270 -19981 -254 -19947
rect 254 -19981 270 -19947
rect -270 -19997 270 -19981
rect -270 -20055 270 -20039
rect -270 -20089 -254 -20055
rect 254 -20089 270 -20055
rect -270 -20127 270 -20089
rect -270 -39965 270 -39927
rect -270 -39999 -254 -39965
rect 254 -39999 270 -39965
rect -270 -40015 270 -39999
rect -270 -40073 270 -40057
rect -270 -40107 -254 -40073
rect 254 -40107 270 -40073
rect -270 -40145 270 -40107
rect -270 -59983 270 -59945
rect -270 -60017 -254 -59983
rect 254 -60017 270 -59983
rect -270 -60033 270 -60017
rect -270 -60091 270 -60075
rect -270 -60125 -254 -60091
rect 254 -60125 270 -60091
rect -270 -60163 270 -60125
rect -270 -80001 270 -79963
rect -270 -80035 -254 -80001
rect 254 -80035 270 -80001
rect -270 -80051 270 -80035
<< polycont >>
rect -254 80001 254 80035
rect -254 60091 254 60125
rect -254 59983 254 60017
rect -254 40073 254 40107
rect -254 39965 254 39999
rect -254 20055 254 20089
rect -254 19947 254 19981
rect -254 37 254 71
rect -254 -71 254 -37
rect -254 -19981 254 -19947
rect -254 -20089 254 -20055
rect -254 -39999 254 -39965
rect -254 -40107 254 -40073
rect -254 -60017 254 -59983
rect -254 -60125 254 -60091
rect -254 -80035 254 -80001
<< locali >>
rect -270 80001 -254 80035
rect 254 80001 270 80035
rect -316 79951 -282 79967
rect -316 60159 -282 60175
rect 282 79951 316 79967
rect 282 60159 316 60175
rect -270 60091 -254 60125
rect 254 60091 270 60125
rect -270 59983 -254 60017
rect 254 59983 270 60017
rect -316 59933 -282 59949
rect -316 40141 -282 40157
rect 282 59933 316 59949
rect 282 40141 316 40157
rect -270 40073 -254 40107
rect 254 40073 270 40107
rect -270 39965 -254 39999
rect 254 39965 270 39999
rect -316 39915 -282 39931
rect -316 20123 -282 20139
rect 282 39915 316 39931
rect 282 20123 316 20139
rect -270 20055 -254 20089
rect 254 20055 270 20089
rect -270 19947 -254 19981
rect 254 19947 270 19981
rect -316 19897 -282 19913
rect -316 105 -282 121
rect 282 19897 316 19913
rect 282 105 316 121
rect -270 37 -254 71
rect 254 37 270 71
rect -270 -71 -254 -37
rect 254 -71 270 -37
rect -316 -121 -282 -105
rect -316 -19913 -282 -19897
rect 282 -121 316 -105
rect 282 -19913 316 -19897
rect -270 -19981 -254 -19947
rect 254 -19981 270 -19947
rect -270 -20089 -254 -20055
rect 254 -20089 270 -20055
rect -316 -20139 -282 -20123
rect -316 -39931 -282 -39915
rect 282 -20139 316 -20123
rect 282 -39931 316 -39915
rect -270 -39999 -254 -39965
rect 254 -39999 270 -39965
rect -270 -40107 -254 -40073
rect 254 -40107 270 -40073
rect -316 -40157 -282 -40141
rect -316 -59949 -282 -59933
rect 282 -40157 316 -40141
rect 282 -59949 316 -59933
rect -270 -60017 -254 -59983
rect 254 -60017 270 -59983
rect -270 -60125 -254 -60091
rect 254 -60125 270 -60091
rect -316 -60175 -282 -60159
rect -316 -79967 -282 -79951
rect 282 -60175 316 -60159
rect 282 -79967 316 -79951
rect -270 -80035 -254 -80001
rect 254 -80035 270 -80001
<< viali >>
rect -254 80001 254 80035
rect -316 60175 -282 79951
rect 282 60175 316 79951
rect -254 60091 254 60125
rect -254 59983 254 60017
rect -316 40157 -282 59933
rect 282 40157 316 59933
rect -254 40073 254 40107
rect -254 39965 254 39999
rect -316 20139 -282 39915
rect 282 20139 316 39915
rect -254 20055 254 20089
rect -254 19947 254 19981
rect -316 121 -282 19897
rect 282 121 316 19897
rect -254 37 254 71
rect -254 -71 254 -37
rect -316 -19897 -282 -121
rect 282 -19897 316 -121
rect -254 -19981 254 -19947
rect -254 -20089 254 -20055
rect -316 -39915 -282 -20139
rect 282 -39915 316 -20139
rect -254 -39999 254 -39965
rect -254 -40107 254 -40073
rect -316 -59933 -282 -40157
rect 282 -59933 316 -40157
rect -254 -60017 254 -59983
rect -254 -60125 254 -60091
rect -316 -79951 -282 -60175
rect 282 -79951 316 -60175
rect -254 -80035 254 -80001
<< metal1 >>
rect -266 80035 266 80041
rect -266 80001 -254 80035
rect 254 80001 266 80035
rect -266 79995 266 80001
rect -322 79951 -276 79963
rect -322 60175 -316 79951
rect -282 60175 -276 79951
rect -322 60163 -276 60175
rect 276 79951 322 79963
rect 276 60175 282 79951
rect 316 60175 322 79951
rect 276 60163 322 60175
rect -266 60125 266 60131
rect -266 60091 -254 60125
rect 254 60091 266 60125
rect -266 60085 266 60091
rect -266 60017 266 60023
rect -266 59983 -254 60017
rect 254 59983 266 60017
rect -266 59977 266 59983
rect -322 59933 -276 59945
rect -322 40157 -316 59933
rect -282 40157 -276 59933
rect -322 40145 -276 40157
rect 276 59933 322 59945
rect 276 40157 282 59933
rect 316 40157 322 59933
rect 276 40145 322 40157
rect -266 40107 266 40113
rect -266 40073 -254 40107
rect 254 40073 266 40107
rect -266 40067 266 40073
rect -266 39999 266 40005
rect -266 39965 -254 39999
rect 254 39965 266 39999
rect -266 39959 266 39965
rect -322 39915 -276 39927
rect -322 20139 -316 39915
rect -282 20139 -276 39915
rect -322 20127 -276 20139
rect 276 39915 322 39927
rect 276 20139 282 39915
rect 316 20139 322 39915
rect 276 20127 322 20139
rect -266 20089 266 20095
rect -266 20055 -254 20089
rect 254 20055 266 20089
rect -266 20049 266 20055
rect -266 19981 266 19987
rect -266 19947 -254 19981
rect 254 19947 266 19981
rect -266 19941 266 19947
rect -322 19897 -276 19909
rect -322 121 -316 19897
rect -282 121 -276 19897
rect -322 109 -276 121
rect 276 19897 322 19909
rect 276 121 282 19897
rect 316 121 322 19897
rect 276 109 322 121
rect -266 71 266 77
rect -266 37 -254 71
rect 254 37 266 71
rect -266 31 266 37
rect -266 -37 266 -31
rect -266 -71 -254 -37
rect 254 -71 266 -37
rect -266 -77 266 -71
rect -322 -121 -276 -109
rect -322 -19897 -316 -121
rect -282 -19897 -276 -121
rect -322 -19909 -276 -19897
rect 276 -121 322 -109
rect 276 -19897 282 -121
rect 316 -19897 322 -121
rect 276 -19909 322 -19897
rect -266 -19947 266 -19941
rect -266 -19981 -254 -19947
rect 254 -19981 266 -19947
rect -266 -19987 266 -19981
rect -266 -20055 266 -20049
rect -266 -20089 -254 -20055
rect 254 -20089 266 -20055
rect -266 -20095 266 -20089
rect -322 -20139 -276 -20127
rect -322 -39915 -316 -20139
rect -282 -39915 -276 -20139
rect -322 -39927 -276 -39915
rect 276 -20139 322 -20127
rect 276 -39915 282 -20139
rect 316 -39915 322 -20139
rect 276 -39927 322 -39915
rect -266 -39965 266 -39959
rect -266 -39999 -254 -39965
rect 254 -39999 266 -39965
rect -266 -40005 266 -39999
rect -266 -40073 266 -40067
rect -266 -40107 -254 -40073
rect 254 -40107 266 -40073
rect -266 -40113 266 -40107
rect -322 -40157 -276 -40145
rect -322 -59933 -316 -40157
rect -282 -59933 -276 -40157
rect -322 -59945 -276 -59933
rect 276 -40157 322 -40145
rect 276 -59933 282 -40157
rect 316 -59933 322 -40157
rect 276 -59945 322 -59933
rect -266 -59983 266 -59977
rect -266 -60017 -254 -59983
rect 254 -60017 266 -59983
rect -266 -60023 266 -60017
rect -266 -60091 266 -60085
rect -266 -60125 -254 -60091
rect 254 -60125 266 -60091
rect -266 -60131 266 -60125
rect -322 -60175 -276 -60163
rect -322 -79951 -316 -60175
rect -282 -79951 -276 -60175
rect -322 -79963 -276 -79951
rect 276 -60175 322 -60163
rect 276 -79951 282 -60175
rect 316 -79951 322 -60175
rect 276 -79963 322 -79951
rect -266 -80001 266 -79995
rect -266 -80035 -254 -80001
rect 254 -80035 266 -80001
rect -266 -80041 266 -80035
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 99.0 l 2.7 m 8 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
