magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect -29 -347 29 -341
<< pwell >>
rect -114 -295 114 357
<< nmos >>
rect -30 -269 30 331
<< ndiff >>
rect -88 286 -30 331
rect -88 252 -76 286
rect -42 252 -30 286
rect -88 218 -30 252
rect -88 184 -76 218
rect -42 184 -30 218
rect -88 150 -30 184
rect -88 116 -76 150
rect -42 116 -30 150
rect -88 82 -30 116
rect -88 48 -76 82
rect -42 48 -30 82
rect -88 14 -30 48
rect -88 -20 -76 14
rect -42 -20 -30 14
rect -88 -54 -30 -20
rect -88 -88 -76 -54
rect -42 -88 -30 -54
rect -88 -122 -30 -88
rect -88 -156 -76 -122
rect -42 -156 -30 -122
rect -88 -190 -30 -156
rect -88 -224 -76 -190
rect -42 -224 -30 -190
rect -88 -269 -30 -224
rect 30 286 88 331
rect 30 252 42 286
rect 76 252 88 286
rect 30 218 88 252
rect 30 184 42 218
rect 76 184 88 218
rect 30 150 88 184
rect 30 116 42 150
rect 76 116 88 150
rect 30 82 88 116
rect 30 48 42 82
rect 76 48 88 82
rect 30 14 88 48
rect 30 -20 42 14
rect 76 -20 88 14
rect 30 -54 88 -20
rect 30 -88 42 -54
rect 76 -88 88 -54
rect 30 -122 88 -88
rect 30 -156 42 -122
rect 76 -156 88 -122
rect 30 -190 88 -156
rect 30 -224 42 -190
rect 76 -224 88 -190
rect 30 -269 88 -224
<< ndiffc >>
rect -76 252 -42 286
rect -76 184 -42 218
rect -76 116 -42 150
rect -76 48 -42 82
rect -76 -20 -42 14
rect -76 -88 -42 -54
rect -76 -156 -42 -122
rect -76 -224 -42 -190
rect 42 252 76 286
rect 42 184 76 218
rect 42 116 76 150
rect 42 48 76 82
rect 42 -20 76 14
rect 42 -88 76 -54
rect 42 -156 76 -122
rect 42 -224 76 -190
<< poly >>
rect -30 331 30 357
rect -30 -291 30 -269
rect -33 -307 33 -291
rect -33 -341 -17 -307
rect 17 -341 33 -307
rect -33 -357 33 -341
<< polycont >>
rect -17 -341 17 -307
<< locali >>
rect -76 300 -42 335
rect -76 228 -42 252
rect -76 156 -42 184
rect -76 84 -42 116
rect -76 14 -42 48
rect -76 -54 -42 -22
rect -76 -122 -42 -94
rect -76 -190 -42 -166
rect -76 -273 -42 -238
rect 42 300 76 335
rect 42 228 76 252
rect 42 156 76 184
rect 42 84 76 116
rect 42 14 76 48
rect 42 -54 76 -22
rect 42 -122 76 -94
rect 42 -190 76 -166
rect 42 -273 76 -238
rect -33 -341 -17 -307
rect 17 -341 33 -307
<< viali >>
rect -76 286 -42 300
rect -76 266 -42 286
rect -76 218 -42 228
rect -76 194 -42 218
rect -76 150 -42 156
rect -76 122 -42 150
rect -76 82 -42 84
rect -76 50 -42 82
rect -76 -20 -42 12
rect -76 -22 -42 -20
rect -76 -88 -42 -60
rect -76 -94 -42 -88
rect -76 -156 -42 -132
rect -76 -166 -42 -156
rect -76 -224 -42 -204
rect -76 -238 -42 -224
rect 42 286 76 300
rect 42 266 76 286
rect 42 218 76 228
rect 42 194 76 218
rect 42 150 76 156
rect 42 122 76 150
rect 42 82 76 84
rect 42 50 76 82
rect 42 -20 76 12
rect 42 -22 76 -20
rect 42 -88 76 -60
rect 42 -94 76 -88
rect 42 -156 76 -132
rect 42 -166 76 -156
rect 42 -224 76 -204
rect 42 -238 76 -224
rect -17 -341 17 -307
<< metal1 >>
rect -82 300 -36 331
rect -82 266 -76 300
rect -42 266 -36 300
rect -82 228 -36 266
rect -82 194 -76 228
rect -42 194 -36 228
rect -82 156 -36 194
rect -82 122 -76 156
rect -42 122 -36 156
rect -82 84 -36 122
rect -82 50 -76 84
rect -42 50 -36 84
rect -82 12 -36 50
rect -82 -22 -76 12
rect -42 -22 -36 12
rect -82 -60 -36 -22
rect -82 -94 -76 -60
rect -42 -94 -36 -60
rect -82 -132 -36 -94
rect -82 -166 -76 -132
rect -42 -166 -36 -132
rect -82 -204 -36 -166
rect -82 -238 -76 -204
rect -42 -238 -36 -204
rect -82 -269 -36 -238
rect 36 300 82 331
rect 36 266 42 300
rect 76 266 82 300
rect 36 228 82 266
rect 36 194 42 228
rect 76 194 82 228
rect 36 156 82 194
rect 36 122 42 156
rect 76 122 82 156
rect 36 84 82 122
rect 36 50 42 84
rect 76 50 82 84
rect 36 12 82 50
rect 36 -22 42 12
rect 76 -22 82 12
rect 36 -60 82 -22
rect 36 -94 42 -60
rect 76 -94 82 -60
rect 36 -132 82 -94
rect 36 -166 42 -132
rect 76 -166 82 -132
rect 36 -204 82 -166
rect 36 -238 42 -204
rect 76 -238 82 -204
rect 36 -269 82 -238
rect -29 -307 29 -301
rect -29 -341 -17 -307
rect 17 -341 29 -307
rect -29 -347 29 -341
<< end >>
