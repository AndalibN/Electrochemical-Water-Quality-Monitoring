magic
tech sky130A
magscale 1 2
timestamp 1666105618
<< nmos >>
rect -50 11071 50 12071
rect -50 9853 50 10853
rect -50 8635 50 9635
rect -50 7417 50 8417
rect -50 6199 50 7199
rect -50 4981 50 5981
rect -50 3763 50 4763
rect -50 2545 50 3545
rect -50 1327 50 2327
rect -50 109 50 1109
rect -50 -1109 50 -109
rect -50 -2327 50 -1327
rect -50 -3545 50 -2545
rect -50 -4763 50 -3763
rect -50 -5981 50 -4981
rect -50 -7199 50 -6199
rect -50 -8417 50 -7417
rect -50 -9635 50 -8635
rect -50 -10853 50 -9853
rect -50 -12071 50 -11071
<< ndiff >>
rect -108 12059 -50 12071
rect -108 11083 -96 12059
rect -62 11083 -50 12059
rect -108 11071 -50 11083
rect 50 12059 108 12071
rect 50 11083 62 12059
rect 96 11083 108 12059
rect 50 11071 108 11083
rect -108 10841 -50 10853
rect -108 9865 -96 10841
rect -62 9865 -50 10841
rect -108 9853 -50 9865
rect 50 10841 108 10853
rect 50 9865 62 10841
rect 96 9865 108 10841
rect 50 9853 108 9865
rect -108 9623 -50 9635
rect -108 8647 -96 9623
rect -62 8647 -50 9623
rect -108 8635 -50 8647
rect 50 9623 108 9635
rect 50 8647 62 9623
rect 96 8647 108 9623
rect 50 8635 108 8647
rect -108 8405 -50 8417
rect -108 7429 -96 8405
rect -62 7429 -50 8405
rect -108 7417 -50 7429
rect 50 8405 108 8417
rect 50 7429 62 8405
rect 96 7429 108 8405
rect 50 7417 108 7429
rect -108 7187 -50 7199
rect -108 6211 -96 7187
rect -62 6211 -50 7187
rect -108 6199 -50 6211
rect 50 7187 108 7199
rect 50 6211 62 7187
rect 96 6211 108 7187
rect 50 6199 108 6211
rect -108 5969 -50 5981
rect -108 4993 -96 5969
rect -62 4993 -50 5969
rect -108 4981 -50 4993
rect 50 5969 108 5981
rect 50 4993 62 5969
rect 96 4993 108 5969
rect 50 4981 108 4993
rect -108 4751 -50 4763
rect -108 3775 -96 4751
rect -62 3775 -50 4751
rect -108 3763 -50 3775
rect 50 4751 108 4763
rect 50 3775 62 4751
rect 96 3775 108 4751
rect 50 3763 108 3775
rect -108 3533 -50 3545
rect -108 2557 -96 3533
rect -62 2557 -50 3533
rect -108 2545 -50 2557
rect 50 3533 108 3545
rect 50 2557 62 3533
rect 96 2557 108 3533
rect 50 2545 108 2557
rect -108 2315 -50 2327
rect -108 1339 -96 2315
rect -62 1339 -50 2315
rect -108 1327 -50 1339
rect 50 2315 108 2327
rect 50 1339 62 2315
rect 96 1339 108 2315
rect 50 1327 108 1339
rect -108 1097 -50 1109
rect -108 121 -96 1097
rect -62 121 -50 1097
rect -108 109 -50 121
rect 50 1097 108 1109
rect 50 121 62 1097
rect 96 121 108 1097
rect 50 109 108 121
rect -108 -121 -50 -109
rect -108 -1097 -96 -121
rect -62 -1097 -50 -121
rect -108 -1109 -50 -1097
rect 50 -121 108 -109
rect 50 -1097 62 -121
rect 96 -1097 108 -121
rect 50 -1109 108 -1097
rect -108 -1339 -50 -1327
rect -108 -2315 -96 -1339
rect -62 -2315 -50 -1339
rect -108 -2327 -50 -2315
rect 50 -1339 108 -1327
rect 50 -2315 62 -1339
rect 96 -2315 108 -1339
rect 50 -2327 108 -2315
rect -108 -2557 -50 -2545
rect -108 -3533 -96 -2557
rect -62 -3533 -50 -2557
rect -108 -3545 -50 -3533
rect 50 -2557 108 -2545
rect 50 -3533 62 -2557
rect 96 -3533 108 -2557
rect 50 -3545 108 -3533
rect -108 -3775 -50 -3763
rect -108 -4751 -96 -3775
rect -62 -4751 -50 -3775
rect -108 -4763 -50 -4751
rect 50 -3775 108 -3763
rect 50 -4751 62 -3775
rect 96 -4751 108 -3775
rect 50 -4763 108 -4751
rect -108 -4993 -50 -4981
rect -108 -5969 -96 -4993
rect -62 -5969 -50 -4993
rect -108 -5981 -50 -5969
rect 50 -4993 108 -4981
rect 50 -5969 62 -4993
rect 96 -5969 108 -4993
rect 50 -5981 108 -5969
rect -108 -6211 -50 -6199
rect -108 -7187 -96 -6211
rect -62 -7187 -50 -6211
rect -108 -7199 -50 -7187
rect 50 -6211 108 -6199
rect 50 -7187 62 -6211
rect 96 -7187 108 -6211
rect 50 -7199 108 -7187
rect -108 -7429 -50 -7417
rect -108 -8405 -96 -7429
rect -62 -8405 -50 -7429
rect -108 -8417 -50 -8405
rect 50 -7429 108 -7417
rect 50 -8405 62 -7429
rect 96 -8405 108 -7429
rect 50 -8417 108 -8405
rect -108 -8647 -50 -8635
rect -108 -9623 -96 -8647
rect -62 -9623 -50 -8647
rect -108 -9635 -50 -9623
rect 50 -8647 108 -8635
rect 50 -9623 62 -8647
rect 96 -9623 108 -8647
rect 50 -9635 108 -9623
rect -108 -9865 -50 -9853
rect -108 -10841 -96 -9865
rect -62 -10841 -50 -9865
rect -108 -10853 -50 -10841
rect 50 -9865 108 -9853
rect 50 -10841 62 -9865
rect 96 -10841 108 -9865
rect 50 -10853 108 -10841
rect -108 -11083 -50 -11071
rect -108 -12059 -96 -11083
rect -62 -12059 -50 -11083
rect -108 -12071 -50 -12059
rect 50 -11083 108 -11071
rect 50 -12059 62 -11083
rect 96 -12059 108 -11083
rect 50 -12071 108 -12059
<< ndiffc >>
rect -96 11083 -62 12059
rect 62 11083 96 12059
rect -96 9865 -62 10841
rect 62 9865 96 10841
rect -96 8647 -62 9623
rect 62 8647 96 9623
rect -96 7429 -62 8405
rect 62 7429 96 8405
rect -96 6211 -62 7187
rect 62 6211 96 7187
rect -96 4993 -62 5969
rect 62 4993 96 5969
rect -96 3775 -62 4751
rect 62 3775 96 4751
rect -96 2557 -62 3533
rect 62 2557 96 3533
rect -96 1339 -62 2315
rect 62 1339 96 2315
rect -96 121 -62 1097
rect 62 121 96 1097
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -96 -2315 -62 -1339
rect 62 -2315 96 -1339
rect -96 -3533 -62 -2557
rect 62 -3533 96 -2557
rect -96 -4751 -62 -3775
rect 62 -4751 96 -3775
rect -96 -5969 -62 -4993
rect 62 -5969 96 -4993
rect -96 -7187 -62 -6211
rect 62 -7187 96 -6211
rect -96 -8405 -62 -7429
rect 62 -8405 96 -7429
rect -96 -9623 -62 -8647
rect 62 -9623 96 -8647
rect -96 -10841 -62 -9865
rect 62 -10841 96 -9865
rect -96 -12059 -62 -11083
rect 62 -12059 96 -11083
<< poly >>
rect -50 12143 50 12159
rect -50 12109 -34 12143
rect 34 12109 50 12143
rect -50 12071 50 12109
rect -50 11033 50 11071
rect -50 10999 -34 11033
rect 34 10999 50 11033
rect -50 10983 50 10999
rect -50 10925 50 10941
rect -50 10891 -34 10925
rect 34 10891 50 10925
rect -50 10853 50 10891
rect -50 9815 50 9853
rect -50 9781 -34 9815
rect 34 9781 50 9815
rect -50 9765 50 9781
rect -50 9707 50 9723
rect -50 9673 -34 9707
rect 34 9673 50 9707
rect -50 9635 50 9673
rect -50 8597 50 8635
rect -50 8563 -34 8597
rect 34 8563 50 8597
rect -50 8547 50 8563
rect -50 8489 50 8505
rect -50 8455 -34 8489
rect 34 8455 50 8489
rect -50 8417 50 8455
rect -50 7379 50 7417
rect -50 7345 -34 7379
rect 34 7345 50 7379
rect -50 7329 50 7345
rect -50 7271 50 7287
rect -50 7237 -34 7271
rect 34 7237 50 7271
rect -50 7199 50 7237
rect -50 6161 50 6199
rect -50 6127 -34 6161
rect 34 6127 50 6161
rect -50 6111 50 6127
rect -50 6053 50 6069
rect -50 6019 -34 6053
rect 34 6019 50 6053
rect -50 5981 50 6019
rect -50 4943 50 4981
rect -50 4909 -34 4943
rect 34 4909 50 4943
rect -50 4893 50 4909
rect -50 4835 50 4851
rect -50 4801 -34 4835
rect 34 4801 50 4835
rect -50 4763 50 4801
rect -50 3725 50 3763
rect -50 3691 -34 3725
rect 34 3691 50 3725
rect -50 3675 50 3691
rect -50 3617 50 3633
rect -50 3583 -34 3617
rect 34 3583 50 3617
rect -50 3545 50 3583
rect -50 2507 50 2545
rect -50 2473 -34 2507
rect 34 2473 50 2507
rect -50 2457 50 2473
rect -50 2399 50 2415
rect -50 2365 -34 2399
rect 34 2365 50 2399
rect -50 2327 50 2365
rect -50 1289 50 1327
rect -50 1255 -34 1289
rect 34 1255 50 1289
rect -50 1239 50 1255
rect -50 1181 50 1197
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -50 1109 50 1147
rect -50 71 50 109
rect -50 37 -34 71
rect 34 37 50 71
rect -50 21 50 37
rect -50 -37 50 -21
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -50 -109 50 -71
rect -50 -1147 50 -1109
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1197 50 -1181
rect -50 -1255 50 -1239
rect -50 -1289 -34 -1255
rect 34 -1289 50 -1255
rect -50 -1327 50 -1289
rect -50 -2365 50 -2327
rect -50 -2399 -34 -2365
rect 34 -2399 50 -2365
rect -50 -2415 50 -2399
rect -50 -2473 50 -2457
rect -50 -2507 -34 -2473
rect 34 -2507 50 -2473
rect -50 -2545 50 -2507
rect -50 -3583 50 -3545
rect -50 -3617 -34 -3583
rect 34 -3617 50 -3583
rect -50 -3633 50 -3617
rect -50 -3691 50 -3675
rect -50 -3725 -34 -3691
rect 34 -3725 50 -3691
rect -50 -3763 50 -3725
rect -50 -4801 50 -4763
rect -50 -4835 -34 -4801
rect 34 -4835 50 -4801
rect -50 -4851 50 -4835
rect -50 -4909 50 -4893
rect -50 -4943 -34 -4909
rect 34 -4943 50 -4909
rect -50 -4981 50 -4943
rect -50 -6019 50 -5981
rect -50 -6053 -34 -6019
rect 34 -6053 50 -6019
rect -50 -6069 50 -6053
rect -50 -6127 50 -6111
rect -50 -6161 -34 -6127
rect 34 -6161 50 -6127
rect -50 -6199 50 -6161
rect -50 -7237 50 -7199
rect -50 -7271 -34 -7237
rect 34 -7271 50 -7237
rect -50 -7287 50 -7271
rect -50 -7345 50 -7329
rect -50 -7379 -34 -7345
rect 34 -7379 50 -7345
rect -50 -7417 50 -7379
rect -50 -8455 50 -8417
rect -50 -8489 -34 -8455
rect 34 -8489 50 -8455
rect -50 -8505 50 -8489
rect -50 -8563 50 -8547
rect -50 -8597 -34 -8563
rect 34 -8597 50 -8563
rect -50 -8635 50 -8597
rect -50 -9673 50 -9635
rect -50 -9707 -34 -9673
rect 34 -9707 50 -9673
rect -50 -9723 50 -9707
rect -50 -9781 50 -9765
rect -50 -9815 -34 -9781
rect 34 -9815 50 -9781
rect -50 -9853 50 -9815
rect -50 -10891 50 -10853
rect -50 -10925 -34 -10891
rect 34 -10925 50 -10891
rect -50 -10941 50 -10925
rect -50 -10999 50 -10983
rect -50 -11033 -34 -10999
rect 34 -11033 50 -10999
rect -50 -11071 50 -11033
rect -50 -12109 50 -12071
rect -50 -12143 -34 -12109
rect 34 -12143 50 -12109
rect -50 -12159 50 -12143
<< polycont >>
rect -34 12109 34 12143
rect -34 10999 34 11033
rect -34 10891 34 10925
rect -34 9781 34 9815
rect -34 9673 34 9707
rect -34 8563 34 8597
rect -34 8455 34 8489
rect -34 7345 34 7379
rect -34 7237 34 7271
rect -34 6127 34 6161
rect -34 6019 34 6053
rect -34 4909 34 4943
rect -34 4801 34 4835
rect -34 3691 34 3725
rect -34 3583 34 3617
rect -34 2473 34 2507
rect -34 2365 34 2399
rect -34 1255 34 1289
rect -34 1147 34 1181
rect -34 37 34 71
rect -34 -71 34 -37
rect -34 -1181 34 -1147
rect -34 -1289 34 -1255
rect -34 -2399 34 -2365
rect -34 -2507 34 -2473
rect -34 -3617 34 -3583
rect -34 -3725 34 -3691
rect -34 -4835 34 -4801
rect -34 -4943 34 -4909
rect -34 -6053 34 -6019
rect -34 -6161 34 -6127
rect -34 -7271 34 -7237
rect -34 -7379 34 -7345
rect -34 -8489 34 -8455
rect -34 -8597 34 -8563
rect -34 -9707 34 -9673
rect -34 -9815 34 -9781
rect -34 -10925 34 -10891
rect -34 -11033 34 -10999
rect -34 -12143 34 -12109
<< locali >>
rect -50 12109 -34 12143
rect 34 12109 50 12143
rect -96 12059 -62 12075
rect -96 11067 -62 11083
rect 62 12059 96 12075
rect 62 11067 96 11083
rect -50 10999 -34 11033
rect 34 10999 50 11033
rect -50 10891 -34 10925
rect 34 10891 50 10925
rect -96 10841 -62 10857
rect -96 9849 -62 9865
rect 62 10841 96 10857
rect 62 9849 96 9865
rect -50 9781 -34 9815
rect 34 9781 50 9815
rect -50 9673 -34 9707
rect 34 9673 50 9707
rect -96 9623 -62 9639
rect -96 8631 -62 8647
rect 62 9623 96 9639
rect 62 8631 96 8647
rect -50 8563 -34 8597
rect 34 8563 50 8597
rect -50 8455 -34 8489
rect 34 8455 50 8489
rect -96 8405 -62 8421
rect -96 7413 -62 7429
rect 62 8405 96 8421
rect 62 7413 96 7429
rect -50 7345 -34 7379
rect 34 7345 50 7379
rect -50 7237 -34 7271
rect 34 7237 50 7271
rect -96 7187 -62 7203
rect -96 6195 -62 6211
rect 62 7187 96 7203
rect 62 6195 96 6211
rect -50 6127 -34 6161
rect 34 6127 50 6161
rect -50 6019 -34 6053
rect 34 6019 50 6053
rect -96 5969 -62 5985
rect -96 4977 -62 4993
rect 62 5969 96 5985
rect 62 4977 96 4993
rect -50 4909 -34 4943
rect 34 4909 50 4943
rect -50 4801 -34 4835
rect 34 4801 50 4835
rect -96 4751 -62 4767
rect -96 3759 -62 3775
rect 62 4751 96 4767
rect 62 3759 96 3775
rect -50 3691 -34 3725
rect 34 3691 50 3725
rect -50 3583 -34 3617
rect 34 3583 50 3617
rect -96 3533 -62 3549
rect -96 2541 -62 2557
rect 62 3533 96 3549
rect 62 2541 96 2557
rect -50 2473 -34 2507
rect 34 2473 50 2507
rect -50 2365 -34 2399
rect 34 2365 50 2399
rect -96 2315 -62 2331
rect -96 1323 -62 1339
rect 62 2315 96 2331
rect 62 1323 96 1339
rect -50 1255 -34 1289
rect 34 1255 50 1289
rect -50 1147 -34 1181
rect 34 1147 50 1181
rect -96 1097 -62 1113
rect -96 105 -62 121
rect 62 1097 96 1113
rect 62 105 96 121
rect -50 37 -34 71
rect 34 37 50 71
rect -50 -71 -34 -37
rect 34 -71 50 -37
rect -96 -121 -62 -105
rect -96 -1113 -62 -1097
rect 62 -121 96 -105
rect 62 -1113 96 -1097
rect -50 -1181 -34 -1147
rect 34 -1181 50 -1147
rect -50 -1289 -34 -1255
rect 34 -1289 50 -1255
rect -96 -1339 -62 -1323
rect -96 -2331 -62 -2315
rect 62 -1339 96 -1323
rect 62 -2331 96 -2315
rect -50 -2399 -34 -2365
rect 34 -2399 50 -2365
rect -50 -2507 -34 -2473
rect 34 -2507 50 -2473
rect -96 -2557 -62 -2541
rect -96 -3549 -62 -3533
rect 62 -2557 96 -2541
rect 62 -3549 96 -3533
rect -50 -3617 -34 -3583
rect 34 -3617 50 -3583
rect -50 -3725 -34 -3691
rect 34 -3725 50 -3691
rect -96 -3775 -62 -3759
rect -96 -4767 -62 -4751
rect 62 -3775 96 -3759
rect 62 -4767 96 -4751
rect -50 -4835 -34 -4801
rect 34 -4835 50 -4801
rect -50 -4943 -34 -4909
rect 34 -4943 50 -4909
rect -96 -4993 -62 -4977
rect -96 -5985 -62 -5969
rect 62 -4993 96 -4977
rect 62 -5985 96 -5969
rect -50 -6053 -34 -6019
rect 34 -6053 50 -6019
rect -50 -6161 -34 -6127
rect 34 -6161 50 -6127
rect -96 -6211 -62 -6195
rect -96 -7203 -62 -7187
rect 62 -6211 96 -6195
rect 62 -7203 96 -7187
rect -50 -7271 -34 -7237
rect 34 -7271 50 -7237
rect -50 -7379 -34 -7345
rect 34 -7379 50 -7345
rect -96 -7429 -62 -7413
rect -96 -8421 -62 -8405
rect 62 -7429 96 -7413
rect 62 -8421 96 -8405
rect -50 -8489 -34 -8455
rect 34 -8489 50 -8455
rect -50 -8597 -34 -8563
rect 34 -8597 50 -8563
rect -96 -8647 -62 -8631
rect -96 -9639 -62 -9623
rect 62 -8647 96 -8631
rect 62 -9639 96 -9623
rect -50 -9707 -34 -9673
rect 34 -9707 50 -9673
rect -50 -9815 -34 -9781
rect 34 -9815 50 -9781
rect -96 -9865 -62 -9849
rect -96 -10857 -62 -10841
rect 62 -9865 96 -9849
rect 62 -10857 96 -10841
rect -50 -10925 -34 -10891
rect 34 -10925 50 -10891
rect -50 -11033 -34 -10999
rect 34 -11033 50 -10999
rect -96 -11083 -62 -11067
rect -96 -12075 -62 -12059
rect 62 -11083 96 -11067
rect 62 -12075 96 -12059
rect -50 -12143 -34 -12109
rect 34 -12143 50 -12109
<< viali >>
rect -34 12109 34 12143
rect -96 11083 -62 12059
rect 62 11083 96 12059
rect -34 10999 34 11033
rect -34 10891 34 10925
rect -96 9865 -62 10841
rect 62 9865 96 10841
rect -34 9781 34 9815
rect -34 9673 34 9707
rect -96 8647 -62 9623
rect 62 8647 96 9623
rect -34 8563 34 8597
rect -34 8455 34 8489
rect -96 7429 -62 8405
rect 62 7429 96 8405
rect -34 7345 34 7379
rect -34 7237 34 7271
rect -96 6211 -62 7187
rect 62 6211 96 7187
rect -34 6127 34 6161
rect -34 6019 34 6053
rect -96 4993 -62 5969
rect 62 4993 96 5969
rect -34 4909 34 4943
rect -34 4801 34 4835
rect -96 3775 -62 4751
rect 62 3775 96 4751
rect -34 3691 34 3725
rect -34 3583 34 3617
rect -96 2557 -62 3533
rect 62 2557 96 3533
rect -34 2473 34 2507
rect -34 2365 34 2399
rect -96 1339 -62 2315
rect 62 1339 96 2315
rect -34 1255 34 1289
rect -34 1147 34 1181
rect -96 121 -62 1097
rect 62 121 96 1097
rect -34 37 34 71
rect -34 -71 34 -37
rect -96 -1097 -62 -121
rect 62 -1097 96 -121
rect -34 -1181 34 -1147
rect -34 -1289 34 -1255
rect -96 -2315 -62 -1339
rect 62 -2315 96 -1339
rect -34 -2399 34 -2365
rect -34 -2507 34 -2473
rect -96 -3533 -62 -2557
rect 62 -3533 96 -2557
rect -34 -3617 34 -3583
rect -34 -3725 34 -3691
rect -96 -4751 -62 -3775
rect 62 -4751 96 -3775
rect -34 -4835 34 -4801
rect -34 -4943 34 -4909
rect -96 -5969 -62 -4993
rect 62 -5969 96 -4993
rect -34 -6053 34 -6019
rect -34 -6161 34 -6127
rect -96 -7187 -62 -6211
rect 62 -7187 96 -6211
rect -34 -7271 34 -7237
rect -34 -7379 34 -7345
rect -96 -8405 -62 -7429
rect 62 -8405 96 -7429
rect -34 -8489 34 -8455
rect -34 -8597 34 -8563
rect -96 -9623 -62 -8647
rect 62 -9623 96 -8647
rect -34 -9707 34 -9673
rect -34 -9815 34 -9781
rect -96 -10841 -62 -9865
rect 62 -10841 96 -9865
rect -34 -10925 34 -10891
rect -34 -11033 34 -10999
rect -96 -12059 -62 -11083
rect 62 -12059 96 -11083
rect -34 -12143 34 -12109
<< metal1 >>
rect -46 12143 46 12149
rect -46 12109 -34 12143
rect 34 12109 46 12143
rect -46 12103 46 12109
rect -102 12059 -56 12071
rect -102 11083 -96 12059
rect -62 11083 -56 12059
rect -102 11071 -56 11083
rect 56 12059 102 12071
rect 56 11083 62 12059
rect 96 11083 102 12059
rect 56 11071 102 11083
rect -46 11033 46 11039
rect -46 10999 -34 11033
rect 34 10999 46 11033
rect -46 10993 46 10999
rect -46 10925 46 10931
rect -46 10891 -34 10925
rect 34 10891 46 10925
rect -46 10885 46 10891
rect -102 10841 -56 10853
rect -102 9865 -96 10841
rect -62 9865 -56 10841
rect -102 9853 -56 9865
rect 56 10841 102 10853
rect 56 9865 62 10841
rect 96 9865 102 10841
rect 56 9853 102 9865
rect -46 9815 46 9821
rect -46 9781 -34 9815
rect 34 9781 46 9815
rect -46 9775 46 9781
rect -46 9707 46 9713
rect -46 9673 -34 9707
rect 34 9673 46 9707
rect -46 9667 46 9673
rect -102 9623 -56 9635
rect -102 8647 -96 9623
rect -62 8647 -56 9623
rect -102 8635 -56 8647
rect 56 9623 102 9635
rect 56 8647 62 9623
rect 96 8647 102 9623
rect 56 8635 102 8647
rect -46 8597 46 8603
rect -46 8563 -34 8597
rect 34 8563 46 8597
rect -46 8557 46 8563
rect -46 8489 46 8495
rect -46 8455 -34 8489
rect 34 8455 46 8489
rect -46 8449 46 8455
rect -102 8405 -56 8417
rect -102 7429 -96 8405
rect -62 7429 -56 8405
rect -102 7417 -56 7429
rect 56 8405 102 8417
rect 56 7429 62 8405
rect 96 7429 102 8405
rect 56 7417 102 7429
rect -46 7379 46 7385
rect -46 7345 -34 7379
rect 34 7345 46 7379
rect -46 7339 46 7345
rect -46 7271 46 7277
rect -46 7237 -34 7271
rect 34 7237 46 7271
rect -46 7231 46 7237
rect -102 7187 -56 7199
rect -102 6211 -96 7187
rect -62 6211 -56 7187
rect -102 6199 -56 6211
rect 56 7187 102 7199
rect 56 6211 62 7187
rect 96 6211 102 7187
rect 56 6199 102 6211
rect -46 6161 46 6167
rect -46 6127 -34 6161
rect 34 6127 46 6161
rect -46 6121 46 6127
rect -46 6053 46 6059
rect -46 6019 -34 6053
rect 34 6019 46 6053
rect -46 6013 46 6019
rect -102 5969 -56 5981
rect -102 4993 -96 5969
rect -62 4993 -56 5969
rect -102 4981 -56 4993
rect 56 5969 102 5981
rect 56 4993 62 5969
rect 96 4993 102 5969
rect 56 4981 102 4993
rect -46 4943 46 4949
rect -46 4909 -34 4943
rect 34 4909 46 4943
rect -46 4903 46 4909
rect -46 4835 46 4841
rect -46 4801 -34 4835
rect 34 4801 46 4835
rect -46 4795 46 4801
rect -102 4751 -56 4763
rect -102 3775 -96 4751
rect -62 3775 -56 4751
rect -102 3763 -56 3775
rect 56 4751 102 4763
rect 56 3775 62 4751
rect 96 3775 102 4751
rect 56 3763 102 3775
rect -46 3725 46 3731
rect -46 3691 -34 3725
rect 34 3691 46 3725
rect -46 3685 46 3691
rect -46 3617 46 3623
rect -46 3583 -34 3617
rect 34 3583 46 3617
rect -46 3577 46 3583
rect -102 3533 -56 3545
rect -102 2557 -96 3533
rect -62 2557 -56 3533
rect -102 2545 -56 2557
rect 56 3533 102 3545
rect 56 2557 62 3533
rect 96 2557 102 3533
rect 56 2545 102 2557
rect -46 2507 46 2513
rect -46 2473 -34 2507
rect 34 2473 46 2507
rect -46 2467 46 2473
rect -46 2399 46 2405
rect -46 2365 -34 2399
rect 34 2365 46 2399
rect -46 2359 46 2365
rect -102 2315 -56 2327
rect -102 1339 -96 2315
rect -62 1339 -56 2315
rect -102 1327 -56 1339
rect 56 2315 102 2327
rect 56 1339 62 2315
rect 96 1339 102 2315
rect 56 1327 102 1339
rect -46 1289 46 1295
rect -46 1255 -34 1289
rect 34 1255 46 1289
rect -46 1249 46 1255
rect -46 1181 46 1187
rect -46 1147 -34 1181
rect 34 1147 46 1181
rect -46 1141 46 1147
rect -102 1097 -56 1109
rect -102 121 -96 1097
rect -62 121 -56 1097
rect -102 109 -56 121
rect 56 1097 102 1109
rect 56 121 62 1097
rect 96 121 102 1097
rect 56 109 102 121
rect -46 71 46 77
rect -46 37 -34 71
rect 34 37 46 71
rect -46 31 46 37
rect -46 -37 46 -31
rect -46 -71 -34 -37
rect 34 -71 46 -37
rect -46 -77 46 -71
rect -102 -121 -56 -109
rect -102 -1097 -96 -121
rect -62 -1097 -56 -121
rect -102 -1109 -56 -1097
rect 56 -121 102 -109
rect 56 -1097 62 -121
rect 96 -1097 102 -121
rect 56 -1109 102 -1097
rect -46 -1147 46 -1141
rect -46 -1181 -34 -1147
rect 34 -1181 46 -1147
rect -46 -1187 46 -1181
rect -46 -1255 46 -1249
rect -46 -1289 -34 -1255
rect 34 -1289 46 -1255
rect -46 -1295 46 -1289
rect -102 -1339 -56 -1327
rect -102 -2315 -96 -1339
rect -62 -2315 -56 -1339
rect -102 -2327 -56 -2315
rect 56 -1339 102 -1327
rect 56 -2315 62 -1339
rect 96 -2315 102 -1339
rect 56 -2327 102 -2315
rect -46 -2365 46 -2359
rect -46 -2399 -34 -2365
rect 34 -2399 46 -2365
rect -46 -2405 46 -2399
rect -46 -2473 46 -2467
rect -46 -2507 -34 -2473
rect 34 -2507 46 -2473
rect -46 -2513 46 -2507
rect -102 -2557 -56 -2545
rect -102 -3533 -96 -2557
rect -62 -3533 -56 -2557
rect -102 -3545 -56 -3533
rect 56 -2557 102 -2545
rect 56 -3533 62 -2557
rect 96 -3533 102 -2557
rect 56 -3545 102 -3533
rect -46 -3583 46 -3577
rect -46 -3617 -34 -3583
rect 34 -3617 46 -3583
rect -46 -3623 46 -3617
rect -46 -3691 46 -3685
rect -46 -3725 -34 -3691
rect 34 -3725 46 -3691
rect -46 -3731 46 -3725
rect -102 -3775 -56 -3763
rect -102 -4751 -96 -3775
rect -62 -4751 -56 -3775
rect -102 -4763 -56 -4751
rect 56 -3775 102 -3763
rect 56 -4751 62 -3775
rect 96 -4751 102 -3775
rect 56 -4763 102 -4751
rect -46 -4801 46 -4795
rect -46 -4835 -34 -4801
rect 34 -4835 46 -4801
rect -46 -4841 46 -4835
rect -46 -4909 46 -4903
rect -46 -4943 -34 -4909
rect 34 -4943 46 -4909
rect -46 -4949 46 -4943
rect -102 -4993 -56 -4981
rect -102 -5969 -96 -4993
rect -62 -5969 -56 -4993
rect -102 -5981 -56 -5969
rect 56 -4993 102 -4981
rect 56 -5969 62 -4993
rect 96 -5969 102 -4993
rect 56 -5981 102 -5969
rect -46 -6019 46 -6013
rect -46 -6053 -34 -6019
rect 34 -6053 46 -6019
rect -46 -6059 46 -6053
rect -46 -6127 46 -6121
rect -46 -6161 -34 -6127
rect 34 -6161 46 -6127
rect -46 -6167 46 -6161
rect -102 -6211 -56 -6199
rect -102 -7187 -96 -6211
rect -62 -7187 -56 -6211
rect -102 -7199 -56 -7187
rect 56 -6211 102 -6199
rect 56 -7187 62 -6211
rect 96 -7187 102 -6211
rect 56 -7199 102 -7187
rect -46 -7237 46 -7231
rect -46 -7271 -34 -7237
rect 34 -7271 46 -7237
rect -46 -7277 46 -7271
rect -46 -7345 46 -7339
rect -46 -7379 -34 -7345
rect 34 -7379 46 -7345
rect -46 -7385 46 -7379
rect -102 -7429 -56 -7417
rect -102 -8405 -96 -7429
rect -62 -8405 -56 -7429
rect -102 -8417 -56 -8405
rect 56 -7429 102 -7417
rect 56 -8405 62 -7429
rect 96 -8405 102 -7429
rect 56 -8417 102 -8405
rect -46 -8455 46 -8449
rect -46 -8489 -34 -8455
rect 34 -8489 46 -8455
rect -46 -8495 46 -8489
rect -46 -8563 46 -8557
rect -46 -8597 -34 -8563
rect 34 -8597 46 -8563
rect -46 -8603 46 -8597
rect -102 -8647 -56 -8635
rect -102 -9623 -96 -8647
rect -62 -9623 -56 -8647
rect -102 -9635 -56 -9623
rect 56 -8647 102 -8635
rect 56 -9623 62 -8647
rect 96 -9623 102 -8647
rect 56 -9635 102 -9623
rect -46 -9673 46 -9667
rect -46 -9707 -34 -9673
rect 34 -9707 46 -9673
rect -46 -9713 46 -9707
rect -46 -9781 46 -9775
rect -46 -9815 -34 -9781
rect 34 -9815 46 -9781
rect -46 -9821 46 -9815
rect -102 -9865 -56 -9853
rect -102 -10841 -96 -9865
rect -62 -10841 -56 -9865
rect -102 -10853 -56 -10841
rect 56 -9865 102 -9853
rect 56 -10841 62 -9865
rect 96 -10841 102 -9865
rect 56 -10853 102 -10841
rect -46 -10891 46 -10885
rect -46 -10925 -34 -10891
rect 34 -10925 46 -10891
rect -46 -10931 46 -10925
rect -46 -10999 46 -10993
rect -46 -11033 -34 -10999
rect 34 -11033 46 -10999
rect -46 -11039 46 -11033
rect -102 -11083 -56 -11071
rect -102 -12059 -96 -11083
rect -62 -12059 -56 -11083
rect -102 -12071 -56 -12059
rect 56 -11083 102 -11071
rect 56 -12059 62 -11083
rect 96 -12059 102 -11083
rect 56 -12071 102 -12059
rect -46 -12109 46 -12103
rect -46 -12143 -34 -12109
rect 34 -12143 46 -12109
rect -46 -12149 46 -12143
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 20 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
