magic
tech sky130A
magscale 1 2
timestamp 1666901446
<< error_p >>
rect -29 845 29 851
rect -29 811 -17 845
rect -29 805 29 811
<< nwell >>
rect -109 -898 109 864
<< pmos >>
rect -15 -836 15 764
<< pdiff >>
rect -73 752 -15 764
rect -73 -824 -61 752
rect -27 -824 -15 752
rect -73 -836 -15 -824
rect 15 752 73 764
rect 15 -824 27 752
rect 61 -824 73 752
rect 15 -836 73 -824
<< pdiffc >>
rect -61 -824 -27 752
rect 27 -824 61 752
<< poly >>
rect -33 845 33 861
rect -33 811 -17 845
rect 17 811 33 845
rect -33 795 33 811
rect -15 764 15 795
rect -15 -862 15 -836
<< polycont >>
rect -17 811 17 845
<< locali >>
rect -33 811 -17 845
rect 17 811 33 845
rect -61 752 -27 768
rect -61 -840 -27 -824
rect 27 752 61 768
rect 27 -840 61 -824
<< viali >>
rect -17 811 17 845
rect -61 -824 -27 752
rect 27 -824 61 752
<< metal1 >>
rect -29 845 29 851
rect -29 811 -17 845
rect 17 811 29 845
rect -29 805 29 811
rect -67 752 -21 764
rect -67 -824 -61 752
rect -27 -824 -21 752
rect -67 -836 -21 -824
rect 21 752 67 764
rect 21 -824 27 752
rect 61 -824 67 752
rect 21 -836 67 -824
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
