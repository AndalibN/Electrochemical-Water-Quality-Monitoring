magic
tech sky130A
magscale 1 2
timestamp 1667402611
<< nwell >>
rect 5406 5880 7632 5882
rect 8288 5880 10228 5882
rect 474 5674 10228 5880
rect 472 5256 10228 5674
rect 472 5248 10230 5256
rect 474 5208 10230 5248
rect 474 5204 2060 5208
rect 3012 5204 10230 5208
rect 474 5194 10230 5204
rect 474 5156 1062 5194
rect 474 5116 1060 5156
rect 520 5034 560 5102
rect 1320 2174 1708 5194
rect 1966 5168 10230 5194
rect 1966 5166 3012 5168
rect 3314 5166 10230 5168
rect 4356 5162 10230 5166
rect 5406 5134 10230 5162
rect 7596 5118 10230 5134
rect 7596 5112 9582 5118
rect 7870 4622 8256 5112
rect 8540 5108 9582 5112
rect 8540 4738 8932 5108
rect 9196 4776 9582 5108
rect 9196 4520 9584 4776
rect 9840 4220 10230 5118
<< nbase >>
rect 2060 5204 3012 5208
<< psubdiff >>
rect 6910 -3598 9628 -3596
rect 13264 -3598 13664 -3596
rect 6910 -3600 10504 -3598
rect 11476 -3600 14238 -3598
rect -1886 -3634 14238 -3600
rect -1886 -3636 11314 -3634
rect -1886 -3838 -1856 -3636
rect -1616 -3646 11314 -3636
rect -1616 -3654 2012 -3646
rect -1616 -3824 -842 -3654
rect -530 -3824 2012 -3654
rect -1616 -3832 2012 -3824
rect 2332 -3648 7540 -3646
rect 2332 -3832 2388 -3648
rect -1616 -3838 2388 -3832
rect -1886 -3840 2388 -3838
rect 2736 -3654 7540 -3648
rect 2736 -3834 6022 -3654
rect 6284 -3834 6426 -3654
rect 2736 -3838 6426 -3834
rect 6698 -3834 6742 -3654
rect 7146 -3834 7540 -3654
rect 6698 -3838 7540 -3834
rect 2736 -3840 7540 -3838
rect -1886 -3842 7540 -3840
rect 8038 -3652 11314 -3646
rect 8038 -3834 9656 -3652
rect 10398 -3834 11314 -3652
rect 11736 -3642 14238 -3634
rect 11736 -3646 13838 -3642
rect 11736 -3834 13030 -3646
rect 13442 -3834 13838 -3646
rect 14164 -3834 14238 -3642
rect 8038 -3842 14238 -3834
rect -1886 -3860 14238 -3842
rect -1886 -3862 -876 -3860
<< nsubdiff >>
rect 2936 5790 10190 5792
rect 510 5746 10190 5790
rect 510 5730 5306 5746
rect 510 5520 520 5730
rect 970 5716 5306 5730
rect 970 5532 2262 5716
rect 2706 5714 5306 5716
rect 2706 5532 3598 5714
rect 970 5528 3598 5532
rect 4050 5528 5306 5714
rect 970 5520 5306 5528
rect 510 5512 5306 5520
rect 5736 5742 10190 5746
rect 5736 5740 9168 5742
rect 5736 5738 7852 5740
rect 5736 5512 7132 5738
rect 510 5504 7132 5512
rect 7562 5504 7852 5738
rect 510 5500 7852 5504
rect 8180 5500 8464 5740
rect 8810 5508 9168 5740
rect 9468 5508 9858 5742
rect 8810 5506 9858 5508
rect 10162 5506 10190 5742
rect 8810 5500 10190 5506
rect 510 5460 10190 5500
rect 2936 5458 4300 5460
rect 7580 5458 10190 5460
<< psubdiffcont >>
rect -1856 -3838 -1616 -3636
rect -842 -3824 -530 -3654
rect 2012 -3832 2332 -3646
rect 2388 -3840 2736 -3648
rect 6022 -3834 6284 -3654
rect 6426 -3838 6698 -3654
rect 6742 -3834 7146 -3654
rect 7540 -3842 8038 -3646
rect 9656 -3834 10398 -3652
rect 11314 -3834 11736 -3634
rect 13030 -3834 13442 -3646
rect 13838 -3834 14164 -3642
<< nsubdiffcont >>
rect 520 5520 970 5730
rect 2262 5532 2706 5716
rect 3598 5528 4050 5714
rect 5306 5512 5736 5746
rect 7132 5504 7562 5738
rect 7852 5500 8180 5740
rect 8464 5500 8810 5740
rect 9168 5508 9468 5742
rect 9858 5506 10162 5742
<< locali >>
rect 520 5746 10180 5760
rect 520 5730 5306 5746
rect 970 5716 5306 5730
rect 970 5532 2262 5716
rect 2706 5714 5306 5716
rect 2706 5532 3598 5714
rect 970 5528 3598 5532
rect 4050 5528 5306 5714
rect 970 5520 5306 5528
rect 520 5512 5306 5520
rect 5736 5742 10180 5746
rect 5736 5740 9168 5742
rect 5736 5738 7852 5740
rect 5736 5512 7132 5738
rect 520 5504 7132 5512
rect 7562 5504 7852 5738
rect 520 5500 7852 5504
rect 8180 5500 8464 5740
rect 8810 5508 9168 5740
rect 9468 5508 9858 5742
rect 8810 5506 9858 5508
rect 10162 5506 10180 5742
rect 8810 5500 10180 5506
rect 520 5490 10180 5500
rect 520 5460 560 5490
rect 522 5202 560 5460
rect 2470 5220 2508 5490
rect 522 5098 558 5202
rect 2472 5086 2506 5220
rect 3820 5204 3858 5490
rect 5452 5228 5490 5490
rect 5676 5488 7564 5490
rect 3820 5108 3854 5204
rect 5456 5082 5490 5228
rect 7514 5230 7552 5488
rect 7912 5456 7952 5490
rect 7912 5256 7950 5456
rect 7514 5084 7548 5230
rect 7912 5224 7952 5256
rect -1140 4706 -520 4774
rect -574 4186 -520 4706
rect 7914 4530 7952 5224
rect 8590 5216 8628 5490
rect 9240 5218 9278 5490
rect 9886 5222 9924 5490
rect 8590 4650 8626 5216
rect 9242 4446 9278 5218
rect 9244 4440 9278 4446
rect 9276 4434 9278 4440
rect 9888 4130 9924 5222
rect 4312 3102 4662 3152
rect 4910 3102 5280 3150
rect 4312 3100 4608 3102
rect 5230 2750 5280 3102
rect 10168 3090 10192 3130
rect 7468 2998 7996 3034
rect 8130 2996 8672 3034
rect 8836 2998 9290 3032
rect 9460 2996 9968 3032
rect 10290 2998 10472 3042
rect 5230 2692 8186 2750
rect 5230 2538 5280 2692
rect 8140 2528 8186 2692
rect 10290 2586 10340 2998
rect 9324 2518 10340 2586
rect 1242 2120 1430 2156
rect -2190 -1660 -2152 1302
rect 1242 1152 1276 2120
rect 6520 1872 6560 2372
rect 6520 1432 6562 1872
rect 3390 1190 3392 1200
rect 1014 1118 1276 1152
rect 1660 1146 2014 1182
rect 968 1012 1372 1048
rect 1920 730 1960 1146
rect 3220 1116 3362 1190
rect 3364 1120 3392 1190
rect 2710 1056 3460 1058
rect 2710 1024 3408 1056
rect 2240 950 2310 1024
rect 3980 950 4040 1024
rect 2240 880 4040 950
rect 4470 844 4544 1140
rect 3220 766 4544 844
rect 1920 690 3510 730
rect 3460 636 3510 690
rect 5000 660 5038 1040
rect 3930 608 5038 660
rect -864 270 -828 466
rect -2190 -1698 -1734 -1660
rect -2190 -1700 -2152 -1698
rect -1802 -2500 -1734 -1698
rect -788 -1874 -744 194
rect 1234 28 1268 454
rect 1630 410 1660 506
rect 3320 490 3354 580
rect 3930 400 3980 608
rect 3814 350 4066 400
rect 1234 -6 1430 28
rect -1800 -3622 -1732 -2500
rect -788 -2512 -742 -1874
rect 2104 -1876 2164 -140
rect 2104 -1880 2168 -1876
rect 6120 -1880 6156 -1404
rect 6520 -1880 6560 1432
rect 6796 -1880 6864 1556
rect 7652 1298 7732 1580
rect 7644 448 7724 730
rect 7642 -400 7722 -118
rect 2106 -2494 2168 -1880
rect -1876 -3624 -872 -3622
rect -788 -3624 -740 -2512
rect 2106 -3624 2170 -2494
rect 6122 -2500 6156 -1880
rect 6522 -2500 6558 -1880
rect 6798 -2500 6864 -1880
rect 7638 -2496 7724 -980
rect 7640 -2500 7724 -2496
rect 6122 -2558 6158 -2500
rect 6120 -3624 6160 -2558
rect 6522 -3624 6562 -2500
rect 6798 -3624 6866 -2500
rect 7640 -3624 7726 -2500
rect 9380 -2680 9420 -1448
rect 8964 -2736 9420 -2680
rect 8958 -3108 9846 -3052
rect 9782 -3544 9846 -3108
rect 10200 -3442 10468 -3396
rect 9782 -3622 9844 -3544
rect 10200 -3546 10258 -3442
rect 10200 -3622 10256 -3546
rect 11462 -3622 11520 -416
rect 11610 -1960 12210 -1956
rect 12428 -1960 12486 -136
rect 13390 -1932 13448 -574
rect 14172 -1580 14238 -706
rect 13954 -1660 14238 -1580
rect 11610 -2010 12486 -1960
rect 13184 -1984 13448 -1932
rect 13390 -1986 13448 -1984
rect 11610 -2012 12210 -2010
rect 11610 -3622 11676 -2012
rect 13132 -2472 13188 -2108
rect 13132 -3622 13186 -2472
rect 13922 -3622 13970 -1968
rect 9598 -3624 10504 -3622
rect 11462 -3624 11958 -3622
rect 12400 -3624 14238 -3622
rect -1876 -3634 14238 -3624
rect -1876 -3636 11314 -3634
rect -1876 -3838 -1856 -3636
rect -1616 -3646 11314 -3636
rect -1616 -3654 2012 -3646
rect -1616 -3824 -842 -3654
rect -530 -3824 2012 -3654
rect -1616 -3832 2012 -3824
rect 2332 -3648 7540 -3646
rect 2332 -3832 2388 -3648
rect -1616 -3838 2388 -3832
rect -1876 -3840 2388 -3838
rect 2736 -3654 7540 -3648
rect 2736 -3834 6022 -3654
rect 6284 -3834 6426 -3654
rect 2736 -3838 6426 -3834
rect 6698 -3834 6742 -3654
rect 7146 -3834 7540 -3654
rect 6698 -3838 7540 -3834
rect 2736 -3840 7540 -3838
rect -1876 -3842 7540 -3840
rect 8038 -3652 11314 -3646
rect 8038 -3834 9656 -3652
rect 10398 -3834 11314 -3652
rect 11736 -3642 14238 -3634
rect 11736 -3646 13838 -3642
rect 11736 -3834 13030 -3646
rect 13442 -3834 13838 -3646
rect 14164 -3834 14238 -3642
rect 8038 -3842 14238 -3834
rect -1876 -3850 14238 -3842
rect -1876 -3852 -872 -3850
<< metal1 >>
rect 520 5460 560 5730
rect 2472 5516 2506 5716
rect 522 5202 560 5460
rect 2470 5220 2508 5516
rect 3820 5500 3854 5714
rect 5456 5524 5490 5746
rect 522 5070 558 5202
rect 2472 5086 2506 5220
rect 3820 5204 3858 5500
rect 5452 5228 5490 5524
rect 3820 5044 3854 5204
rect 5456 5080 5490 5228
rect 7514 5526 7548 5738
rect 7514 5230 7552 5526
rect 7914 5520 7952 5738
rect 7912 5456 7952 5520
rect 8590 5512 8626 5738
rect 9242 5514 9278 5742
rect 9888 5518 9924 5738
rect 7912 5256 7950 5456
rect 7514 5080 7548 5230
rect 7912 5224 7952 5256
rect -1140 4706 -520 4774
rect -574 4186 -520 4706
rect 7914 4530 7952 5224
rect 8590 5216 8628 5512
rect 9240 5218 9278 5514
rect 9886 5222 9924 5518
rect 8590 4650 8626 5216
rect 9242 4446 9278 5218
rect 9244 4440 9278 4446
rect 9276 4434 9278 4440
rect 9888 4130 9924 5222
rect 4312 3102 4662 3152
rect 8166 3150 8230 3170
rect 4910 3102 5280 3150
rect 4312 3100 4608 3102
rect -580 3040 -510 3046
rect -580 2976 -570 3040
rect -518 2976 -510 3040
rect -580 2966 -510 2976
rect 4278 2882 4312 2930
rect 5230 2750 5280 3102
rect 8166 3098 8172 3150
rect 8224 3098 8230 3150
rect 8166 3092 8230 3098
rect 8840 3152 8900 3158
rect 8840 3100 8848 3152
rect 8840 3090 8900 3100
rect 9492 3152 9552 3160
rect 9492 3100 9500 3152
rect 9492 3090 9552 3100
rect 10136 3142 10202 3144
rect 10136 3090 10144 3142
rect 10196 3090 10202 3142
rect 10136 3080 10202 3090
rect 5610 3052 5680 3060
rect 5610 3000 5620 3052
rect 5672 3000 5680 3052
rect 5610 2990 5680 3000
rect 7468 2998 7996 3034
rect 8130 2996 8672 3034
rect 8802 2998 9320 3032
rect 9460 2996 9968 3032
rect 10290 2998 10472 3042
rect 5230 2692 8186 2750
rect 5230 2538 5280 2692
rect 7550 2592 7620 2600
rect 7550 2536 7558 2592
rect 7610 2536 7620 2592
rect 7550 2530 7620 2536
rect 8140 2528 8186 2692
rect 10290 2586 10340 2998
rect 9324 2518 10340 2586
rect 1242 2120 1598 2156
rect -2190 -1660 -2152 1302
rect 1242 1152 1276 2120
rect 6520 1872 6560 2372
rect 6520 1432 6562 1872
rect 8900 1632 8992 1660
rect 3390 1190 3392 1200
rect 980 1118 1276 1152
rect 1626 1146 2048 1184
rect 3220 1180 3362 1190
rect 584 1014 1406 1048
rect 1368 1010 1402 1014
rect 1362 934 1408 950
rect 1362 928 1420 934
rect 1414 876 1420 928
rect 1362 842 1408 876
rect 1920 730 1960 1146
rect 3220 1128 3230 1180
rect 3300 1128 3362 1180
rect 3220 1116 3362 1128
rect 3364 1120 3392 1190
rect 3570 1074 3670 1080
rect 2240 1054 2320 1056
rect 2240 950 2310 1054
rect 2706 1024 3468 1058
rect 3570 1016 3584 1074
rect 3656 1016 3670 1074
rect 4152 1072 4240 1078
rect 3570 1010 3670 1016
rect 3580 1008 3662 1010
rect 3980 950 4040 1052
rect 4152 1020 4166 1072
rect 4222 1020 4240 1072
rect 4152 1008 4240 1020
rect 2240 942 4040 950
rect 2240 890 2250 942
rect 2310 890 4040 942
rect 2240 880 4040 890
rect 4470 844 4544 1140
rect 3220 836 4544 844
rect 3220 774 3234 836
rect 3306 774 4544 836
rect 3220 766 4544 774
rect 1618 712 1680 720
rect 1618 660 1626 712
rect 1678 660 1680 712
rect 1920 690 3510 730
rect 1618 652 1680 660
rect 3460 636 3510 690
rect 5000 660 5038 1040
rect 3930 608 5038 660
rect 3320 550 3354 580
rect 3300 542 3368 550
rect -864 270 -828 466
rect -746 226 -744 228
rect -2190 -1698 -1734 -1660
rect -2190 -1700 -2152 -1698
rect -1802 -2500 -1734 -1698
rect -788 -1874 -744 226
rect 1234 28 1268 454
rect 1630 410 1660 506
rect 3300 490 3310 542
rect 3362 490 3368 542
rect 3300 482 3368 490
rect 3782 482 3814 522
rect 3930 400 3980 608
rect 4150 512 4252 514
rect 4150 460 4168 512
rect 4240 460 4252 512
rect 4150 450 4252 460
rect 3814 350 4066 400
rect 1616 180 1690 192
rect 1616 110 1624 180
rect 1676 110 1690 180
rect 1616 88 1690 110
rect 1234 -6 1430 28
rect -1800 -3836 -1732 -2500
rect -788 -2512 -742 -1874
rect 2104 -1876 2164 -140
rect 2104 -1880 2168 -1876
rect 6120 -1880 6156 -1404
rect 6520 -1880 6560 1432
rect 6796 -1880 6864 1556
rect 7652 1298 7732 1580
rect 8900 1560 8920 1632
rect 8972 1560 8992 1632
rect 8900 1542 8992 1560
rect 12158 1322 12278 1334
rect 12158 1238 12170 1322
rect 12258 1238 12278 1322
rect 12158 1230 12176 1238
rect 12244 1230 12278 1238
rect 12158 1216 12278 1230
rect 13110 894 13216 898
rect 13104 892 13216 894
rect 13104 820 13118 892
rect 13110 812 13118 820
rect 13206 812 13216 892
rect 13110 804 13216 812
rect 7644 448 7724 730
rect 13900 724 13988 726
rect 13900 670 13910 724
rect 13980 670 13988 724
rect 13900 664 13988 670
rect 7642 -400 7722 -118
rect 2106 -2494 2168 -1880
rect -788 -3726 -740 -2512
rect 2106 -3822 2170 -2494
rect 6122 -2500 6156 -1880
rect 6522 -2500 6558 -1880
rect 6798 -2500 6864 -1880
rect 7638 -2496 7724 -980
rect 7640 -2500 7724 -2496
rect 6122 -2558 6158 -2500
rect 2490 -3732 2632 -3696
rect 2490 -3814 2522 -3732
rect 2584 -3814 2632 -3732
rect 6120 -3744 6160 -2558
rect 2490 -3832 2632 -3814
rect 6522 -3834 6562 -2500
rect 6798 -3784 6866 -2500
rect 6934 -3676 7076 -3654
rect 6934 -3758 6966 -3676
rect 7028 -3758 7076 -3676
rect 6934 -3776 7076 -3758
rect 7640 -3826 7726 -2500
rect 9380 -2680 9420 -1448
rect 8964 -2736 9420 -2680
rect 8958 -3108 9846 -3052
rect 9782 -3544 9846 -3108
rect 10200 -3442 10468 -3396
rect 7766 -3712 7904 -3690
rect 7766 -3794 7798 -3712
rect 7860 -3794 7904 -3712
rect 9782 -3778 9844 -3544
rect 10200 -3546 10258 -3442
rect 7766 -3812 7904 -3794
rect 10200 -3808 10256 -3546
rect 11462 -3766 11520 -416
rect 11610 -1960 12210 -1956
rect 12428 -1960 12486 -136
rect 13390 -1932 13448 -574
rect 14172 -1580 14238 -706
rect 13954 -1660 14238 -1580
rect 11610 -2010 12486 -1960
rect 13184 -1984 13448 -1932
rect 13390 -1986 13448 -1984
rect 11610 -2012 12210 -2010
rect 11610 -3776 11676 -2012
rect 13132 -2472 13188 -2108
rect 13132 -3814 13186 -2472
rect 13922 -3814 13970 -1968
<< via1 >>
rect -570 2976 -518 3040
rect 8172 3098 8224 3150
rect 8848 3100 8900 3152
rect 9500 3100 9552 3152
rect 10144 3090 10196 3142
rect 5620 3000 5672 3052
rect 7558 2536 7610 2592
rect 7114 1806 7218 1912
rect 7960 1808 8058 1914
rect 1362 876 1414 928
rect 3230 1128 3300 1180
rect 3584 1016 3656 1074
rect 4166 1020 4222 1072
rect 2250 890 2310 942
rect 3234 774 3306 836
rect 1626 660 1678 712
rect 3310 490 3362 542
rect 4168 460 4240 512
rect 1624 110 1676 180
rect 2334 94 2434 190
rect 8920 1560 8972 1632
rect 12170 1238 12258 1322
rect 12176 1230 12244 1238
rect 7108 958 7210 1060
rect 7954 962 8052 1068
rect 13118 812 13206 892
rect 13910 670 13980 724
rect 7108 106 7210 208
rect 7954 106 8052 212
rect 7112 -734 7214 -632
rect 7954 -732 8056 -630
rect 2522 -3814 2584 -3732
rect 6966 -3758 7028 -3676
rect 7798 -3794 7860 -3712
<< metal2 >>
rect 8164 3150 8330 3160
rect 8164 3098 8172 3150
rect 8224 3098 8330 3150
rect 8164 3092 8330 3098
rect 5610 3052 5680 3060
rect -580 3040 -510 3050
rect -580 2976 -570 3040
rect -518 2976 -510 3040
rect -580 722 -510 2976
rect 5610 3000 5620 3052
rect 5672 3000 5680 3052
rect 5610 2920 5680 3000
rect 4382 2880 5680 2920
rect 3220 1180 3310 1190
rect 2966 1102 3120 1180
rect 3050 950 3120 1102
rect 1362 948 3120 950
rect 3220 1128 3230 1180
rect 3300 1128 3310 1180
rect 1362 942 3122 948
rect 1362 928 2250 942
rect 1414 890 2250 928
rect 2310 890 3122 942
rect 1414 876 3122 890
rect 1362 846 3122 876
rect 1362 842 3050 846
rect -580 712 1682 722
rect -580 660 1626 712
rect 1678 660 1682 712
rect -580 650 1682 660
rect 3220 926 3310 1128
rect 3560 1074 3680 1090
rect 3560 1016 3584 1074
rect 3656 1016 3680 1074
rect 3220 836 3312 926
rect 3220 774 3234 836
rect 3306 774 3312 836
rect 3220 766 3312 774
rect 3560 800 3680 1016
rect 4150 1072 4240 1078
rect 4150 1020 4166 1072
rect 4222 1020 4240 1072
rect 4150 970 4240 1020
rect 4382 970 4420 2880
rect 7550 2592 7630 2600
rect 7550 2536 7558 2592
rect 7610 2536 7630 2592
rect 7550 2400 7630 2536
rect 7102 2350 7630 2400
rect 8290 2424 8330 3092
rect 8840 3152 9030 3160
rect 8840 3100 8848 3152
rect 8900 3100 9030 3152
rect 8840 3090 9030 3100
rect 9492 3152 9680 3160
rect 9492 3100 9500 3152
rect 9552 3100 9680 3152
rect 10286 3150 10390 3152
rect 9492 3090 9680 3100
rect 8990 2770 9030 3090
rect 9640 2900 9680 3090
rect 10136 3142 10390 3150
rect 10136 3090 10144 3142
rect 10196 3090 10390 3142
rect 10136 3080 10390 3090
rect 9640 2860 10160 2900
rect 8990 2730 10020 2770
rect 8290 2382 8650 2424
rect 7102 1920 7222 2350
rect 8574 2156 8650 2382
rect 8574 2054 9012 2156
rect 8570 2052 9012 2054
rect 8570 2038 8690 2052
rect 8570 1956 8582 2038
rect 8670 1956 8690 2038
rect 8570 1934 8690 1956
rect 7102 1912 7226 1920
rect 7102 1806 7114 1912
rect 7218 1806 7226 1912
rect 7102 1798 7226 1806
rect 4150 930 4420 970
rect 7100 1796 7226 1798
rect 7942 1914 8072 1926
rect 7942 1808 7960 1914
rect 8058 1808 8072 1914
rect 7100 1060 7224 1796
rect 7100 958 7108 1060
rect 7210 958 7224 1060
rect 7100 942 7224 958
rect 3560 740 4260 800
rect 3926 738 4260 740
rect 3120 542 3368 550
rect 3120 490 3310 542
rect 3362 490 3368 542
rect 3120 480 3368 490
rect 4150 512 4260 738
rect 4150 460 4168 512
rect 4240 460 4260 512
rect 4150 450 4260 460
rect 7102 208 7224 942
rect 2322 190 2444 198
rect 1616 180 2334 190
rect 1616 110 1624 180
rect 1676 110 2334 180
rect 1616 94 2334 110
rect 2434 94 2444 190
rect 1616 88 2444 94
rect 2322 80 2444 88
rect 7102 106 7108 208
rect 7210 106 7224 208
rect 7102 -616 7224 106
rect 7942 1068 8072 1808
rect 8890 1632 9012 2052
rect 8890 1560 8920 1632
rect 8972 1560 9012 1632
rect 8890 1542 9012 1560
rect 9980 1262 10020 2730
rect 10120 1452 10160 2860
rect 10346 1570 10390 3080
rect 10346 1530 13610 1570
rect 10346 1528 10390 1530
rect 12328 1452 12872 1454
rect 10120 1408 12872 1452
rect 10120 1406 10160 1408
rect 12158 1322 12278 1334
rect 12158 1262 12170 1322
rect 9980 1238 12170 1262
rect 12258 1238 12278 1322
rect 9980 1230 12176 1238
rect 12244 1230 12278 1238
rect 9980 1220 12278 1230
rect 12158 1216 12278 1220
rect 7942 962 7954 1068
rect 8052 962 8072 1068
rect 7942 212 8072 962
rect 12778 1210 12872 1408
rect 12778 922 12870 1210
rect 12778 900 13198 922
rect 12778 892 13220 900
rect 12778 832 13118 892
rect 13102 810 13118 832
rect 13206 810 13220 892
rect 13106 788 13220 810
rect 13500 752 13610 1530
rect 13890 752 14000 754
rect 13500 744 14002 752
rect 13500 662 13900 744
rect 13988 662 14002 744
rect 13500 644 14002 662
rect 13888 642 14002 644
rect 7942 106 7954 212
rect 8052 106 8072 212
rect 7942 -616 8072 106
rect 7100 -630 8072 -616
rect 7100 -632 7954 -630
rect 7100 -734 7112 -632
rect 7214 -732 7954 -632
rect 8056 -732 8072 -630
rect 7214 -734 8072 -732
rect 7100 -750 8072 -734
rect 6952 -3676 7038 -3666
rect 2508 -3732 2594 -3722
rect 2508 -3814 2522 -3732
rect 2584 -3814 2594 -3732
rect 6952 -3758 6966 -3676
rect 7028 -3758 7038 -3676
rect 6952 -3768 7038 -3758
rect 7784 -3712 7870 -3702
rect 7784 -3794 7798 -3712
rect 7860 -3794 7870 -3712
rect 7784 -3804 7870 -3794
rect 2508 -3824 2594 -3814
<< rmetal2 >>
rect 3050 550 3122 846
rect 3050 480 3120 550
<< via2 >>
rect 8582 1956 8670 2038
rect 12170 1238 12258 1320
rect 13118 812 13206 892
rect 13118 810 13206 812
rect 13900 724 13988 744
rect 13900 670 13910 724
rect 13910 670 13980 724
rect 13980 670 13988 724
rect 13900 662 13988 670
rect 2522 -3814 2582 -3732
rect 6966 -3758 7026 -3676
rect 7798 -3794 7858 -3712
<< metal3 >>
rect 8572 2040 8684 2046
rect 8572 1956 8582 2040
rect 8670 1956 8684 2040
rect 8572 1944 8684 1956
rect 12160 1322 12272 1328
rect 12160 1238 12170 1322
rect 12258 1238 12272 1322
rect 12160 1226 12272 1238
rect 13108 894 13220 900
rect 13108 810 13118 894
rect 13206 810 13220 894
rect 13108 798 13220 810
rect 13890 746 14002 752
rect 13890 662 13900 746
rect 13988 662 14002 746
rect 13890 650 14002 662
rect 6946 -3676 7044 -3664
rect 2502 -3732 2600 -3720
rect 2502 -3814 2522 -3732
rect 2582 -3814 2600 -3732
rect 6946 -3758 6966 -3676
rect 7026 -3758 7044 -3676
rect 6946 -3766 7044 -3758
rect 7778 -3712 7876 -3700
rect 7778 -3794 7798 -3712
rect 7858 -3794 7876 -3712
rect 7778 -3802 7876 -3794
rect 2502 -3822 2600 -3814
<< via3 >>
rect 8582 2038 8670 2040
rect 8582 1956 8670 2038
rect 12170 1320 12258 1322
rect 12170 1238 12258 1320
rect 13118 892 13206 894
rect 13118 810 13206 892
rect 13900 744 13988 746
rect 13900 662 13988 744
<< metal4 >>
rect 8572 2040 8684 2046
rect 8572 1956 8582 2040
rect 8670 1956 8684 2040
rect 8572 1948 8684 1956
rect 8570 1858 8684 1948
rect 13978 1858 14200 2120
rect 8570 1798 14200 1858
rect 6962 254 7030 1716
rect 7812 1164 7872 1720
rect 14280 1328 14530 1612
rect 12158 1322 14530 1328
rect 12158 1238 12170 1322
rect 12258 1238 14530 1322
rect 12158 1216 14530 1238
rect 14970 920 15220 1244
rect 13106 894 15220 920
rect 7806 306 7866 862
rect 13106 810 13118 894
rect 13206 860 15220 894
rect 13206 858 13810 860
rect 13206 810 13220 858
rect 13106 788 13220 810
rect 13888 746 14002 752
rect 13888 662 13900 746
rect 13988 702 14002 746
rect 15462 702 15700 956
rect 13988 662 15700 702
rect 13888 642 15700 662
rect 6960 252 7030 254
rect 2510 -640 2592 2
rect 2508 -1278 2590 -640
rect 2506 -2500 2592 -1278
rect 6960 -2500 7028 252
rect 7806 -538 7866 18
rect 7800 -1254 7864 -824
rect 7800 -1876 7866 -1254
rect 2508 -3824 2594 -2500
rect 6960 -2506 7030 -2500
rect 7800 -2506 7868 -1876
rect 6962 -3654 7030 -2506
rect 7802 -2546 7868 -2506
rect 7802 -3594 7870 -2546
rect 6952 -3768 7038 -3654
rect 7802 -3684 7868 -3594
rect 7802 -3686 7870 -3684
rect 7794 -3690 7870 -3686
rect 7784 -3804 7870 -3690
use 298k  R1
timestamp 1666627716
transform 1 0 6899 0 1 335
box 0 0 1 1
use 52k  R2
timestamp 1666627716
transform 1 0 6895 0 1 335
box 0 0 1 1
use 485k  R3
timestamp 1666627716
transform 1 0 6896 0 1 335
box 0 0 1 1
use 520k  R4
timestamp 1666627716
transform 1 0 6897 0 1 335
box 0 0 1 1
use 520k  R5
timestamp 1666627716
transform 1 0 6898 0 1 335
box 0 0 1 1
use 295k  R6
timestamp 1666627716
transform 1 0 8517 0 1 176
box 0 0 1 1
use 298k  R7
timestamp 1666627716
transform 1 0 8518 0 1 176
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_C6T788  XM6
timestamp 1666968066
transform 1 0 6502 0 1 4044
box -1094 -1064 1094 1098
use sky130_fd_pr__pfet_01v8_E8XWE6  XM7
timestamp 1666896002
transform 1 0 4066 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__nfet_01v8_VYYYB6  XM8
timestamp 1666901352
transform 1 0 3568 0 1 -387
box -258 -1057 258 1057
use sky130_fd_pr__nfet_01v8_VJC34T  XM10
timestamp 1666903823
transform 1 0 5110 0 1 -543
box -1058 -1057 1058 1057
use sky130_fd_pr__pfet_01v8_ANL9FS  XM11
timestamp 1667046312
transform 1 0 8062 0 1 3784
box -194 -804 194 838
use sky130_fd_pr__pfet_01v8_E8XWA6  XM12
timestamp 1666810850
transform 1 0 2260 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_4QVNZ8  XM13
timestamp 1667048966
transform 1 0 8737 0 1 3843
box -194 -864 194 898
use sky130_fd_pr__pfet_01v8_AN68VM  XM15
timestamp 1667053331
transform 1 0 10034 0 1 3582
box -194 -604 194 638
use sky130_fd_pr__pfet_01v8_6ECZVM  XM16
timestamp 1667053331
transform 1 0 9389 0 1 3733
box -194 -754 194 788
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ1 pdk/open_pdks/share/pdk/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1653785680
transform 1 0 1986 0 1 -258
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ2
timestamp 1653785680
transform 1 0 6768 0 1 1458
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ3
timestamp 1653785680
transform 1 0 6762 0 1 610
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ4
timestamp 1653785680
transform 1 0 6762 0 1 -242
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ5
timestamp 1653785680
transform 1 0 6766 0 1 -1080
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ6
timestamp 1653785680
transform 1 0 7608 0 1 -1078
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ7
timestamp 1653785680
transform 1 0 7608 0 1 -242
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ8
timestamp 1653785680
transform 1 0 7608 0 1 614
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  XQ10
timestamp 1653785680
transform 1 0 7612 0 1 1462
box 0 0 796 796
use res52_504  res52_504_0
timestamp 1667019087
transform 0 -1 7886 1 0 2528
box -202 0 74 2664
use res54_789k  res54_789k_0
timestamp 1667400688
transform -1 0 10486 0 -1 3662
box -3806 2918 -3420 5662
use res63_92k  res63_92k_0
timestamp 1667400564
transform -1 0 9706 0 -1 3838
box -3806 2918 -3420 6106
use res298k  res298k_0
timestamp 1667400309
transform -1 0 8744 0 -1 4252
box -3806 2918 -3420 6312
use res484_3K  res484_3K_0
timestamp 1667399187
transform -1 0 8984 0 -1 1656
box -654 0 74 4764
use res517_512K  res517_512K_0
timestamp 1667019531
transform 1 0 -1806 0 1 -1726
box -608 0 710 6864
use res517_512K  res517_512K_1
timestamp 1667019531
transform -1 0 11154 0 -1 3418
box -608 0 710 6864
use sky130_fd_pr__nfet_01v8_7ZFCMD  sky130_fd_pr__nfet_01v8_7ZFCMD_0
timestamp 1666810850
transform 1 0 188 0 1 366
box -1058 -188 1058 188
use sky130_fd_pr__nfet_01v8_VYYYF6  sky130_fd_pr__nfet_01v8_VYYYF6_0
timestamp 1666903823
transform 1 0 4790 0 1 2061
box -258 -1057 258 1057
use sky130_fd_pr__pfet_01v8_A42UEE  sky130_fd_pr__pfet_01v8_A42UEE_0
timestamp 1666810850
transform 1 0 768 0 1 3058
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_0
timestamp 1666810850
transform 1 0 2718 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_E8XWA6  sky130_fd_pr__pfet_01v8_E8XWA6_1
timestamp 1666810850
transform 1 0 3608 0 1 3068
box -294 -2064 294 2098
use sky130_fd_pr__pfet_01v8_GGSNBJ  sky130_fd_pr__pfet_01v8_GGSNBJ_0
timestamp 1666797418
transform 1 0 1514 0 1 1074
box -194 -1100 194 1100
use sky130_fd_pr__res_high_po_0p35_XUGN4V  sky130_fd_pr__res_high_po_0p35_XUGN4V_1
timestamp 1667332169
transform 0 -1 8763 1 0 2553
box -37 -627 37 627
use sky130_fd_pr__res_high_po_0p35_XUGN4V  sky130_fd_pr__res_high_po_0p35_XUGN4V_2
timestamp 1667332169
transform 1 0 -545 0 1 3597
box -37 -627 37 627
<< end >>
