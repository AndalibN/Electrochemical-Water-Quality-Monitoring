magic
tech sky130A
timestamp 1667443396
<< pwell >>
rect -198 -1505 198 1505
<< nmos >>
rect -100 -1400 100 1400
<< ndiff >>
rect -129 1394 -100 1400
rect -129 -1394 -123 1394
rect -106 -1394 -100 1394
rect -129 -1400 -100 -1394
rect 100 1394 129 1400
rect 100 -1394 106 1394
rect 123 -1394 129 1394
rect 100 -1400 129 -1394
<< ndiffc >>
rect -123 -1394 -106 1394
rect 106 -1394 123 1394
<< psubdiff >>
rect -180 1470 -132 1487
rect 132 1470 180 1487
rect -180 1439 -163 1470
rect 163 1439 180 1470
rect -180 -1470 -163 -1439
rect 163 -1470 180 -1439
rect -180 -1487 -132 -1470
rect 132 -1487 180 -1470
<< psubdiffcont >>
rect -132 1470 132 1487
rect -180 -1439 -163 1439
rect 163 -1439 180 1439
rect -132 -1487 132 -1470
<< poly >>
rect -100 1436 100 1444
rect -100 1419 -92 1436
rect 92 1419 100 1436
rect -100 1400 100 1419
rect -100 -1419 100 -1400
rect -100 -1436 -92 -1419
rect 92 -1436 100 -1419
rect -100 -1444 100 -1436
<< polycont >>
rect -92 1419 92 1436
rect -92 -1436 92 -1419
<< locali >>
rect -180 1470 -132 1487
rect 132 1470 180 1487
rect -180 1439 -163 1470
rect 163 1439 180 1470
rect -100 1419 -92 1436
rect 92 1419 100 1436
rect -123 1394 -106 1402
rect -123 -1402 -106 -1394
rect 106 1394 123 1402
rect 106 -1402 123 -1394
rect -100 -1436 -92 -1419
rect 92 -1436 100 -1419
rect -180 -1470 -163 -1439
rect 163 -1470 180 -1439
rect -180 -1487 -132 -1470
rect 132 -1487 180 -1470
<< viali >>
rect -92 1419 92 1436
rect -123 -1394 -106 1394
rect 106 -1394 123 1394
rect -92 -1436 92 -1419
<< metal1 >>
rect -98 1436 98 1439
rect -98 1419 -92 1436
rect 92 1419 98 1436
rect -98 1416 98 1419
rect -126 1394 -103 1400
rect -126 -1394 -123 1394
rect -106 -1394 -103 1394
rect -126 -1400 -103 -1394
rect 103 1394 126 1400
rect 103 -1394 106 1394
rect 123 -1394 126 1394
rect 103 -1400 126 -1394
rect -98 -1419 98 -1416
rect -98 -1436 -92 -1419
rect 92 -1436 98 -1419
rect -98 -1439 98 -1436
<< properties >>
string FIXED_BBOX -171 -1478 171 1478
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 28.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
