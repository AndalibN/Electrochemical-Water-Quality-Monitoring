magic
tech sky130A
magscale 1 2
timestamp 1666812247
<< error_p >>
rect -227 975 -163 981
rect -97 975 -33 981
rect 33 975 97 981
rect 163 975 227 981
rect -227 941 -215 975
rect -97 941 -85 975
rect 33 941 45 975
rect 163 941 175 975
rect -227 935 -163 941
rect -97 935 -33 941
rect 33 935 97 941
rect 163 935 227 941
rect -227 -941 -163 -935
rect -97 -941 -33 -935
rect 33 -941 97 -935
rect 163 -941 227 -935
rect -227 -975 -215 -941
rect -97 -975 -85 -941
rect 33 -975 45 -941
rect 163 -975 175 -941
rect -227 -981 -163 -975
rect -97 -981 -33 -975
rect 33 -981 97 -975
rect 163 -981 227 -975
<< nmos >>
rect -231 -903 -159 903
rect -101 -903 -29 903
rect 29 -903 101 903
rect 159 -903 231 903
<< ndiff >>
rect -289 891 -231 903
rect -289 -891 -277 891
rect -243 -891 -231 891
rect -289 -903 -231 -891
rect -159 891 -101 903
rect -159 -891 -147 891
rect -113 -891 -101 891
rect -159 -903 -101 -891
rect -29 891 29 903
rect -29 -891 -17 891
rect 17 -891 29 891
rect -29 -903 29 -891
rect 101 891 159 903
rect 101 -891 113 891
rect 147 -891 159 891
rect 101 -903 159 -891
rect 231 891 289 903
rect 231 -891 243 891
rect 277 -891 289 891
rect 231 -903 289 -891
<< ndiffc >>
rect -277 -891 -243 891
rect -147 -891 -113 891
rect -17 -891 17 891
rect 113 -891 147 891
rect 243 -891 277 891
<< poly >>
rect -231 975 -159 991
rect -231 941 -215 975
rect -175 941 -159 975
rect -231 903 -159 941
rect -101 975 -29 991
rect -101 941 -85 975
rect -45 941 -29 975
rect -101 903 -29 941
rect 29 975 101 991
rect 29 941 45 975
rect 85 941 101 975
rect 29 903 101 941
rect 159 975 231 991
rect 159 941 175 975
rect 215 941 231 975
rect 159 903 231 941
rect -231 -941 -159 -903
rect -231 -975 -215 -941
rect -175 -975 -159 -941
rect -231 -991 -159 -975
rect -101 -941 -29 -903
rect -101 -975 -85 -941
rect -45 -975 -29 -941
rect -101 -991 -29 -975
rect 29 -941 101 -903
rect 29 -975 45 -941
rect 85 -975 101 -941
rect 29 -991 101 -975
rect 159 -941 231 -903
rect 159 -975 175 -941
rect 215 -975 231 -941
rect 159 -991 231 -975
<< polycont >>
rect -215 941 -175 975
rect -85 941 -45 975
rect 45 941 85 975
rect 175 941 215 975
rect -215 -975 -175 -941
rect -85 -975 -45 -941
rect 45 -975 85 -941
rect 175 -975 215 -941
<< locali >>
rect -231 941 -215 975
rect -175 941 -159 975
rect -101 941 -85 975
rect -45 941 -29 975
rect 29 941 45 975
rect 85 941 101 975
rect 159 941 175 975
rect 215 941 231 975
rect -277 891 -243 907
rect -277 -907 -243 -891
rect -147 891 -113 907
rect -147 -907 -113 -891
rect -17 891 17 907
rect -17 -907 17 -891
rect 113 891 147 907
rect 113 -907 147 -891
rect 243 891 277 907
rect 243 -907 277 -891
rect -231 -975 -215 -941
rect -175 -975 -159 -941
rect -101 -975 -85 -941
rect -45 -975 -29 -941
rect 29 -975 45 -941
rect 85 -975 101 -941
rect 159 -975 175 -941
rect 215 -975 231 -941
<< viali >>
rect -215 941 -175 975
rect -85 941 -45 975
rect 45 941 85 975
rect 175 941 215 975
rect -277 -891 -243 891
rect -147 -891 -113 891
rect -17 -891 17 891
rect 113 -891 147 891
rect 243 -891 277 891
rect -215 -975 -175 -941
rect -85 -975 -45 -941
rect 45 -975 85 -941
rect 175 -975 215 -941
<< metal1 >>
rect -227 975 -163 981
rect -227 941 -215 975
rect -175 941 -163 975
rect -227 935 -163 941
rect -97 975 -33 981
rect -97 941 -85 975
rect -45 941 -33 975
rect -97 935 -33 941
rect 33 975 97 981
rect 33 941 45 975
rect 85 941 97 975
rect 33 935 97 941
rect 163 975 227 981
rect 163 941 175 975
rect 215 941 227 975
rect 163 935 227 941
rect -283 891 -237 903
rect -283 -891 -277 891
rect -243 -891 -237 891
rect -283 -903 -237 -891
rect -153 891 -107 903
rect -153 -891 -147 891
rect -113 -891 -107 891
rect -153 -903 -107 -891
rect -23 891 23 903
rect -23 -891 -17 891
rect 17 -891 23 891
rect -23 -903 23 -891
rect 107 891 153 903
rect 107 -891 113 891
rect 147 -891 153 891
rect 107 -903 153 -891
rect 237 891 283 903
rect 237 -891 243 891
rect 277 -891 283 891
rect 237 -903 283 -891
rect -227 -941 -163 -935
rect -227 -975 -215 -941
rect -175 -975 -163 -941
rect -227 -981 -163 -975
rect -97 -941 -33 -935
rect -97 -975 -85 -941
rect -45 -975 -33 -941
rect -97 -981 -33 -975
rect 33 -941 97 -935
rect 33 -975 45 -941
rect 85 -975 97 -941
rect 33 -981 97 -975
rect 163 -941 227 -935
rect 163 -975 175 -941
rect 215 -975 227 -941
rect 163 -981 227 -975
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 9.03 l 0.361 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
