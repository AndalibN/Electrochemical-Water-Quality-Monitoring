magic
tech sky130A
magscale 1 2
timestamp 1666902736
<< pwell >>
rect -396 -1179 396 1179
<< nmos >>
rect -200 -969 200 1031
<< ndiff >>
rect -258 1019 -200 1031
rect -258 -957 -246 1019
rect -212 -957 -200 1019
rect -258 -969 -200 -957
rect 200 1019 258 1031
rect 200 -957 212 1019
rect 246 -957 258 1019
rect 200 -969 258 -957
<< ndiffc >>
rect -246 -957 -212 1019
rect 212 -957 246 1019
<< psubdiff >>
rect -360 1109 -264 1143
rect 264 1109 360 1143
rect -360 1047 -326 1109
rect 326 1047 360 1109
rect -360 -1109 -326 -1047
rect 326 -1109 360 -1047
rect -360 -1143 -264 -1109
rect 264 -1143 360 -1109
<< psubdiffcont >>
rect -264 1109 264 1143
rect -360 -1047 -326 1047
rect 326 -1047 360 1047
rect -264 -1143 264 -1109
<< poly >>
rect -200 1031 200 1057
rect -200 -1007 200 -969
rect -200 -1041 -184 -1007
rect 184 -1041 200 -1007
rect -200 -1057 200 -1041
<< polycont >>
rect -184 -1041 184 -1007
<< locali >>
rect -280 1109 -264 1143
rect 264 1109 280 1143
rect -360 1047 -326 1063
rect 326 1047 360 1063
rect -246 1019 -212 1035
rect -246 -973 -212 -957
rect 212 1019 246 1035
rect 212 -973 246 -957
rect -200 -1041 -184 -1007
rect 184 -1041 200 -1007
rect -360 -1063 -326 -1047
rect 326 -1063 360 -1047
rect -280 -1143 -264 -1109
rect 264 -1143 280 -1109
<< viali >>
rect -246 -957 -212 1019
rect 212 -957 246 1019
rect -184 -1041 184 -1007
<< metal1 >>
rect -252 1019 -206 1031
rect -252 -957 -246 1019
rect -212 -957 -206 1019
rect -252 -969 -206 -957
rect 206 1019 252 1031
rect 206 -957 212 1019
rect 246 -957 252 1019
rect 206 -969 252 -957
rect -196 -1007 196 -1001
rect -196 -1041 -184 -1007
rect 184 -1041 196 -1007
rect -196 -1047 196 -1041
<< properties >>
string FIXED_BBOX -343 -1126 343 1126
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
