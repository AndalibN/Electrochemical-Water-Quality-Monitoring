magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -277 1878 -213 1884
rect -277 1844 -262 1878
rect -277 1838 -213 1844
<< pwell >>
rect -365 -1832 315 1832
<< nmos >>
rect -281 -1806 -209 1806
rect -101 -1806 -29 1806
rect 29 -1806 101 1806
rect 159 -1806 231 1806
<< ndiff >>
rect -339 1785 -281 1806
rect -339 1751 -327 1785
rect -293 1751 -281 1785
rect -339 1717 -281 1751
rect -339 1683 -327 1717
rect -293 1683 -281 1717
rect -339 1649 -281 1683
rect -339 1615 -327 1649
rect -293 1615 -281 1649
rect -339 1581 -281 1615
rect -339 1547 -327 1581
rect -293 1547 -281 1581
rect -339 1513 -281 1547
rect -339 1479 -327 1513
rect -293 1479 -281 1513
rect -339 1445 -281 1479
rect -339 1411 -327 1445
rect -293 1411 -281 1445
rect -339 1377 -281 1411
rect -339 1343 -327 1377
rect -293 1343 -281 1377
rect -339 1309 -281 1343
rect -339 1275 -327 1309
rect -293 1275 -281 1309
rect -339 1241 -281 1275
rect -339 1207 -327 1241
rect -293 1207 -281 1241
rect -339 1173 -281 1207
rect -339 1139 -327 1173
rect -293 1139 -281 1173
rect -339 1105 -281 1139
rect -339 1071 -327 1105
rect -293 1071 -281 1105
rect -339 1037 -281 1071
rect -339 1003 -327 1037
rect -293 1003 -281 1037
rect -339 969 -281 1003
rect -339 935 -327 969
rect -293 935 -281 969
rect -339 901 -281 935
rect -339 867 -327 901
rect -293 867 -281 901
rect -339 833 -281 867
rect -339 799 -327 833
rect -293 799 -281 833
rect -339 765 -281 799
rect -339 731 -327 765
rect -293 731 -281 765
rect -339 697 -281 731
rect -339 663 -327 697
rect -293 663 -281 697
rect -339 629 -281 663
rect -339 595 -327 629
rect -293 595 -281 629
rect -339 561 -281 595
rect -339 527 -327 561
rect -293 527 -281 561
rect -339 493 -281 527
rect -339 459 -327 493
rect -293 459 -281 493
rect -339 425 -281 459
rect -339 391 -327 425
rect -293 391 -281 425
rect -339 357 -281 391
rect -339 323 -327 357
rect -293 323 -281 357
rect -339 289 -281 323
rect -339 255 -327 289
rect -293 255 -281 289
rect -339 221 -281 255
rect -339 187 -327 221
rect -293 187 -281 221
rect -339 153 -281 187
rect -339 119 -327 153
rect -293 119 -281 153
rect -339 85 -281 119
rect -339 51 -327 85
rect -293 51 -281 85
rect -339 17 -281 51
rect -339 -17 -327 17
rect -293 -17 -281 17
rect -339 -51 -281 -17
rect -339 -85 -327 -51
rect -293 -85 -281 -51
rect -339 -119 -281 -85
rect -339 -153 -327 -119
rect -293 -153 -281 -119
rect -339 -187 -281 -153
rect -339 -221 -327 -187
rect -293 -221 -281 -187
rect -339 -255 -281 -221
rect -339 -289 -327 -255
rect -293 -289 -281 -255
rect -339 -323 -281 -289
rect -339 -357 -327 -323
rect -293 -357 -281 -323
rect -339 -391 -281 -357
rect -339 -425 -327 -391
rect -293 -425 -281 -391
rect -339 -459 -281 -425
rect -339 -493 -327 -459
rect -293 -493 -281 -459
rect -339 -527 -281 -493
rect -339 -561 -327 -527
rect -293 -561 -281 -527
rect -339 -595 -281 -561
rect -339 -629 -327 -595
rect -293 -629 -281 -595
rect -339 -663 -281 -629
rect -339 -697 -327 -663
rect -293 -697 -281 -663
rect -339 -731 -281 -697
rect -339 -765 -327 -731
rect -293 -765 -281 -731
rect -339 -799 -281 -765
rect -339 -833 -327 -799
rect -293 -833 -281 -799
rect -339 -867 -281 -833
rect -339 -901 -327 -867
rect -293 -901 -281 -867
rect -339 -935 -281 -901
rect -339 -969 -327 -935
rect -293 -969 -281 -935
rect -339 -1003 -281 -969
rect -339 -1037 -327 -1003
rect -293 -1037 -281 -1003
rect -339 -1071 -281 -1037
rect -339 -1105 -327 -1071
rect -293 -1105 -281 -1071
rect -339 -1139 -281 -1105
rect -339 -1173 -327 -1139
rect -293 -1173 -281 -1139
rect -339 -1207 -281 -1173
rect -339 -1241 -327 -1207
rect -293 -1241 -281 -1207
rect -339 -1275 -281 -1241
rect -339 -1309 -327 -1275
rect -293 -1309 -281 -1275
rect -339 -1343 -281 -1309
rect -339 -1377 -327 -1343
rect -293 -1377 -281 -1343
rect -339 -1411 -281 -1377
rect -339 -1445 -327 -1411
rect -293 -1445 -281 -1411
rect -339 -1479 -281 -1445
rect -339 -1513 -327 -1479
rect -293 -1513 -281 -1479
rect -339 -1547 -281 -1513
rect -339 -1581 -327 -1547
rect -293 -1581 -281 -1547
rect -339 -1615 -281 -1581
rect -339 -1649 -327 -1615
rect -293 -1649 -281 -1615
rect -339 -1683 -281 -1649
rect -339 -1717 -327 -1683
rect -293 -1717 -281 -1683
rect -339 -1751 -281 -1717
rect -339 -1785 -327 -1751
rect -293 -1785 -281 -1751
rect -339 -1806 -281 -1785
rect -209 1785 -101 1806
rect -209 1751 -172 1785
rect -138 1751 -101 1785
rect -209 1717 -101 1751
rect -209 1683 -172 1717
rect -138 1683 -101 1717
rect -209 1649 -101 1683
rect -209 1615 -172 1649
rect -138 1615 -101 1649
rect -209 1581 -101 1615
rect -209 1547 -172 1581
rect -138 1547 -101 1581
rect -209 1513 -101 1547
rect -209 1479 -172 1513
rect -138 1479 -101 1513
rect -209 1445 -101 1479
rect -209 1411 -172 1445
rect -138 1411 -101 1445
rect -209 1377 -101 1411
rect -209 1343 -172 1377
rect -138 1343 -101 1377
rect -209 1309 -101 1343
rect -209 1275 -172 1309
rect -138 1275 -101 1309
rect -209 1241 -101 1275
rect -209 1207 -172 1241
rect -138 1207 -101 1241
rect -209 1173 -101 1207
rect -209 1139 -172 1173
rect -138 1139 -101 1173
rect -209 1105 -101 1139
rect -209 1071 -172 1105
rect -138 1071 -101 1105
rect -209 1037 -101 1071
rect -209 1003 -172 1037
rect -138 1003 -101 1037
rect -209 969 -101 1003
rect -209 935 -172 969
rect -138 935 -101 969
rect -209 901 -101 935
rect -209 867 -172 901
rect -138 867 -101 901
rect -209 833 -101 867
rect -209 799 -172 833
rect -138 799 -101 833
rect -209 765 -101 799
rect -209 731 -172 765
rect -138 731 -101 765
rect -209 697 -101 731
rect -209 663 -172 697
rect -138 663 -101 697
rect -209 629 -101 663
rect -209 595 -172 629
rect -138 595 -101 629
rect -209 561 -101 595
rect -209 527 -172 561
rect -138 527 -101 561
rect -209 493 -101 527
rect -209 459 -172 493
rect -138 459 -101 493
rect -209 425 -101 459
rect -209 391 -172 425
rect -138 391 -101 425
rect -209 357 -101 391
rect -209 323 -172 357
rect -138 323 -101 357
rect -209 289 -101 323
rect -209 255 -172 289
rect -138 255 -101 289
rect -209 221 -101 255
rect -209 187 -172 221
rect -138 187 -101 221
rect -209 153 -101 187
rect -209 119 -172 153
rect -138 119 -101 153
rect -209 85 -101 119
rect -209 51 -172 85
rect -138 51 -101 85
rect -209 17 -101 51
rect -209 -17 -172 17
rect -138 -17 -101 17
rect -209 -51 -101 -17
rect -209 -85 -172 -51
rect -138 -85 -101 -51
rect -209 -119 -101 -85
rect -209 -153 -172 -119
rect -138 -153 -101 -119
rect -209 -187 -101 -153
rect -209 -221 -172 -187
rect -138 -221 -101 -187
rect -209 -255 -101 -221
rect -209 -289 -172 -255
rect -138 -289 -101 -255
rect -209 -323 -101 -289
rect -209 -357 -172 -323
rect -138 -357 -101 -323
rect -209 -391 -101 -357
rect -209 -425 -172 -391
rect -138 -425 -101 -391
rect -209 -459 -101 -425
rect -209 -493 -172 -459
rect -138 -493 -101 -459
rect -209 -527 -101 -493
rect -209 -561 -172 -527
rect -138 -561 -101 -527
rect -209 -595 -101 -561
rect -209 -629 -172 -595
rect -138 -629 -101 -595
rect -209 -663 -101 -629
rect -209 -697 -172 -663
rect -138 -697 -101 -663
rect -209 -731 -101 -697
rect -209 -765 -172 -731
rect -138 -765 -101 -731
rect -209 -799 -101 -765
rect -209 -833 -172 -799
rect -138 -833 -101 -799
rect -209 -867 -101 -833
rect -209 -901 -172 -867
rect -138 -901 -101 -867
rect -209 -935 -101 -901
rect -209 -969 -172 -935
rect -138 -969 -101 -935
rect -209 -1003 -101 -969
rect -209 -1037 -172 -1003
rect -138 -1037 -101 -1003
rect -209 -1071 -101 -1037
rect -209 -1105 -172 -1071
rect -138 -1105 -101 -1071
rect -209 -1139 -101 -1105
rect -209 -1173 -172 -1139
rect -138 -1173 -101 -1139
rect -209 -1207 -101 -1173
rect -209 -1241 -172 -1207
rect -138 -1241 -101 -1207
rect -209 -1275 -101 -1241
rect -209 -1309 -172 -1275
rect -138 -1309 -101 -1275
rect -209 -1343 -101 -1309
rect -209 -1377 -172 -1343
rect -138 -1377 -101 -1343
rect -209 -1411 -101 -1377
rect -209 -1445 -172 -1411
rect -138 -1445 -101 -1411
rect -209 -1479 -101 -1445
rect -209 -1513 -172 -1479
rect -138 -1513 -101 -1479
rect -209 -1547 -101 -1513
rect -209 -1581 -172 -1547
rect -138 -1581 -101 -1547
rect -209 -1615 -101 -1581
rect -209 -1649 -172 -1615
rect -138 -1649 -101 -1615
rect -209 -1683 -101 -1649
rect -209 -1717 -172 -1683
rect -138 -1717 -101 -1683
rect -209 -1751 -101 -1717
rect -209 -1785 -172 -1751
rect -138 -1785 -101 -1751
rect -209 -1806 -101 -1785
rect -29 1785 29 1806
rect -29 1751 -17 1785
rect 17 1751 29 1785
rect -29 1717 29 1751
rect -29 1683 -17 1717
rect 17 1683 29 1717
rect -29 1649 29 1683
rect -29 1615 -17 1649
rect 17 1615 29 1649
rect -29 1581 29 1615
rect -29 1547 -17 1581
rect 17 1547 29 1581
rect -29 1513 29 1547
rect -29 1479 -17 1513
rect 17 1479 29 1513
rect -29 1445 29 1479
rect -29 1411 -17 1445
rect 17 1411 29 1445
rect -29 1377 29 1411
rect -29 1343 -17 1377
rect 17 1343 29 1377
rect -29 1309 29 1343
rect -29 1275 -17 1309
rect 17 1275 29 1309
rect -29 1241 29 1275
rect -29 1207 -17 1241
rect 17 1207 29 1241
rect -29 1173 29 1207
rect -29 1139 -17 1173
rect 17 1139 29 1173
rect -29 1105 29 1139
rect -29 1071 -17 1105
rect 17 1071 29 1105
rect -29 1037 29 1071
rect -29 1003 -17 1037
rect 17 1003 29 1037
rect -29 969 29 1003
rect -29 935 -17 969
rect 17 935 29 969
rect -29 901 29 935
rect -29 867 -17 901
rect 17 867 29 901
rect -29 833 29 867
rect -29 799 -17 833
rect 17 799 29 833
rect -29 765 29 799
rect -29 731 -17 765
rect 17 731 29 765
rect -29 697 29 731
rect -29 663 -17 697
rect 17 663 29 697
rect -29 629 29 663
rect -29 595 -17 629
rect 17 595 29 629
rect -29 561 29 595
rect -29 527 -17 561
rect 17 527 29 561
rect -29 493 29 527
rect -29 459 -17 493
rect 17 459 29 493
rect -29 425 29 459
rect -29 391 -17 425
rect 17 391 29 425
rect -29 357 29 391
rect -29 323 -17 357
rect 17 323 29 357
rect -29 289 29 323
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -323 29 -289
rect -29 -357 -17 -323
rect 17 -357 29 -323
rect -29 -391 29 -357
rect -29 -425 -17 -391
rect 17 -425 29 -391
rect -29 -459 29 -425
rect -29 -493 -17 -459
rect 17 -493 29 -459
rect -29 -527 29 -493
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -595 29 -561
rect -29 -629 -17 -595
rect 17 -629 29 -595
rect -29 -663 29 -629
rect -29 -697 -17 -663
rect 17 -697 29 -663
rect -29 -731 29 -697
rect -29 -765 -17 -731
rect 17 -765 29 -731
rect -29 -799 29 -765
rect -29 -833 -17 -799
rect 17 -833 29 -799
rect -29 -867 29 -833
rect -29 -901 -17 -867
rect 17 -901 29 -867
rect -29 -935 29 -901
rect -29 -969 -17 -935
rect 17 -969 29 -935
rect -29 -1003 29 -969
rect -29 -1037 -17 -1003
rect 17 -1037 29 -1003
rect -29 -1071 29 -1037
rect -29 -1105 -17 -1071
rect 17 -1105 29 -1071
rect -29 -1139 29 -1105
rect -29 -1173 -17 -1139
rect 17 -1173 29 -1139
rect -29 -1207 29 -1173
rect -29 -1241 -17 -1207
rect 17 -1241 29 -1207
rect -29 -1275 29 -1241
rect -29 -1309 -17 -1275
rect 17 -1309 29 -1275
rect -29 -1343 29 -1309
rect -29 -1377 -17 -1343
rect 17 -1377 29 -1343
rect -29 -1411 29 -1377
rect -29 -1445 -17 -1411
rect 17 -1445 29 -1411
rect -29 -1479 29 -1445
rect -29 -1513 -17 -1479
rect 17 -1513 29 -1479
rect -29 -1547 29 -1513
rect -29 -1581 -17 -1547
rect 17 -1581 29 -1547
rect -29 -1615 29 -1581
rect -29 -1649 -17 -1615
rect 17 -1649 29 -1615
rect -29 -1683 29 -1649
rect -29 -1717 -17 -1683
rect 17 -1717 29 -1683
rect -29 -1751 29 -1717
rect -29 -1785 -17 -1751
rect 17 -1785 29 -1751
rect -29 -1806 29 -1785
rect 101 1785 159 1806
rect 101 1751 113 1785
rect 147 1751 159 1785
rect 101 1717 159 1751
rect 101 1683 113 1717
rect 147 1683 159 1717
rect 101 1649 159 1683
rect 101 1615 113 1649
rect 147 1615 159 1649
rect 101 1581 159 1615
rect 101 1547 113 1581
rect 147 1547 159 1581
rect 101 1513 159 1547
rect 101 1479 113 1513
rect 147 1479 159 1513
rect 101 1445 159 1479
rect 101 1411 113 1445
rect 147 1411 159 1445
rect 101 1377 159 1411
rect 101 1343 113 1377
rect 147 1343 159 1377
rect 101 1309 159 1343
rect 101 1275 113 1309
rect 147 1275 159 1309
rect 101 1241 159 1275
rect 101 1207 113 1241
rect 147 1207 159 1241
rect 101 1173 159 1207
rect 101 1139 113 1173
rect 147 1139 159 1173
rect 101 1105 159 1139
rect 101 1071 113 1105
rect 147 1071 159 1105
rect 101 1037 159 1071
rect 101 1003 113 1037
rect 147 1003 159 1037
rect 101 969 159 1003
rect 101 935 113 969
rect 147 935 159 969
rect 101 901 159 935
rect 101 867 113 901
rect 147 867 159 901
rect 101 833 159 867
rect 101 799 113 833
rect 147 799 159 833
rect 101 765 159 799
rect 101 731 113 765
rect 147 731 159 765
rect 101 697 159 731
rect 101 663 113 697
rect 147 663 159 697
rect 101 629 159 663
rect 101 595 113 629
rect 147 595 159 629
rect 101 561 159 595
rect 101 527 113 561
rect 147 527 159 561
rect 101 493 159 527
rect 101 459 113 493
rect 147 459 159 493
rect 101 425 159 459
rect 101 391 113 425
rect 147 391 159 425
rect 101 357 159 391
rect 101 323 113 357
rect 147 323 159 357
rect 101 289 159 323
rect 101 255 113 289
rect 147 255 159 289
rect 101 221 159 255
rect 101 187 113 221
rect 147 187 159 221
rect 101 153 159 187
rect 101 119 113 153
rect 147 119 159 153
rect 101 85 159 119
rect 101 51 113 85
rect 147 51 159 85
rect 101 17 159 51
rect 101 -17 113 17
rect 147 -17 159 17
rect 101 -51 159 -17
rect 101 -85 113 -51
rect 147 -85 159 -51
rect 101 -119 159 -85
rect 101 -153 113 -119
rect 147 -153 159 -119
rect 101 -187 159 -153
rect 101 -221 113 -187
rect 147 -221 159 -187
rect 101 -255 159 -221
rect 101 -289 113 -255
rect 147 -289 159 -255
rect 101 -323 159 -289
rect 101 -357 113 -323
rect 147 -357 159 -323
rect 101 -391 159 -357
rect 101 -425 113 -391
rect 147 -425 159 -391
rect 101 -459 159 -425
rect 101 -493 113 -459
rect 147 -493 159 -459
rect 101 -527 159 -493
rect 101 -561 113 -527
rect 147 -561 159 -527
rect 101 -595 159 -561
rect 101 -629 113 -595
rect 147 -629 159 -595
rect 101 -663 159 -629
rect 101 -697 113 -663
rect 147 -697 159 -663
rect 101 -731 159 -697
rect 101 -765 113 -731
rect 147 -765 159 -731
rect 101 -799 159 -765
rect 101 -833 113 -799
rect 147 -833 159 -799
rect 101 -867 159 -833
rect 101 -901 113 -867
rect 147 -901 159 -867
rect 101 -935 159 -901
rect 101 -969 113 -935
rect 147 -969 159 -935
rect 101 -1003 159 -969
rect 101 -1037 113 -1003
rect 147 -1037 159 -1003
rect 101 -1071 159 -1037
rect 101 -1105 113 -1071
rect 147 -1105 159 -1071
rect 101 -1139 159 -1105
rect 101 -1173 113 -1139
rect 147 -1173 159 -1139
rect 101 -1207 159 -1173
rect 101 -1241 113 -1207
rect 147 -1241 159 -1207
rect 101 -1275 159 -1241
rect 101 -1309 113 -1275
rect 147 -1309 159 -1275
rect 101 -1343 159 -1309
rect 101 -1377 113 -1343
rect 147 -1377 159 -1343
rect 101 -1411 159 -1377
rect 101 -1445 113 -1411
rect 147 -1445 159 -1411
rect 101 -1479 159 -1445
rect 101 -1513 113 -1479
rect 147 -1513 159 -1479
rect 101 -1547 159 -1513
rect 101 -1581 113 -1547
rect 147 -1581 159 -1547
rect 101 -1615 159 -1581
rect 101 -1649 113 -1615
rect 147 -1649 159 -1615
rect 101 -1683 159 -1649
rect 101 -1717 113 -1683
rect 147 -1717 159 -1683
rect 101 -1751 159 -1717
rect 101 -1785 113 -1751
rect 147 -1785 159 -1751
rect 101 -1806 159 -1785
rect 231 1785 289 1806
rect 231 1751 243 1785
rect 277 1751 289 1785
rect 231 1717 289 1751
rect 231 1683 243 1717
rect 277 1683 289 1717
rect 231 1649 289 1683
rect 231 1615 243 1649
rect 277 1615 289 1649
rect 231 1581 289 1615
rect 231 1547 243 1581
rect 277 1547 289 1581
rect 231 1513 289 1547
rect 231 1479 243 1513
rect 277 1479 289 1513
rect 231 1445 289 1479
rect 231 1411 243 1445
rect 277 1411 289 1445
rect 231 1377 289 1411
rect 231 1343 243 1377
rect 277 1343 289 1377
rect 231 1309 289 1343
rect 231 1275 243 1309
rect 277 1275 289 1309
rect 231 1241 289 1275
rect 231 1207 243 1241
rect 277 1207 289 1241
rect 231 1173 289 1207
rect 231 1139 243 1173
rect 277 1139 289 1173
rect 231 1105 289 1139
rect 231 1071 243 1105
rect 277 1071 289 1105
rect 231 1037 289 1071
rect 231 1003 243 1037
rect 277 1003 289 1037
rect 231 969 289 1003
rect 231 935 243 969
rect 277 935 289 969
rect 231 901 289 935
rect 231 867 243 901
rect 277 867 289 901
rect 231 833 289 867
rect 231 799 243 833
rect 277 799 289 833
rect 231 765 289 799
rect 231 731 243 765
rect 277 731 289 765
rect 231 697 289 731
rect 231 663 243 697
rect 277 663 289 697
rect 231 629 289 663
rect 231 595 243 629
rect 277 595 289 629
rect 231 561 289 595
rect 231 527 243 561
rect 277 527 289 561
rect 231 493 289 527
rect 231 459 243 493
rect 277 459 289 493
rect 231 425 289 459
rect 231 391 243 425
rect 277 391 289 425
rect 231 357 289 391
rect 231 323 243 357
rect 277 323 289 357
rect 231 289 289 323
rect 231 255 243 289
rect 277 255 289 289
rect 231 221 289 255
rect 231 187 243 221
rect 277 187 289 221
rect 231 153 289 187
rect 231 119 243 153
rect 277 119 289 153
rect 231 85 289 119
rect 231 51 243 85
rect 277 51 289 85
rect 231 17 289 51
rect 231 -17 243 17
rect 277 -17 289 17
rect 231 -51 289 -17
rect 231 -85 243 -51
rect 277 -85 289 -51
rect 231 -119 289 -85
rect 231 -153 243 -119
rect 277 -153 289 -119
rect 231 -187 289 -153
rect 231 -221 243 -187
rect 277 -221 289 -187
rect 231 -255 289 -221
rect 231 -289 243 -255
rect 277 -289 289 -255
rect 231 -323 289 -289
rect 231 -357 243 -323
rect 277 -357 289 -323
rect 231 -391 289 -357
rect 231 -425 243 -391
rect 277 -425 289 -391
rect 231 -459 289 -425
rect 231 -493 243 -459
rect 277 -493 289 -459
rect 231 -527 289 -493
rect 231 -561 243 -527
rect 277 -561 289 -527
rect 231 -595 289 -561
rect 231 -629 243 -595
rect 277 -629 289 -595
rect 231 -663 289 -629
rect 231 -697 243 -663
rect 277 -697 289 -663
rect 231 -731 289 -697
rect 231 -765 243 -731
rect 277 -765 289 -731
rect 231 -799 289 -765
rect 231 -833 243 -799
rect 277 -833 289 -799
rect 231 -867 289 -833
rect 231 -901 243 -867
rect 277 -901 289 -867
rect 231 -935 289 -901
rect 231 -969 243 -935
rect 277 -969 289 -935
rect 231 -1003 289 -969
rect 231 -1037 243 -1003
rect 277 -1037 289 -1003
rect 231 -1071 289 -1037
rect 231 -1105 243 -1071
rect 277 -1105 289 -1071
rect 231 -1139 289 -1105
rect 231 -1173 243 -1139
rect 277 -1173 289 -1139
rect 231 -1207 289 -1173
rect 231 -1241 243 -1207
rect 277 -1241 289 -1207
rect 231 -1275 289 -1241
rect 231 -1309 243 -1275
rect 277 -1309 289 -1275
rect 231 -1343 289 -1309
rect 231 -1377 243 -1343
rect 277 -1377 289 -1343
rect 231 -1411 289 -1377
rect 231 -1445 243 -1411
rect 277 -1445 289 -1411
rect 231 -1479 289 -1445
rect 231 -1513 243 -1479
rect 277 -1513 289 -1479
rect 231 -1547 289 -1513
rect 231 -1581 243 -1547
rect 277 -1581 289 -1547
rect 231 -1615 289 -1581
rect 231 -1649 243 -1615
rect 277 -1649 289 -1615
rect 231 -1683 289 -1649
rect 231 -1717 243 -1683
rect 277 -1717 289 -1683
rect 231 -1751 289 -1717
rect 231 -1785 243 -1751
rect 277 -1785 289 -1751
rect 231 -1806 289 -1785
<< ndiffc >>
rect -327 1751 -293 1785
rect -327 1683 -293 1717
rect -327 1615 -293 1649
rect -327 1547 -293 1581
rect -327 1479 -293 1513
rect -327 1411 -293 1445
rect -327 1343 -293 1377
rect -327 1275 -293 1309
rect -327 1207 -293 1241
rect -327 1139 -293 1173
rect -327 1071 -293 1105
rect -327 1003 -293 1037
rect -327 935 -293 969
rect -327 867 -293 901
rect -327 799 -293 833
rect -327 731 -293 765
rect -327 663 -293 697
rect -327 595 -293 629
rect -327 527 -293 561
rect -327 459 -293 493
rect -327 391 -293 425
rect -327 323 -293 357
rect -327 255 -293 289
rect -327 187 -293 221
rect -327 119 -293 153
rect -327 51 -293 85
rect -327 -17 -293 17
rect -327 -85 -293 -51
rect -327 -153 -293 -119
rect -327 -221 -293 -187
rect -327 -289 -293 -255
rect -327 -357 -293 -323
rect -327 -425 -293 -391
rect -327 -493 -293 -459
rect -327 -561 -293 -527
rect -327 -629 -293 -595
rect -327 -697 -293 -663
rect -327 -765 -293 -731
rect -327 -833 -293 -799
rect -327 -901 -293 -867
rect -327 -969 -293 -935
rect -327 -1037 -293 -1003
rect -327 -1105 -293 -1071
rect -327 -1173 -293 -1139
rect -327 -1241 -293 -1207
rect -327 -1309 -293 -1275
rect -327 -1377 -293 -1343
rect -327 -1445 -293 -1411
rect -327 -1513 -293 -1479
rect -327 -1581 -293 -1547
rect -327 -1649 -293 -1615
rect -327 -1717 -293 -1683
rect -327 -1785 -293 -1751
rect -172 1751 -138 1785
rect -172 1683 -138 1717
rect -172 1615 -138 1649
rect -172 1547 -138 1581
rect -172 1479 -138 1513
rect -172 1411 -138 1445
rect -172 1343 -138 1377
rect -172 1275 -138 1309
rect -172 1207 -138 1241
rect -172 1139 -138 1173
rect -172 1071 -138 1105
rect -172 1003 -138 1037
rect -172 935 -138 969
rect -172 867 -138 901
rect -172 799 -138 833
rect -172 731 -138 765
rect -172 663 -138 697
rect -172 595 -138 629
rect -172 527 -138 561
rect -172 459 -138 493
rect -172 391 -138 425
rect -172 323 -138 357
rect -172 255 -138 289
rect -172 187 -138 221
rect -172 119 -138 153
rect -172 51 -138 85
rect -172 -17 -138 17
rect -172 -85 -138 -51
rect -172 -153 -138 -119
rect -172 -221 -138 -187
rect -172 -289 -138 -255
rect -172 -357 -138 -323
rect -172 -425 -138 -391
rect -172 -493 -138 -459
rect -172 -561 -138 -527
rect -172 -629 -138 -595
rect -172 -697 -138 -663
rect -172 -765 -138 -731
rect -172 -833 -138 -799
rect -172 -901 -138 -867
rect -172 -969 -138 -935
rect -172 -1037 -138 -1003
rect -172 -1105 -138 -1071
rect -172 -1173 -138 -1139
rect -172 -1241 -138 -1207
rect -172 -1309 -138 -1275
rect -172 -1377 -138 -1343
rect -172 -1445 -138 -1411
rect -172 -1513 -138 -1479
rect -172 -1581 -138 -1547
rect -172 -1649 -138 -1615
rect -172 -1717 -138 -1683
rect -172 -1785 -138 -1751
rect -17 1751 17 1785
rect -17 1683 17 1717
rect -17 1615 17 1649
rect -17 1547 17 1581
rect -17 1479 17 1513
rect -17 1411 17 1445
rect -17 1343 17 1377
rect -17 1275 17 1309
rect -17 1207 17 1241
rect -17 1139 17 1173
rect -17 1071 17 1105
rect -17 1003 17 1037
rect -17 935 17 969
rect -17 867 17 901
rect -17 799 17 833
rect -17 731 17 765
rect -17 663 17 697
rect -17 595 17 629
rect -17 527 17 561
rect -17 459 17 493
rect -17 391 17 425
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect -17 -425 17 -391
rect -17 -493 17 -459
rect -17 -561 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -663
rect -17 -765 17 -731
rect -17 -833 17 -799
rect -17 -901 17 -867
rect -17 -969 17 -935
rect -17 -1037 17 -1003
rect -17 -1105 17 -1071
rect -17 -1173 17 -1139
rect -17 -1241 17 -1207
rect -17 -1309 17 -1275
rect -17 -1377 17 -1343
rect -17 -1445 17 -1411
rect -17 -1513 17 -1479
rect -17 -1581 17 -1547
rect -17 -1649 17 -1615
rect -17 -1717 17 -1683
rect -17 -1785 17 -1751
rect 113 1751 147 1785
rect 113 1683 147 1717
rect 113 1615 147 1649
rect 113 1547 147 1581
rect 113 1479 147 1513
rect 113 1411 147 1445
rect 113 1343 147 1377
rect 113 1275 147 1309
rect 113 1207 147 1241
rect 113 1139 147 1173
rect 113 1071 147 1105
rect 113 1003 147 1037
rect 113 935 147 969
rect 113 867 147 901
rect 113 799 147 833
rect 113 731 147 765
rect 113 663 147 697
rect 113 595 147 629
rect 113 527 147 561
rect 113 459 147 493
rect 113 391 147 425
rect 113 323 147 357
rect 113 255 147 289
rect 113 187 147 221
rect 113 119 147 153
rect 113 51 147 85
rect 113 -17 147 17
rect 113 -85 147 -51
rect 113 -153 147 -119
rect 113 -221 147 -187
rect 113 -289 147 -255
rect 113 -357 147 -323
rect 113 -425 147 -391
rect 113 -493 147 -459
rect 113 -561 147 -527
rect 113 -629 147 -595
rect 113 -697 147 -663
rect 113 -765 147 -731
rect 113 -833 147 -799
rect 113 -901 147 -867
rect 113 -969 147 -935
rect 113 -1037 147 -1003
rect 113 -1105 147 -1071
rect 113 -1173 147 -1139
rect 113 -1241 147 -1207
rect 113 -1309 147 -1275
rect 113 -1377 147 -1343
rect 113 -1445 147 -1411
rect 113 -1513 147 -1479
rect 113 -1581 147 -1547
rect 113 -1649 147 -1615
rect 113 -1717 147 -1683
rect 113 -1785 147 -1751
rect 243 1751 277 1785
rect 243 1683 277 1717
rect 243 1615 277 1649
rect 243 1547 277 1581
rect 243 1479 277 1513
rect 243 1411 277 1445
rect 243 1343 277 1377
rect 243 1275 277 1309
rect 243 1207 277 1241
rect 243 1139 277 1173
rect 243 1071 277 1105
rect 243 1003 277 1037
rect 243 935 277 969
rect 243 867 277 901
rect 243 799 277 833
rect 243 731 277 765
rect 243 663 277 697
rect 243 595 277 629
rect 243 527 277 561
rect 243 459 277 493
rect 243 391 277 425
rect 243 323 277 357
rect 243 255 277 289
rect 243 187 277 221
rect 243 119 277 153
rect 243 51 277 85
rect 243 -17 277 17
rect 243 -85 277 -51
rect 243 -153 277 -119
rect 243 -221 277 -187
rect 243 -289 277 -255
rect 243 -357 277 -323
rect 243 -425 277 -391
rect 243 -493 277 -459
rect 243 -561 277 -527
rect 243 -629 277 -595
rect 243 -697 277 -663
rect 243 -765 277 -731
rect 243 -833 277 -799
rect 243 -901 277 -867
rect 243 -969 277 -935
rect 243 -1037 277 -1003
rect 243 -1105 277 -1071
rect 243 -1173 277 -1139
rect 243 -1241 277 -1207
rect 243 -1309 277 -1275
rect 243 -1377 277 -1343
rect 243 -1445 277 -1411
rect 243 -1513 277 -1479
rect 243 -1581 277 -1547
rect 243 -1649 277 -1615
rect 243 -1717 277 -1683
rect 243 -1785 277 -1751
<< poly >>
rect -281 1878 -209 1894
rect -281 1844 -262 1878
rect -228 1844 -209 1878
rect -281 1806 -209 1844
rect -101 1838 101 1894
rect -101 1806 -29 1838
rect 29 1806 101 1838
rect 159 1806 231 1838
rect -281 -1837 -209 -1806
rect -101 -1837 -29 -1806
rect -281 -1893 -29 -1837
rect 29 -1837 101 -1806
rect 159 -1837 231 -1806
rect 29 -1893 231 -1837
<< polycont >>
rect -262 1844 -228 1878
<< locali >>
rect -281 1844 -262 1878
rect -228 1844 -209 1878
rect -327 1785 -293 1810
rect -327 1717 -293 1747
rect -327 1649 -293 1675
rect -327 1581 -293 1603
rect -327 1513 -293 1531
rect -327 1445 -293 1459
rect -327 1377 -293 1387
rect -327 1309 -293 1315
rect -327 1241 -293 1243
rect -327 1205 -293 1207
rect -327 1133 -293 1139
rect -327 1061 -293 1071
rect -327 989 -293 1003
rect -327 917 -293 935
rect -327 845 -293 867
rect -327 773 -293 799
rect -327 701 -293 731
rect -327 629 -293 663
rect -327 561 -293 595
rect -327 493 -293 523
rect -327 425 -293 451
rect -327 357 -293 379
rect -327 289 -293 307
rect -327 221 -293 235
rect -327 153 -293 163
rect -327 85 -293 91
rect -327 17 -293 19
rect -327 -19 -293 -17
rect -327 -91 -293 -85
rect -327 -163 -293 -153
rect -327 -235 -293 -221
rect -327 -307 -293 -289
rect -327 -379 -293 -357
rect -327 -451 -293 -425
rect -327 -523 -293 -493
rect -327 -595 -293 -561
rect -327 -663 -293 -629
rect -327 -731 -293 -701
rect -327 -799 -293 -773
rect -327 -867 -293 -845
rect -327 -935 -293 -917
rect -327 -1003 -293 -989
rect -327 -1071 -293 -1061
rect -327 -1139 -293 -1133
rect -327 -1207 -293 -1205
rect -327 -1243 -293 -1241
rect -327 -1315 -293 -1309
rect -327 -1387 -293 -1377
rect -327 -1459 -293 -1445
rect -327 -1531 -293 -1513
rect -327 -1603 -293 -1581
rect -327 -1675 -293 -1649
rect -327 -1747 -293 -1717
rect -327 -1810 -293 -1785
rect -197 1785 -113 1810
rect -197 1747 -172 1785
rect -138 1747 -113 1785
rect -197 1717 -113 1747
rect -197 1675 -172 1717
rect -138 1675 -113 1717
rect -197 1649 -113 1675
rect -197 1603 -172 1649
rect -138 1603 -113 1649
rect -197 1581 -113 1603
rect -197 1531 -172 1581
rect -138 1531 -113 1581
rect -197 1513 -113 1531
rect -197 1459 -172 1513
rect -138 1459 -113 1513
rect -197 1445 -113 1459
rect -197 1387 -172 1445
rect -138 1387 -113 1445
rect -197 1377 -113 1387
rect -197 1315 -172 1377
rect -138 1315 -113 1377
rect -197 1309 -113 1315
rect -197 1243 -172 1309
rect -138 1243 -113 1309
rect -197 1241 -113 1243
rect -197 1207 -172 1241
rect -138 1207 -113 1241
rect -197 1205 -113 1207
rect -197 1139 -172 1205
rect -138 1139 -113 1205
rect -197 1133 -113 1139
rect -197 1071 -172 1133
rect -138 1071 -113 1133
rect -197 1061 -113 1071
rect -197 1003 -172 1061
rect -138 1003 -113 1061
rect -197 989 -113 1003
rect -197 935 -172 989
rect -138 935 -113 989
rect -197 917 -113 935
rect -197 867 -172 917
rect -138 867 -113 917
rect -197 845 -113 867
rect -197 799 -172 845
rect -138 799 -113 845
rect -197 773 -113 799
rect -197 731 -172 773
rect -138 731 -113 773
rect -197 701 -113 731
rect -197 663 -172 701
rect -138 663 -113 701
rect -197 629 -113 663
rect -197 595 -172 629
rect -138 595 -113 629
rect -197 561 -113 595
rect -197 523 -172 561
rect -138 523 -113 561
rect -197 493 -113 523
rect -197 451 -172 493
rect -138 451 -113 493
rect -197 425 -113 451
rect -197 379 -172 425
rect -138 379 -113 425
rect -197 357 -113 379
rect -197 307 -172 357
rect -138 307 -113 357
rect -197 289 -113 307
rect -197 235 -172 289
rect -138 235 -113 289
rect -197 221 -113 235
rect -197 163 -172 221
rect -138 163 -113 221
rect -197 153 -113 163
rect -197 91 -172 153
rect -138 91 -113 153
rect -197 85 -113 91
rect -197 19 -172 85
rect -138 19 -113 85
rect -197 17 -113 19
rect -197 -17 -172 17
rect -138 -17 -113 17
rect -197 -19 -113 -17
rect -197 -85 -172 -19
rect -138 -85 -113 -19
rect -197 -91 -113 -85
rect -197 -153 -172 -91
rect -138 -153 -113 -91
rect -197 -163 -113 -153
rect -197 -221 -172 -163
rect -138 -221 -113 -163
rect -197 -235 -113 -221
rect -197 -289 -172 -235
rect -138 -289 -113 -235
rect -197 -307 -113 -289
rect -197 -357 -172 -307
rect -138 -357 -113 -307
rect -197 -379 -113 -357
rect -197 -425 -172 -379
rect -138 -425 -113 -379
rect -197 -451 -113 -425
rect -197 -493 -172 -451
rect -138 -493 -113 -451
rect -197 -523 -113 -493
rect -197 -561 -172 -523
rect -138 -561 -113 -523
rect -197 -595 -113 -561
rect -197 -629 -172 -595
rect -138 -629 -113 -595
rect -197 -663 -113 -629
rect -197 -701 -172 -663
rect -138 -701 -113 -663
rect -197 -731 -113 -701
rect -197 -773 -172 -731
rect -138 -773 -113 -731
rect -197 -799 -113 -773
rect -197 -845 -172 -799
rect -138 -845 -113 -799
rect -197 -867 -113 -845
rect -197 -917 -172 -867
rect -138 -917 -113 -867
rect -197 -935 -113 -917
rect -197 -989 -172 -935
rect -138 -989 -113 -935
rect -197 -1003 -113 -989
rect -197 -1061 -172 -1003
rect -138 -1061 -113 -1003
rect -197 -1071 -113 -1061
rect -197 -1133 -172 -1071
rect -138 -1133 -113 -1071
rect -197 -1139 -113 -1133
rect -197 -1205 -172 -1139
rect -138 -1205 -113 -1139
rect -197 -1207 -113 -1205
rect -197 -1241 -172 -1207
rect -138 -1241 -113 -1207
rect -197 -1243 -113 -1241
rect -197 -1309 -172 -1243
rect -138 -1309 -113 -1243
rect -197 -1315 -113 -1309
rect -197 -1377 -172 -1315
rect -138 -1377 -113 -1315
rect -197 -1387 -113 -1377
rect -197 -1445 -172 -1387
rect -138 -1445 -113 -1387
rect -197 -1459 -113 -1445
rect -197 -1513 -172 -1459
rect -138 -1513 -113 -1459
rect -197 -1531 -113 -1513
rect -197 -1581 -172 -1531
rect -138 -1581 -113 -1531
rect -197 -1603 -113 -1581
rect -197 -1649 -172 -1603
rect -138 -1649 -113 -1603
rect -197 -1675 -113 -1649
rect -197 -1717 -172 -1675
rect -138 -1717 -113 -1675
rect -197 -1747 -113 -1717
rect -197 -1785 -172 -1747
rect -138 -1785 -113 -1747
rect -197 -1810 -113 -1785
rect -17 1785 17 1810
rect -17 1717 17 1747
rect -17 1649 17 1675
rect -17 1581 17 1603
rect -17 1513 17 1531
rect -17 1445 17 1459
rect -17 1377 17 1387
rect -17 1309 17 1315
rect -17 1241 17 1243
rect -17 1205 17 1207
rect -17 1133 17 1139
rect -17 1061 17 1071
rect -17 989 17 1003
rect -17 917 17 935
rect -17 845 17 867
rect -17 773 17 799
rect -17 701 17 731
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 523
rect -17 425 17 451
rect -17 357 17 379
rect -17 289 17 307
rect -17 221 17 235
rect -17 153 17 163
rect -17 85 17 91
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -91 17 -85
rect -17 -163 17 -153
rect -17 -235 17 -221
rect -17 -307 17 -289
rect -17 -379 17 -357
rect -17 -451 17 -425
rect -17 -523 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect -17 -731 17 -701
rect -17 -799 17 -773
rect -17 -867 17 -845
rect -17 -935 17 -917
rect -17 -1003 17 -989
rect -17 -1071 17 -1061
rect -17 -1139 17 -1133
rect -17 -1207 17 -1205
rect -17 -1243 17 -1241
rect -17 -1315 17 -1309
rect -17 -1387 17 -1377
rect -17 -1459 17 -1445
rect -17 -1531 17 -1513
rect -17 -1603 17 -1581
rect -17 -1675 17 -1649
rect -17 -1747 17 -1717
rect -17 -1810 17 -1785
rect 113 1785 147 1810
rect 113 1717 147 1747
rect 113 1649 147 1675
rect 113 1581 147 1603
rect 113 1513 147 1531
rect 113 1445 147 1459
rect 113 1377 147 1387
rect 113 1309 147 1315
rect 113 1241 147 1243
rect 113 1205 147 1207
rect 113 1133 147 1139
rect 113 1061 147 1071
rect 113 989 147 1003
rect 113 917 147 935
rect 113 845 147 867
rect 113 773 147 799
rect 113 701 147 731
rect 113 629 147 663
rect 113 561 147 595
rect 113 493 147 523
rect 113 425 147 451
rect 113 357 147 379
rect 113 289 147 307
rect 113 221 147 235
rect 113 153 147 163
rect 113 85 147 91
rect 113 17 147 19
rect 113 -19 147 -17
rect 113 -91 147 -85
rect 113 -163 147 -153
rect 113 -235 147 -221
rect 113 -307 147 -289
rect 113 -379 147 -357
rect 113 -451 147 -425
rect 113 -523 147 -493
rect 113 -595 147 -561
rect 113 -663 147 -629
rect 113 -731 147 -701
rect 113 -799 147 -773
rect 113 -867 147 -845
rect 113 -935 147 -917
rect 113 -1003 147 -989
rect 113 -1071 147 -1061
rect 113 -1139 147 -1133
rect 113 -1207 147 -1205
rect 113 -1243 147 -1241
rect 113 -1315 147 -1309
rect 113 -1387 147 -1377
rect 113 -1459 147 -1445
rect 113 -1531 147 -1513
rect 113 -1603 147 -1581
rect 113 -1675 147 -1649
rect 113 -1747 147 -1717
rect 113 -1810 147 -1785
rect 243 1785 277 1810
rect 243 1717 277 1747
rect 243 1649 277 1675
rect 243 1581 277 1603
rect 243 1513 277 1531
rect 243 1445 277 1459
rect 243 1377 277 1387
rect 243 1309 277 1315
rect 243 1241 277 1243
rect 243 1205 277 1207
rect 243 1133 277 1139
rect 243 1061 277 1071
rect 243 989 277 1003
rect 243 917 277 935
rect 243 845 277 867
rect 243 773 277 799
rect 243 701 277 731
rect 243 629 277 663
rect 243 561 277 595
rect 243 493 277 523
rect 243 425 277 451
rect 243 357 277 379
rect 243 289 277 307
rect 243 221 277 235
rect 243 153 277 163
rect 243 85 277 91
rect 243 17 277 19
rect 243 -19 277 -17
rect 243 -91 277 -85
rect 243 -163 277 -153
rect 243 -235 277 -221
rect 243 -307 277 -289
rect 243 -379 277 -357
rect 243 -451 277 -425
rect 243 -523 277 -493
rect 243 -595 277 -561
rect 243 -663 277 -629
rect 243 -731 277 -701
rect 243 -799 277 -773
rect 243 -867 277 -845
rect 243 -935 277 -917
rect 243 -1003 277 -989
rect 243 -1071 277 -1061
rect 243 -1139 277 -1133
rect 243 -1207 277 -1205
rect 243 -1243 277 -1241
rect 243 -1315 277 -1309
rect 243 -1387 277 -1377
rect 243 -1459 277 -1445
rect 243 -1531 277 -1513
rect 243 -1603 277 -1581
rect 243 -1675 277 -1649
rect 243 -1747 277 -1717
rect 243 -1810 277 -1785
<< viali >>
rect -262 1844 -228 1878
rect -327 1751 -293 1781
rect -327 1747 -293 1751
rect -327 1683 -293 1709
rect -327 1675 -293 1683
rect -327 1615 -293 1637
rect -327 1603 -293 1615
rect -327 1547 -293 1565
rect -327 1531 -293 1547
rect -327 1479 -293 1493
rect -327 1459 -293 1479
rect -327 1411 -293 1421
rect -327 1387 -293 1411
rect -327 1343 -293 1349
rect -327 1315 -293 1343
rect -327 1275 -293 1277
rect -327 1243 -293 1275
rect -327 1173 -293 1205
rect -327 1171 -293 1173
rect -327 1105 -293 1133
rect -327 1099 -293 1105
rect -327 1037 -293 1061
rect -327 1027 -293 1037
rect -327 969 -293 989
rect -327 955 -293 969
rect -327 901 -293 917
rect -327 883 -293 901
rect -327 833 -293 845
rect -327 811 -293 833
rect -327 765 -293 773
rect -327 739 -293 765
rect -327 697 -293 701
rect -327 667 -293 697
rect -327 595 -293 629
rect -327 527 -293 557
rect -327 523 -293 527
rect -327 459 -293 485
rect -327 451 -293 459
rect -327 391 -293 413
rect -327 379 -293 391
rect -327 323 -293 341
rect -327 307 -293 323
rect -327 255 -293 269
rect -327 235 -293 255
rect -327 187 -293 197
rect -327 163 -293 187
rect -327 119 -293 125
rect -327 91 -293 119
rect -327 51 -293 53
rect -327 19 -293 51
rect -327 -51 -293 -19
rect -327 -53 -293 -51
rect -327 -119 -293 -91
rect -327 -125 -293 -119
rect -327 -187 -293 -163
rect -327 -197 -293 -187
rect -327 -255 -293 -235
rect -327 -269 -293 -255
rect -327 -323 -293 -307
rect -327 -341 -293 -323
rect -327 -391 -293 -379
rect -327 -413 -293 -391
rect -327 -459 -293 -451
rect -327 -485 -293 -459
rect -327 -527 -293 -523
rect -327 -557 -293 -527
rect -327 -629 -293 -595
rect -327 -697 -293 -667
rect -327 -701 -293 -697
rect -327 -765 -293 -739
rect -327 -773 -293 -765
rect -327 -833 -293 -811
rect -327 -845 -293 -833
rect -327 -901 -293 -883
rect -327 -917 -293 -901
rect -327 -969 -293 -955
rect -327 -989 -293 -969
rect -327 -1037 -293 -1027
rect -327 -1061 -293 -1037
rect -327 -1105 -293 -1099
rect -327 -1133 -293 -1105
rect -327 -1173 -293 -1171
rect -327 -1205 -293 -1173
rect -327 -1275 -293 -1243
rect -327 -1277 -293 -1275
rect -327 -1343 -293 -1315
rect -327 -1349 -293 -1343
rect -327 -1411 -293 -1387
rect -327 -1421 -293 -1411
rect -327 -1479 -293 -1459
rect -327 -1493 -293 -1479
rect -327 -1547 -293 -1531
rect -327 -1565 -293 -1547
rect -327 -1615 -293 -1603
rect -327 -1637 -293 -1615
rect -327 -1683 -293 -1675
rect -327 -1709 -293 -1683
rect -327 -1751 -293 -1747
rect -327 -1781 -293 -1751
rect -172 1751 -138 1781
rect -172 1747 -138 1751
rect -172 1683 -138 1709
rect -172 1675 -138 1683
rect -172 1615 -138 1637
rect -172 1603 -138 1615
rect -172 1547 -138 1565
rect -172 1531 -138 1547
rect -172 1479 -138 1493
rect -172 1459 -138 1479
rect -172 1411 -138 1421
rect -172 1387 -138 1411
rect -172 1343 -138 1349
rect -172 1315 -138 1343
rect -172 1275 -138 1277
rect -172 1243 -138 1275
rect -172 1173 -138 1205
rect -172 1171 -138 1173
rect -172 1105 -138 1133
rect -172 1099 -138 1105
rect -172 1037 -138 1061
rect -172 1027 -138 1037
rect -172 969 -138 989
rect -172 955 -138 969
rect -172 901 -138 917
rect -172 883 -138 901
rect -172 833 -138 845
rect -172 811 -138 833
rect -172 765 -138 773
rect -172 739 -138 765
rect -172 697 -138 701
rect -172 667 -138 697
rect -172 595 -138 629
rect -172 527 -138 557
rect -172 523 -138 527
rect -172 459 -138 485
rect -172 451 -138 459
rect -172 391 -138 413
rect -172 379 -138 391
rect -172 323 -138 341
rect -172 307 -138 323
rect -172 255 -138 269
rect -172 235 -138 255
rect -172 187 -138 197
rect -172 163 -138 187
rect -172 119 -138 125
rect -172 91 -138 119
rect -172 51 -138 53
rect -172 19 -138 51
rect -172 -51 -138 -19
rect -172 -53 -138 -51
rect -172 -119 -138 -91
rect -172 -125 -138 -119
rect -172 -187 -138 -163
rect -172 -197 -138 -187
rect -172 -255 -138 -235
rect -172 -269 -138 -255
rect -172 -323 -138 -307
rect -172 -341 -138 -323
rect -172 -391 -138 -379
rect -172 -413 -138 -391
rect -172 -459 -138 -451
rect -172 -485 -138 -459
rect -172 -527 -138 -523
rect -172 -557 -138 -527
rect -172 -629 -138 -595
rect -172 -697 -138 -667
rect -172 -701 -138 -697
rect -172 -765 -138 -739
rect -172 -773 -138 -765
rect -172 -833 -138 -811
rect -172 -845 -138 -833
rect -172 -901 -138 -883
rect -172 -917 -138 -901
rect -172 -969 -138 -955
rect -172 -989 -138 -969
rect -172 -1037 -138 -1027
rect -172 -1061 -138 -1037
rect -172 -1105 -138 -1099
rect -172 -1133 -138 -1105
rect -172 -1173 -138 -1171
rect -172 -1205 -138 -1173
rect -172 -1275 -138 -1243
rect -172 -1277 -138 -1275
rect -172 -1343 -138 -1315
rect -172 -1349 -138 -1343
rect -172 -1411 -138 -1387
rect -172 -1421 -138 -1411
rect -172 -1479 -138 -1459
rect -172 -1493 -138 -1479
rect -172 -1547 -138 -1531
rect -172 -1565 -138 -1547
rect -172 -1615 -138 -1603
rect -172 -1637 -138 -1615
rect -172 -1683 -138 -1675
rect -172 -1709 -138 -1683
rect -172 -1751 -138 -1747
rect -172 -1781 -138 -1751
rect -17 1751 17 1781
rect -17 1747 17 1751
rect -17 1683 17 1709
rect -17 1675 17 1683
rect -17 1615 17 1637
rect -17 1603 17 1615
rect -17 1547 17 1565
rect -17 1531 17 1547
rect -17 1479 17 1493
rect -17 1459 17 1479
rect -17 1411 17 1421
rect -17 1387 17 1411
rect -17 1343 17 1349
rect -17 1315 17 1343
rect -17 1275 17 1277
rect -17 1243 17 1275
rect -17 1173 17 1205
rect -17 1171 17 1173
rect -17 1105 17 1133
rect -17 1099 17 1105
rect -17 1037 17 1061
rect -17 1027 17 1037
rect -17 969 17 989
rect -17 955 17 969
rect -17 901 17 917
rect -17 883 17 901
rect -17 833 17 845
rect -17 811 17 833
rect -17 765 17 773
rect -17 739 17 765
rect -17 697 17 701
rect -17 667 17 697
rect -17 595 17 629
rect -17 527 17 557
rect -17 523 17 527
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect -17 -527 17 -523
rect -17 -557 17 -527
rect -17 -629 17 -595
rect -17 -697 17 -667
rect -17 -701 17 -697
rect -17 -765 17 -739
rect -17 -773 17 -765
rect -17 -833 17 -811
rect -17 -845 17 -833
rect -17 -901 17 -883
rect -17 -917 17 -901
rect -17 -969 17 -955
rect -17 -989 17 -969
rect -17 -1037 17 -1027
rect -17 -1061 17 -1037
rect -17 -1105 17 -1099
rect -17 -1133 17 -1105
rect -17 -1173 17 -1171
rect -17 -1205 17 -1173
rect -17 -1275 17 -1243
rect -17 -1277 17 -1275
rect -17 -1343 17 -1315
rect -17 -1349 17 -1343
rect -17 -1411 17 -1387
rect -17 -1421 17 -1411
rect -17 -1479 17 -1459
rect -17 -1493 17 -1479
rect -17 -1547 17 -1531
rect -17 -1565 17 -1547
rect -17 -1615 17 -1603
rect -17 -1637 17 -1615
rect -17 -1683 17 -1675
rect -17 -1709 17 -1683
rect -17 -1751 17 -1747
rect -17 -1781 17 -1751
rect 113 1751 147 1781
rect 113 1747 147 1751
rect 113 1683 147 1709
rect 113 1675 147 1683
rect 113 1615 147 1637
rect 113 1603 147 1615
rect 113 1547 147 1565
rect 113 1531 147 1547
rect 113 1479 147 1493
rect 113 1459 147 1479
rect 113 1411 147 1421
rect 113 1387 147 1411
rect 113 1343 147 1349
rect 113 1315 147 1343
rect 113 1275 147 1277
rect 113 1243 147 1275
rect 113 1173 147 1205
rect 113 1171 147 1173
rect 113 1105 147 1133
rect 113 1099 147 1105
rect 113 1037 147 1061
rect 113 1027 147 1037
rect 113 969 147 989
rect 113 955 147 969
rect 113 901 147 917
rect 113 883 147 901
rect 113 833 147 845
rect 113 811 147 833
rect 113 765 147 773
rect 113 739 147 765
rect 113 697 147 701
rect 113 667 147 697
rect 113 595 147 629
rect 113 527 147 557
rect 113 523 147 527
rect 113 459 147 485
rect 113 451 147 459
rect 113 391 147 413
rect 113 379 147 391
rect 113 323 147 341
rect 113 307 147 323
rect 113 255 147 269
rect 113 235 147 255
rect 113 187 147 197
rect 113 163 147 187
rect 113 119 147 125
rect 113 91 147 119
rect 113 51 147 53
rect 113 19 147 51
rect 113 -51 147 -19
rect 113 -53 147 -51
rect 113 -119 147 -91
rect 113 -125 147 -119
rect 113 -187 147 -163
rect 113 -197 147 -187
rect 113 -255 147 -235
rect 113 -269 147 -255
rect 113 -323 147 -307
rect 113 -341 147 -323
rect 113 -391 147 -379
rect 113 -413 147 -391
rect 113 -459 147 -451
rect 113 -485 147 -459
rect 113 -527 147 -523
rect 113 -557 147 -527
rect 113 -629 147 -595
rect 113 -697 147 -667
rect 113 -701 147 -697
rect 113 -765 147 -739
rect 113 -773 147 -765
rect 113 -833 147 -811
rect 113 -845 147 -833
rect 113 -901 147 -883
rect 113 -917 147 -901
rect 113 -969 147 -955
rect 113 -989 147 -969
rect 113 -1037 147 -1027
rect 113 -1061 147 -1037
rect 113 -1105 147 -1099
rect 113 -1133 147 -1105
rect 113 -1173 147 -1171
rect 113 -1205 147 -1173
rect 113 -1275 147 -1243
rect 113 -1277 147 -1275
rect 113 -1343 147 -1315
rect 113 -1349 147 -1343
rect 113 -1411 147 -1387
rect 113 -1421 147 -1411
rect 113 -1479 147 -1459
rect 113 -1493 147 -1479
rect 113 -1547 147 -1531
rect 113 -1565 147 -1547
rect 113 -1615 147 -1603
rect 113 -1637 147 -1615
rect 113 -1683 147 -1675
rect 113 -1709 147 -1683
rect 113 -1751 147 -1747
rect 113 -1781 147 -1751
rect 243 1751 277 1781
rect 243 1747 277 1751
rect 243 1683 277 1709
rect 243 1675 277 1683
rect 243 1615 277 1637
rect 243 1603 277 1615
rect 243 1547 277 1565
rect 243 1531 277 1547
rect 243 1479 277 1493
rect 243 1459 277 1479
rect 243 1411 277 1421
rect 243 1387 277 1411
rect 243 1343 277 1349
rect 243 1315 277 1343
rect 243 1275 277 1277
rect 243 1243 277 1275
rect 243 1173 277 1205
rect 243 1171 277 1173
rect 243 1105 277 1133
rect 243 1099 277 1105
rect 243 1037 277 1061
rect 243 1027 277 1037
rect 243 969 277 989
rect 243 955 277 969
rect 243 901 277 917
rect 243 883 277 901
rect 243 833 277 845
rect 243 811 277 833
rect 243 765 277 773
rect 243 739 277 765
rect 243 697 277 701
rect 243 667 277 697
rect 243 595 277 629
rect 243 527 277 557
rect 243 523 277 527
rect 243 459 277 485
rect 243 451 277 459
rect 243 391 277 413
rect 243 379 277 391
rect 243 323 277 341
rect 243 307 277 323
rect 243 255 277 269
rect 243 235 277 255
rect 243 187 277 197
rect 243 163 277 187
rect 243 119 277 125
rect 243 91 277 119
rect 243 51 277 53
rect 243 19 277 51
rect 243 -51 277 -19
rect 243 -53 277 -51
rect 243 -119 277 -91
rect 243 -125 277 -119
rect 243 -187 277 -163
rect 243 -197 277 -187
rect 243 -255 277 -235
rect 243 -269 277 -255
rect 243 -323 277 -307
rect 243 -341 277 -323
rect 243 -391 277 -379
rect 243 -413 277 -391
rect 243 -459 277 -451
rect 243 -485 277 -459
rect 243 -527 277 -523
rect 243 -557 277 -527
rect 243 -629 277 -595
rect 243 -697 277 -667
rect 243 -701 277 -697
rect 243 -765 277 -739
rect 243 -773 277 -765
rect 243 -833 277 -811
rect 243 -845 277 -833
rect 243 -901 277 -883
rect 243 -917 277 -901
rect 243 -969 277 -955
rect 243 -989 277 -969
rect 243 -1037 277 -1027
rect 243 -1061 277 -1037
rect 243 -1105 277 -1099
rect 243 -1133 277 -1105
rect 243 -1173 277 -1171
rect 243 -1205 277 -1173
rect 243 -1275 277 -1243
rect 243 -1277 277 -1275
rect 243 -1343 277 -1315
rect 243 -1349 277 -1343
rect 243 -1411 277 -1387
rect 243 -1421 277 -1411
rect 243 -1479 277 -1459
rect 243 -1493 277 -1479
rect 243 -1547 277 -1531
rect 243 -1565 277 -1547
rect 243 -1615 277 -1603
rect 243 -1637 277 -1615
rect 243 -1683 277 -1675
rect 243 -1709 277 -1683
rect 243 -1751 277 -1747
rect 243 -1781 277 -1751
<< metal1 >>
rect -277 1878 -213 1884
rect -277 1844 -262 1878
rect -228 1844 -213 1878
rect -277 1838 -213 1844
rect -333 1781 -287 1806
rect -333 1747 -327 1781
rect -293 1747 -287 1781
rect -333 1709 -287 1747
rect -333 1675 -327 1709
rect -293 1675 -287 1709
rect -333 1637 -287 1675
rect -333 1603 -327 1637
rect -293 1603 -287 1637
rect -333 1565 -287 1603
rect -333 1531 -327 1565
rect -293 1531 -287 1565
rect -333 1493 -287 1531
rect -333 1459 -327 1493
rect -293 1459 -287 1493
rect -333 1421 -287 1459
rect -333 1387 -327 1421
rect -293 1387 -287 1421
rect -333 1349 -287 1387
rect -333 1315 -327 1349
rect -293 1315 -287 1349
rect -333 1277 -287 1315
rect -333 1243 -327 1277
rect -293 1243 -287 1277
rect -333 1205 -287 1243
rect -333 1171 -327 1205
rect -293 1171 -287 1205
rect -333 1133 -287 1171
rect -333 1099 -327 1133
rect -293 1099 -287 1133
rect -333 1061 -287 1099
rect -333 1027 -327 1061
rect -293 1027 -287 1061
rect -333 989 -287 1027
rect -333 955 -327 989
rect -293 955 -287 989
rect -333 917 -287 955
rect -333 883 -327 917
rect -293 883 -287 917
rect -333 845 -287 883
rect -333 811 -327 845
rect -293 811 -287 845
rect -333 773 -287 811
rect -333 739 -327 773
rect -293 739 -287 773
rect -333 701 -287 739
rect -333 667 -327 701
rect -293 667 -287 701
rect -333 629 -287 667
rect -333 595 -327 629
rect -293 595 -287 629
rect -333 557 -287 595
rect -333 523 -327 557
rect -293 523 -287 557
rect -333 485 -287 523
rect -333 451 -327 485
rect -293 451 -287 485
rect -333 413 -287 451
rect -333 379 -327 413
rect -293 379 -287 413
rect -333 341 -287 379
rect -333 307 -327 341
rect -293 307 -287 341
rect -333 269 -287 307
rect -333 235 -327 269
rect -293 235 -287 269
rect -333 197 -287 235
rect -333 163 -327 197
rect -293 163 -287 197
rect -333 125 -287 163
rect -333 91 -327 125
rect -293 91 -287 125
rect -333 53 -287 91
rect -333 19 -327 53
rect -293 19 -287 53
rect -333 -19 -287 19
rect -333 -53 -327 -19
rect -293 -53 -287 -19
rect -333 -91 -287 -53
rect -333 -125 -327 -91
rect -293 -125 -287 -91
rect -333 -163 -287 -125
rect -333 -197 -327 -163
rect -293 -197 -287 -163
rect -333 -235 -287 -197
rect -333 -269 -327 -235
rect -293 -269 -287 -235
rect -333 -307 -287 -269
rect -333 -341 -327 -307
rect -293 -341 -287 -307
rect -333 -379 -287 -341
rect -333 -413 -327 -379
rect -293 -413 -287 -379
rect -333 -451 -287 -413
rect -333 -485 -327 -451
rect -293 -485 -287 -451
rect -333 -523 -287 -485
rect -333 -557 -327 -523
rect -293 -557 -287 -523
rect -333 -595 -287 -557
rect -333 -629 -327 -595
rect -293 -629 -287 -595
rect -333 -667 -287 -629
rect -333 -701 -327 -667
rect -293 -701 -287 -667
rect -333 -739 -287 -701
rect -333 -773 -327 -739
rect -293 -773 -287 -739
rect -333 -811 -287 -773
rect -333 -845 -327 -811
rect -293 -845 -287 -811
rect -333 -883 -287 -845
rect -333 -917 -327 -883
rect -293 -917 -287 -883
rect -333 -955 -287 -917
rect -333 -989 -327 -955
rect -293 -989 -287 -955
rect -333 -1027 -287 -989
rect -333 -1061 -327 -1027
rect -293 -1061 -287 -1027
rect -333 -1099 -287 -1061
rect -333 -1133 -327 -1099
rect -293 -1133 -287 -1099
rect -333 -1171 -287 -1133
rect -333 -1205 -327 -1171
rect -293 -1205 -287 -1171
rect -333 -1243 -287 -1205
rect -333 -1277 -327 -1243
rect -293 -1277 -287 -1243
rect -333 -1315 -287 -1277
rect -333 -1349 -327 -1315
rect -293 -1349 -287 -1315
rect -333 -1387 -287 -1349
rect -333 -1421 -327 -1387
rect -293 -1421 -287 -1387
rect -333 -1459 -287 -1421
rect -333 -1493 -327 -1459
rect -293 -1493 -287 -1459
rect -333 -1531 -287 -1493
rect -333 -1565 -327 -1531
rect -293 -1565 -287 -1531
rect -333 -1603 -287 -1565
rect -333 -1637 -327 -1603
rect -293 -1637 -287 -1603
rect -333 -1675 -287 -1637
rect -333 -1709 -327 -1675
rect -293 -1709 -287 -1675
rect -333 -1747 -287 -1709
rect -333 -1781 -327 -1747
rect -293 -1781 -287 -1747
rect -333 -1806 -287 -1781
rect -203 1781 -107 1806
rect -203 1747 -172 1781
rect -138 1747 -107 1781
rect -203 1709 -107 1747
rect -203 1675 -172 1709
rect -138 1675 -107 1709
rect -203 1637 -107 1675
rect -203 1603 -172 1637
rect -138 1603 -107 1637
rect -203 1565 -107 1603
rect -203 1531 -172 1565
rect -138 1531 -107 1565
rect -203 1493 -107 1531
rect -203 1459 -172 1493
rect -138 1459 -107 1493
rect -203 1421 -107 1459
rect -203 1387 -172 1421
rect -138 1387 -107 1421
rect -203 1349 -107 1387
rect -203 1315 -172 1349
rect -138 1315 -107 1349
rect -203 1277 -107 1315
rect -203 1243 -172 1277
rect -138 1243 -107 1277
rect -203 1205 -107 1243
rect -203 1171 -172 1205
rect -138 1171 -107 1205
rect -203 1133 -107 1171
rect -203 1099 -172 1133
rect -138 1099 -107 1133
rect -203 1061 -107 1099
rect -203 1027 -172 1061
rect -138 1027 -107 1061
rect -203 989 -107 1027
rect -203 955 -172 989
rect -138 955 -107 989
rect -203 917 -107 955
rect -203 883 -172 917
rect -138 883 -107 917
rect -203 845 -107 883
rect -203 811 -172 845
rect -138 811 -107 845
rect -203 773 -107 811
rect -203 739 -172 773
rect -138 739 -107 773
rect -203 701 -107 739
rect -203 667 -172 701
rect -138 667 -107 701
rect -203 629 -107 667
rect -203 595 -172 629
rect -138 595 -107 629
rect -203 557 -107 595
rect -203 523 -172 557
rect -138 523 -107 557
rect -203 485 -107 523
rect -203 451 -172 485
rect -138 451 -107 485
rect -203 413 -107 451
rect -203 379 -172 413
rect -138 379 -107 413
rect -203 341 -107 379
rect -203 307 -172 341
rect -138 307 -107 341
rect -203 269 -107 307
rect -203 235 -172 269
rect -138 235 -107 269
rect -203 197 -107 235
rect -203 163 -172 197
rect -138 163 -107 197
rect -203 125 -107 163
rect -203 91 -172 125
rect -138 91 -107 125
rect -203 53 -107 91
rect -203 19 -172 53
rect -138 19 -107 53
rect -203 -19 -107 19
rect -203 -53 -172 -19
rect -138 -53 -107 -19
rect -203 -91 -107 -53
rect -203 -125 -172 -91
rect -138 -125 -107 -91
rect -203 -163 -107 -125
rect -203 -197 -172 -163
rect -138 -197 -107 -163
rect -203 -235 -107 -197
rect -203 -269 -172 -235
rect -138 -269 -107 -235
rect -203 -307 -107 -269
rect -203 -341 -172 -307
rect -138 -341 -107 -307
rect -203 -379 -107 -341
rect -203 -413 -172 -379
rect -138 -413 -107 -379
rect -203 -451 -107 -413
rect -203 -485 -172 -451
rect -138 -485 -107 -451
rect -203 -523 -107 -485
rect -203 -557 -172 -523
rect -138 -557 -107 -523
rect -203 -595 -107 -557
rect -203 -629 -172 -595
rect -138 -629 -107 -595
rect -203 -667 -107 -629
rect -203 -701 -172 -667
rect -138 -701 -107 -667
rect -203 -739 -107 -701
rect -203 -773 -172 -739
rect -138 -773 -107 -739
rect -203 -811 -107 -773
rect -203 -845 -172 -811
rect -138 -845 -107 -811
rect -203 -883 -107 -845
rect -203 -917 -172 -883
rect -138 -917 -107 -883
rect -203 -955 -107 -917
rect -203 -989 -172 -955
rect -138 -989 -107 -955
rect -203 -1027 -107 -989
rect -203 -1061 -172 -1027
rect -138 -1061 -107 -1027
rect -203 -1099 -107 -1061
rect -203 -1133 -172 -1099
rect -138 -1133 -107 -1099
rect -203 -1171 -107 -1133
rect -203 -1205 -172 -1171
rect -138 -1205 -107 -1171
rect -203 -1243 -107 -1205
rect -203 -1277 -172 -1243
rect -138 -1277 -107 -1243
rect -203 -1315 -107 -1277
rect -203 -1349 -172 -1315
rect -138 -1349 -107 -1315
rect -203 -1387 -107 -1349
rect -203 -1421 -172 -1387
rect -138 -1421 -107 -1387
rect -203 -1459 -107 -1421
rect -203 -1493 -172 -1459
rect -138 -1493 -107 -1459
rect -203 -1531 -107 -1493
rect -203 -1565 -172 -1531
rect -138 -1565 -107 -1531
rect -203 -1603 -107 -1565
rect -203 -1637 -172 -1603
rect -138 -1637 -107 -1603
rect -203 -1675 -107 -1637
rect -203 -1709 -172 -1675
rect -138 -1709 -107 -1675
rect -203 -1747 -107 -1709
rect -203 -1781 -172 -1747
rect -138 -1781 -107 -1747
rect -203 -1806 -107 -1781
rect -23 1781 23 1806
rect -23 1747 -17 1781
rect 17 1747 23 1781
rect -23 1709 23 1747
rect -23 1675 -17 1709
rect 17 1675 23 1709
rect -23 1637 23 1675
rect -23 1603 -17 1637
rect 17 1603 23 1637
rect -23 1565 23 1603
rect -23 1531 -17 1565
rect 17 1531 23 1565
rect -23 1493 23 1531
rect -23 1459 -17 1493
rect 17 1459 23 1493
rect -23 1421 23 1459
rect -23 1387 -17 1421
rect 17 1387 23 1421
rect -23 1349 23 1387
rect -23 1315 -17 1349
rect 17 1315 23 1349
rect -23 1277 23 1315
rect -23 1243 -17 1277
rect 17 1243 23 1277
rect -23 1205 23 1243
rect -23 1171 -17 1205
rect 17 1171 23 1205
rect -23 1133 23 1171
rect -23 1099 -17 1133
rect 17 1099 23 1133
rect -23 1061 23 1099
rect -23 1027 -17 1061
rect 17 1027 23 1061
rect -23 989 23 1027
rect -23 955 -17 989
rect 17 955 23 989
rect -23 917 23 955
rect -23 883 -17 917
rect 17 883 23 917
rect -23 845 23 883
rect -23 811 -17 845
rect 17 811 23 845
rect -23 773 23 811
rect -23 739 -17 773
rect 17 739 23 773
rect -23 701 23 739
rect -23 667 -17 701
rect 17 667 23 701
rect -23 629 23 667
rect -23 595 -17 629
rect 17 595 23 629
rect -23 557 23 595
rect -23 523 -17 557
rect 17 523 23 557
rect -23 485 23 523
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -523 23 -485
rect -23 -557 -17 -523
rect 17 -557 23 -523
rect -23 -595 23 -557
rect -23 -629 -17 -595
rect 17 -629 23 -595
rect -23 -667 23 -629
rect -23 -701 -17 -667
rect 17 -701 23 -667
rect -23 -739 23 -701
rect -23 -773 -17 -739
rect 17 -773 23 -739
rect -23 -811 23 -773
rect -23 -845 -17 -811
rect 17 -845 23 -811
rect -23 -883 23 -845
rect -23 -917 -17 -883
rect 17 -917 23 -883
rect -23 -955 23 -917
rect -23 -989 -17 -955
rect 17 -989 23 -955
rect -23 -1027 23 -989
rect -23 -1061 -17 -1027
rect 17 -1061 23 -1027
rect -23 -1099 23 -1061
rect -23 -1133 -17 -1099
rect 17 -1133 23 -1099
rect -23 -1171 23 -1133
rect -23 -1205 -17 -1171
rect 17 -1205 23 -1171
rect -23 -1243 23 -1205
rect -23 -1277 -17 -1243
rect 17 -1277 23 -1243
rect -23 -1315 23 -1277
rect -23 -1349 -17 -1315
rect 17 -1349 23 -1315
rect -23 -1387 23 -1349
rect -23 -1421 -17 -1387
rect 17 -1421 23 -1387
rect -23 -1459 23 -1421
rect -23 -1493 -17 -1459
rect 17 -1493 23 -1459
rect -23 -1531 23 -1493
rect -23 -1565 -17 -1531
rect 17 -1565 23 -1531
rect -23 -1603 23 -1565
rect -23 -1637 -17 -1603
rect 17 -1637 23 -1603
rect -23 -1675 23 -1637
rect -23 -1709 -17 -1675
rect 17 -1709 23 -1675
rect -23 -1747 23 -1709
rect -23 -1781 -17 -1747
rect 17 -1781 23 -1747
rect -23 -1806 23 -1781
rect 107 1781 153 1806
rect 107 1747 113 1781
rect 147 1747 153 1781
rect 107 1709 153 1747
rect 107 1675 113 1709
rect 147 1675 153 1709
rect 107 1637 153 1675
rect 107 1603 113 1637
rect 147 1603 153 1637
rect 107 1565 153 1603
rect 107 1531 113 1565
rect 147 1531 153 1565
rect 107 1493 153 1531
rect 107 1459 113 1493
rect 147 1459 153 1493
rect 107 1421 153 1459
rect 107 1387 113 1421
rect 147 1387 153 1421
rect 107 1349 153 1387
rect 107 1315 113 1349
rect 147 1315 153 1349
rect 107 1277 153 1315
rect 107 1243 113 1277
rect 147 1243 153 1277
rect 107 1205 153 1243
rect 107 1171 113 1205
rect 147 1171 153 1205
rect 107 1133 153 1171
rect 107 1099 113 1133
rect 147 1099 153 1133
rect 107 1061 153 1099
rect 107 1027 113 1061
rect 147 1027 153 1061
rect 107 989 153 1027
rect 107 955 113 989
rect 147 955 153 989
rect 107 917 153 955
rect 107 883 113 917
rect 147 883 153 917
rect 107 845 153 883
rect 107 811 113 845
rect 147 811 153 845
rect 107 773 153 811
rect 107 739 113 773
rect 147 739 153 773
rect 107 701 153 739
rect 107 667 113 701
rect 147 667 153 701
rect 107 629 153 667
rect 107 595 113 629
rect 147 595 153 629
rect 107 557 153 595
rect 107 523 113 557
rect 147 523 153 557
rect 107 485 153 523
rect 107 451 113 485
rect 147 451 153 485
rect 107 413 153 451
rect 107 379 113 413
rect 147 379 153 413
rect 107 341 153 379
rect 107 307 113 341
rect 147 307 153 341
rect 107 269 153 307
rect 107 235 113 269
rect 147 235 153 269
rect 107 197 153 235
rect 107 163 113 197
rect 147 163 153 197
rect 107 125 153 163
rect 107 91 113 125
rect 147 91 153 125
rect 107 53 153 91
rect 107 19 113 53
rect 147 19 153 53
rect 107 -19 153 19
rect 107 -53 113 -19
rect 147 -53 153 -19
rect 107 -91 153 -53
rect 107 -125 113 -91
rect 147 -125 153 -91
rect 107 -163 153 -125
rect 107 -197 113 -163
rect 147 -197 153 -163
rect 107 -235 153 -197
rect 107 -269 113 -235
rect 147 -269 153 -235
rect 107 -307 153 -269
rect 107 -341 113 -307
rect 147 -341 153 -307
rect 107 -379 153 -341
rect 107 -413 113 -379
rect 147 -413 153 -379
rect 107 -451 153 -413
rect 107 -485 113 -451
rect 147 -485 153 -451
rect 107 -523 153 -485
rect 107 -557 113 -523
rect 147 -557 153 -523
rect 107 -595 153 -557
rect 107 -629 113 -595
rect 147 -629 153 -595
rect 107 -667 153 -629
rect 107 -701 113 -667
rect 147 -701 153 -667
rect 107 -739 153 -701
rect 107 -773 113 -739
rect 147 -773 153 -739
rect 107 -811 153 -773
rect 107 -845 113 -811
rect 147 -845 153 -811
rect 107 -883 153 -845
rect 107 -917 113 -883
rect 147 -917 153 -883
rect 107 -955 153 -917
rect 107 -989 113 -955
rect 147 -989 153 -955
rect 107 -1027 153 -989
rect 107 -1061 113 -1027
rect 147 -1061 153 -1027
rect 107 -1099 153 -1061
rect 107 -1133 113 -1099
rect 147 -1133 153 -1099
rect 107 -1171 153 -1133
rect 107 -1205 113 -1171
rect 147 -1205 153 -1171
rect 107 -1243 153 -1205
rect 107 -1277 113 -1243
rect 147 -1277 153 -1243
rect 107 -1315 153 -1277
rect 107 -1349 113 -1315
rect 147 -1349 153 -1315
rect 107 -1387 153 -1349
rect 107 -1421 113 -1387
rect 147 -1421 153 -1387
rect 107 -1459 153 -1421
rect 107 -1493 113 -1459
rect 147 -1493 153 -1459
rect 107 -1531 153 -1493
rect 107 -1565 113 -1531
rect 147 -1565 153 -1531
rect 107 -1603 153 -1565
rect 107 -1637 113 -1603
rect 147 -1637 153 -1603
rect 107 -1675 153 -1637
rect 107 -1709 113 -1675
rect 147 -1709 153 -1675
rect 107 -1747 153 -1709
rect 107 -1781 113 -1747
rect 147 -1781 153 -1747
rect 107 -1806 153 -1781
rect 237 1781 283 1806
rect 237 1747 243 1781
rect 277 1747 283 1781
rect 237 1709 283 1747
rect 237 1675 243 1709
rect 277 1675 283 1709
rect 237 1637 283 1675
rect 237 1603 243 1637
rect 277 1603 283 1637
rect 237 1565 283 1603
rect 237 1531 243 1565
rect 277 1531 283 1565
rect 237 1493 283 1531
rect 237 1459 243 1493
rect 277 1459 283 1493
rect 237 1421 283 1459
rect 237 1387 243 1421
rect 277 1387 283 1421
rect 237 1349 283 1387
rect 237 1315 243 1349
rect 277 1315 283 1349
rect 237 1277 283 1315
rect 237 1243 243 1277
rect 277 1243 283 1277
rect 237 1205 283 1243
rect 237 1171 243 1205
rect 277 1171 283 1205
rect 237 1133 283 1171
rect 237 1099 243 1133
rect 277 1099 283 1133
rect 237 1061 283 1099
rect 237 1027 243 1061
rect 277 1027 283 1061
rect 237 989 283 1027
rect 237 955 243 989
rect 277 955 283 989
rect 237 917 283 955
rect 237 883 243 917
rect 277 883 283 917
rect 237 845 283 883
rect 237 811 243 845
rect 277 811 283 845
rect 237 773 283 811
rect 237 739 243 773
rect 277 739 283 773
rect 237 701 283 739
rect 237 667 243 701
rect 277 667 283 701
rect 237 629 283 667
rect 237 595 243 629
rect 277 595 283 629
rect 237 557 283 595
rect 237 523 243 557
rect 277 523 283 557
rect 237 485 283 523
rect 237 451 243 485
rect 277 451 283 485
rect 237 413 283 451
rect 237 379 243 413
rect 277 379 283 413
rect 237 341 283 379
rect 237 307 243 341
rect 277 307 283 341
rect 237 269 283 307
rect 237 235 243 269
rect 277 235 283 269
rect 237 197 283 235
rect 237 163 243 197
rect 277 163 283 197
rect 237 125 283 163
rect 237 91 243 125
rect 277 91 283 125
rect 237 53 283 91
rect 237 19 243 53
rect 277 19 283 53
rect 237 -19 283 19
rect 237 -53 243 -19
rect 277 -53 283 -19
rect 237 -91 283 -53
rect 237 -125 243 -91
rect 277 -125 283 -91
rect 237 -163 283 -125
rect 237 -197 243 -163
rect 277 -197 283 -163
rect 237 -235 283 -197
rect 237 -269 243 -235
rect 277 -269 283 -235
rect 237 -307 283 -269
rect 237 -341 243 -307
rect 277 -341 283 -307
rect 237 -379 283 -341
rect 237 -413 243 -379
rect 277 -413 283 -379
rect 237 -451 283 -413
rect 237 -485 243 -451
rect 277 -485 283 -451
rect 237 -523 283 -485
rect 237 -557 243 -523
rect 277 -557 283 -523
rect 237 -595 283 -557
rect 237 -629 243 -595
rect 277 -629 283 -595
rect 237 -667 283 -629
rect 237 -701 243 -667
rect 277 -701 283 -667
rect 237 -739 283 -701
rect 237 -773 243 -739
rect 277 -773 283 -739
rect 237 -811 283 -773
rect 237 -845 243 -811
rect 277 -845 283 -811
rect 237 -883 283 -845
rect 237 -917 243 -883
rect 277 -917 283 -883
rect 237 -955 283 -917
rect 237 -989 243 -955
rect 277 -989 283 -955
rect 237 -1027 283 -989
rect 237 -1061 243 -1027
rect 277 -1061 283 -1027
rect 237 -1099 283 -1061
rect 237 -1133 243 -1099
rect 277 -1133 283 -1099
rect 237 -1171 283 -1133
rect 237 -1205 243 -1171
rect 277 -1205 283 -1171
rect 237 -1243 283 -1205
rect 237 -1277 243 -1243
rect 277 -1277 283 -1243
rect 237 -1315 283 -1277
rect 237 -1349 243 -1315
rect 277 -1349 283 -1315
rect 237 -1387 283 -1349
rect 237 -1421 243 -1387
rect 277 -1421 283 -1387
rect 237 -1459 283 -1421
rect 237 -1493 243 -1459
rect 277 -1493 283 -1459
rect 237 -1531 283 -1493
rect 237 -1565 243 -1531
rect 277 -1565 283 -1531
rect 237 -1603 283 -1565
rect 237 -1637 243 -1603
rect 277 -1637 283 -1603
rect 237 -1675 283 -1637
rect 237 -1709 243 -1675
rect 277 -1709 283 -1675
rect 237 -1747 283 -1709
rect 237 -1781 243 -1747
rect 277 -1781 283 -1747
rect 237 -1806 283 -1781
<< end >>
