magic
tech sky130A
magscale 1 2
timestamp 1667951016
<< error_p >>
rect -29 341 29 347
rect -29 307 -17 341
rect -29 301 29 307
<< nmos >>
rect -30 -331 30 269
<< ndiff >>
rect -88 257 -30 269
rect -88 -319 -76 257
rect -42 -319 -30 257
rect -88 -331 -30 -319
rect 30 257 88 269
rect 30 -319 42 257
rect 76 -319 88 257
rect 30 -331 88 -319
<< ndiffc >>
rect -76 -319 -42 257
rect 42 -319 76 257
<< poly >>
rect -33 341 33 357
rect -33 307 -17 341
rect 17 307 33 341
rect -33 291 33 307
rect -30 269 30 291
rect -30 -357 30 -331
<< polycont >>
rect -17 307 17 341
<< locali >>
rect -33 307 -17 341
rect 17 307 33 341
rect -76 257 -42 273
rect -76 -335 -42 -319
rect 42 257 76 273
rect 42 -335 76 -319
<< viali >>
rect -17 307 17 341
rect -76 -319 -42 257
rect 42 -319 76 257
<< metal1 >>
rect -29 341 29 347
rect -29 307 -17 341
rect 17 307 29 341
rect -29 301 29 307
rect -82 257 -36 269
rect -82 -319 -76 257
rect -42 -319 -36 257
rect -82 -331 -36 -319
rect 36 257 82 269
rect 36 -319 42 257
rect 76 -319 82 257
rect 36 -331 82 -319
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
