magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< error_p >>
rect -594 18 594 236
<< nwell >>
rect -594 18 594 418
rect -594 -418 594 -18
<< pmos >>
rect -500 118 500 318
rect -500 -318 500 -118
<< pdiff >>
rect -558 306 -500 318
rect -558 130 -546 306
rect -512 130 -500 306
rect -558 118 -500 130
rect 500 306 558 318
rect 500 130 512 306
rect 546 130 558 306
rect 500 118 558 130
rect -558 -130 -500 -118
rect -558 -306 -546 -130
rect -512 -306 -500 -130
rect -558 -318 -500 -306
rect 500 -130 558 -118
rect 500 -306 512 -130
rect 546 -306 558 -130
rect 500 -318 558 -306
<< pdiffc >>
rect -546 130 -512 306
rect 512 130 546 306
rect -546 -306 -512 -130
rect 512 -306 546 -130
<< poly >>
rect -500 399 500 415
rect -500 365 -484 399
rect 484 365 500 399
rect -500 318 500 365
rect -500 71 500 118
rect -500 37 -484 71
rect 484 37 500 71
rect -500 21 500 37
rect -500 -37 500 -21
rect -500 -71 -484 -37
rect 484 -71 500 -37
rect -500 -118 500 -71
rect -500 -365 500 -318
rect -500 -399 -484 -365
rect 484 -399 500 -365
rect -500 -415 500 -399
<< polycont >>
rect -484 365 484 399
rect -484 37 484 71
rect -484 -71 484 -37
rect -484 -399 484 -365
<< locali >>
rect -500 365 -484 399
rect 484 365 500 399
rect -546 306 -512 322
rect -546 114 -512 130
rect 512 306 546 322
rect 512 114 546 130
rect -500 37 -484 71
rect 484 37 500 71
rect -500 -71 -484 -37
rect 484 -71 500 -37
rect -546 -130 -512 -114
rect -546 -322 -512 -306
rect 512 -130 546 -114
rect 512 -322 546 -306
rect -500 -399 -484 -365
rect 484 -399 500 -365
<< viali >>
rect -484 365 484 399
rect -546 130 -512 306
rect 512 130 546 306
rect -484 37 484 71
rect -484 -71 484 -37
rect -546 -306 -512 -130
rect 512 -306 546 -130
rect -484 -399 484 -365
<< metal1 >>
rect -496 399 496 405
rect -496 365 -484 399
rect 484 365 496 399
rect -496 359 496 365
rect -552 306 -506 318
rect -552 130 -546 306
rect -512 130 -506 306
rect -552 118 -506 130
rect 506 306 552 318
rect 506 130 512 306
rect 546 130 552 306
rect 506 118 552 130
rect -496 71 496 77
rect -496 37 -484 71
rect 484 37 496 71
rect -496 31 496 37
rect -496 -37 496 -31
rect -496 -71 -484 -37
rect 484 -71 496 -37
rect -496 -77 496 -71
rect -552 -130 -506 -118
rect -552 -306 -546 -130
rect -512 -306 -506 -130
rect -552 -318 -506 -306
rect 506 -130 552 -118
rect 506 -306 512 -130
rect 546 -306 552 -130
rect 506 -318 552 -306
rect -496 -365 496 -359
rect -496 -399 -484 -365
rect 484 -399 496 -365
rect -496 -405 496 -399
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 5.0 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
