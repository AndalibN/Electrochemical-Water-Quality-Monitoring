magic
tech sky130A
timestamp 1669661075
<< nwell >>
rect -160 330 1819 1085
rect -159 263 1819 330
<< psubdiff >>
rect -25 79 1726 93
rect -25 45 77 79
rect 1615 45 1726 79
rect -25 36 1726 45
rect -25 -592 -9 36
rect 57 30 1726 36
rect 57 20 1645 30
rect 57 -10 71 20
rect 57 -592 72 -10
rect 1631 -592 1645 20
rect -27 -596 1645 -592
rect 1699 20 1726 30
rect 1699 -596 1721 20
rect -27 -604 1721 -596
rect -27 -614 1719 -604
rect -27 -676 57 -614
rect 1649 -676 1719 -614
rect -27 -697 1719 -676
<< nsubdiff >>
rect -29 1027 1729 1046
rect -29 953 -18 1027
rect 1693 953 1729 1027
rect -29 932 1729 953
rect -29 931 65 932
rect -29 362 -22 931
rect 49 362 65 931
rect 1636 392 1654 932
rect 1707 392 1729 932
rect 1636 378 1729 392
rect -29 347 65 362
rect 1635 372 1729 378
rect 1635 347 1731 372
rect -31 334 1732 347
rect -31 299 62 334
rect 1649 299 1732 334
rect -31 285 1732 299
<< psubdiffcont >>
rect 77 45 1615 79
rect -9 -592 57 36
rect 1645 -596 1699 30
rect 57 -676 1649 -614
<< nsubdiffcont >>
rect -18 953 1693 1027
rect -22 362 49 931
rect 1654 392 1707 932
rect 62 299 1649 334
<< poly >>
rect 401 887 664 902
rect 221 843 343 870
rect 401 843 431 887
rect 634 868 664 887
rect 693 889 962 904
rect 693 843 723 889
rect 932 851 962 889
rect 221 833 251 843
rect 224 508 242 575
rect 190 494 242 508
rect 190 468 203 494
rect 230 468 242 494
rect 190 456 242 468
rect 135 -95 190 -83
rect 135 -124 148 -95
rect 180 -99 190 -95
rect 180 -123 253 -99
rect 180 -124 190 -123
rect 135 -137 190 -124
rect 230 -174 252 -123
rect 232 -519 247 -371
rect 408 -517 423 -484
rect 694 -517 713 -484
rect 408 -518 713 -517
rect 1001 -518 1018 -486
rect 408 -519 1018 -518
rect 232 -538 1018 -519
rect 419 -539 713 -538
<< polycont >>
rect 203 468 230 494
rect 148 -124 180 -95
<< locali >>
rect -25 1027 1718 1039
rect -25 953 -18 1027
rect 1693 953 1718 1027
rect -25 950 1718 953
rect -27 943 1718 950
rect -27 931 60 943
rect -27 362 -22 931
rect 49 362 60 931
rect 1644 932 1715 943
rect 194 496 236 502
rect 194 467 200 496
rect 232 467 236 496
rect 194 460 236 467
rect 1644 392 1654 932
rect 1707 392 1715 932
rect 1644 383 1715 392
rect -27 344 60 362
rect 1642 344 1715 383
rect -27 334 1715 344
rect -27 299 62 334
rect 1649 328 1715 334
rect 1649 299 1713 328
rect -27 292 1713 299
rect -16 86 1709 89
rect -19 79 1710 86
rect -19 45 77 79
rect 1615 45 1710 79
rect -19 36 1710 45
rect -19 -592 -9 36
rect 57 30 1710 36
rect 57 28 1645 30
rect 57 -592 64 28
rect 139 -92 188 -86
rect 139 -126 145 -92
rect 183 -126 188 -92
rect 139 -132 188 -126
rect -19 -606 64 -592
rect 1637 -596 1645 28
rect 1699 -596 1710 30
rect 1637 -606 1710 -596
rect -19 -612 1710 -606
rect -19 -614 1706 -612
rect -19 -676 57 -614
rect 1649 -676 1706 -614
rect -19 -686 1706 -676
rect -10 -689 1706 -686
<< viali >>
rect 194 974 218 996
rect 374 976 398 998
rect 666 977 690 999
rect 966 979 990 1001
rect 1262 975 1286 994
rect 1448 975 1468 992
rect 200 494 232 496
rect 200 468 203 494
rect 203 468 230 494
rect 230 468 232 494
rect 200 467 232 468
rect 145 -95 183 -92
rect 145 -124 148 -95
rect 148 -124 180 -95
rect 180 -124 183 -95
rect 145 -126 183 -124
rect 197 -647 216 -629
rect 374 -654 398 -635
rect 669 -647 690 -629
rect 966 -642 987 -622
<< metal1 >>
rect 187 996 225 1004
rect 187 974 194 996
rect 218 974 225 996
rect 187 965 225 974
rect 367 998 405 1006
rect 367 976 374 998
rect 398 976 405 998
rect 367 967 405 976
rect 659 999 697 1007
rect 659 977 666 999
rect 690 977 697 999
rect 659 968 697 977
rect 959 1001 997 1009
rect 959 979 966 1001
rect 990 979 997 1001
rect 959 970 997 979
rect 1256 994 1293 1000
rect 1256 975 1262 994
rect 1286 975 1293 994
rect 1256 970 1293 975
rect 1442 992 1474 996
rect 1442 975 1448 992
rect 1468 975 1474 992
rect 195 820 218 965
rect 375 829 398 967
rect 437 869 573 883
rect 437 827 454 869
rect 555 829 573 869
rect 667 830 690 968
rect 965 908 988 970
rect 729 871 865 885
rect 729 828 746 871
rect 847 828 865 871
rect 965 829 989 908
rect 1027 878 1165 893
rect 1027 827 1046 878
rect 1145 827 1165 878
rect 1267 843 1284 970
rect 1442 969 1474 975
rect 1450 848 1467 969
rect 268 582 277 584
rect 192 498 240 506
rect 192 496 243 498
rect 260 496 277 582
rect 192 467 200 496
rect 232 474 277 496
rect 318 490 335 530
rect 437 490 454 534
rect 318 475 454 490
rect 611 493 627 534
rect 729 493 747 532
rect 611 476 747 493
rect 909 491 926 532
rect 1027 491 1044 532
rect 909 475 1045 491
rect 1209 479 1225 498
rect 1391 483 1408 502
rect 1391 482 1477 483
rect 232 469 243 474
rect 232 467 240 469
rect 192 459 240 467
rect -140 -95 -57 -68
rect 136 -92 189 -84
rect 136 -94 145 -92
rect 51 -95 145 -94
rect -140 -124 145 -95
rect -140 -152 -57 -124
rect 136 -126 145 -124
rect 183 -126 189 -92
rect 136 -135 189 -126
rect 260 -184 277 474
rect 1209 465 1343 479
rect 1391 467 1527 482
rect 1391 466 1477 467
rect 376 223 441 240
rect 376 192 393 223
rect 426 216 441 223
rect 1176 226 1241 243
rect 1176 216 1193 226
rect 426 196 470 216
rect 513 196 762 216
rect 426 192 441 196
rect 807 194 1061 215
rect 1101 195 1193 216
rect 1226 216 1241 226
rect 1226 195 1305 216
rect 1628 215 1683 235
rect 1101 193 1196 195
rect 376 176 395 192
rect 420 176 441 192
rect 1176 179 1196 193
rect 1216 193 1305 195
rect 1338 193 1495 214
rect 1526 194 1683 215
rect 1216 179 1241 193
rect 1628 181 1683 194
rect 1468 -228 1469 -215
rect 395 -238 397 -229
rect 200 -623 216 -359
rect 189 -629 225 -623
rect 380 -626 397 -472
rect 672 -624 689 -474
rect 969 -615 985 -474
rect 960 -622 995 -615
rect 189 -647 197 -629
rect 216 -647 225 -629
rect 189 -655 225 -647
rect 367 -635 408 -626
rect 367 -654 374 -635
rect 398 -654 408 -635
rect 662 -629 699 -624
rect 662 -647 669 -629
rect 690 -647 699 -629
rect 960 -642 966 -622
rect 987 -642 995 -622
rect 960 -647 995 -642
rect 662 -653 699 -647
rect 367 -661 408 -654
<< via1 >>
rect 393 192 426 223
rect 1193 195 1226 226
<< metal2 >>
rect 1199 241 1221 243
rect 399 238 421 240
rect 378 223 439 238
rect 378 192 393 223
rect 426 192 439 223
rect 378 177 439 192
rect 1178 226 1239 241
rect 1178 195 1193 226
rect 1226 195 1239 226
rect 1178 180 1239 195
rect 394 155 419 177
rect 1195 155 1218 180
rect 393 134 1218 155
use inv  inv_0
timestamp 1669661075
transform 1 0 1184 0 1 460
box 0 -1128 183 415
use inv  inv_1
timestamp 1669661075
transform 1 0 1367 0 1 465
box 0 -1128 183 415
use sky130_fd_pr__nfet_01v8_7R257D  sky130_fd_pr__nfet_01v8_7R257D_0
timestamp 1669522153
transform 1 0 240 0 1 -273
box -57 -103 57 103
use sky130_fd_pr__pfet_01v8_GRHA7T  sky130_fd_pr__pfet_01v8_GRHA7T_0
timestamp 1669522153
transform 1 0 236 0 1 700
box -62 -151 62 151
use stage  stage_0
timestamp 1669661075
transform 1 0 295 0 1 499
box 0 -988 301 382
use stage  stage_1
timestamp 1669661075
transform 1 0 587 0 1 499
box 0 -988 301 382
use stage  stage_2
timestamp 1669661075
transform 1 0 885 0 1 498
box 0 -988 301 382
<< labels >>
rlabel nwell -10 960 1683 1018 7 VDD
port 1 w
rlabel metal1 1637 187 1673 226 7 Out
port 2 w
rlabel psubdiffcont 67 -670 1639 -617 7 gnd
port 3 w
rlabel metal1 -128 -142 -66 -79 7 In
port 4 w
<< end >>
