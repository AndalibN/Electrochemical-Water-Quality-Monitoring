magic
tech sky130A
magscale 1 2
timestamp 1666406900
<< error_p >>
rect -29 -788 29 -782
rect -29 -822 -17 -788
rect -29 -828 29 -822
<< nmos >>
rect -30 -750 30 750
<< ndiff >>
rect -88 738 -30 750
rect -88 -738 -76 738
rect -42 -738 -30 738
rect -88 -750 -30 -738
rect 30 738 88 750
rect 30 -738 42 738
rect 76 -738 88 738
rect 30 -750 88 -738
<< ndiffc >>
rect -76 -738 -42 738
rect 42 -738 76 738
<< poly >>
rect -30 750 30 838
rect -30 -772 30 -750
rect -33 -788 33 -772
rect -33 -822 -17 -788
rect 17 -822 33 -788
rect -33 -838 33 -822
<< polycont >>
rect -17 -822 17 -788
<< locali >>
rect -76 738 -42 754
rect -76 -754 -42 -738
rect 42 738 76 754
rect 42 -754 76 -738
rect -33 -822 -17 -788
rect 17 -822 33 -788
<< viali >>
rect -76 -738 -42 738
rect 42 -738 76 738
rect -17 -822 17 -788
<< metal1 >>
rect -82 738 -36 750
rect -82 -738 -76 738
rect -42 -738 -36 738
rect -82 -750 -36 -738
rect 36 738 82 750
rect 36 -738 42 738
rect 76 -738 82 738
rect 36 -750 82 -738
rect -29 -788 29 -782
rect -29 -822 -17 -788
rect 17 -822 29 -788
rect -29 -828 29 -822
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 7.5 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
