magic
tech sky130A
magscale 1 2
timestamp 1666815934
<< error_p >>
rect -29 739 29 745
rect -29 705 -17 739
rect -29 699 29 705
rect -29 -705 29 -699
rect -29 -739 -17 -705
rect -29 -745 29 -739
<< pwell >>
rect -226 -877 226 877
<< nmos >>
rect -30 -667 30 667
<< ndiff >>
rect -88 655 -30 667
rect -88 -655 -76 655
rect -42 -655 -30 655
rect -88 -667 -30 -655
rect 30 655 88 667
rect 30 -655 42 655
rect 76 -655 88 655
rect 30 -667 88 -655
<< ndiffc >>
rect -76 -655 -42 655
rect 42 -655 76 655
<< psubdiff >>
rect -190 807 -94 841
rect 94 807 190 841
rect -190 745 -156 807
rect 156 745 190 807
rect -190 -807 -156 -745
rect 156 -807 190 -745
rect -190 -841 -94 -807
rect 94 -841 190 -807
<< psubdiffcont >>
rect -94 807 94 841
rect -190 -745 -156 745
rect 156 -745 190 745
rect -94 -841 94 -807
<< poly >>
rect -33 739 33 755
rect -33 705 -17 739
rect 17 705 33 739
rect -33 689 33 705
rect -30 667 30 689
rect -30 -689 30 -667
rect -33 -705 33 -689
rect -33 -739 -17 -705
rect 17 -739 33 -705
rect -33 -755 33 -739
<< polycont >>
rect -17 705 17 739
rect -17 -739 17 -705
<< locali >>
rect -190 807 -94 841
rect 94 807 190 841
rect -190 745 -156 807
rect 156 745 190 807
rect -33 705 -17 739
rect 17 705 33 739
rect -76 655 -42 671
rect -76 -671 -42 -655
rect 42 655 76 671
rect 42 -671 76 -655
rect -33 -739 -17 -705
rect 17 -739 33 -705
rect -190 -807 -156 -745
rect 156 -807 190 -745
rect -190 -841 -94 -807
rect 94 -841 190 -807
<< viali >>
rect -17 705 17 739
rect -76 -655 -42 655
rect 42 -655 76 655
rect -17 -739 17 -705
<< metal1 >>
rect -29 739 29 745
rect -29 705 -17 739
rect 17 705 29 739
rect -29 699 29 705
rect -82 655 -36 667
rect -82 -655 -76 655
rect -42 -655 -36 655
rect -82 -667 -36 -655
rect 36 655 82 667
rect 36 -655 42 655
rect 76 -655 82 655
rect 36 -667 82 -655
rect -29 -705 29 -699
rect -29 -739 -17 -705
rect 17 -739 29 -705
rect -29 -745 29 -739
<< properties >>
string FIXED_BBOX -173 -824 173 824
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.67 l 0.3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
