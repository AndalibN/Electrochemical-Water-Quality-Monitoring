magic
tech sky130a
timestamp 1668788242
<< checkpaint >>
rect 0 0 2850 3000
use diffind_sam_bk diffind_sam_bk_1
timestamp 1668788242
transform 1 0 1750 0 1 700
box -1750 -700 1100 2300
<< end >>
