magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -294 -2064 294 2098
<< pmos >>
rect -200 -1964 200 2036
<< pdiff >>
rect -258 1991 -200 2036
rect -258 1957 -246 1991
rect -212 1957 -200 1991
rect -258 1923 -200 1957
rect -258 1889 -246 1923
rect -212 1889 -200 1923
rect -258 1855 -200 1889
rect -258 1821 -246 1855
rect -212 1821 -200 1855
rect -258 1787 -200 1821
rect -258 1753 -246 1787
rect -212 1753 -200 1787
rect -258 1719 -200 1753
rect -258 1685 -246 1719
rect -212 1685 -200 1719
rect -258 1651 -200 1685
rect -258 1617 -246 1651
rect -212 1617 -200 1651
rect -258 1583 -200 1617
rect -258 1549 -246 1583
rect -212 1549 -200 1583
rect -258 1515 -200 1549
rect -258 1481 -246 1515
rect -212 1481 -200 1515
rect -258 1447 -200 1481
rect -258 1413 -246 1447
rect -212 1413 -200 1447
rect -258 1379 -200 1413
rect -258 1345 -246 1379
rect -212 1345 -200 1379
rect -258 1311 -200 1345
rect -258 1277 -246 1311
rect -212 1277 -200 1311
rect -258 1243 -200 1277
rect -258 1209 -246 1243
rect -212 1209 -200 1243
rect -258 1175 -200 1209
rect -258 1141 -246 1175
rect -212 1141 -200 1175
rect -258 1107 -200 1141
rect -258 1073 -246 1107
rect -212 1073 -200 1107
rect -258 1039 -200 1073
rect -258 1005 -246 1039
rect -212 1005 -200 1039
rect -258 971 -200 1005
rect -258 937 -246 971
rect -212 937 -200 971
rect -258 903 -200 937
rect -258 869 -246 903
rect -212 869 -200 903
rect -258 835 -200 869
rect -258 801 -246 835
rect -212 801 -200 835
rect -258 767 -200 801
rect -258 733 -246 767
rect -212 733 -200 767
rect -258 699 -200 733
rect -258 665 -246 699
rect -212 665 -200 699
rect -258 631 -200 665
rect -258 597 -246 631
rect -212 597 -200 631
rect -258 563 -200 597
rect -258 529 -246 563
rect -212 529 -200 563
rect -258 495 -200 529
rect -258 461 -246 495
rect -212 461 -200 495
rect -258 427 -200 461
rect -258 393 -246 427
rect -212 393 -200 427
rect -258 359 -200 393
rect -258 325 -246 359
rect -212 325 -200 359
rect -258 291 -200 325
rect -258 257 -246 291
rect -212 257 -200 291
rect -258 223 -200 257
rect -258 189 -246 223
rect -212 189 -200 223
rect -258 155 -200 189
rect -258 121 -246 155
rect -212 121 -200 155
rect -258 87 -200 121
rect -258 53 -246 87
rect -212 53 -200 87
rect -258 19 -200 53
rect -258 -15 -246 19
rect -212 -15 -200 19
rect -258 -49 -200 -15
rect -258 -83 -246 -49
rect -212 -83 -200 -49
rect -258 -117 -200 -83
rect -258 -151 -246 -117
rect -212 -151 -200 -117
rect -258 -185 -200 -151
rect -258 -219 -246 -185
rect -212 -219 -200 -185
rect -258 -253 -200 -219
rect -258 -287 -246 -253
rect -212 -287 -200 -253
rect -258 -321 -200 -287
rect -258 -355 -246 -321
rect -212 -355 -200 -321
rect -258 -389 -200 -355
rect -258 -423 -246 -389
rect -212 -423 -200 -389
rect -258 -457 -200 -423
rect -258 -491 -246 -457
rect -212 -491 -200 -457
rect -258 -525 -200 -491
rect -258 -559 -246 -525
rect -212 -559 -200 -525
rect -258 -593 -200 -559
rect -258 -627 -246 -593
rect -212 -627 -200 -593
rect -258 -661 -200 -627
rect -258 -695 -246 -661
rect -212 -695 -200 -661
rect -258 -729 -200 -695
rect -258 -763 -246 -729
rect -212 -763 -200 -729
rect -258 -797 -200 -763
rect -258 -831 -246 -797
rect -212 -831 -200 -797
rect -258 -865 -200 -831
rect -258 -899 -246 -865
rect -212 -899 -200 -865
rect -258 -933 -200 -899
rect -258 -967 -246 -933
rect -212 -967 -200 -933
rect -258 -1001 -200 -967
rect -258 -1035 -246 -1001
rect -212 -1035 -200 -1001
rect -258 -1069 -200 -1035
rect -258 -1103 -246 -1069
rect -212 -1103 -200 -1069
rect -258 -1137 -200 -1103
rect -258 -1171 -246 -1137
rect -212 -1171 -200 -1137
rect -258 -1205 -200 -1171
rect -258 -1239 -246 -1205
rect -212 -1239 -200 -1205
rect -258 -1273 -200 -1239
rect -258 -1307 -246 -1273
rect -212 -1307 -200 -1273
rect -258 -1341 -200 -1307
rect -258 -1375 -246 -1341
rect -212 -1375 -200 -1341
rect -258 -1409 -200 -1375
rect -258 -1443 -246 -1409
rect -212 -1443 -200 -1409
rect -258 -1477 -200 -1443
rect -258 -1511 -246 -1477
rect -212 -1511 -200 -1477
rect -258 -1545 -200 -1511
rect -258 -1579 -246 -1545
rect -212 -1579 -200 -1545
rect -258 -1613 -200 -1579
rect -258 -1647 -246 -1613
rect -212 -1647 -200 -1613
rect -258 -1681 -200 -1647
rect -258 -1715 -246 -1681
rect -212 -1715 -200 -1681
rect -258 -1749 -200 -1715
rect -258 -1783 -246 -1749
rect -212 -1783 -200 -1749
rect -258 -1817 -200 -1783
rect -258 -1851 -246 -1817
rect -212 -1851 -200 -1817
rect -258 -1885 -200 -1851
rect -258 -1919 -246 -1885
rect -212 -1919 -200 -1885
rect -258 -1964 -200 -1919
rect 200 1991 258 2036
rect 200 1957 212 1991
rect 246 1957 258 1991
rect 200 1923 258 1957
rect 200 1889 212 1923
rect 246 1889 258 1923
rect 200 1855 258 1889
rect 200 1821 212 1855
rect 246 1821 258 1855
rect 200 1787 258 1821
rect 200 1753 212 1787
rect 246 1753 258 1787
rect 200 1719 258 1753
rect 200 1685 212 1719
rect 246 1685 258 1719
rect 200 1651 258 1685
rect 200 1617 212 1651
rect 246 1617 258 1651
rect 200 1583 258 1617
rect 200 1549 212 1583
rect 246 1549 258 1583
rect 200 1515 258 1549
rect 200 1481 212 1515
rect 246 1481 258 1515
rect 200 1447 258 1481
rect 200 1413 212 1447
rect 246 1413 258 1447
rect 200 1379 258 1413
rect 200 1345 212 1379
rect 246 1345 258 1379
rect 200 1311 258 1345
rect 200 1277 212 1311
rect 246 1277 258 1311
rect 200 1243 258 1277
rect 200 1209 212 1243
rect 246 1209 258 1243
rect 200 1175 258 1209
rect 200 1141 212 1175
rect 246 1141 258 1175
rect 200 1107 258 1141
rect 200 1073 212 1107
rect 246 1073 258 1107
rect 200 1039 258 1073
rect 200 1005 212 1039
rect 246 1005 258 1039
rect 200 971 258 1005
rect 200 937 212 971
rect 246 937 258 971
rect 200 903 258 937
rect 200 869 212 903
rect 246 869 258 903
rect 200 835 258 869
rect 200 801 212 835
rect 246 801 258 835
rect 200 767 258 801
rect 200 733 212 767
rect 246 733 258 767
rect 200 699 258 733
rect 200 665 212 699
rect 246 665 258 699
rect 200 631 258 665
rect 200 597 212 631
rect 246 597 258 631
rect 200 563 258 597
rect 200 529 212 563
rect 246 529 258 563
rect 200 495 258 529
rect 200 461 212 495
rect 246 461 258 495
rect 200 427 258 461
rect 200 393 212 427
rect 246 393 258 427
rect 200 359 258 393
rect 200 325 212 359
rect 246 325 258 359
rect 200 291 258 325
rect 200 257 212 291
rect 246 257 258 291
rect 200 223 258 257
rect 200 189 212 223
rect 246 189 258 223
rect 200 155 258 189
rect 200 121 212 155
rect 246 121 258 155
rect 200 87 258 121
rect 200 53 212 87
rect 246 53 258 87
rect 200 19 258 53
rect 200 -15 212 19
rect 246 -15 258 19
rect 200 -49 258 -15
rect 200 -83 212 -49
rect 246 -83 258 -49
rect 200 -117 258 -83
rect 200 -151 212 -117
rect 246 -151 258 -117
rect 200 -185 258 -151
rect 200 -219 212 -185
rect 246 -219 258 -185
rect 200 -253 258 -219
rect 200 -287 212 -253
rect 246 -287 258 -253
rect 200 -321 258 -287
rect 200 -355 212 -321
rect 246 -355 258 -321
rect 200 -389 258 -355
rect 200 -423 212 -389
rect 246 -423 258 -389
rect 200 -457 258 -423
rect 200 -491 212 -457
rect 246 -491 258 -457
rect 200 -525 258 -491
rect 200 -559 212 -525
rect 246 -559 258 -525
rect 200 -593 258 -559
rect 200 -627 212 -593
rect 246 -627 258 -593
rect 200 -661 258 -627
rect 200 -695 212 -661
rect 246 -695 258 -661
rect 200 -729 258 -695
rect 200 -763 212 -729
rect 246 -763 258 -729
rect 200 -797 258 -763
rect 200 -831 212 -797
rect 246 -831 258 -797
rect 200 -865 258 -831
rect 200 -899 212 -865
rect 246 -899 258 -865
rect 200 -933 258 -899
rect 200 -967 212 -933
rect 246 -967 258 -933
rect 200 -1001 258 -967
rect 200 -1035 212 -1001
rect 246 -1035 258 -1001
rect 200 -1069 258 -1035
rect 200 -1103 212 -1069
rect 246 -1103 258 -1069
rect 200 -1137 258 -1103
rect 200 -1171 212 -1137
rect 246 -1171 258 -1137
rect 200 -1205 258 -1171
rect 200 -1239 212 -1205
rect 246 -1239 258 -1205
rect 200 -1273 258 -1239
rect 200 -1307 212 -1273
rect 246 -1307 258 -1273
rect 200 -1341 258 -1307
rect 200 -1375 212 -1341
rect 246 -1375 258 -1341
rect 200 -1409 258 -1375
rect 200 -1443 212 -1409
rect 246 -1443 258 -1409
rect 200 -1477 258 -1443
rect 200 -1511 212 -1477
rect 246 -1511 258 -1477
rect 200 -1545 258 -1511
rect 200 -1579 212 -1545
rect 246 -1579 258 -1545
rect 200 -1613 258 -1579
rect 200 -1647 212 -1613
rect 246 -1647 258 -1613
rect 200 -1681 258 -1647
rect 200 -1715 212 -1681
rect 246 -1715 258 -1681
rect 200 -1749 258 -1715
rect 200 -1783 212 -1749
rect 246 -1783 258 -1749
rect 200 -1817 258 -1783
rect 200 -1851 212 -1817
rect 246 -1851 258 -1817
rect 200 -1885 258 -1851
rect 200 -1919 212 -1885
rect 246 -1919 258 -1885
rect 200 -1964 258 -1919
<< pdiffc >>
rect -246 1957 -212 1991
rect -246 1889 -212 1923
rect -246 1821 -212 1855
rect -246 1753 -212 1787
rect -246 1685 -212 1719
rect -246 1617 -212 1651
rect -246 1549 -212 1583
rect -246 1481 -212 1515
rect -246 1413 -212 1447
rect -246 1345 -212 1379
rect -246 1277 -212 1311
rect -246 1209 -212 1243
rect -246 1141 -212 1175
rect -246 1073 -212 1107
rect -246 1005 -212 1039
rect -246 937 -212 971
rect -246 869 -212 903
rect -246 801 -212 835
rect -246 733 -212 767
rect -246 665 -212 699
rect -246 597 -212 631
rect -246 529 -212 563
rect -246 461 -212 495
rect -246 393 -212 427
rect -246 325 -212 359
rect -246 257 -212 291
rect -246 189 -212 223
rect -246 121 -212 155
rect -246 53 -212 87
rect -246 -15 -212 19
rect -246 -83 -212 -49
rect -246 -151 -212 -117
rect -246 -219 -212 -185
rect -246 -287 -212 -253
rect -246 -355 -212 -321
rect -246 -423 -212 -389
rect -246 -491 -212 -457
rect -246 -559 -212 -525
rect -246 -627 -212 -593
rect -246 -695 -212 -661
rect -246 -763 -212 -729
rect -246 -831 -212 -797
rect -246 -899 -212 -865
rect -246 -967 -212 -933
rect -246 -1035 -212 -1001
rect -246 -1103 -212 -1069
rect -246 -1171 -212 -1137
rect -246 -1239 -212 -1205
rect -246 -1307 -212 -1273
rect -246 -1375 -212 -1341
rect -246 -1443 -212 -1409
rect -246 -1511 -212 -1477
rect -246 -1579 -212 -1545
rect -246 -1647 -212 -1613
rect -246 -1715 -212 -1681
rect -246 -1783 -212 -1749
rect -246 -1851 -212 -1817
rect -246 -1919 -212 -1885
rect 212 1957 246 1991
rect 212 1889 246 1923
rect 212 1821 246 1855
rect 212 1753 246 1787
rect 212 1685 246 1719
rect 212 1617 246 1651
rect 212 1549 246 1583
rect 212 1481 246 1515
rect 212 1413 246 1447
rect 212 1345 246 1379
rect 212 1277 246 1311
rect 212 1209 246 1243
rect 212 1141 246 1175
rect 212 1073 246 1107
rect 212 1005 246 1039
rect 212 937 246 971
rect 212 869 246 903
rect 212 801 246 835
rect 212 733 246 767
rect 212 665 246 699
rect 212 597 246 631
rect 212 529 246 563
rect 212 461 246 495
rect 212 393 246 427
rect 212 325 246 359
rect 212 257 246 291
rect 212 189 246 223
rect 212 121 246 155
rect 212 53 246 87
rect 212 -15 246 19
rect 212 -83 246 -49
rect 212 -151 246 -117
rect 212 -219 246 -185
rect 212 -287 246 -253
rect 212 -355 246 -321
rect 212 -423 246 -389
rect 212 -491 246 -457
rect 212 -559 246 -525
rect 212 -627 246 -593
rect 212 -695 246 -661
rect 212 -763 246 -729
rect 212 -831 246 -797
rect 212 -899 246 -865
rect 212 -967 246 -933
rect 212 -1035 246 -1001
rect 212 -1103 246 -1069
rect 212 -1171 246 -1137
rect 212 -1239 246 -1205
rect 212 -1307 246 -1273
rect 212 -1375 246 -1341
rect 212 -1443 246 -1409
rect 212 -1511 246 -1477
rect 212 -1579 246 -1545
rect 212 -1647 246 -1613
rect 212 -1715 246 -1681
rect 212 -1783 246 -1749
rect 212 -1851 246 -1817
rect 212 -1919 246 -1885
<< poly >>
rect -200 2036 200 2062
rect -200 -2011 200 -1964
rect -200 -2045 -153 -2011
rect -119 -2045 -85 -2011
rect -51 -2045 -17 -2011
rect 17 -2045 51 -2011
rect 85 -2045 119 -2011
rect 153 -2045 200 -2011
rect -200 -2061 200 -2045
<< polycont >>
rect -153 -2045 -119 -2011
rect -85 -2045 -51 -2011
rect -17 -2045 17 -2011
rect 51 -2045 85 -2011
rect 119 -2045 153 -2011
<< locali >>
rect -246 1997 -212 2040
rect -246 1925 -212 1957
rect -246 1855 -212 1889
rect -246 1787 -212 1819
rect -246 1719 -212 1747
rect -246 1651 -212 1675
rect -246 1583 -212 1603
rect -246 1515 -212 1531
rect -246 1447 -212 1459
rect -246 1379 -212 1387
rect -246 1311 -212 1315
rect -246 1205 -212 1209
rect -246 1133 -212 1141
rect -246 1061 -212 1073
rect -246 989 -212 1005
rect -246 917 -212 937
rect -246 845 -212 869
rect -246 773 -212 801
rect -246 701 -212 733
rect -246 631 -212 665
rect -246 563 -212 595
rect -246 495 -212 523
rect -246 427 -212 451
rect -246 359 -212 379
rect -246 291 -212 307
rect -246 223 -212 235
rect -246 155 -212 163
rect -246 87 -212 91
rect -246 -19 -212 -15
rect -246 -91 -212 -83
rect -246 -163 -212 -151
rect -246 -235 -212 -219
rect -246 -307 -212 -287
rect -246 -379 -212 -355
rect -246 -451 -212 -423
rect -246 -523 -212 -491
rect -246 -593 -212 -559
rect -246 -661 -212 -629
rect -246 -729 -212 -701
rect -246 -797 -212 -773
rect -246 -865 -212 -845
rect -246 -933 -212 -917
rect -246 -1001 -212 -989
rect -246 -1069 -212 -1061
rect -246 -1137 -212 -1133
rect -246 -1243 -212 -1239
rect -246 -1315 -212 -1307
rect -246 -1387 -212 -1375
rect -246 -1459 -212 -1443
rect -246 -1531 -212 -1511
rect -246 -1603 -212 -1579
rect -246 -1675 -212 -1647
rect -246 -1747 -212 -1715
rect -246 -1817 -212 -1783
rect -246 -1885 -212 -1853
rect -246 -1968 -212 -1925
rect 212 1997 246 2040
rect 212 1925 246 1957
rect 212 1855 246 1889
rect 212 1787 246 1819
rect 212 1719 246 1747
rect 212 1651 246 1675
rect 212 1583 246 1603
rect 212 1515 246 1531
rect 212 1447 246 1459
rect 212 1379 246 1387
rect 212 1311 246 1315
rect 212 1205 246 1209
rect 212 1133 246 1141
rect 212 1061 246 1073
rect 212 989 246 1005
rect 212 917 246 937
rect 212 845 246 869
rect 212 773 246 801
rect 212 701 246 733
rect 212 631 246 665
rect 212 563 246 595
rect 212 495 246 523
rect 212 427 246 451
rect 212 359 246 379
rect 212 291 246 307
rect 212 223 246 235
rect 212 155 246 163
rect 212 87 246 91
rect 212 -19 246 -15
rect 212 -91 246 -83
rect 212 -163 246 -151
rect 212 -235 246 -219
rect 212 -307 246 -287
rect 212 -379 246 -355
rect 212 -451 246 -423
rect 212 -523 246 -491
rect 212 -593 246 -559
rect 212 -661 246 -629
rect 212 -729 246 -701
rect 212 -797 246 -773
rect 212 -865 246 -845
rect 212 -933 246 -917
rect 212 -1001 246 -989
rect 212 -1069 246 -1061
rect 212 -1137 246 -1133
rect 212 -1243 246 -1239
rect 212 -1315 246 -1307
rect 212 -1387 246 -1375
rect 212 -1459 246 -1443
rect 212 -1531 246 -1511
rect 212 -1603 246 -1579
rect 212 -1675 246 -1647
rect 212 -1747 246 -1715
rect 212 -1817 246 -1783
rect 212 -1885 246 -1853
rect 212 -1968 246 -1925
rect -200 -2045 -161 -2011
rect -119 -2045 -89 -2011
rect -51 -2045 -17 -2011
rect 17 -2045 51 -2011
rect 89 -2045 119 -2011
rect 161 -2045 200 -2011
<< viali >>
rect -246 1991 -212 1997
rect -246 1963 -212 1991
rect -246 1923 -212 1925
rect -246 1891 -212 1923
rect -246 1821 -212 1853
rect -246 1819 -212 1821
rect -246 1753 -212 1781
rect -246 1747 -212 1753
rect -246 1685 -212 1709
rect -246 1675 -212 1685
rect -246 1617 -212 1637
rect -246 1603 -212 1617
rect -246 1549 -212 1565
rect -246 1531 -212 1549
rect -246 1481 -212 1493
rect -246 1459 -212 1481
rect -246 1413 -212 1421
rect -246 1387 -212 1413
rect -246 1345 -212 1349
rect -246 1315 -212 1345
rect -246 1243 -212 1277
rect -246 1175 -212 1205
rect -246 1171 -212 1175
rect -246 1107 -212 1133
rect -246 1099 -212 1107
rect -246 1039 -212 1061
rect -246 1027 -212 1039
rect -246 971 -212 989
rect -246 955 -212 971
rect -246 903 -212 917
rect -246 883 -212 903
rect -246 835 -212 845
rect -246 811 -212 835
rect -246 767 -212 773
rect -246 739 -212 767
rect -246 699 -212 701
rect -246 667 -212 699
rect -246 597 -212 629
rect -246 595 -212 597
rect -246 529 -212 557
rect -246 523 -212 529
rect -246 461 -212 485
rect -246 451 -212 461
rect -246 393 -212 413
rect -246 379 -212 393
rect -246 325 -212 341
rect -246 307 -212 325
rect -246 257 -212 269
rect -246 235 -212 257
rect -246 189 -212 197
rect -246 163 -212 189
rect -246 121 -212 125
rect -246 91 -212 121
rect -246 19 -212 53
rect -246 -49 -212 -19
rect -246 -53 -212 -49
rect -246 -117 -212 -91
rect -246 -125 -212 -117
rect -246 -185 -212 -163
rect -246 -197 -212 -185
rect -246 -253 -212 -235
rect -246 -269 -212 -253
rect -246 -321 -212 -307
rect -246 -341 -212 -321
rect -246 -389 -212 -379
rect -246 -413 -212 -389
rect -246 -457 -212 -451
rect -246 -485 -212 -457
rect -246 -525 -212 -523
rect -246 -557 -212 -525
rect -246 -627 -212 -595
rect -246 -629 -212 -627
rect -246 -695 -212 -667
rect -246 -701 -212 -695
rect -246 -763 -212 -739
rect -246 -773 -212 -763
rect -246 -831 -212 -811
rect -246 -845 -212 -831
rect -246 -899 -212 -883
rect -246 -917 -212 -899
rect -246 -967 -212 -955
rect -246 -989 -212 -967
rect -246 -1035 -212 -1027
rect -246 -1061 -212 -1035
rect -246 -1103 -212 -1099
rect -246 -1133 -212 -1103
rect -246 -1205 -212 -1171
rect -246 -1273 -212 -1243
rect -246 -1277 -212 -1273
rect -246 -1341 -212 -1315
rect -246 -1349 -212 -1341
rect -246 -1409 -212 -1387
rect -246 -1421 -212 -1409
rect -246 -1477 -212 -1459
rect -246 -1493 -212 -1477
rect -246 -1545 -212 -1531
rect -246 -1565 -212 -1545
rect -246 -1613 -212 -1603
rect -246 -1637 -212 -1613
rect -246 -1681 -212 -1675
rect -246 -1709 -212 -1681
rect -246 -1749 -212 -1747
rect -246 -1781 -212 -1749
rect -246 -1851 -212 -1819
rect -246 -1853 -212 -1851
rect -246 -1919 -212 -1891
rect -246 -1925 -212 -1919
rect 212 1991 246 1997
rect 212 1963 246 1991
rect 212 1923 246 1925
rect 212 1891 246 1923
rect 212 1821 246 1853
rect 212 1819 246 1821
rect 212 1753 246 1781
rect 212 1747 246 1753
rect 212 1685 246 1709
rect 212 1675 246 1685
rect 212 1617 246 1637
rect 212 1603 246 1617
rect 212 1549 246 1565
rect 212 1531 246 1549
rect 212 1481 246 1493
rect 212 1459 246 1481
rect 212 1413 246 1421
rect 212 1387 246 1413
rect 212 1345 246 1349
rect 212 1315 246 1345
rect 212 1243 246 1277
rect 212 1175 246 1205
rect 212 1171 246 1175
rect 212 1107 246 1133
rect 212 1099 246 1107
rect 212 1039 246 1061
rect 212 1027 246 1039
rect 212 971 246 989
rect 212 955 246 971
rect 212 903 246 917
rect 212 883 246 903
rect 212 835 246 845
rect 212 811 246 835
rect 212 767 246 773
rect 212 739 246 767
rect 212 699 246 701
rect 212 667 246 699
rect 212 597 246 629
rect 212 595 246 597
rect 212 529 246 557
rect 212 523 246 529
rect 212 461 246 485
rect 212 451 246 461
rect 212 393 246 413
rect 212 379 246 393
rect 212 325 246 341
rect 212 307 246 325
rect 212 257 246 269
rect 212 235 246 257
rect 212 189 246 197
rect 212 163 246 189
rect 212 121 246 125
rect 212 91 246 121
rect 212 19 246 53
rect 212 -49 246 -19
rect 212 -53 246 -49
rect 212 -117 246 -91
rect 212 -125 246 -117
rect 212 -185 246 -163
rect 212 -197 246 -185
rect 212 -253 246 -235
rect 212 -269 246 -253
rect 212 -321 246 -307
rect 212 -341 246 -321
rect 212 -389 246 -379
rect 212 -413 246 -389
rect 212 -457 246 -451
rect 212 -485 246 -457
rect 212 -525 246 -523
rect 212 -557 246 -525
rect 212 -627 246 -595
rect 212 -629 246 -627
rect 212 -695 246 -667
rect 212 -701 246 -695
rect 212 -763 246 -739
rect 212 -773 246 -763
rect 212 -831 246 -811
rect 212 -845 246 -831
rect 212 -899 246 -883
rect 212 -917 246 -899
rect 212 -967 246 -955
rect 212 -989 246 -967
rect 212 -1035 246 -1027
rect 212 -1061 246 -1035
rect 212 -1103 246 -1099
rect 212 -1133 246 -1103
rect 212 -1205 246 -1171
rect 212 -1273 246 -1243
rect 212 -1277 246 -1273
rect 212 -1341 246 -1315
rect 212 -1349 246 -1341
rect 212 -1409 246 -1387
rect 212 -1421 246 -1409
rect 212 -1477 246 -1459
rect 212 -1493 246 -1477
rect 212 -1545 246 -1531
rect 212 -1565 246 -1545
rect 212 -1613 246 -1603
rect 212 -1637 246 -1613
rect 212 -1681 246 -1675
rect 212 -1709 246 -1681
rect 212 -1749 246 -1747
rect 212 -1781 246 -1749
rect 212 -1851 246 -1819
rect 212 -1853 246 -1851
rect 212 -1919 246 -1891
rect 212 -1925 246 -1919
rect -161 -2045 -153 -2011
rect -153 -2045 -127 -2011
rect -89 -2045 -85 -2011
rect -85 -2045 -55 -2011
rect -17 -2045 17 -2011
rect 55 -2045 85 -2011
rect 85 -2045 89 -2011
rect 127 -2045 153 -2011
rect 153 -2045 161 -2011
<< metal1 >>
rect -252 1997 -206 2036
rect -252 1963 -246 1997
rect -212 1963 -206 1997
rect -252 1925 -206 1963
rect -252 1891 -246 1925
rect -212 1891 -206 1925
rect -252 1853 -206 1891
rect -252 1819 -246 1853
rect -212 1819 -206 1853
rect -252 1781 -206 1819
rect -252 1747 -246 1781
rect -212 1747 -206 1781
rect -252 1709 -206 1747
rect -252 1675 -246 1709
rect -212 1675 -206 1709
rect -252 1637 -206 1675
rect -252 1603 -246 1637
rect -212 1603 -206 1637
rect -252 1565 -206 1603
rect -252 1531 -246 1565
rect -212 1531 -206 1565
rect -252 1493 -206 1531
rect -252 1459 -246 1493
rect -212 1459 -206 1493
rect -252 1421 -206 1459
rect -252 1387 -246 1421
rect -212 1387 -206 1421
rect -252 1349 -206 1387
rect -252 1315 -246 1349
rect -212 1315 -206 1349
rect -252 1277 -206 1315
rect -252 1243 -246 1277
rect -212 1243 -206 1277
rect -252 1205 -206 1243
rect -252 1171 -246 1205
rect -212 1171 -206 1205
rect -252 1133 -206 1171
rect -252 1099 -246 1133
rect -212 1099 -206 1133
rect -252 1061 -206 1099
rect -252 1027 -246 1061
rect -212 1027 -206 1061
rect -252 989 -206 1027
rect -252 955 -246 989
rect -212 955 -206 989
rect -252 917 -206 955
rect -252 883 -246 917
rect -212 883 -206 917
rect -252 845 -206 883
rect -252 811 -246 845
rect -212 811 -206 845
rect -252 773 -206 811
rect -252 739 -246 773
rect -212 739 -206 773
rect -252 701 -206 739
rect -252 667 -246 701
rect -212 667 -206 701
rect -252 629 -206 667
rect -252 595 -246 629
rect -212 595 -206 629
rect -252 557 -206 595
rect -252 523 -246 557
rect -212 523 -206 557
rect -252 485 -206 523
rect -252 451 -246 485
rect -212 451 -206 485
rect -252 413 -206 451
rect -252 379 -246 413
rect -212 379 -206 413
rect -252 341 -206 379
rect -252 307 -246 341
rect -212 307 -206 341
rect -252 269 -206 307
rect -252 235 -246 269
rect -212 235 -206 269
rect -252 197 -206 235
rect -252 163 -246 197
rect -212 163 -206 197
rect -252 125 -206 163
rect -252 91 -246 125
rect -212 91 -206 125
rect -252 53 -206 91
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -91 -206 -53
rect -252 -125 -246 -91
rect -212 -125 -206 -91
rect -252 -163 -206 -125
rect -252 -197 -246 -163
rect -212 -197 -206 -163
rect -252 -235 -206 -197
rect -252 -269 -246 -235
rect -212 -269 -206 -235
rect -252 -307 -206 -269
rect -252 -341 -246 -307
rect -212 -341 -206 -307
rect -252 -379 -206 -341
rect -252 -413 -246 -379
rect -212 -413 -206 -379
rect -252 -451 -206 -413
rect -252 -485 -246 -451
rect -212 -485 -206 -451
rect -252 -523 -206 -485
rect -252 -557 -246 -523
rect -212 -557 -206 -523
rect -252 -595 -206 -557
rect -252 -629 -246 -595
rect -212 -629 -206 -595
rect -252 -667 -206 -629
rect -252 -701 -246 -667
rect -212 -701 -206 -667
rect -252 -739 -206 -701
rect -252 -773 -246 -739
rect -212 -773 -206 -739
rect -252 -811 -206 -773
rect -252 -845 -246 -811
rect -212 -845 -206 -811
rect -252 -883 -206 -845
rect -252 -917 -246 -883
rect -212 -917 -206 -883
rect -252 -955 -206 -917
rect -252 -989 -246 -955
rect -212 -989 -206 -955
rect -252 -1027 -206 -989
rect -252 -1061 -246 -1027
rect -212 -1061 -206 -1027
rect -252 -1099 -206 -1061
rect -252 -1133 -246 -1099
rect -212 -1133 -206 -1099
rect -252 -1171 -206 -1133
rect -252 -1205 -246 -1171
rect -212 -1205 -206 -1171
rect -252 -1243 -206 -1205
rect -252 -1277 -246 -1243
rect -212 -1277 -206 -1243
rect -252 -1315 -206 -1277
rect -252 -1349 -246 -1315
rect -212 -1349 -206 -1315
rect -252 -1387 -206 -1349
rect -252 -1421 -246 -1387
rect -212 -1421 -206 -1387
rect -252 -1459 -206 -1421
rect -252 -1493 -246 -1459
rect -212 -1493 -206 -1459
rect -252 -1531 -206 -1493
rect -252 -1565 -246 -1531
rect -212 -1565 -206 -1531
rect -252 -1603 -206 -1565
rect -252 -1637 -246 -1603
rect -212 -1637 -206 -1603
rect -252 -1675 -206 -1637
rect -252 -1709 -246 -1675
rect -212 -1709 -206 -1675
rect -252 -1747 -206 -1709
rect -252 -1781 -246 -1747
rect -212 -1781 -206 -1747
rect -252 -1819 -206 -1781
rect -252 -1853 -246 -1819
rect -212 -1853 -206 -1819
rect -252 -1891 -206 -1853
rect -252 -1925 -246 -1891
rect -212 -1925 -206 -1891
rect -252 -1964 -206 -1925
rect 206 1997 252 2036
rect 206 1963 212 1997
rect 246 1963 252 1997
rect 206 1925 252 1963
rect 206 1891 212 1925
rect 246 1891 252 1925
rect 206 1853 252 1891
rect 206 1819 212 1853
rect 246 1819 252 1853
rect 206 1781 252 1819
rect 206 1747 212 1781
rect 246 1747 252 1781
rect 206 1709 252 1747
rect 206 1675 212 1709
rect 246 1675 252 1709
rect 206 1637 252 1675
rect 206 1603 212 1637
rect 246 1603 252 1637
rect 206 1565 252 1603
rect 206 1531 212 1565
rect 246 1531 252 1565
rect 206 1493 252 1531
rect 206 1459 212 1493
rect 246 1459 252 1493
rect 206 1421 252 1459
rect 206 1387 212 1421
rect 246 1387 252 1421
rect 206 1349 252 1387
rect 206 1315 212 1349
rect 246 1315 252 1349
rect 206 1277 252 1315
rect 206 1243 212 1277
rect 246 1243 252 1277
rect 206 1205 252 1243
rect 206 1171 212 1205
rect 246 1171 252 1205
rect 206 1133 252 1171
rect 206 1099 212 1133
rect 246 1099 252 1133
rect 206 1061 252 1099
rect 206 1027 212 1061
rect 246 1027 252 1061
rect 206 989 252 1027
rect 206 955 212 989
rect 246 955 252 989
rect 206 917 252 955
rect 206 883 212 917
rect 246 883 252 917
rect 206 845 252 883
rect 206 811 212 845
rect 246 811 252 845
rect 206 773 252 811
rect 206 739 212 773
rect 246 739 252 773
rect 206 701 252 739
rect 206 667 212 701
rect 246 667 252 701
rect 206 629 252 667
rect 206 595 212 629
rect 246 595 252 629
rect 206 557 252 595
rect 206 523 212 557
rect 246 523 252 557
rect 206 485 252 523
rect 206 451 212 485
rect 246 451 252 485
rect 206 413 252 451
rect 206 379 212 413
rect 246 379 252 413
rect 206 341 252 379
rect 206 307 212 341
rect 246 307 252 341
rect 206 269 252 307
rect 206 235 212 269
rect 246 235 252 269
rect 206 197 252 235
rect 206 163 212 197
rect 246 163 252 197
rect 206 125 252 163
rect 206 91 212 125
rect 246 91 252 125
rect 206 53 252 91
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -91 252 -53
rect 206 -125 212 -91
rect 246 -125 252 -91
rect 206 -163 252 -125
rect 206 -197 212 -163
rect 246 -197 252 -163
rect 206 -235 252 -197
rect 206 -269 212 -235
rect 246 -269 252 -235
rect 206 -307 252 -269
rect 206 -341 212 -307
rect 246 -341 252 -307
rect 206 -379 252 -341
rect 206 -413 212 -379
rect 246 -413 252 -379
rect 206 -451 252 -413
rect 206 -485 212 -451
rect 246 -485 252 -451
rect 206 -523 252 -485
rect 206 -557 212 -523
rect 246 -557 252 -523
rect 206 -595 252 -557
rect 206 -629 212 -595
rect 246 -629 252 -595
rect 206 -667 252 -629
rect 206 -701 212 -667
rect 246 -701 252 -667
rect 206 -739 252 -701
rect 206 -773 212 -739
rect 246 -773 252 -739
rect 206 -811 252 -773
rect 206 -845 212 -811
rect 246 -845 252 -811
rect 206 -883 252 -845
rect 206 -917 212 -883
rect 246 -917 252 -883
rect 206 -955 252 -917
rect 206 -989 212 -955
rect 246 -989 252 -955
rect 206 -1027 252 -989
rect 206 -1061 212 -1027
rect 246 -1061 252 -1027
rect 206 -1099 252 -1061
rect 206 -1133 212 -1099
rect 246 -1133 252 -1099
rect 206 -1171 252 -1133
rect 206 -1205 212 -1171
rect 246 -1205 252 -1171
rect 206 -1243 252 -1205
rect 206 -1277 212 -1243
rect 246 -1277 252 -1243
rect 206 -1315 252 -1277
rect 206 -1349 212 -1315
rect 246 -1349 252 -1315
rect 206 -1387 252 -1349
rect 206 -1421 212 -1387
rect 246 -1421 252 -1387
rect 206 -1459 252 -1421
rect 206 -1493 212 -1459
rect 246 -1493 252 -1459
rect 206 -1531 252 -1493
rect 206 -1565 212 -1531
rect 246 -1565 252 -1531
rect 206 -1603 252 -1565
rect 206 -1637 212 -1603
rect 246 -1637 252 -1603
rect 206 -1675 252 -1637
rect 206 -1709 212 -1675
rect 246 -1709 252 -1675
rect 206 -1747 252 -1709
rect 206 -1781 212 -1747
rect 246 -1781 252 -1747
rect 206 -1819 252 -1781
rect 206 -1853 212 -1819
rect 246 -1853 252 -1819
rect 206 -1891 252 -1853
rect 206 -1925 212 -1891
rect 246 -1925 252 -1891
rect 206 -1964 252 -1925
rect -196 -2011 196 -2005
rect -196 -2045 -161 -2011
rect -127 -2045 -89 -2011
rect -55 -2045 -17 -2011
rect 17 -2045 55 -2011
rect 89 -2045 127 -2011
rect 161 -2045 196 -2011
rect -196 -2051 196 -2045
<< end >>
