magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< nwell >>
rect -109 -290 109 276
<< pmos >>
rect -15 -228 15 156
<< pdiff >>
rect -73 117 -15 156
rect -73 83 -61 117
rect -27 83 -15 117
rect -73 49 -15 83
rect -73 15 -61 49
rect -27 15 -15 49
rect -73 -19 -15 15
rect -73 -53 -61 -19
rect -27 -53 -15 -19
rect -73 -87 -15 -53
rect -73 -121 -61 -87
rect -27 -121 -15 -87
rect -73 -155 -15 -121
rect -73 -189 -61 -155
rect -27 -189 -15 -155
rect -73 -228 -15 -189
rect 15 117 73 156
rect 15 83 27 117
rect 61 83 73 117
rect 15 49 73 83
rect 15 15 27 49
rect 61 15 73 49
rect 15 -19 73 15
rect 15 -53 27 -19
rect 61 -53 73 -19
rect 15 -87 73 -53
rect 15 -121 27 -87
rect 61 -121 73 -87
rect 15 -155 73 -121
rect 15 -189 27 -155
rect 61 -189 73 -155
rect 15 -228 73 -189
<< pdiffc >>
rect -61 83 -27 117
rect -61 15 -27 49
rect -61 -53 -27 -19
rect -61 -121 -27 -87
rect -61 -189 -27 -155
rect 27 83 61 117
rect 27 15 61 49
rect 27 -53 61 -19
rect 27 -121 61 -87
rect 27 -189 61 -155
<< poly >>
rect -66 257 0 273
rect -66 223 -50 257
rect -16 223 0 257
rect -66 220 0 223
rect -66 207 15 220
rect -37 190 15 207
rect -15 156 15 190
rect -15 -254 15 -228
<< polycont >>
rect -50 223 -16 257
<< locali >>
rect -66 223 -50 257
rect -16 223 0 257
rect -61 125 -27 160
rect -61 53 -27 83
rect -61 -19 -27 15
rect -61 -87 -27 -53
rect -61 -155 -27 -125
rect -61 -232 -27 -197
rect 27 125 61 160
rect 27 53 61 83
rect 27 -19 61 15
rect 27 -87 61 -53
rect 27 -155 61 -125
rect 27 -232 61 -197
<< viali >>
rect -50 223 -16 257
rect -61 117 -27 125
rect -61 91 -27 117
rect -61 49 -27 53
rect -61 19 -27 49
rect -61 -53 -27 -19
rect -61 -121 -27 -91
rect -61 -125 -27 -121
rect -61 -189 -27 -163
rect -61 -197 -27 -189
rect 27 117 61 125
rect 27 91 61 117
rect 27 49 61 53
rect 27 19 61 49
rect 27 -53 61 -19
rect 27 -121 61 -91
rect 27 -125 61 -121
rect 27 -189 61 -163
rect 27 -197 61 -189
<< metal1 >>
rect -64 257 -2 268
rect -64 223 -50 257
rect -16 223 -2 257
rect -64 214 -2 223
rect -67 125 -21 156
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -163 -21 -125
rect -67 -197 -61 -163
rect -27 -197 -21 -163
rect -67 -228 -21 -197
rect 21 125 67 156
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -163 67 -125
rect 21 -197 27 -163
rect 61 -197 67 -163
rect 21 -228 67 -197
<< end >>
