magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< error_p >>
rect -88 -971 -30 -965
rect 30 -971 88 -965
rect -88 -1005 -76 -971
rect 30 -1005 42 -971
rect -88 -1011 -30 -1005
rect 30 -1011 88 -1005
<< nwell >>
rect -183 -1024 183 1058
<< pmos >>
rect -89 -924 -29 996
rect 29 -924 89 996
<< pdiff >>
rect -147 971 -89 996
rect -147 937 -135 971
rect -101 937 -89 971
rect -147 903 -89 937
rect -147 869 -135 903
rect -101 869 -89 903
rect -147 835 -89 869
rect -147 801 -135 835
rect -101 801 -89 835
rect -147 767 -89 801
rect -147 733 -135 767
rect -101 733 -89 767
rect -147 699 -89 733
rect -147 665 -135 699
rect -101 665 -89 699
rect -147 631 -89 665
rect -147 597 -135 631
rect -101 597 -89 631
rect -147 563 -89 597
rect -147 529 -135 563
rect -101 529 -89 563
rect -147 495 -89 529
rect -147 461 -135 495
rect -101 461 -89 495
rect -147 427 -89 461
rect -147 393 -135 427
rect -101 393 -89 427
rect -147 359 -89 393
rect -147 325 -135 359
rect -101 325 -89 359
rect -147 291 -89 325
rect -147 257 -135 291
rect -101 257 -89 291
rect -147 223 -89 257
rect -147 189 -135 223
rect -101 189 -89 223
rect -147 155 -89 189
rect -147 121 -135 155
rect -101 121 -89 155
rect -147 87 -89 121
rect -147 53 -135 87
rect -101 53 -89 87
rect -147 19 -89 53
rect -147 -15 -135 19
rect -101 -15 -89 19
rect -147 -49 -89 -15
rect -147 -83 -135 -49
rect -101 -83 -89 -49
rect -147 -117 -89 -83
rect -147 -151 -135 -117
rect -101 -151 -89 -117
rect -147 -185 -89 -151
rect -147 -219 -135 -185
rect -101 -219 -89 -185
rect -147 -253 -89 -219
rect -147 -287 -135 -253
rect -101 -287 -89 -253
rect -147 -321 -89 -287
rect -147 -355 -135 -321
rect -101 -355 -89 -321
rect -147 -389 -89 -355
rect -147 -423 -135 -389
rect -101 -423 -89 -389
rect -147 -457 -89 -423
rect -147 -491 -135 -457
rect -101 -491 -89 -457
rect -147 -525 -89 -491
rect -147 -559 -135 -525
rect -101 -559 -89 -525
rect -147 -593 -89 -559
rect -147 -627 -135 -593
rect -101 -627 -89 -593
rect -147 -661 -89 -627
rect -147 -695 -135 -661
rect -101 -695 -89 -661
rect -147 -729 -89 -695
rect -147 -763 -135 -729
rect -101 -763 -89 -729
rect -147 -797 -89 -763
rect -147 -831 -135 -797
rect -101 -831 -89 -797
rect -147 -865 -89 -831
rect -147 -899 -135 -865
rect -101 -899 -89 -865
rect -147 -924 -89 -899
rect -29 971 29 996
rect -29 937 -17 971
rect 17 937 29 971
rect -29 903 29 937
rect -29 869 -17 903
rect 17 869 29 903
rect -29 835 29 869
rect -29 801 -17 835
rect 17 801 29 835
rect -29 767 29 801
rect -29 733 -17 767
rect 17 733 29 767
rect -29 699 29 733
rect -29 665 -17 699
rect 17 665 29 699
rect -29 631 29 665
rect -29 597 -17 631
rect 17 597 29 631
rect -29 563 29 597
rect -29 529 -17 563
rect 17 529 29 563
rect -29 495 29 529
rect -29 461 -17 495
rect 17 461 29 495
rect -29 427 29 461
rect -29 393 -17 427
rect 17 393 29 427
rect -29 359 29 393
rect -29 325 -17 359
rect 17 325 29 359
rect -29 291 29 325
rect -29 257 -17 291
rect 17 257 29 291
rect -29 223 29 257
rect -29 189 -17 223
rect 17 189 29 223
rect -29 155 29 189
rect -29 121 -17 155
rect 17 121 29 155
rect -29 87 29 121
rect -29 53 -17 87
rect 17 53 29 87
rect -29 19 29 53
rect -29 -15 -17 19
rect 17 -15 29 19
rect -29 -49 29 -15
rect -29 -83 -17 -49
rect 17 -83 29 -49
rect -29 -117 29 -83
rect -29 -151 -17 -117
rect 17 -151 29 -117
rect -29 -185 29 -151
rect -29 -219 -17 -185
rect 17 -219 29 -185
rect -29 -253 29 -219
rect -29 -287 -17 -253
rect 17 -287 29 -253
rect -29 -321 29 -287
rect -29 -355 -17 -321
rect 17 -355 29 -321
rect -29 -389 29 -355
rect -29 -423 -17 -389
rect 17 -423 29 -389
rect -29 -457 29 -423
rect -29 -491 -17 -457
rect 17 -491 29 -457
rect -29 -525 29 -491
rect -29 -559 -17 -525
rect 17 -559 29 -525
rect -29 -593 29 -559
rect -29 -627 -17 -593
rect 17 -627 29 -593
rect -29 -661 29 -627
rect -29 -695 -17 -661
rect 17 -695 29 -661
rect -29 -729 29 -695
rect -29 -763 -17 -729
rect 17 -763 29 -729
rect -29 -797 29 -763
rect -29 -831 -17 -797
rect 17 -831 29 -797
rect -29 -865 29 -831
rect -29 -899 -17 -865
rect 17 -899 29 -865
rect -29 -924 29 -899
rect 89 971 147 996
rect 89 937 101 971
rect 135 937 147 971
rect 89 903 147 937
rect 89 869 101 903
rect 135 869 147 903
rect 89 835 147 869
rect 89 801 101 835
rect 135 801 147 835
rect 89 767 147 801
rect 89 733 101 767
rect 135 733 147 767
rect 89 699 147 733
rect 89 665 101 699
rect 135 665 147 699
rect 89 631 147 665
rect 89 597 101 631
rect 135 597 147 631
rect 89 563 147 597
rect 89 529 101 563
rect 135 529 147 563
rect 89 495 147 529
rect 89 461 101 495
rect 135 461 147 495
rect 89 427 147 461
rect 89 393 101 427
rect 135 393 147 427
rect 89 359 147 393
rect 89 325 101 359
rect 135 325 147 359
rect 89 291 147 325
rect 89 257 101 291
rect 135 257 147 291
rect 89 223 147 257
rect 89 189 101 223
rect 135 189 147 223
rect 89 155 147 189
rect 89 121 101 155
rect 135 121 147 155
rect 89 87 147 121
rect 89 53 101 87
rect 135 53 147 87
rect 89 19 147 53
rect 89 -15 101 19
rect 135 -15 147 19
rect 89 -49 147 -15
rect 89 -83 101 -49
rect 135 -83 147 -49
rect 89 -117 147 -83
rect 89 -151 101 -117
rect 135 -151 147 -117
rect 89 -185 147 -151
rect 89 -219 101 -185
rect 135 -219 147 -185
rect 89 -253 147 -219
rect 89 -287 101 -253
rect 135 -287 147 -253
rect 89 -321 147 -287
rect 89 -355 101 -321
rect 135 -355 147 -321
rect 89 -389 147 -355
rect 89 -423 101 -389
rect 135 -423 147 -389
rect 89 -457 147 -423
rect 89 -491 101 -457
rect 135 -491 147 -457
rect 89 -525 147 -491
rect 89 -559 101 -525
rect 135 -559 147 -525
rect 89 -593 147 -559
rect 89 -627 101 -593
rect 135 -627 147 -593
rect 89 -661 147 -627
rect 89 -695 101 -661
rect 135 -695 147 -661
rect 89 -729 147 -695
rect 89 -763 101 -729
rect 135 -763 147 -729
rect 89 -797 147 -763
rect 89 -831 101 -797
rect 135 -831 147 -797
rect 89 -865 147 -831
rect 89 -899 101 -865
rect 135 -899 147 -865
rect 89 -924 147 -899
<< pdiffc >>
rect -135 937 -101 971
rect -135 869 -101 903
rect -135 801 -101 835
rect -135 733 -101 767
rect -135 665 -101 699
rect -135 597 -101 631
rect -135 529 -101 563
rect -135 461 -101 495
rect -135 393 -101 427
rect -135 325 -101 359
rect -135 257 -101 291
rect -135 189 -101 223
rect -135 121 -101 155
rect -135 53 -101 87
rect -135 -15 -101 19
rect -135 -83 -101 -49
rect -135 -151 -101 -117
rect -135 -219 -101 -185
rect -135 -287 -101 -253
rect -135 -355 -101 -321
rect -135 -423 -101 -389
rect -135 -491 -101 -457
rect -135 -559 -101 -525
rect -135 -627 -101 -593
rect -135 -695 -101 -661
rect -135 -763 -101 -729
rect -135 -831 -101 -797
rect -135 -899 -101 -865
rect -17 937 17 971
rect -17 869 17 903
rect -17 801 17 835
rect -17 733 17 767
rect -17 665 17 699
rect -17 597 17 631
rect -17 529 17 563
rect -17 461 17 495
rect -17 393 17 427
rect -17 325 17 359
rect -17 257 17 291
rect -17 189 17 223
rect -17 121 17 155
rect -17 53 17 87
rect -17 -15 17 19
rect -17 -83 17 -49
rect -17 -151 17 -117
rect -17 -219 17 -185
rect -17 -287 17 -253
rect -17 -355 17 -321
rect -17 -423 17 -389
rect -17 -491 17 -457
rect -17 -559 17 -525
rect -17 -627 17 -593
rect -17 -695 17 -661
rect -17 -763 17 -729
rect -17 -831 17 -797
rect -17 -899 17 -865
rect 101 937 135 971
rect 101 869 135 903
rect 101 801 135 835
rect 101 733 135 767
rect 101 665 135 699
rect 101 597 135 631
rect 101 529 135 563
rect 101 461 135 495
rect 101 393 135 427
rect 101 325 135 359
rect 101 257 135 291
rect 101 189 135 223
rect 101 121 135 155
rect 101 53 135 87
rect 101 -15 135 19
rect 101 -83 135 -49
rect 101 -151 135 -117
rect 101 -219 135 -185
rect 101 -287 135 -253
rect 101 -355 135 -321
rect 101 -423 135 -389
rect 101 -491 135 -457
rect 101 -559 135 -525
rect 101 -627 135 -593
rect 101 -695 135 -661
rect 101 -763 135 -729
rect 101 -831 135 -797
rect 101 -899 135 -865
<< poly >>
rect -89 1011 89 1056
rect -89 996 -29 1011
rect 29 996 89 1011
rect -89 -955 -29 -924
rect 29 -955 89 -924
rect -92 -971 -26 -955
rect -92 -1005 -76 -971
rect -42 -1005 -26 -971
rect -92 -1021 -26 -1005
rect 26 -971 92 -955
rect 26 -1005 42 -971
rect 76 -1005 92 -971
rect 26 -1021 92 -1005
<< polycont >>
rect -76 -1005 -42 -971
rect 42 -1005 76 -971
<< locali >>
rect -135 971 -101 1000
rect -135 903 -101 919
rect -135 835 -101 847
rect -135 767 -101 775
rect -135 699 -101 703
rect -135 593 -101 597
rect -135 521 -101 529
rect -135 449 -101 461
rect -135 377 -101 393
rect -135 305 -101 325
rect -135 233 -101 257
rect -135 161 -101 189
rect -135 89 -101 121
rect -135 19 -101 53
rect -135 -49 -101 -17
rect -135 -117 -101 -89
rect -135 -185 -101 -161
rect -135 -253 -101 -233
rect -135 -321 -101 -305
rect -135 -389 -101 -377
rect -135 -457 -101 -449
rect -135 -525 -101 -521
rect -135 -631 -101 -627
rect -135 -703 -101 -695
rect -135 -775 -101 -763
rect -135 -847 -101 -831
rect -135 -928 -101 -899
rect -17 971 17 1000
rect -17 903 17 919
rect -17 835 17 847
rect -17 767 17 775
rect -17 699 17 703
rect -17 593 17 597
rect -17 521 17 529
rect -17 449 17 461
rect -17 377 17 393
rect -17 305 17 325
rect -17 233 17 257
rect -17 161 17 189
rect -17 89 17 121
rect -17 19 17 53
rect -17 -49 17 -17
rect -17 -117 17 -89
rect -17 -185 17 -161
rect -17 -253 17 -233
rect -17 -321 17 -305
rect -17 -389 17 -377
rect -17 -457 17 -449
rect -17 -525 17 -521
rect -17 -631 17 -627
rect -17 -703 17 -695
rect -17 -775 17 -763
rect -17 -847 17 -831
rect -17 -928 17 -899
rect 101 971 135 1000
rect 101 903 135 919
rect 101 835 135 847
rect 101 767 135 775
rect 101 699 135 703
rect 101 593 135 597
rect 101 521 135 529
rect 101 449 135 461
rect 101 377 135 393
rect 101 305 135 325
rect 101 233 135 257
rect 101 161 135 189
rect 101 89 135 121
rect 101 19 135 53
rect 101 -49 135 -17
rect 101 -117 135 -89
rect 101 -185 135 -161
rect 101 -253 135 -233
rect 101 -321 135 -305
rect 101 -389 135 -377
rect 101 -457 135 -449
rect 101 -525 135 -521
rect 101 -631 135 -627
rect 101 -703 135 -695
rect 101 -775 135 -763
rect 101 -847 135 -831
rect 101 -928 135 -899
rect -92 -1005 -76 -971
rect -42 -1005 -26 -971
rect 26 -1005 42 -971
rect 76 -1005 92 -971
<< viali >>
rect -135 937 -101 953
rect -135 919 -101 937
rect -135 869 -101 881
rect -135 847 -101 869
rect -135 801 -101 809
rect -135 775 -101 801
rect -135 733 -101 737
rect -135 703 -101 733
rect -135 631 -101 665
rect -135 563 -101 593
rect -135 559 -101 563
rect -135 495 -101 521
rect -135 487 -101 495
rect -135 427 -101 449
rect -135 415 -101 427
rect -135 359 -101 377
rect -135 343 -101 359
rect -135 291 -101 305
rect -135 271 -101 291
rect -135 223 -101 233
rect -135 199 -101 223
rect -135 155 -101 161
rect -135 127 -101 155
rect -135 87 -101 89
rect -135 55 -101 87
rect -135 -15 -101 17
rect -135 -17 -101 -15
rect -135 -83 -101 -55
rect -135 -89 -101 -83
rect -135 -151 -101 -127
rect -135 -161 -101 -151
rect -135 -219 -101 -199
rect -135 -233 -101 -219
rect -135 -287 -101 -271
rect -135 -305 -101 -287
rect -135 -355 -101 -343
rect -135 -377 -101 -355
rect -135 -423 -101 -415
rect -135 -449 -101 -423
rect -135 -491 -101 -487
rect -135 -521 -101 -491
rect -135 -593 -101 -559
rect -135 -661 -101 -631
rect -135 -665 -101 -661
rect -135 -729 -101 -703
rect -135 -737 -101 -729
rect -135 -797 -101 -775
rect -135 -809 -101 -797
rect -135 -865 -101 -847
rect -135 -881 -101 -865
rect -17 937 17 953
rect -17 919 17 937
rect -17 869 17 881
rect -17 847 17 869
rect -17 801 17 809
rect -17 775 17 801
rect -17 733 17 737
rect -17 703 17 733
rect -17 631 17 665
rect -17 563 17 593
rect -17 559 17 563
rect -17 495 17 521
rect -17 487 17 495
rect -17 427 17 449
rect -17 415 17 427
rect -17 359 17 377
rect -17 343 17 359
rect -17 291 17 305
rect -17 271 17 291
rect -17 223 17 233
rect -17 199 17 223
rect -17 155 17 161
rect -17 127 17 155
rect -17 87 17 89
rect -17 55 17 87
rect -17 -15 17 17
rect -17 -17 17 -15
rect -17 -83 17 -55
rect -17 -89 17 -83
rect -17 -151 17 -127
rect -17 -161 17 -151
rect -17 -219 17 -199
rect -17 -233 17 -219
rect -17 -287 17 -271
rect -17 -305 17 -287
rect -17 -355 17 -343
rect -17 -377 17 -355
rect -17 -423 17 -415
rect -17 -449 17 -423
rect -17 -491 17 -487
rect -17 -521 17 -491
rect -17 -593 17 -559
rect -17 -661 17 -631
rect -17 -665 17 -661
rect -17 -729 17 -703
rect -17 -737 17 -729
rect -17 -797 17 -775
rect -17 -809 17 -797
rect -17 -865 17 -847
rect -17 -881 17 -865
rect 101 937 135 953
rect 101 919 135 937
rect 101 869 135 881
rect 101 847 135 869
rect 101 801 135 809
rect 101 775 135 801
rect 101 733 135 737
rect 101 703 135 733
rect 101 631 135 665
rect 101 563 135 593
rect 101 559 135 563
rect 101 495 135 521
rect 101 487 135 495
rect 101 427 135 449
rect 101 415 135 427
rect 101 359 135 377
rect 101 343 135 359
rect 101 291 135 305
rect 101 271 135 291
rect 101 223 135 233
rect 101 199 135 223
rect 101 155 135 161
rect 101 127 135 155
rect 101 87 135 89
rect 101 55 135 87
rect 101 -15 135 17
rect 101 -17 135 -15
rect 101 -83 135 -55
rect 101 -89 135 -83
rect 101 -151 135 -127
rect 101 -161 135 -151
rect 101 -219 135 -199
rect 101 -233 135 -219
rect 101 -287 135 -271
rect 101 -305 135 -287
rect 101 -355 135 -343
rect 101 -377 135 -355
rect 101 -423 135 -415
rect 101 -449 135 -423
rect 101 -491 135 -487
rect 101 -521 135 -491
rect 101 -593 135 -559
rect 101 -661 135 -631
rect 101 -665 135 -661
rect 101 -729 135 -703
rect 101 -737 135 -729
rect 101 -797 135 -775
rect 101 -809 135 -797
rect 101 -865 135 -847
rect 101 -881 135 -865
rect -76 -1005 -42 -971
rect 42 -1005 76 -971
<< metal1 >>
rect -141 953 -95 996
rect -141 919 -135 953
rect -101 919 -95 953
rect -141 881 -95 919
rect -141 847 -135 881
rect -101 847 -95 881
rect -141 809 -95 847
rect -141 775 -135 809
rect -101 775 -95 809
rect -141 737 -95 775
rect -141 703 -135 737
rect -101 703 -95 737
rect -141 665 -95 703
rect -141 631 -135 665
rect -101 631 -95 665
rect -141 593 -95 631
rect -141 559 -135 593
rect -101 559 -95 593
rect -141 521 -95 559
rect -141 487 -135 521
rect -101 487 -95 521
rect -141 449 -95 487
rect -141 415 -135 449
rect -101 415 -95 449
rect -141 377 -95 415
rect -141 343 -135 377
rect -101 343 -95 377
rect -141 305 -95 343
rect -141 271 -135 305
rect -101 271 -95 305
rect -141 233 -95 271
rect -141 199 -135 233
rect -101 199 -95 233
rect -141 161 -95 199
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -199 -95 -161
rect -141 -233 -135 -199
rect -101 -233 -95 -199
rect -141 -271 -95 -233
rect -141 -305 -135 -271
rect -101 -305 -95 -271
rect -141 -343 -95 -305
rect -141 -377 -135 -343
rect -101 -377 -95 -343
rect -141 -415 -95 -377
rect -141 -449 -135 -415
rect -101 -449 -95 -415
rect -141 -487 -95 -449
rect -141 -521 -135 -487
rect -101 -521 -95 -487
rect -141 -559 -95 -521
rect -141 -593 -135 -559
rect -101 -593 -95 -559
rect -141 -631 -95 -593
rect -141 -665 -135 -631
rect -101 -665 -95 -631
rect -141 -703 -95 -665
rect -141 -737 -135 -703
rect -101 -737 -95 -703
rect -141 -775 -95 -737
rect -141 -809 -135 -775
rect -101 -809 -95 -775
rect -141 -847 -95 -809
rect -141 -881 -135 -847
rect -101 -881 -95 -847
rect -141 -924 -95 -881
rect -23 953 23 996
rect -23 919 -17 953
rect 17 919 23 953
rect -23 881 23 919
rect -23 847 -17 881
rect 17 847 23 881
rect -23 809 23 847
rect -23 775 -17 809
rect 17 775 23 809
rect -23 737 23 775
rect -23 703 -17 737
rect 17 703 23 737
rect -23 665 23 703
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -703 23 -665
rect -23 -737 -17 -703
rect 17 -737 23 -703
rect -23 -775 23 -737
rect -23 -809 -17 -775
rect 17 -809 23 -775
rect -23 -847 23 -809
rect -23 -881 -17 -847
rect 17 -881 23 -847
rect -23 -924 23 -881
rect 95 953 141 996
rect 95 919 101 953
rect 135 919 141 953
rect 95 881 141 919
rect 95 847 101 881
rect 135 847 141 881
rect 95 809 141 847
rect 95 775 101 809
rect 135 775 141 809
rect 95 737 141 775
rect 95 703 101 737
rect 135 703 141 737
rect 95 665 141 703
rect 95 631 101 665
rect 135 631 141 665
rect 95 593 141 631
rect 95 559 101 593
rect 135 559 141 593
rect 95 521 141 559
rect 95 487 101 521
rect 135 487 141 521
rect 95 449 141 487
rect 95 415 101 449
rect 135 415 141 449
rect 95 377 141 415
rect 95 343 101 377
rect 135 343 141 377
rect 95 305 141 343
rect 95 271 101 305
rect 135 271 141 305
rect 95 233 141 271
rect 95 199 101 233
rect 135 199 141 233
rect 95 161 141 199
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -199 141 -161
rect 95 -233 101 -199
rect 135 -233 141 -199
rect 95 -271 141 -233
rect 95 -305 101 -271
rect 135 -305 141 -271
rect 95 -343 141 -305
rect 95 -377 101 -343
rect 135 -377 141 -343
rect 95 -415 141 -377
rect 95 -449 101 -415
rect 135 -449 141 -415
rect 95 -487 141 -449
rect 95 -521 101 -487
rect 135 -521 141 -487
rect 95 -559 141 -521
rect 95 -593 101 -559
rect 135 -593 141 -559
rect 95 -631 141 -593
rect 95 -665 101 -631
rect 135 -665 141 -631
rect 95 -703 141 -665
rect 95 -737 101 -703
rect 135 -737 141 -703
rect 95 -775 141 -737
rect 95 -809 101 -775
rect 135 -809 141 -775
rect 95 -847 141 -809
rect 95 -881 101 -847
rect 135 -881 141 -847
rect 95 -924 141 -881
rect -88 -971 -30 -965
rect -88 -1005 -76 -971
rect -42 -1005 -30 -971
rect -88 -1011 -30 -1005
rect 30 -971 88 -965
rect 30 -1005 42 -971
rect 76 -1005 88 -971
rect 30 -1011 88 -1005
<< end >>
