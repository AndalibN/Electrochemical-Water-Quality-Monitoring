magic
tech sky130A
magscale 1 2
timestamp 1669522153
<< pwell >>
rect -424 2444 -120 3856
<< psubdiff >>
rect -398 3779 -146 3830
rect -398 2521 -391 3779
rect -153 2521 -146 3779
rect -398 2470 -146 2521
<< psubdiffcont >>
rect -391 2521 -153 3779
<< locali >>
rect -398 3779 -146 3822
rect -398 2521 -391 3779
rect -153 2521 -146 3779
rect -398 2478 -146 2521
use sky130_fd_pr__res_xhigh_po_0p35_57VM9D  sky130_fd_pr__res_xhigh_po_0p35_57VM9D_0
timestamp 1669522153
transform 1 0 37 0 1 2889
box -35 -2889 35 2889
<< labels >>
rlabel locali s -302 3098 -302 3098 4 gnd
port 1 nsew
<< end >>
