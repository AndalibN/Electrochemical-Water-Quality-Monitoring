magic
tech sky130A
magscale 1 2
timestamp 1667254537
<< error_p >>
rect -274 1331 -216 1337
rect -78 1331 -20 1337
rect 118 1331 176 1337
rect 314 1331 372 1337
rect -274 1297 -262 1331
rect -78 1297 -66 1331
rect 118 1297 130 1331
rect 314 1297 326 1331
rect -274 1291 -216 1297
rect -78 1291 -20 1297
rect 118 1291 176 1297
rect 314 1291 372 1297
rect -372 -1297 -314 -1291
rect -176 -1297 -118 -1291
rect 20 -1297 78 -1291
rect 216 -1297 274 -1291
rect -372 -1331 -360 -1297
rect -176 -1331 -164 -1297
rect 20 -1331 32 -1297
rect 216 -1331 228 -1297
rect -372 -1337 -314 -1331
rect -176 -1337 -118 -1331
rect 20 -1337 78 -1331
rect 216 -1337 274 -1331
<< nwell >>
rect -359 1312 457 1350
rect -457 -1312 457 1312
rect -457 -1350 359 -1312
<< pmos >>
rect -363 -1250 -323 1250
rect -265 -1250 -225 1250
rect -167 -1250 -127 1250
rect -69 -1250 -29 1250
rect 29 -1250 69 1250
rect 127 -1250 167 1250
rect 225 -1250 265 1250
rect 323 -1250 363 1250
<< pdiff >>
rect -421 1238 -363 1250
rect -421 -1238 -409 1238
rect -375 -1238 -363 1238
rect -421 -1250 -363 -1238
rect -323 1238 -265 1250
rect -323 -1238 -311 1238
rect -277 -1238 -265 1238
rect -323 -1250 -265 -1238
rect -225 1238 -167 1250
rect -225 -1238 -213 1238
rect -179 -1238 -167 1238
rect -225 -1250 -167 -1238
rect -127 1238 -69 1250
rect -127 -1238 -115 1238
rect -81 -1238 -69 1238
rect -127 -1250 -69 -1238
rect -29 1238 29 1250
rect -29 -1238 -17 1238
rect 17 -1238 29 1238
rect -29 -1250 29 -1238
rect 69 1238 127 1250
rect 69 -1238 81 1238
rect 115 -1238 127 1238
rect 69 -1250 127 -1238
rect 167 1238 225 1250
rect 167 -1238 179 1238
rect 213 -1238 225 1238
rect 167 -1250 225 -1238
rect 265 1238 323 1250
rect 265 -1238 277 1238
rect 311 -1238 323 1238
rect 265 -1250 323 -1238
rect 363 1238 421 1250
rect 363 -1238 375 1238
rect 409 -1238 421 1238
rect 363 -1250 421 -1238
<< pdiffc >>
rect -409 -1238 -375 1238
rect -311 -1238 -277 1238
rect -213 -1238 -179 1238
rect -115 -1238 -81 1238
rect -17 -1238 17 1238
rect 81 -1238 115 1238
rect 179 -1238 213 1238
rect 277 -1238 311 1238
rect 375 -1238 409 1238
<< poly >>
rect -278 1331 -212 1347
rect -278 1297 -262 1331
rect -228 1297 -212 1331
rect -278 1281 -212 1297
rect -82 1331 -16 1347
rect -82 1297 -66 1331
rect -32 1297 -16 1331
rect -82 1281 -16 1297
rect 114 1331 180 1347
rect 114 1297 130 1331
rect 164 1297 180 1331
rect 114 1281 180 1297
rect 310 1331 376 1347
rect 310 1297 326 1331
rect 360 1297 376 1331
rect 310 1281 376 1297
rect -363 1250 -323 1276
rect -265 1250 -225 1281
rect -167 1250 -127 1276
rect -69 1250 -29 1281
rect 29 1250 69 1276
rect 127 1250 167 1281
rect 225 1250 265 1276
rect 323 1250 363 1281
rect -363 -1281 -323 -1250
rect -265 -1276 -225 -1250
rect -167 -1281 -127 -1250
rect -69 -1276 -29 -1250
rect 29 -1281 69 -1250
rect 127 -1276 167 -1250
rect 225 -1281 265 -1250
rect 323 -1276 363 -1250
rect -376 -1297 -310 -1281
rect -376 -1331 -360 -1297
rect -326 -1331 -310 -1297
rect -376 -1347 -310 -1331
rect -180 -1297 -114 -1281
rect -180 -1331 -164 -1297
rect -130 -1331 -114 -1297
rect -180 -1347 -114 -1331
rect 16 -1297 82 -1281
rect 16 -1331 32 -1297
rect 66 -1331 82 -1297
rect 16 -1347 82 -1331
rect 212 -1297 278 -1281
rect 212 -1331 228 -1297
rect 262 -1331 278 -1297
rect 212 -1347 278 -1331
<< polycont >>
rect -262 1297 -228 1331
rect -66 1297 -32 1331
rect 130 1297 164 1331
rect 326 1297 360 1331
rect -360 -1331 -326 -1297
rect -164 -1331 -130 -1297
rect 32 -1331 66 -1297
rect 228 -1331 262 -1297
<< locali >>
rect -278 1297 -262 1331
rect -228 1297 -212 1331
rect -82 1297 -66 1331
rect -32 1297 -16 1331
rect 114 1297 130 1331
rect 164 1297 180 1331
rect 310 1297 326 1331
rect 360 1297 376 1331
rect -409 1238 -375 1254
rect -409 -1254 -375 -1238
rect -311 1238 -277 1254
rect -311 -1254 -277 -1238
rect -213 1238 -179 1254
rect -213 -1254 -179 -1238
rect -115 1238 -81 1254
rect -115 -1254 -81 -1238
rect -17 1238 17 1254
rect -17 -1254 17 -1238
rect 81 1238 115 1254
rect 81 -1254 115 -1238
rect 179 1238 213 1254
rect 179 -1254 213 -1238
rect 277 1238 311 1254
rect 277 -1254 311 -1238
rect 375 1238 409 1254
rect 375 -1254 409 -1238
rect -376 -1331 -360 -1297
rect -326 -1331 -310 -1297
rect -180 -1331 -164 -1297
rect -130 -1331 -114 -1297
rect 16 -1331 32 -1297
rect 66 -1331 82 -1297
rect 212 -1331 228 -1297
rect 262 -1331 278 -1297
<< viali >>
rect -262 1297 -228 1331
rect -66 1297 -32 1331
rect 130 1297 164 1331
rect 326 1297 360 1331
rect -409 -1238 -375 1238
rect -311 -1238 -277 1238
rect -213 -1238 -179 1238
rect -115 -1238 -81 1238
rect -17 -1238 17 1238
rect 81 -1238 115 1238
rect 179 -1238 213 1238
rect 277 -1238 311 1238
rect 375 -1238 409 1238
rect -360 -1331 -326 -1297
rect -164 -1331 -130 -1297
rect 32 -1331 66 -1297
rect 228 -1331 262 -1297
<< metal1 >>
rect -274 1331 -216 1337
rect -274 1297 -262 1331
rect -228 1297 -216 1331
rect -274 1291 -216 1297
rect -78 1331 -20 1337
rect -78 1297 -66 1331
rect -32 1297 -20 1331
rect -78 1291 -20 1297
rect 118 1331 176 1337
rect 118 1297 130 1331
rect 164 1297 176 1331
rect 118 1291 176 1297
rect 314 1331 372 1337
rect 314 1297 326 1331
rect 360 1297 372 1331
rect 314 1291 372 1297
rect -415 1238 -369 1250
rect -415 -1238 -409 1238
rect -375 -1238 -369 1238
rect -415 -1250 -369 -1238
rect -317 1238 -271 1250
rect -317 -1238 -311 1238
rect -277 -1238 -271 1238
rect -317 -1250 -271 -1238
rect -219 1238 -173 1250
rect -219 -1238 -213 1238
rect -179 -1238 -173 1238
rect -219 -1250 -173 -1238
rect -121 1238 -75 1250
rect -121 -1238 -115 1238
rect -81 -1238 -75 1238
rect -121 -1250 -75 -1238
rect -23 1238 23 1250
rect -23 -1238 -17 1238
rect 17 -1238 23 1238
rect -23 -1250 23 -1238
rect 75 1238 121 1250
rect 75 -1238 81 1238
rect 115 -1238 121 1238
rect 75 -1250 121 -1238
rect 173 1238 219 1250
rect 173 -1238 179 1238
rect 213 -1238 219 1238
rect 173 -1250 219 -1238
rect 271 1238 317 1250
rect 271 -1238 277 1238
rect 311 -1238 317 1238
rect 271 -1250 317 -1238
rect 369 1238 415 1250
rect 369 -1238 375 1238
rect 409 -1238 415 1238
rect 369 -1250 415 -1238
rect -372 -1297 -314 -1291
rect -372 -1331 -360 -1297
rect -326 -1331 -314 -1297
rect -372 -1337 -314 -1331
rect -176 -1297 -118 -1291
rect -176 -1331 -164 -1297
rect -130 -1331 -118 -1297
rect -176 -1337 -118 -1331
rect 20 -1297 78 -1291
rect 20 -1331 32 -1297
rect 66 -1331 78 -1297
rect 20 -1337 78 -1331
rect 216 -1297 274 -1291
rect 216 -1331 228 -1297
rect 262 -1331 274 -1297
rect 216 -1337 274 -1331
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 12.5 l 0.2 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
