magic
tech sky130A
magscale 1 2
timestamp 1662642932
<< error_p >>
rect -31 -222 31 -216
rect -31 -256 -19 -222
rect -31 -262 31 -256
<< nwell >>
rect -129 -275 129 275
<< pmos >>
rect -35 -175 35 175
<< pdiff >>
rect -93 163 -35 175
rect -93 -163 -81 163
rect -47 -163 -35 163
rect -93 -175 -35 -163
rect 35 163 93 175
rect 35 -163 47 163
rect 81 -163 93 163
rect 35 -175 93 -163
<< pdiffc >>
rect -81 -163 -47 163
rect 47 -163 81 163
<< poly >>
rect -35 175 35 201
rect -35 -222 35 -175
rect -35 -256 -19 -222
rect 19 -256 35 -222
rect -35 -272 35 -256
<< polycont >>
rect -19 -256 19 -222
<< locali >>
rect -81 163 -47 179
rect -81 -179 -47 -163
rect 47 163 81 179
rect 47 -179 81 -163
rect -35 -256 -19 -222
rect 19 -256 35 -222
<< viali >>
rect -81 -163 -47 163
rect 47 -163 81 163
rect -19 -256 19 -222
<< metal1 >>
rect -87 163 -41 175
rect -87 -163 -81 163
rect -47 -163 -41 163
rect -87 -175 -41 -163
rect 41 163 87 175
rect 41 -163 47 163
rect 81 -163 87 163
rect 41 -175 87 -163
rect -31 -222 31 -216
rect -31 -256 -19 -222
rect 19 -256 31 -222
rect -31 -262 31 -256
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.75 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
