magic
tech sky130A
magscale 1 2
timestamp 1667267346
<< error_s >>
rect -7270 8160 -7006 8334
rect -8197 7885 -8139 7891
rect -8001 7885 -7943 7891
rect -7805 7885 -7747 7891
rect -7609 7885 -7551 7891
rect -7413 7885 -7355 7891
rect -8197 7851 -8185 7885
rect -8001 7851 -7989 7885
rect -7805 7851 -7793 7885
rect -7609 7851 -7597 7885
rect -7413 7851 -7401 7885
rect -8197 7845 -8139 7851
rect -8001 7845 -7943 7851
rect -7805 7845 -7747 7851
rect -7609 7845 -7551 7851
rect -7413 7845 -7355 7851
rect -8295 5757 -8237 5763
rect -8099 5757 -8041 5763
rect -7903 5757 -7845 5763
rect -7707 5757 -7649 5763
rect -7511 5757 -7453 5763
rect -8295 5723 -8283 5757
rect -8099 5723 -8087 5757
rect -7903 5723 -7891 5757
rect -7707 5723 -7695 5757
rect -7511 5723 -7499 5757
rect -8295 5717 -8237 5723
rect -8099 5717 -8041 5723
rect -7903 5717 -7845 5723
rect -7707 5717 -7649 5723
rect -7511 5717 -7453 5723
<< nwell >>
rect -8380 8180 -4280 9020
rect -8380 8160 -5640 8180
rect -8380 8080 -7270 8160
rect -8380 5700 -7260 8080
rect -6040 6600 -5640 8160
rect -5820 6100 -5640 6600
use sky130_fd_pr__nfet_01v8_8AGWK6  XM4
timestamp 1667254537
transform 1 0 -6401 0 1 6348
box -187 -1088 187 1088
use sky130_fd_pr__nfet_01v8_JTEWKG  XM5
timestamp 1667254537
transform 1 0 -6822 0 1 6354
box -108 -1088 108 1088
use sky130_fd_pr__pfet_01v8_XP5NZ5  XM6
timestamp 1667254537
transform 1 0 -5896 0 1 7700
box -144 -1100 144 1100
use sky130_fd_pr__pfet_01v8_NMFWVH  XM7
timestamp 1667254537
transform 1 0 -4975 0 1 7456
box -697 -1350 697 1350
use sky130_fd_pr__nfet_01v8_JXHLW7  XM8
timestamp 1667254537
transform 1 0 -5005 0 1 4638
box -661 -1338 661 1338
use sky130_fd_pr__pfet_01v8_SK7ZVM  XM9
timestamp 1667266911
transform 1 0 -7251 0 1 8500
box -1123 -300 1123 300
use sky130_fd_pr__nfet_01v8_69FTK7  XM10
timestamp 1667254537
transform 1 0 -6402 0 1 7888
box -258 -188 258 188
use sky130_fd_pr__cap_mim_m3_1_A5GGR2  sky130_fd_pr__cap_mim_m3_1_A5GGR2_0
timestamp 1667266911
transform 1 0 -2931 0 1 7427
box -1249 -1199 1248 1199
use sky130_fd_pr__pfet_01v8_NDY9L5  sky130_fd_pr__pfet_01v8_NDY9L5_0
timestamp 1667265963
transform 1 0 -7825 0 1 6804
box -555 -1100 555 1100
<< end >>
