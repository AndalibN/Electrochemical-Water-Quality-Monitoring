magic
tech sky130A
magscale 1 2
timestamp 1666625676
<< error_p >>
rect -353 586 -283 730
rect -35 586 35 730
rect 283 586 353 730
rect -353 -482 -283 -338
rect -35 -482 35 -338
rect 283 -482 353 -338
<< xpolycontact >>
rect -353 1118 -283 1550
rect -353 586 -283 1018
rect -35 1118 35 1550
rect -35 586 35 1018
rect 283 1118 353 1550
rect 283 586 353 1018
rect -353 50 -283 482
rect -353 -482 -283 -50
rect -35 50 35 482
rect -35 -482 35 -50
rect 283 50 353 482
rect 283 -482 353 -50
rect -353 -1018 -283 -586
rect -353 -1550 -283 -1118
rect -35 -1018 35 -586
rect -35 -1550 35 -1118
rect 283 -1018 353 -586
rect 283 -1550 353 -1118
<< xpolyres >>
rect -353 1018 -283 1118
rect -35 1018 35 1118
rect 283 1018 353 1118
rect -353 -50 -283 50
rect -35 -50 35 50
rect 283 -50 353 50
rect -353 -1118 -283 -1018
rect -35 -1118 35 -1018
rect 283 -1118 353 -1018
<< viali >>
rect -337 1135 -299 1532
rect -19 1135 19 1532
rect 299 1135 337 1532
rect -337 604 -299 1001
rect -19 604 19 1001
rect 299 604 337 1001
rect -337 67 -299 464
rect -19 67 19 464
rect 299 67 337 464
rect -337 -464 -299 -67
rect -19 -464 19 -67
rect 299 -464 337 -67
rect -337 -1001 -299 -604
rect -19 -1001 19 -604
rect 299 -1001 337 -604
rect -337 -1532 -299 -1135
rect -19 -1532 19 -1135
rect 299 -1532 337 -1135
<< metal1 >>
rect -343 1532 -293 1544
rect -343 1135 -337 1532
rect -299 1135 -293 1532
rect -343 1123 -293 1135
rect -25 1532 25 1544
rect -25 1135 -19 1532
rect 19 1135 25 1532
rect -25 1123 25 1135
rect 293 1532 343 1544
rect 293 1135 299 1532
rect 337 1135 343 1532
rect 293 1123 343 1135
rect -343 1001 -293 1013
rect -343 604 -337 1001
rect -299 604 -293 1001
rect -343 592 -293 604
rect -25 1001 25 1013
rect -25 604 -19 1001
rect 19 604 25 1001
rect -25 592 25 604
rect 293 1001 343 1013
rect 293 604 299 1001
rect 337 604 343 1001
rect 293 592 343 604
rect -343 464 -293 476
rect -343 67 -337 464
rect -299 67 -293 464
rect -343 55 -293 67
rect -25 464 25 476
rect -25 67 -19 464
rect 19 67 25 464
rect -25 55 25 67
rect 293 464 343 476
rect 293 67 299 464
rect 337 67 343 464
rect 293 55 343 67
rect -343 -67 -293 -55
rect -343 -464 -337 -67
rect -299 -464 -293 -67
rect -343 -476 -293 -464
rect -25 -67 25 -55
rect -25 -464 -19 -67
rect 19 -464 25 -67
rect -25 -476 25 -464
rect 293 -67 343 -55
rect 293 -464 299 -67
rect 337 -464 343 -67
rect 293 -476 343 -464
rect -343 -604 -293 -592
rect -343 -1001 -337 -604
rect -299 -1001 -293 -604
rect -343 -1013 -293 -1001
rect -25 -604 25 -592
rect -25 -1001 -19 -604
rect 19 -1001 25 -604
rect -25 -1013 25 -1001
rect 293 -604 343 -592
rect 293 -1001 299 -604
rect 337 -1001 343 -604
rect 293 -1013 343 -1001
rect -343 -1135 -293 -1123
rect -343 -1532 -337 -1135
rect -299 -1532 -293 -1135
rect -343 -1544 -293 -1532
rect -25 -1135 25 -1123
rect -25 -1532 -19 -1135
rect 19 -1532 25 -1135
rect -25 -1544 25 -1532
rect 293 -1135 343 -1123
rect 293 -1532 299 -1135
rect 337 -1532 343 -1135
rect 293 -1544 343 -1532
<< res0p35 >>
rect -355 1016 -281 1120
rect -37 1016 37 1120
rect 281 1016 355 1120
rect -355 -52 -281 52
rect -37 -52 37 52
rect 281 -52 355 52
rect -355 -1120 -281 -1016
rect -37 -1120 37 -1016
rect 281 -1120 355 -1016
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.5 m 3 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 3.932k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
